* NGSPICE file created from lpopamp_slice_.ext - technology: sky130A

.subckt lpopamp_slice_ im ip o avdd avss en enb bpa bpb bnb bna xp ypm ypp zpm zpp
+ xn ynm ynp znm znp vsub
X0 a_13000_n800# ip ypp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1 a_21550_n1650# bnb a_23200_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X2 ypp zpp a_22900_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X3 a_28450_5000# bpa a_28300_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X4 a_27250_n1650# znp a_27100_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X5 a_26350_4350# bpa a_26200_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X6 a_25150_3050# bpa a_25000_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X7 a_100_3050# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X8 a_18100_900# znp avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X9 a_4000_n800# en bna avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X10 ynm im xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X11 a_28150_50# znp a_28000_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X12 a_1150_n1650# bnb a_5800_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X13 a_25000_50# znp a_24850_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X14 a_8200_50# bna a_8050_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X15 a_28600_5000# bpa a_28450_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X16 a_20050_3050# bpa a_19900_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X17 a_26500_4350# bpa a_26350_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X18 a_13300_n1650# im xn avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X19 a_25300_5000# bpb a_25150_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X20 a_17200_n1650# znp a_17050_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X21 a_19900_50# znp a_19750_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X22 xp ip ynp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X23 a_23200_4350# zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X24 a_13450_3050# zpp a_13300_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X25 a_8200_3700# bpa a_8050_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X26 avdd bpa bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X27 a_4300_n1650# en a_1150_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X28 a_8200_n1650# bna a_8050_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X29 a_17650_n800# znp a_17500_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X30 a_14050_5000# zpp a_13900_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X31 a_550_3050# bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X32 avdd zpp a_11800_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X33 xn im a_14200_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X34 bna enb avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=3.5 ps=15 w=7 l=1
X35 avdd bpa bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X36 a_4450_3050# bpa a_4300_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X37 xn ip a_12400_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X38 ynm im xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X39 a_550_3050# bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X40 a_13600_3050# zpp a_13450_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X41 a_20050_n1650# znp a_19900_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X42 bpa bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X43 a_8650_n800# bna a_8500_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X44 a_550_3050# bpb a_4900_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X45 a_550_3050# bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X46 a_1150_n1650# bnb a_5200_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X47 a_550_3050# bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X48 a_17800_n800# znp a_17650_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X49 a_7900_3050# bpa a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X50 a_27850_3700# bpb znp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X51 a_14500_n800# bna xn avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X52 a_10900_5000# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X53 a_4600_3050# bpa a_4450_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X54 avdd zpp a_24400_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X55 a_11200_n800# bna a_11050_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X56 a_23500_n1650# bna a_21550_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X57 xn bna a_11800_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X58 a_27400_n1650# znp a_27250_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X59 bpb bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X60 a_21250_3700# zpp a_21100_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X61 a_23800_900# bna a_23650_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X62 zpp bnb a_22300_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X63 a_8800_n800# bna a_8650_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X64 a_21250_900# bna a_21100_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X65 a_2500_50# bnb a_1150_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X66 a_17350_50# znp a_17200_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X67 a_5500_n800# bnb a_1150_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X68 bpa enb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X69 a_2200_n800# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X70 a_4900_900# bnb a_1150_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X71 a_28000_3700# bpb a_27850_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X72 a_16000_900# znp a_15850_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X73 a_100_4350# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X74 a_1150_n1650# bnb a_2200_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X75 a_24700_3700# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X76 ypm im a_13300_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X77 a_25300_900# znp a_25150_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X78 zpp zpp a_21250_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X79 a_10150_n1650# bna a_10000_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X80 a_18250_3050# bpa a_18100_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X81 bpa en avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=2.5 ps=11 w=5 l=1
X82 a_20050_4350# bpa a_19900_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X83 ypp zpp a_20800_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X84 a_6400_900# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X85 xp im ynm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X86 a_1150_n1650# bna a_1000_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X87 a_27250_50# znp a_27100_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X88 a_17500_900# znp a_17350_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X89 xp ip ynp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X90 bnb bnb a_4900_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X91 ynm znp a_19000_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X92 a_7300_50# bna a_1150_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X93 avdd zpp a_15400_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X94 avdd bpa bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X95 a_13450_4350# zpp a_13300_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X96 a_12250_5000# zpp a_12100_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X97 avdd bpa bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X98 a_18400_3050# bpa a_18250_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X99 a_21850_n800# bnb a_21700_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X100 a_19000_50# znp a_18850_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X101 a_15100_3050# zpp ypm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X102 avdd bpa bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X103 a_250_n1650# bna a_100_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X104 a_550_3050# bpb a_6700_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X105 a_550_3050# enb bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X106 ynm im xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X107 a_4450_4350# bpa a_4300_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X108 ynm im xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X109 a_550_3050# bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X110 a_19300_n800# znp ynm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X111 a_550_3050# bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X112 a_15700_5000# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X113 a_13600_4350# zpp a_13450_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X114 bpa bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X115 a_12400_5000# zpp a_12250_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X116 bpa enb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X117 bpa bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X118 a_11650_50# bna a_11500_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X119 a_22000_n800# bnb a_21850_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X120 avss znp a_20200_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X121 a_9850_50# bna a_9700_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X122 a_24250_n1650# bna a_24100_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X123 bpa bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X124 a_7900_4350# bpa a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X125 a_28150_n1650# znp a_28000_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X126 a_6700_5000# bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X127 a_4600_4350# bpa a_4450_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X128 bpb bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X129 bpb bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X130 a_26200_3700# bpa a_25150_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X131 a_10300_n1650# bna a_10150_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X132 a_21550_n1650# bna a_21400_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X133 a_14200_n1650# im ypm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X134 a_1600_50# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X135 a_18100_n1650# znp avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X136 a_25750_3050# bpb znp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X137 a_16450_50# znp a_16300_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X138 a_20650_900# bna a_20500_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X139 avdd zpp a_22300_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X140 ypm zpp a_14800_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X141 a_1300_n1650# bnb a_1150_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X142 a_11650_3700# zpp a_11500_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X143 a_18250_4350# bpa a_18100_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X144 a_5200_n1650# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X145 a_9100_n1650# bna a_8950_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X146 znp znp a_26500_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X147 ypp zpp a_22900_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X148 a_1150_n1650# bnb a_1600_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X149 ypp zpp a_20800_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X150 a_21550_n1650# bnb a_23200_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X151 ypp ip a_12700_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X152 a_550_3050# bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X153 a_24700_900# znp avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X154 a_25900_3050# bpb a_25750_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X155 a_400_n1650# bna a_250_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X156 avdd bpa bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X157 a_17050_n1650# znp a_16900_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X158 a_550_3050# bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X159 a_250_n800# bna a_100_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X160 a_22150_900# bnb a_22000_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X161 a_22600_3050# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X162 a_26350_50# znp a_26200_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X163 a_18400_4350# bpa a_18250_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X164 a_11800_3700# zpp a_11650_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X165 ynm im xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X166 a_6400_50# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X167 a_15100_4350# zpp ypm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X168 a_5800_900# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X169 a_16900_900# znp ynp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X170 a_26800_n800# znp znp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X171 a_8050_n1650# bna a_7900_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X172 bnb bnb a_3100_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X173 xn im a_14200_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X174 a_23500_n800# bna a_21550_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X175 a_20500_n1650# bna avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X176 a_26200_900# znp a_26050_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X177 a_20200_n800# znp a_20050_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X178 a_24400_n1650# bna a_24250_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X179 bpa bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X180 a_28300_n1650# znp a_28150_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X181 a_400_n800# bna a_250_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X182 bpb bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X183 a_8200_5000# bpa a_8050_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X184 bpa enb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X185 a_7300_900# bna a_1150_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X186 a_18400_900# znp a_18250_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X187 avss bna a_10600_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X188 a_8950_50# bna a_8800_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X189 a_28000_50# znp a_27850_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X190 xp ip ynp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X191 a_25150_3050# bpa a_27100_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X192 xp ip ynp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X193 avdd zpp a_13000_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X194 a_27850_5000# bpb znp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X195 a_25750_4350# bpb znp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X196 a_28150_n800# znp a_28000_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X197 avdd zpp a_24400_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X198 a_850_50# bna a_700_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X199 avdd zpp a_22300_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X200 a_20650_50# bna a_20500_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X201 a_21250_5000# zpp a_21100_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X202 a_550_3050# bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X203 a_27400_3050# bpb a_25150_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X204 a_19900_3700# bpa xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X205 avss bna a_15400_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X206 avdd bpa a_4000_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X207 a_24100_3050# zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X208 ynp ip xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X209 a_13300_3700# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X210 a_28000_5000# bpb a_27850_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X211 a_25900_4350# bpb a_25750_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X212 a_28300_n800# znp a_28150_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X213 a_24700_5000# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X214 a_22600_4350# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X215 zpp zpp a_21250_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X216 a_12850_3050# zpp a_12700_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X217 bpb bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X218 a_4300_3700# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X219 a_21250_n1650# bna a_21100_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X220 bpa en avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=2.5 ps=11 w=5 l=1
X221 a_25150_n1650# znp a_25000_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X222 a_25450_50# znp a_25300_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X223 a_17050_n800# znp a_16900_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X224 a_21550_n1650# bna a_21400_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X225 xn im a_13600_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X226 a_5500_50# bnb a_1150_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X227 a_3850_3050# bpa a_3700_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X228 a_10450_n800# bna a_10300_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X229 avdd en bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X230 a_13000_3050# zpp a_12850_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X231 bnb bnb a_2500_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X232 a_8050_n800# bna a_7900_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X233 xn im a_13600_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X234 a_11200_n1650# bna a_11050_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X235 a_25600_900# znp a_25450_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X236 a_1150_n1650# en a_4600_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X237 a_15100_n1650# bna a_14950_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X238 bnb bnb a_1300_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X239 a_13900_n800# im xn avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X240 a_4000_3050# bpa a_3850_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X241 ypp zpp a_23800_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X242 a_10600_n800# bna a_10450_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X243 a_2200_n1650# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X244 a_6700_900# bnb a_1150_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X245 a_25150_3050# bpa a_27100_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X246 a_17800_900# znp a_17650_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X247 a_20650_3700# zpp a_20500_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X248 a_12100_50# ip xn avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X249 a_8050_50# bna a_7900_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X250 a_6100_n1650# bnb a_1150_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X251 a_550_3050# bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X252 a_1150_n1650# en a_4000_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X253 a_15250_900# bna a_15100_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X254 a_27100_900# znp a_26950_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X255 a_4900_n800# bnb a_1150_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X256 a_18100_3700# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X257 a_1600_n800# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X258 ypm im a_13900_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X259 avss znp a_17800_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X260 a_8200_900# bna a_8050_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X261 a_20800_3700# zpp a_20650_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X262 a_27400_4350# bpb a_25150_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X263 a_19300_900# znp ynm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X264 a_26200_5000# bpa a_25150_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X265 a_17650_3050# bpa a_17500_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X266 bpb bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X267 a_24100_4350# zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X268 bnb bnb a_4900_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X269 a_8950_n1650# bna a_8800_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X270 avdd zpp a_14200_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X271 bpa bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X272 a_21400_n1650# bna a_21250_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X273 a_14650_50# bna a_14500_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X274 a_25300_n1650# znp a_25150_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X275 a_18550_n800# znp a_18400_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X276 ypm zpp a_14800_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X277 a_400_900# bna a_250_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X278 avdd bpa bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X279 a_12850_4350# zpp a_12700_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X280 a_15250_n800# bna a_15100_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X281 a_11650_5000# zpp a_11500_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X282 a_550_3050# bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X283 a_17800_3050# bpa a_17650_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X284 a_14500_3050# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X285 a_11200_3050# zpp a_11050_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X286 bpb bna a_9400_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X287 a_550_3050# bpb a_4900_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X288 a_3850_4350# bpa a_3700_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X289 avdd en bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X290 bnb bnb a_6100_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X291 a_550_3050# bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X292 a_18700_n800# znp a_18550_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X293 avss bna a_24400_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X294 bpa bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X295 a_13000_4350# zpp a_12850_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X296 avdd bpa a_28600_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.5 pd=11 as=1.25 ps=5.5 w=5 l=1
X297 a_15400_n800# bna a_15250_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X298 a_4600_50# en bna avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X299 a_11800_5000# zpp a_11650_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X300 a_19450_50# znp a_19300_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X301 bpb bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X302 a_12100_n800# ip xn avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X303 a_25450_3700# bpb a_25300_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X304 a_20950_900# bna a_20800_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X305 bpa enb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X306 a_22150_3700# zpp a_22000_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X307 a_9700_n800# bna bpb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X308 a_4000_4350# bpa a_3850_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X309 a_6400_n800# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X310 bpb bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X311 bnb bnb a_1900_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X312 a_3100_n800# bnb a_1150_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X313 a_25000_900# znp a_24850_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X314 znp bpb a_25450_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X315 zpp bnb a_22300_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X316 a_22300_3700# zpp a_22150_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X317 a_11200_50# bna a_11050_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X318 xp im ynm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X319 a_9400_50# bna a_9250_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X320 a_1150_n1650# bnb a_3400_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X321 a_14650_900# bna a_14500_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X322 ypp zpp a_21700_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X323 xp ip ynp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X324 a_26500_900# znp a_26350_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X325 a_17650_4350# bpa a_17500_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X326 a_11050_3700# zpp a_10900_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X327 a_22150_n1650# bnb a_22000_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X328 xp ip ynp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X329 avdd zpp a_14200_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X330 a_26050_n800# znp a_25900_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X331 avdd zpp a_13000_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X332 ynp ip xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X333 a_22750_n800# bnb a_22600_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X334 a_7600_900# bna a_7450_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X335 a_18700_900# znp a_18550_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X336 a_21100_50# bna a_20950_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X337 a_8650_4350# bpa bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X338 xn im a_13600_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X339 a_16150_900# znp a_16000_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X340 a_550_3050# enb bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X341 a_22000_3050# zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X342 a_550_3050# bpb a_6700_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X343 a_550_3050# bpb a_4900_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X344 a_19900_5000# bpa xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X345 a_17800_4350# bpa a_17650_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X346 avdd bpa a_4000_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X347 ynp ip xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X348 a_12100_n1650# ip xn avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X349 a_14500_4350# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X350 a_13300_5000# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X351 a_11200_4350# zpp a_11050_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X352 a_22900_n800# bnb a_22750_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X353 a_9100_900# bna a_8950_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X354 a_3100_n1650# bnb a_1150_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X355 bpa bpa a_8650_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X356 a_6700_5000# bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X357 a_4900_4350# bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X358 a_4300_5000# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X359 a_23650_50# bna a_23500_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X360 bpa enb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X361 a_11050_n1650# bna a_10900_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X362 a_3700_50# en a_1150_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X363 a_18550_50# znp a_18400_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X364 a_27100_3700# bpa a_26950_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X365 a_14950_n1650# bna a_14800_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X366 a_18850_n1650# znp a_18700_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X367 bnb bnb a_1900_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X368 avdd bpa a_26500_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X369 a_1150_n1650# bnb a_5800_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X370 a_23350_3050# zpp a_23200_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X371 a_15850_3700# bpa a_15700_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X372 a_9850_n1650# bna a_9700_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X373 xp im ynm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X374 ypp zpp a_12400_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X375 a_22300_n1650# bnb a_22150_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X376 a_26200_n1650# znp a_26050_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X377 a_250_3050# bpa a_100_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X378 ynp znp a_27400_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X379 a_28450_50# znp a_28300_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X380 ypp zpp a_23800_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X381 a_10300_50# bna a_10150_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X382 ypp zpp a_21700_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X383 a_21850_900# bnb a_21700_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X384 a_24250_n800# bna a_24100_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X385 a_20650_5000# zpp a_20500_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X386 a_8500_50# bna avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X387 a_550_3050# bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X388 a_550_3050# bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X389 a_26800_3050# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X390 a_550_3050# bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X391 a_16000_3700# bpa a_15850_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X392 zpp zpp a_23350_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X393 a_12700_3700# zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X394 ynp ip xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X395 a_1150_n1650# bnb a_2800_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X396 a_20200_3050# bpa a_20050_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X397 a_18100_5000# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X398 ypm im a_13900_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X399 a_400_3050# bpa a_250_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X400 a_27700_n800# znp ynp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X401 a_25900_900# znp ynp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X402 a_22000_4350# zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X403 a_24400_n800# bna a_24250_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X404 a_21550_n1650# bnb a_23200_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X405 a_1150_n1650# bna a_1000_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X406 a_20800_5000# zpp a_20650_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X407 bpb bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X408 bpb bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X409 a_400_50# bna a_250_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X410 a_21100_n800# bna a_20950_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X411 a_20200_50# znp a_20050_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X412 a_3700_3700# bpa a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X413 ypp ip a_12700_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X414 a_7000_900# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X415 bpa bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X416 a_15100_50# bna a_14950_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X417 bna enb avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X418 bna en a_4300_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X419 avss bna a_15400_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X420 a_27400_900# znp a_27250_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X421 a_19000_n1650# znp a_18850_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X422 a_8500_900# bna avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X423 a_19600_900# znp a_19450_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X424 a_25150_3050# bpb a_28000_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X425 avss enb bna avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X426 a_10000_n1650# bna a_9850_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X427 a_22750_50# bnb a_22600_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X428 xp im ynm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X429 a_2800_50# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X430 a_17650_50# znp a_17500_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X431 avdd bpa a_28600_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.5 pd=11 as=1.25 ps=5.5 w=5 l=1
X432 avdd bpa a_26500_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X433 a_25450_5000# bpb a_25300_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X434 a_23350_4350# zpp a_23200_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X435 a_700_900# bna a_550_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X436 a_22150_5000# zpp a_22000_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X437 avdd bpa a_8200_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X438 a_28300_3050# bpa a_25150_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X439 a_250_4350# bpa a_100_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X440 a_17500_3700# bpa xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X441 a_14200_3700# zpp a_14050_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X442 a_26800_4350# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X443 znp bpb a_25450_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X444 ynp znp a_27400_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X445 xp im ynm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X446 zpp zpp a_23350_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X447 a_7600_50# bna a_7450_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X448 a_22300_5000# zpp a_22150_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X449 ypm zpp a_13600_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X450 bpa bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X451 a_20200_4350# bpa a_20050_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X452 a_400_4350# bpa a_250_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X453 avdd bpa bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X454 bpb bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X455 avss znp a_17800_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X456 a_8050_3050# bpa a_7900_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X457 a_14650_n800# bna a_14500_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X458 a_11050_5000# zpp a_10900_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X459 a_550_3050# bpa a_4600_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X460 a_11350_n800# bna a_11200_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X461 bna enb avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X462 a_550_3050# bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X463 xn bna a_11800_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X464 a_13900_3050# zpp ypm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X465 a_15850_n1650# znp a_15700_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X466 a_22750_900# bnb a_22600_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X467 bpa bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X468 a_8950_n800# bna a_8800_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X469 a_19750_n1650# znp a_19600_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X470 xn bna a_11800_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X471 a_550_3050# enb bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X472 bnb bnb a_5500_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X473 a_14200_50# im ypm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X474 a_1150_n1650# bnb a_2200_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X475 a_1150_n1650# bnb a_2800_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X476 a_14800_n800# bna a_14650_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X477 bnb bnb a_6700_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X478 bna en a_3700_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X479 bpb bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X480 a_24850_3700# bpa a_24700_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X481 a_11500_n800# bna a_11350_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X482 a_14950_900# bna a_14800_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X483 a_25150_3050# bpb a_28000_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X484 bpb bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X485 a_21550_3700# zpp zpp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X486 a_23200_n1650# bnb a_23050_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X487 a_26800_900# znp znp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X488 a_27100_n1650# znp a_26950_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X489 a_24250_900# bna a_24100_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X490 a_5800_n800# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X491 a_21850_50# bnb a_21700_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X492 a_2500_n800# bnb a_1150_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X493 a_7900_900# bna a_7750_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X494 a_19000_900# znp a_18850_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X495 a_24100_50# bna a_23950_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X496 a_1900_50# bnb a_1150_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X497 a_1150_n1650# bnb a_5200_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X498 a_25000_3700# bpa a_24850_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X499 ynp znp a_16600_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X500 a_16450_900# znp a_16300_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X501 a_28300_4350# bpa a_25150_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X502 a_28300_900# znp a_28150_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X503 a_21700_3700# zpp a_21550_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X504 a_27100_5000# bpa a_26950_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X505 xp bpa a_18400_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X506 a_26050_n1650# znp a_25900_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X507 a_15250_3050# zpp a_15100_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X508 a_9400_900# bna a_9250_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X509 xp im ynm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X510 a_19450_n800# znp a_19300_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X511 a_15850_5000# bpa a_15700_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X512 avdd bpa bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X513 ypm zpp a_13600_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X514 a_16150_n800# znp a_16000_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X515 ypp zpp a_12400_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X516 a_550_3050# enb bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X517 avdd bpa bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X518 ynm im xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X519 avss enb bna avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X520 znp znp a_26500_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X521 a_6700_50# bnb a_1150_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X522 a_15400_3050# zpp a_15250_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X523 a_16000_n1650# znp a_15850_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X524 bna enb avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X525 a_8050_4350# bpa a_7900_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X526 a_12100_3050# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X527 a_19900_n1650# znp a_19750_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X528 a_550_3050# bpb a_6700_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X529 a_550_3050# bpa a_4600_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X530 a_1150_n1650# bnb a_7000_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X531 a_550_3050# bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X532 a_19600_n800# znp a_19450_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X533 a_550_3050# bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X534 a_16000_5000# bpa a_15850_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X535 a_13900_4350# zpp ypm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X536 bpa bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X537 a_16300_n800# znp a_16150_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X538 a_7000_n1650# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X539 a_12700_5000# zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X540 bpa enb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X541 bpa bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X542 a_26350_3700# bpa a_26200_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X543 bpb bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X544 a_6700_5000# bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X545 a_11050_50# bna a_10900_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X546 a_4900_4350# bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X547 a_7300_n800# bna a_1150_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X548 a_3700_5000# bpa a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X549 a_13300_50# im xn avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X550 bpb bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X551 a_26500_3700# bpa a_26350_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X552 a_23200_3700# zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X553 a_10300_900# bna a_10150_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X554 a_25150_3050# bpb a_25900_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X555 a_23650_900# bna a_23500_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X556 a_1150_n1650# en a_4000_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X557 a_22750_3050# zpp a_22600_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X558 a_20950_50# bna a_20800_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X559 avdd zpp a_11800_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X560 xp bpa a_18400_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X561 a_23200_50# bnb a_23050_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X562 xp im ynm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X563 a_15850_50# znp a_15700_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X564 a_15250_4350# zpp a_15100_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X565 a_26950_n800# znp a_26800_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X566 a_18100_50# znp avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X567 a_1150_n1650# en a_4600_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X568 a_23650_n800# bna a_23500_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X569 a_15850_900# znp a_15700_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X570 a_27700_900# znp ynp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X571 avss znp a_20200_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X572 avdd bpa bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X573 a_550_3050# bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X574 ypp ip a_12700_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X575 a_550_n800# bna a_400_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X576 a_25150_900# znp a_25000_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X577 a_22900_3050# zpp a_22750_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X578 avdd bpa a_8200_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X579 a_550_3050# enb bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X580 ynp znp a_16600_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X581 ynm im xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X582 a_17500_5000# bpa xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X583 a_15400_4350# zpp a_15250_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X584 a_8800_900# bna a_8650_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X585 a_19900_900# znp a_19750_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X586 a_14200_5000# zpp a_14050_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X587 a_12100_4350# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X588 bna en a_3700_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X589 bnb bnb a_6100_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X590 ynp znp a_25600_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X591 a_17350_900# znp a_17200_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X592 a_23800_n800# bna a_23650_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X593 a_7750_n1650# bna a_7600_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X594 a_5800_50# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X595 a_20500_n800# bna avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X596 a_20200_n1650# znp a_20050_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X597 bpa bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X598 a_700_n800# bna a_550_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X599 a_24100_n1650# bna a_23950_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X600 bpa bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X601 bpa enb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X602 a_4900_5000# bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X603 a_100_3700# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X604 a_1000_900# bna a_850_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X605 bpb bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X606 a_20050_3700# bpa a_19900_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X607 a_23050_n1650# bnb a_22900_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X608 a_27550_3050# bpb a_27400_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X609 a_12400_50# ip ypp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X610 a_26950_n1650# znp a_26800_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X611 xp ip ynp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X612 a_24250_3050# zpp a_24100_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X613 a_13450_3700# zpp a_13300_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X614 avdd bpa bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X615 a_25150_3050# bpb a_25900_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X616 a_28450_n800# znp a_28300_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X617 a_24850_5000# bpa a_24700_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X618 a_22750_4350# zpp a_22600_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X619 a_25150_n800# znp a_25000_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X620 a_21550_5000# zpp zpp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X621 a_100_n1650# bna avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X622 a_550_3050# bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X623 znp bpb a_27550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X624 a_4450_3700# bpa a_4300_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X625 a_13000_n1650# ip ypp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X626 a_24400_3050# zpp a_24250_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X627 ynm im xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X628 bnb bnb a_3100_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X629 a_16900_n1650# znp ynp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X630 a_550_3050# bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X631 a_21100_3050# zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X632 a_13600_3700# zpp a_13450_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X633 a_22300_50# bnb a_22150_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X634 a_23050_900# bnb a_22900_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X635 bpa bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X636 a_14950_50# bna a_14800_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X637 a_28600_n800# znp a_28450_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X638 a_25000_5000# bpa a_24850_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X639 a_17200_50# znp a_17050_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X640 bpa en avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X641 a_4000_n1650# en bna avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X642 a_22900_4350# zpp a_22750_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X643 a_25300_n800# znp a_25150_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X644 a_7900_n1650# bna a_7750_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X645 a_21700_5000# zpp a_21550_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X646 a_7900_3700# bpa a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X647 a_4600_3700# bpa a_4450_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X648 a_11200_900# bna a_11050_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X649 bpb bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X650 avss bna a_24400_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X651 ypm im a_13900_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X652 avss bna a_10600_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X653 avdd en bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X654 a_24850_50# znp a_24700_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X655 a_27100_50# znp a_26950_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X656 a_4900_50# bnb a_1150_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X657 bnb bnb a_5500_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X658 a_19750_50# znp a_19600_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X659 ynp znp a_16600_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X660 a_28600_900# znp a_28450_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X661 avss enb bna avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X662 bnb bnb a_4900_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X663 a_18250_3700# bpa a_18100_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X664 a_1150_n1650# bnb a_1600_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X665 a_10900_n800# bna avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X666 a_9700_900# bna bpb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X667 a_27550_4350# bpb a_27400_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X668 ypp zpp a_20800_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X669 a_26350_5000# bpa a_26200_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X670 a_1150_n1650# bnb a_7000_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X671 a_24250_4350# zpp a_24100_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X672 a_18250_900# znp a_18100_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X673 avdd bpa bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X674 a_11500_50# bna a_11350_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X675 a_18400_3700# bpa a_18250_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X676 a_1900_n800# bnb a_1150_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X677 a_9700_50# bna bpb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X678 a_15100_3700# zpp ypm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X679 xn im a_13600_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X680 a_17650_n1650# znp a_17500_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X681 znp bpb a_27550_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X682 a_26500_5000# bpa a_26350_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X683 avdd bpa a_17800_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X684 a_24400_4350# zpp a_24250_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X685 a_23200_5000# zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X686 a_14650_3050# zpp a_14500_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X687 bpa bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X688 a_21100_4350# zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X689 a_1150_n1650# en a_4600_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X690 a_8650_n1650# bna a_8500_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X691 ypp zpp a_11200_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X692 bpa enb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X693 a_1150_n1650# bnb a_2200_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X694 bpa en avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X695 a_21100_n1650# bna a_20950_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X696 a_18850_n800# znp a_18700_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X697 a_21400_50# bna a_21250_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X698 avdd bpa bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X699 avss bna a_15400_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X700 ypm im a_13900_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X701 avdd zpp a_11800_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X702 a_16300_50# znp a_16150_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X703 a_550_3050# bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X704 ypp ip a_12100_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X705 a_550_3050# enb bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X706 a_14800_3050# zpp a_14650_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X707 a_11500_3050# zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X708 a_9850_n800# bna a_9700_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X709 avdd en bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X710 a_1150_n1650# bnb a_6400_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X711 a_550_3050# bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X712 a_19000_n800# znp a_18850_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X713 a_10600_900# bna a_10450_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X714 bnb bnb a_3100_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X715 a_15700_n800# znp avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X716 a_23950_n1650# bna a_23800_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X717 a_27850_n1650# znp a_27700_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X718 bpb bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X719 a_25750_3700# bpb znp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X720 a_12400_n800# ip ypp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X721 a_23950_900# bna a_23800_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X722 a_1150_n1650# bnb a_7000_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X723 a_23950_50# bna a_23800_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X724 bpb bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X725 avdd zpp a_22300_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X726 a_26200_50# znp a_26050_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X727 a_4000_50# en bna avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X728 a_10000_n800# bna a_9850_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X729 a_18850_50# znp a_18700_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X730 a_6700_n800# bnb a_1150_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X731 bnb bnb a_4900_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X732 a_12100_900# ip xn avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X733 a_3400_n800# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X734 a_28000_900# znp a_27850_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X735 a_100_5000# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X736 a_13900_n1650# im xn avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X737 a_25900_3700# bpb a_25750_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X738 a_25450_900# znp a_25300_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X739 a_17800_n1650# znp a_17650_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X740 a_22600_3700# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X741 xp ip ynp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X742 xp bpa a_16000_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X743 a_4900_n1650# bnb a_1150_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X744 a_1150_n1650# bnb a_6400_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X745 a_8800_n1650# bna a_8650_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X746 avss znp a_28600_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=3.5 pd=15 as=1.75 ps=7.5 w=7 l=1
X747 a_17650_900# znp a_17500_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X748 a_10600_50# bna a_10450_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X749 a_20050_5000# bpa a_19900_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X750 avdd bpa a_17800_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X751 a_8800_50# bna a_8650_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X752 xp ip ynp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X753 a_14650_4350# zpp a_14500_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X754 a_13450_5000# zpp a_13300_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X755 a_550_3050# bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X756 ypp zpp a_11200_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X757 ynp ip xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X758 a_23050_n800# bnb a_22900_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X759 avdd bpa bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X760 ynp ip xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X761 avdd bpa bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X762 ynm znp a_19000_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X763 a_550_3050# bpb a_6700_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X764 a_550_3050# bpb a_4900_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X765 bnb bnb a_1300_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X766 a_4450_5000# bpa a_4300_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X767 a_700_50# bna a_550_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X768 ynm im xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X769 a_20500_50# bna avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X770 a_550_3050# enb bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X771 a_14800_4350# zpp a_14650_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X772 a_550_3050# bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X773 a_17200_n800# znp a_17050_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X774 a_13600_5000# zpp a_13450_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X775 a_28000_n1650# znp a_27850_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X776 bpb bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X777 a_25150_3050# bpa a_27100_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X778 a_11500_4350# zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X779 a_15400_50# bna a_15250_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X780 bpa bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X781 a_250_900# bna a_100_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X782 a_7900_5000# bpa a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X783 a_4900_4350# bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X784 a_8200_n800# bna a_8050_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X785 a_4600_5000# bpa a_4450_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X786 bpb bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X787 bpb bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X788 a_27400_3700# bpb a_25150_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X789 avss bna a_10600_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X790 bnb bnb a_6100_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X791 a_23050_50# bnb a_22900_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X792 a_24100_3700# zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X793 a_14650_n1650# bna a_14500_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X794 a_25300_50# znp a_25150_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X795 a_18550_n1650# znp a_18400_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X796 avss znp a_17800_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X797 a_26950_3050# bpa a_26800_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X798 a_1150_n1650# bnb a_1600_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X799 a_23650_3050# zpp zpp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X800 bnb bnb a_5500_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X801 xp ip ynp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X802 avdd bpa a_20200_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X803 a_12850_3700# zpp a_12700_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X804 bpb bna a_9400_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X805 a_18250_5000# bpa a_18100_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X806 a_11500_900# bna a_11350_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X807 a_550_3050# bpa a_400_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X808 xp bpa a_16000_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X809 a_27850_n800# znp a_27700_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X810 a_24850_900# znp a_24700_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X811 avss bna a_24400_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X812 ypp zpp a_20800_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X813 a_850_n1650# bna a_700_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X814 a_21250_n800# bna a_21100_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X815 a_3850_3700# bpa a_3700_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X816 avdd en bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X817 a_27850_50# znp a_27700_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X818 a_23800_3050# zpp a_23650_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X819 avdd bpa bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X820 a_550_3050# bpb a_6700_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X821 a_13000_3700# zpp a_12850_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X822 ynp ip xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X823 a_7900_50# bna a_7750_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X824 a_1150_n1650# bnb a_5800_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X825 a_20500_3050# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X826 a_18400_5000# bpa a_18250_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X827 a_17050_900# znp a_16900_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X828 bpb bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X829 ynp ip xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X830 a_28000_n800# znp a_27850_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X831 avss enb bna avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X832 a_15100_5000# zpp ypm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X833 a_20950_n1650# bna a_20800_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X834 a_24700_n800# znp avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X835 a_24850_n1650# znp a_24700_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X836 a_26350_900# znp a_26200_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X837 avss znp a_28600_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=3.5 pd=15 as=1.75 ps=7.5 w=7 l=1
X838 a_21400_n800# bna a_21250_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X839 a_4000_3700# bpa a_3850_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X840 a_10000_900# bna a_9850_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X841 bpa bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X842 a_6700_4350# bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X843 bna enb avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=3.5 ps=15 w=7 l=1
X844 a_7450_900# bna a_7300_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X845 bpa enb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X846 a_18550_900# znp a_18400_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X847 a_14500_50# bna xn avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X848 a_10900_n1650# bna avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X849 a_14800_n1650# bna a_14650_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X850 a_18700_n1650# znp a_18550_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X851 a_28450_3050# bpa a_28300_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X852 a_1900_n1650# bnb a_1150_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X853 a_25150_3050# bpa a_25000_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X854 a_17650_3700# bpa a_17500_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X855 a_5800_n1650# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X856 avdd zpp a_14200_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X857 a_9700_n1650# bna bpb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X858 a_26950_4350# bpa a_26800_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X859 a_1150_n1650# bnb a_5200_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X860 a_25750_5000# bpb znp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X861 a_24400_50# bna a_24250_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X862 a_23650_4350# zpp zpp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X863 avdd zpp a_22300_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X864 a_1000_n1650# bna a_850_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X865 a_17050_50# znp a_16900_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X866 avdd bpa bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X867 avdd bpa a_20200_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X868 a_28600_3050# bpa a_28450_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X869 a_19300_50# znp ynm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X870 a_550_3050# bpa a_400_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X871 a_550_3050# bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X872 a_25300_3050# bpb a_25150_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X873 a_17800_3700# bpa a_17650_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X874 a_14500_3700# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X875 a_11200_3700# zpp a_11050_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X876 a_25900_5000# bpb a_25750_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X877 a_23800_4350# zpp a_23650_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X878 a_10900_900# bna avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X879 a_26200_n800# znp a_26050_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X880 a_25000_n1650# znp a_24850_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X881 a_22600_5000# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X882 a_14050_3050# zpp a_13900_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X883 bpa bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X884 a_20500_4350# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X885 bpb bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X886 avdd bpa bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X887 a_20200_900# znp a_20050_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X888 bpb bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X889 a_26950_50# znp a_26800_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X890 bpa enb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X891 a_7000_50# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X892 bna enb avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=3.5 ps=15 w=7 l=1
X893 a_14950_n800# bna a_14800_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X894 a_550_3050# bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X895 a_1300_900# bnb a_1150_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X896 a_11650_n800# bna a_11500_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X897 a_12400_900# ip ypp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X898 a_550_3050# bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X899 a_11650_n1650# bna a_11500_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X900 ynp znp a_25600_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X901 a_10900_3050# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X902 avss bna a_15400_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X903 a_1150_n1650# bnb a_5800_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X904 a_19450_n1650# znp a_19300_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X905 xp im ynm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X906 bnb bnb a_2500_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X907 bnb bnb a_2500_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X908 bnb bnb a_6700_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X909 a_11800_n800# bna a_11650_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X910 a_1150_n1650# bnb a_6400_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X911 avss znp a_17800_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X912 a_13600_50# im ypm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X913 a_28450_4350# bpa a_28300_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X914 bpa enb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X915 ypp zpp a_21700_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X916 a_25150_3050# bpa a_27100_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X917 a_25150_3050# bpa a_25000_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X918 a_27250_900# znp a_27100_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X919 ynp ip xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X920 a_2800_n800# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X921 avss bna a_8200_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X922 a_19450_900# znp a_19300_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X923 a_28600_4350# bpa a_28450_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X924 bna en a_4300_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X925 a_22000_3700# zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X926 a_27400_5000# bpb a_25150_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X927 xp im ynm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X928 a_25300_4350# bpb a_25150_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X929 a_23500_50# bna a_21550_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X930 a_24100_5000# zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X931 avdd zpp a_15400_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X932 a_21850_n1650# bnb a_21700_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X933 ynp znp a_25600_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X934 a_18400_50# znp a_18250_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X935 a_12250_3050# zpp a_12100_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X936 a_550_900# bna a_400_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X937 a_19750_n800# znp a_19600_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X938 avdd bpa bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X939 a_14050_4350# zpp a_13900_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X940 a_16450_n800# znp a_16300_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X941 a_12850_5000# zpp a_12700_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X942 a_550_3050# enb bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X943 avdd bpa bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X944 xn ip a_13000_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X945 ynm im xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X946 a_550_3050# bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X947 a_15700_3050# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X948 avss enb bna avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X949 a_11800_n1650# bna a_11650_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X950 a_12400_3050# zpp a_12250_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X951 a_15700_n1650# znp avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X952 a_26050_50# znp a_25900_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X953 a_9250_50# bna a_9100_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X954 a_550_3050# bpb a_4900_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X955 a_7450_n800# bna a_7300_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X956 a_3850_5000# bpa a_3700_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X957 a_19900_n800# znp a_19750_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X958 a_19600_n1650# znp a_19450_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X959 a_28300_50# znp a_28150_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X960 avdd en bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X961 a_550_3050# bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X962 a_1150_n1650# en a_4000_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X963 bpa bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X964 a_16600_n800# znp a_16450_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X965 a_13000_5000# zpp a_12850_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X966 a_2800_n1650# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X967 bpb bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X968 a_10900_4350# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X969 avdd bpa a_26500_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X970 a_13300_n800# im xn avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X971 a_6700_n1650# bnb a_1150_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X972 bpb bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X973 a_23350_3700# zpp a_23200_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X974 a_11800_900# bna a_11650_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X975 a_250_3700# bpa a_100_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X976 a_7600_n800# bna a_7450_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X977 a_4000_5000# bpa a_3850_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X978 a_21100_900# bna a_20950_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X979 bpa enb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X980 a_4300_n800# en a_1150_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X981 a_26800_3700# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X982 a_12700_50# ip xn avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X983 zpp zpp a_23350_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X984 a_2200_900# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X985 a_20200_3700# bpa a_20050_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X986 a_13300_900# im xn avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X987 a_22000_n1650# bnb a_21850_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X988 a_400_3700# bpa a_250_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X989 a_25900_n1650# znp ynp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X990 znp znp a_26500_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X991 ypp zpp a_22900_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X992 xp im ynm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X993 a_17650_5000# bpa a_17500_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X994 avdd zpp a_15400_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X995 avdd zpp a_14200_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X996 a_1150_n1650# bnb a_3400_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X997 a_12250_4350# zpp a_12100_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X998 a_7750_900# bna a_7600_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X999 a_23950_n800# bna a_23800_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1000 a_18850_900# znp a_18700_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1001 a_22600_50# bnb zpp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1002 ynm im xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1003 a_20650_n800# bna a_20500_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1004 avdd bpa bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1005 a_850_n800# bna a_700_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1006 a_17500_50# znp a_17350_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1007 a_28150_900# znp a_28000_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1008 a_8650_5000# bpa bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1009 a_550_3050# enb bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1010 ynm im xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1011 xn ip a_12400_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1012 a_550_3050# bpb a_4900_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1013 a_550_3050# bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1014 a_17800_5000# bpa a_17650_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1015 a_16450_n1650# znp a_16300_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1016 a_15700_4350# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1017 a_18100_n800# znp avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1018 a_14500_5000# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1019 a_8200_3050# bpa a_8050_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1020 a_12400_4350# zpp a_12250_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1021 a_9250_900# bna a_9100_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1022 a_25150_3050# bpb a_28000_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1023 a_11200_5000# zpp a_11050_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1024 a_1150_n1650# bnb a_3400_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1025 a_20800_n800# bna a_20650_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1026 a_7450_n1650# bna a_7300_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1027 bpa bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1028 a_1000_n800# bna a_850_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1029 a_10150_50# bna a_10000_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1030 bpa bpa a_8650_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1031 avss bna a_8200_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1032 a_6700_4350# bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1033 a_9100_n800# bna a_8950_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1034 a_4900_5000# bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1035 a_27400_50# znp a_27250_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1036 bpb bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1037 bpa enb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1038 a_20050_50# znp a_19900_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1039 a_28300_3700# bpa a_25150_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1040 a_27850_3050# bpb znp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1041 a_250_50# bna a_100_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1042 xp im ynm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1043 a_22750_n1650# bnb a_22600_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1044 avdd zpp a_24400_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1045 znp znp a_26500_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1046 a_21250_3050# zpp a_21100_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1047 ypm zpp a_13600_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1048 xp im ynm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1049 a_20500_900# bna avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1050 avdd bpa bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1051 a_11800_50# bna a_11650_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1052 avss znp a_28600_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=3.5 pd=15 as=1.75 ps=7.5 w=7 l=1
X1053 a_10000_50# bna a_9850_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1054 ypp zpp a_22900_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1055 a_25450_n800# znp a_25300_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1056 ypp zpp a_21700_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1057 a_8050_3700# bpa a_7900_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1058 a_28000_3050# bpb a_27850_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1059 a_22150_n800# bnb a_22000_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1060 a_1600_900# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1061 a_12700_900# ip xn avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1062 a_550_3050# bpa a_4600_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1063 a_24700_3050# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1064 a_10150_900# bna a_10000_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1065 a_550_3050# bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1066 a_12700_n1650# ip xn avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1067 zpp zpp a_21250_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1068 a_13900_3700# zpp ypm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1069 ynp ip xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1070 a_16600_n1650# znp a_16450_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1071 a_26050_900# znp a_25900_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1072 bpa bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1073 ynm im xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1074 bnb bnb a_2500_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1075 bpa en avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=2.5 ps=11 w=5 l=1
X1076 a_25600_n800# znp a_25450_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1077 a_22000_5000# zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1078 a_21700_50# bnb a_21550_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1079 a_3700_n1650# en a_1150_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1080 a_22300_n800# bnb a_22150_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1081 a_7600_n1650# bna a_7450_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1082 a_3100_900# bnb a_1150_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1083 bpb bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1084 a_16600_50# znp a_16450_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1085 a_14200_900# im ypm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1086 a_8200_4350# bpa a_8050_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1087 bpb bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1088 ynp znp a_27400_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1089 a_11050_n800# bna a_10900_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1090 a_8650_900# bna a_8500_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1091 a_19750_900# znp a_19600_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1092 a_7450_50# bna a_7300_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1093 a_26500_50# znp a_26350_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1094 xp bpa a_18400_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1095 bnb bnb a_1900_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1096 a_22900_n1650# bnb a_22750_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1097 a_26800_n1650# znp znp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1098 a_15250_3700# zpp a_15100_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1099 avss enb bna avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1100 a_27850_4350# bpb znp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1101 a_850_900# bna a_700_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1102 avdd bpa a_26500_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1103 avdd zpp a_24400_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1104 a_23350_5000# zpp a_23200_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1105 avdd bpa bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1106 a_21250_4350# zpp a_21100_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1107 a_550_3050# enb bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1108 ynm im xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1109 a_250_5000# bpa a_100_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1110 a_26200_3050# bpa a_25150_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1111 a_15400_3700# zpp a_15250_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1112 a_12100_3700# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1113 ypm im a_13300_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1114 a_28000_4350# bpb a_27850_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1115 a_10900_50# bna avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1116 a_26800_5000# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1117 a_17350_n1650# znp a_17200_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1118 a_24700_4350# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1119 a_27100_n800# znp a_26950_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1120 zpp zpp a_23350_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1121 ypm zpp a_14800_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1122 bpa bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1123 zpp zpp a_21250_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1124 a_20200_5000# bpa a_20050_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1125 a_11650_3050# zpp a_11500_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1126 bpa enb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1127 a_400_5000# bpa a_250_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1128 bna en a_4300_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1129 a_100_900# bna avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1130 bpa en avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=2.5 ps=11 w=5 l=1
X1131 avss bna a_8200_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1132 bpb bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1133 a_15850_n800# znp a_15700_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1134 a_550_3050# bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1135 xn ip a_12400_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1136 a_1150_n1650# bnb a_1600_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1137 a_21400_900# bna a_21250_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1138 a_1000_50# bna a_850_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1139 a_550_3050# bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1140 a_20800_50# bna a_20650_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1141 a_11800_3050# zpp a_11650_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1142 a_15700_50# znp avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1143 bnb bnb a_6700_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1144 a_2500_900# bnb a_1150_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1145 a_13600_900# im ypm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1146 a_1150_n1650# bnb a_3400_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1147 a_16000_n800# znp a_15850_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1148 a_25150_3050# bpb a_25900_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1149 a_12700_n800# ip xn avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1150 a_23650_n1650# bna a_23500_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1151 a_26950_900# znp a_26800_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1152 ynp znp a_27400_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1153 bpb bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1154 a_22750_3700# zpp a_22600_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1155 a_25150_3050# bpb a_28000_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1156 a_7000_n800# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1157 a_1150_n1650# bnb a_6400_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1158 a_8050_900# bna a_7900_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1159 a_25600_50# znp a_25450_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1160 a_15100_900# bna a_14950_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1161 a_3700_n800# en a_1150_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1162 a_28450_900# znp a_28300_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1163 a_13600_n1650# im ypm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1164 a_100_50# bna avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1165 a_22900_3700# zpp a_22750_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1166 a_28300_5000# bpa a_25150_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1167 a_17500_n1650# znp a_17350_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1168 xp ip ynp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1169 a_26200_4350# bpa a_25150_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1170 xp ip ynp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1171 bpb bna a_9400_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1172 avdd zpp a_13000_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1173 a_4600_n1650# en bna avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1174 a_8500_n1650# bna avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1175 xn ip a_13000_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1176 xp im ynm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1177 ypm zpp a_14800_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1178 a_17350_n800# znp a_17200_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1179 ypm zpp a_13600_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1180 a_550_3050# bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1181 a_11650_4350# zpp a_11500_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1182 a_19900_3050# bpa xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1183 avdd bpa bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1184 avdd bpa a_4000_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1185 ynp ip xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1186 a_13300_3050# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1187 a_8050_5000# bpa a_7900_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1188 a_550_3050# bpb a_4900_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1189 avss bna a_8200_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1190 a_550_3050# bpa a_4600_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1191 a_550_3050# bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1192 a_550_3050# bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1193 a_17500_n800# znp a_17350_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1194 a_13900_5000# zpp ypm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1195 bpb bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1196 a_27550_3700# bpb a_27400_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1197 a_11800_4350# zpp a_11650_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1198 a_14200_n800# im ypm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1199 a_23800_n1650# bna a_23650_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1200 bpa bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1201 a_27700_n1650# znp ynp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1202 a_3100_50# bnb a_1150_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1203 a_4300_3050# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1204 a_24250_3700# zpp a_24100_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1205 a_20800_900# bna a_20650_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1206 a_14800_50# bna a_14650_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1207 a_8500_n800# bna avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1208 a_4900_5000# bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1209 bpb bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1210 a_5200_n800# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1211 bpb bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1212 a_1900_900# bnb a_1150_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1213 znp bpb a_27550_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1214 a_13000_900# ip ypp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1215 a_24400_3700# zpp a_24250_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1216 a_10450_900# bna a_10300_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1217 a_10450_n1650# bna a_10300_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1218 a_21100_3700# zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1219 a_22300_900# bnb a_22150_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1220 xn im a_14200_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1221 a_18250_n1650# znp a_18100_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1222 bnb bnb a_5500_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1223 ypp zpp a_23800_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1224 bpa en avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1225 a_24700_50# znp avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1226 bnb bnb a_1300_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1227 xp ip ynp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1228 a_20650_3050# zpp a_20500_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1229 a_3400_900# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1230 a_1150_n1650# bnb a_5200_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1231 xp bpa a_18400_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1232 a_19600_50# znp a_19450_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1233 a_14500_900# bna xn avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1234 a_550_3050# bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1235 xp ip ynp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1236 a_9250_n1650# bna a_9100_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1237 a_15250_5000# zpp a_15100_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1238 avdd zpp a_13000_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1239 a_27850_900# znp a_27700_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1240 a_24850_n800# znp a_24700_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1241 a_18100_3050# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1242 a_21550_n1650# bna a_21400_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1243 a_550_n1650# bna a_400_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1244 avdd en bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1245 avdd bpa bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1246 a_550_3050# bpb a_6700_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1247 a_19900_4350# bpa xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1248 a_8950_900# bna a_8800_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1249 a_20800_3050# zpp a_20650_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1250 a_550_3050# enb bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1251 avdd bpa a_4000_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1252 ynm im xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1253 ypp ip a_12100_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1254 a_20050_900# znp a_19900_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1255 bpb bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1256 ynp ip xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1257 a_15400_5000# zpp a_15250_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1258 a_13300_4350# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1259 bpa bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1260 a_25000_n800# znp a_24850_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1261 a_12100_5000# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1262 a_20650_n1650# bna a_20500_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1263 a_21700_n800# bnb a_21550_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1264 avss bna a_24400_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1265 a_28450_n1650# znp a_28300_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1266 bpa bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1267 a_6700_4350# bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1268 bpa enb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1269 a_4300_4350# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1270 bpb bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1271 a_22150_50# bnb a_22000_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1272 a_2200_50# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1273 a_10600_n1650# bna a_10450_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1274 a_14500_n1650# bna xn avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1275 a_18400_n1650# znp a_18250_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1276 a_13900_50# im xn avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1277 avdd bpa a_28600_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.5 pd=11 as=1.25 ps=5.5 w=5 l=1
X1278 a_25450_3050# bpb a_25300_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1279 avdd bpa a_17800_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1280 a_1600_n1650# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1281 a_14650_3700# zpp a_14500_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1282 a_22150_3050# zpp a_22000_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1283 a_5500_n1650# bnb a_1150_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1284 ypp zpp a_11200_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1285 a_9400_n1650# bna a_9250_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1286 a_25150_3050# bpb a_25900_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1287 ypp zpp a_23800_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1288 a_26350_n800# znp a_26200_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1289 a_22750_5000# zpp a_22600_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1290 avdd bpa bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1291 a_20650_4350# zpp a_20500_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1292 a_550_3050# bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1293 a_700_n1650# bna a_550_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1294 a_1150_n1650# en a_4600_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1295 a_550_3050# bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1296 a_21700_900# bnb a_21550_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1297 znp bpb a_25450_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1298 a_23800_50# bna a_23650_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1299 a_550_3050# enb bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1300 a_22300_3050# zpp a_22150_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1301 a_14800_3700# zpp a_14650_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1302 a_18100_4350# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1303 a_18700_50# znp a_18550_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1304 a_11500_3700# zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1305 a_2800_900# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1306 a_13900_900# im xn avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1307 a_26500_n800# znp a_26350_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1308 a_20800_n1650# bna a_20650_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1309 a_22900_5000# zpp a_22750_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1310 a_20800_4350# zpp a_20650_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1311 a_11350_900# bna a_11200_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1312 a_23200_n800# bnb a_23050_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1313 a_24700_n1650# znp avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1314 a_11050_3050# zpp a_10900_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1315 bpb bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1316 a_28600_n1650# znp a_28450_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1317 a_23200_900# bnb a_23050_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1318 bpb bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1319 bpb bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1320 bpa bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1321 a_11350_50# bna a_11200_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1322 bpb bna a_9400_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1323 a_4300_900# en a_1150_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1324 xn bna a_11800_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1325 a_28600_50# znp a_28450_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1326 a_15400_900# bna a_15250_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1327 a_550_3050# enb bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1328 avss znp a_28600_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=3.5 pd=15 as=1.75 ps=7.5 w=7 l=1
X1329 bna enb avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1330 a_11350_n1650# bna a_11200_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1331 a_15250_n1650# bna a_15100_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1332 xp ip ynp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1333 a_1150_n1650# bnb a_2800_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1334 ynm znp a_19000_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1335 xp bpa a_16000_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1336 a_9850_900# bna a_9700_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1337 a_21250_50# bna a_21100_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1338 a_1150_n1650# bnb a_2200_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1339 avdd bpa a_28600_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=2.5 pd=11 as=1.25 ps=5.5 w=5 l=1
X1340 bnb bnb a_6100_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1341 a_1300_50# bnb a_1150_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1342 a_27550_5000# bpb a_27400_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1343 a_25450_4350# bpb a_25300_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1344 a_16150_50# znp a_16000_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1345 a_24250_5000# zpp a_24100_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1346 a_22150_4350# zpp a_22000_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1347 a_13000_50# ip ypp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1348 a_550_3050# bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1349 a_27100_3050# bpa a_26950_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1350 ynp ip xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1351 ynp ip xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1352 a_100_n800# bna avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1353 znp bpb a_27550_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1354 znp bpb a_25450_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1355 a_24400_5000# zpp a_24250_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1356 a_15850_3050# bpa a_15700_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1357 a_22300_4350# zpp a_22150_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1358 a_21100_5000# zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1359 bna en a_3700_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1360 ypp zpp a_12400_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1361 bpb bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1362 a_21550_n1650# bna a_21400_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1363 a_25450_n1650# znp a_25300_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1364 a_6100_50# bnb a_1150_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1365 a_22900_50# bnb a_22750_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1366 bpa en avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1367 a_20050_n800# znp a_19900_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1368 ynp znp a_16600_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1369 a_17800_50# znp a_17650_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1370 a_550_3050# bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1371 a_11050_4350# zpp a_10900_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1372 ypm im a_13300_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1373 a_550_3050# bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1374 a_10150_n800# bna a_10000_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1375 a_16000_3050# bpa a_15850_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1376 a_12700_3050# zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1377 a_11500_n1650# bna a_11350_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1378 a_7750_n800# bna a_7600_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1379 avss bna a_10600_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1380 avdd en bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1381 a_15400_n1650# bna a_15250_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1382 a_550_3050# enb bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1383 a_22600_900# bnb zpp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1384 bna en a_4300_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1385 a_19300_n1650# znp ynm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1386 a_16900_n800# znp ynp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1387 a_10450_50# bna a_10300_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1388 a_8650_50# bna a_8500_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1389 a_1150_n1650# bna a_1000_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1390 bpb bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1391 a_26950_3700# bpa a_26800_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1392 a_13600_n800# im ypm avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1393 a_2500_n1650# bnb a_1150_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1394 a_27700_50# znp ynp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1395 a_3700_3050# bpa a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1396 a_23650_3700# zpp zpp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1397 a_10300_n800# bna a_10150_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1398 a_6400_n1650# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1399 a_3700_900# en a_1150_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1400 a_14800_900# bna a_14650_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1401 avdd bpa a_20200_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1402 a_550_3050# bpa a_400_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1403 a_1150_n1650# bna a_1000_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1404 ypp ip a_12100_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1405 a_7900_n800# bna a_7750_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1406 a_24100_900# bna a_23950_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1407 a_4600_n800# en bna avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1408 a_1300_n800# bnb a_1150_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1409 a_550_50# bna a_400_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1410 avss znp a_20200_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1411 a_23800_3700# zpp a_23650_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1412 a_5200_900# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1413 a_20500_3700# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1414 a_27100_4350# bpa a_26950_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1415 a_15250_50# bna a_15100_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1416 a_16300_900# znp a_16150_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1417 xp im ynm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1418 bpb bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1419 a_21700_n1650# bnb a_21550_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1420 a_25600_n1650# znp a_25450_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1421 avdd bpa a_17800_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1422 a_15850_4350# bpa a_15700_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1423 a_18250_n800# znp a_18100_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1424 a_14650_5000# zpp a_14500_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1425 ypp zpp a_12400_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1426 avdd bpa a_8200_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1427 ypp zpp a_11200_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1428 a_17500_3050# bpa xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1429 a_20950_n800# bna a_20800_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1430 a_25150_50# znp a_25000_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1431 a_14200_3050# zpp a_14050_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1432 a_1150_n1650# bnb a_2800_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1433 avdd bpa bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1434 a_550_3050# bpb a_6700_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1435 a_5200_50# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1436 a_9250_n800# bna a_9100_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1437 a_22000_50# bnb a_21850_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1438 a_550_3050# bpb a_4900_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1439 a_550_3050# bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1440 a_16000_4350# bpa a_15850_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1441 ypp ip a_12100_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1442 a_550_3050# enb bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1443 a_18400_n800# znp a_18250_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1444 a_16900_50# znp ynp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1445 a_16150_n1650# znp a_16000_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1446 a_14800_5000# zpp a_14650_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1447 bpa bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1448 a_12700_4350# zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1449 a_28450_3700# bpa a_28300_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1450 a_15100_n800# bna a_14950_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1451 a_11500_5000# zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1452 bpb bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1453 a_25150_3050# bpa a_25000_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1454 bnb bnb a_3100_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1455 a_1150_n1650# bnb a_7000_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1456 a_6700_4350# bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1457 a_9400_n800# bna a_9250_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1458 a_4900_5000# bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1459 a_3700_4350# bpa a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1460 a_6100_n800# bnb a_1150_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1461 bpb bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1462 a_7750_50# bna a_7600_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1463 a_28600_3700# bpa a_28450_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1464 a_22000_900# bnb a_21850_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1465 a_26800_50# znp znp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1466 a_25300_3700# bpb a_25150_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1467 avss enb bna avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1468 a_24850_3050# bpa a_24700_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1469 a_11650_900# bna a_11500_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1470 a_14050_3700# zpp a_13900_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1471 zpp bnb a_22300_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1472 a_21550_3050# zpp zpp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1473 xp ip ynp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1474 a_23500_900# bna a_21550_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1475 xp im ynm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1476 a_26350_n1650# znp a_26200_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1477 avdd bpa bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1478 xp bpa a_16000_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1479 ynp znp a_25600_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1480 xn im a_14200_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1481 zpp bnb a_22300_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1482 a_4600_900# en bna avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1483 a_15700_900# znp avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1484 a_550_3050# bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1485 a_25000_3050# bpa a_24850_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1486 avdd bpa a_8200_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1487 xn ip a_13000_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1488 a_550_3050# bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1489 a_21700_3050# zpp a_21550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1490 a_550_3050# bpb a_6700_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1491 bna enb avss avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=3.5 ps=15 w=7 l=1
X1492 ynp ip xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1493 a_10900_3700# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1494 a_17500_4350# bpa xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1495 a_12400_n1650# ip ypp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1496 ynp ip xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1497 a_16300_n1650# znp a_16150_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1498 a_14200_4350# zpp a_14050_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1499 a_25900_n800# znp ynp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1500 a_22600_n800# bnb zpp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1501 a_6100_900# bnb a_1150_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1502 a_3400_n1650# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1503 a_24250_50# bna a_24100_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1504 a_17200_900# znp a_17050_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1505 bnb bnb a_1900_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1506 a_7300_n1650# bna a_1150_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1507 bpa enb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1508 bpa bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1509 a_4300_50# en a_1150_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1510 a_6700_5000# bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1511 ynm znp a_19000_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1512 a_4900_4350# bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1513 a_16000_50# znp a_15850_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1514 a_26350_3050# bpa a_26200_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1515 xp im ynm avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1516 avdd zpp a_15400_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1517 a_22600_n1650# bnb zpp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1518 bnb bnb a_6700_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1519 a_26500_n1650# znp a_26350_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1520 a_12250_3700# zpp a_12100_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1521 a_9100_50# bna a_8950_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1522 a_25900_50# znp ynp avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1523 a_26950_5000# bpa a_26800_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1524 a_24850_4350# bpa a_24700_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1525 a_27250_n800# znp a_27100_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1526 a_23650_5000# zpp zpp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1527 avdd bpa bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1528 a_21550_4350# zpp zpp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1529 avdd bpa a_20200_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1530 a_550_3050# enb bpa avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1531 a_550_3050# bpa a_400_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1532 a_26500_3050# bpa a_26350_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1533 ynm im xp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1534 a_550_3050# bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1535 a_15700_3700# bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1536 a_23200_3050# zpp ypp avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1537 a_12400_3700# zpp a_12250_3700# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1538 a_11050_900# bna a_10900_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1539 xn ip a_13000_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1540 a_25000_4350# bpa a_24850_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1541 a_27400_n800# znp a_27250_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1542 a_22900_900# bnb a_22750_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1543 ypm im a_13300_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1544 a_23800_5000# zpp a_23650_5000# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1545 bpa bpa avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1546 a_21700_4350# zpp a_21550_4350# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1547 a_24100_n800# bna a_23950_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1548 avss znp a_20200_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1549 a_20500_5000# zpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1550 avdd zpp a_11800_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1551 bpb bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1552 bpb bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1553 bpb bpb a_550_3050# avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1554 a_1150_n1650# en a_4000_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1555 a_4000_900# en bna avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1556 bnb bnb a_1300_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1557 xn ip a_12400_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1558 ypp ip a_12700_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1559 a_24400_900# bna a_24250_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1560 a_550_3050# bpb bpb avdd sky130_fd_pr__pfet_g5v0d10v5 ad=1.25 pd=5.5 as=1.25 ps=5.5 w=5 l=1
X1561 a_21550_n1650# bnb a_23200_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1562 a_3400_50# bnb bnb avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1563 a_5500_900# bnb a_1150_n1650# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1564 a_18250_50# znp a_18100_50# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1565 a_16600_900# znp a_16450_900# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1566 bna en a_3700_n800# avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
X1567 avss enb bna avss sky130_fd_pr__nfet_g5v0d10v5 ad=1.75 pd=7.5 as=1.75 ps=7.5 w=7 l=1
.ends

