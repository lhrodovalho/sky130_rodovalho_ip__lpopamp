magic
tech sky130A
timestamp 1711497604
<< error_p >>
rect 28800 1850 28833 1883
rect 28767 1800 28833 1850
rect 28800 1767 28833 1800
rect 28800 -1850 28833 -1817
rect 28767 -1900 28833 -1850
rect 28800 -1933 28833 -1900
rect 28350 -2000 28800 -1950
<< dnwell >>
rect -850 -1950 28800 1900
<< nwell >>
rect -700 2900 32150 5650
rect -900 1750 28800 1950
rect -900 -1800 -700 1750
rect -900 -2000 28800 -1800
<< mvnmos >>
rect -600 900 -500 1600
rect -450 900 -350 1600
rect -300 900 -200 1600
rect -150 900 -50 1600
rect 0 900 100 1600
rect 150 900 250 1600
rect 300 900 400 1600
rect 450 900 550 1600
rect 600 900 700 1600
rect 750 900 850 1600
rect 900 900 1000 1600
rect 1050 900 1150 1600
rect 1200 900 1300 1600
rect 1350 900 1450 1600
rect 1500 900 1600 1600
rect 1650 900 1750 1600
rect 1800 900 1900 1600
rect 1950 900 2050 1600
rect 2100 900 2200 1600
rect 2250 900 2350 1600
rect 2400 900 2500 1600
rect 2550 900 2650 1600
rect 2700 900 2800 1600
rect 2850 900 2950 1600
rect 3000 900 3100 1600
rect 3150 900 3250 1600
rect 3300 900 3400 1600
rect 3450 900 3550 1600
rect 3600 900 3700 1600
rect 3750 900 3850 1600
rect 3900 900 4000 1600
rect 4050 900 4150 1600
rect 4200 900 4300 1600
rect 4350 900 4450 1600
rect 4500 900 4600 1600
rect 4650 900 4750 1600
rect 4800 900 4900 1600
rect 4950 900 5050 1600
rect 5100 900 5200 1600
rect 5250 900 5350 1600
rect 5400 900 5500 1600
rect 5550 900 5650 1600
rect 5700 900 5800 1600
rect 5850 900 5950 1600
rect 6000 900 6100 1600
rect 6150 900 6250 1600
rect 6300 900 6400 1600
rect 6450 900 6550 1600
rect 6600 900 6700 1600
rect 6750 900 6850 1600
rect 6900 900 7000 1600
rect 7050 900 7150 1600
rect 7200 900 7300 1600
rect 7350 900 7450 1600
rect 7500 900 7600 1600
rect 7650 900 7750 1600
rect 7800 900 7900 1600
rect 7950 900 8050 1600
rect 8100 900 8200 1600
rect 8250 900 8350 1600
rect 8400 900 8500 1600
rect 8550 900 8650 1600
rect 8700 900 8800 1600
rect 8850 900 8950 1600
rect 9000 900 9100 1600
rect 9150 900 9250 1600
rect 9300 900 9400 1600
rect 9450 900 9550 1600
rect 9600 900 9700 1600
rect 9750 900 9850 1600
rect 9900 900 10000 1600
rect 10050 900 10150 1600
rect 10200 900 10300 1600
rect 10350 900 10450 1600
rect 10500 900 10600 1600
rect 10650 900 10750 1600
rect 10800 900 10900 1600
rect 10950 900 11050 1600
rect 11100 900 11200 1600
rect 11250 900 11350 1600
rect 11400 900 11500 1600
rect 11550 900 11650 1600
rect 11700 900 11800 1600
rect 11850 900 11950 1600
rect 12000 900 12100 1600
rect 12150 900 12250 1600
rect 12300 900 12400 1600
rect 12450 900 12550 1600
rect 12600 900 12700 1600
rect 12750 900 12850 1600
rect 12900 900 13000 1600
rect 13050 900 13150 1600
rect 13200 900 13300 1600
rect 13350 900 13450 1600
rect 13500 900 13600 1600
rect 13650 900 13750 1600
rect 13800 900 13900 1600
rect 13950 900 14050 1600
rect 14100 900 14200 1600
rect 14250 900 14350 1600
rect 14400 900 14500 1600
rect 14550 900 14650 1600
rect 14700 900 14800 1600
rect 14850 900 14950 1600
rect 15000 900 15100 1600
rect 15150 900 15250 1600
rect 15300 900 15400 1600
rect 15450 900 15550 1600
rect 15600 900 15700 1600
rect 15750 900 15850 1600
rect 15900 900 16000 1600
rect 16050 900 16150 1600
rect 16200 900 16300 1600
rect 16350 900 16450 1600
rect 16500 900 16600 1600
rect 16650 900 16750 1600
rect 16800 900 16900 1600
rect 16950 900 17050 1600
rect 17100 900 17200 1600
rect 17250 900 17350 1600
rect 17400 900 17500 1600
rect 17550 900 17650 1600
rect 17700 900 17800 1600
rect 17850 900 17950 1600
rect 18000 900 18100 1600
rect 18150 900 18250 1600
rect 18300 900 18400 1600
rect 18450 900 18550 1600
rect 18600 900 18700 1600
rect 18750 900 18850 1600
rect 18900 900 19000 1600
rect 19050 900 19150 1600
rect 19200 900 19300 1600
rect 19350 900 19450 1600
rect 19500 900 19600 1600
rect 19650 900 19750 1600
rect 19800 900 19900 1600
rect 19950 900 20050 1600
rect 20100 900 20200 1600
rect 20250 900 20350 1600
rect 20400 900 20500 1600
rect 20550 900 20650 1600
rect 20700 900 20800 1600
rect 20850 900 20950 1600
rect 21000 900 21100 1600
rect 21150 900 21250 1600
rect 21300 900 21400 1600
rect 21450 900 21550 1600
rect 21600 900 21700 1600
rect 21750 900 21850 1600
rect 21900 900 22000 1600
rect 22050 900 22150 1600
rect 22200 900 22300 1600
rect 22350 900 22450 1600
rect 22500 900 22600 1600
rect 22650 900 22750 1600
rect 22800 900 22900 1600
rect 22950 900 23050 1600
rect 23100 900 23200 1600
rect 23250 900 23350 1600
rect 23400 900 23500 1600
rect 23550 900 23650 1600
rect 23700 900 23800 1600
rect 23850 900 23950 1600
rect 24000 900 24100 1600
rect 24150 900 24250 1600
rect 24300 900 24400 1600
rect 24450 900 24550 1600
rect 24600 900 24700 1600
rect 24750 900 24850 1600
rect 24900 900 25000 1600
rect 25050 900 25150 1600
rect 25200 900 25300 1600
rect 25350 900 25450 1600
rect 25500 900 25600 1600
rect 25650 900 25750 1600
rect 25800 900 25900 1600
rect 25950 900 26050 1600
rect 26100 900 26200 1600
rect 26250 900 26350 1600
rect 26400 900 26500 1600
rect 26550 900 26650 1600
rect 26700 900 26800 1600
rect 26850 900 26950 1600
rect 27000 900 27100 1600
rect 27150 900 27250 1600
rect 27300 900 27400 1600
rect 27450 900 27550 1600
rect 27600 900 27700 1600
rect 27750 900 27850 1600
rect 27900 900 28000 1600
rect 28050 900 28150 1600
rect 28200 900 28300 1600
rect 28350 900 28450 1600
rect 28500 900 28600 1600
rect 28650 900 28750 1600
rect -600 50 -500 750
rect -450 50 -350 750
rect -300 50 -200 750
rect -150 50 -50 750
rect 0 50 100 750
rect 150 50 250 750
rect 300 50 400 750
rect 450 50 550 750
rect 600 50 700 750
rect 750 50 850 750
rect 900 50 1000 750
rect 1050 50 1150 750
rect 1200 50 1300 750
rect 1350 50 1450 750
rect 1500 50 1600 750
rect 1650 50 1750 750
rect 1800 50 1900 750
rect 1950 50 2050 750
rect 2100 50 2200 750
rect 2250 50 2350 750
rect 2400 50 2500 750
rect 2550 50 2650 750
rect 2700 50 2800 750
rect 2850 50 2950 750
rect 3000 50 3100 750
rect 3150 50 3250 750
rect 3300 50 3400 750
rect 3450 50 3550 750
rect 3600 50 3700 750
rect 3750 50 3850 750
rect 3900 50 4000 750
rect 4050 50 4150 750
rect 4200 50 4300 750
rect 4350 50 4450 750
rect 4500 50 4600 750
rect 4650 50 4750 750
rect 4800 50 4900 750
rect 4950 50 5050 750
rect 5100 50 5200 750
rect 5250 50 5350 750
rect 5400 50 5500 750
rect 5550 50 5650 750
rect 5700 50 5800 750
rect 5850 50 5950 750
rect 6000 50 6100 750
rect 6150 50 6250 750
rect 6300 50 6400 750
rect 6450 50 6550 750
rect 6600 50 6700 750
rect 6750 50 6850 750
rect 6900 50 7000 750
rect 7050 50 7150 750
rect 7200 50 7300 750
rect 7350 50 7450 750
rect 7500 50 7600 750
rect 7650 50 7750 750
rect 7800 50 7900 750
rect 7950 50 8050 750
rect 8100 50 8200 750
rect 8250 50 8350 750
rect 8400 50 8500 750
rect 8550 50 8650 750
rect 8700 50 8800 750
rect 8850 50 8950 750
rect 9000 50 9100 750
rect 9150 50 9250 750
rect 9300 50 9400 750
rect 9450 50 9550 750
rect 9600 50 9700 750
rect 9750 50 9850 750
rect 9900 50 10000 750
rect 10050 50 10150 750
rect 10200 50 10300 750
rect 10350 50 10450 750
rect 10500 50 10600 750
rect 10650 50 10750 750
rect 10800 50 10900 750
rect 10950 50 11050 750
rect 11100 50 11200 750
rect 11250 50 11350 750
rect 11400 50 11500 750
rect 11550 50 11650 750
rect 11700 50 11800 750
rect 11850 50 11950 750
rect 12000 50 12100 750
rect 12150 50 12250 750
rect 12300 50 12400 750
rect 12450 50 12550 750
rect 12600 50 12700 750
rect 12750 50 12850 750
rect 12900 50 13000 750
rect 13050 50 13150 750
rect 13200 50 13300 750
rect 13350 50 13450 750
rect 13500 50 13600 750
rect 13650 50 13750 750
rect 13800 50 13900 750
rect 13950 50 14050 750
rect 14100 50 14200 750
rect 14250 50 14350 750
rect 14400 50 14500 750
rect 14550 50 14650 750
rect 14700 50 14800 750
rect 14850 50 14950 750
rect 15000 50 15100 750
rect 15150 50 15250 750
rect 15300 50 15400 750
rect 15450 50 15550 750
rect 15600 50 15700 750
rect 15750 50 15850 750
rect 15900 50 16000 750
rect 16050 50 16150 750
rect 16200 50 16300 750
rect 16350 50 16450 750
rect 16500 50 16600 750
rect 16650 50 16750 750
rect 16800 50 16900 750
rect 16950 50 17050 750
rect 17100 50 17200 750
rect 17250 50 17350 750
rect 17400 50 17500 750
rect 17550 50 17650 750
rect 17700 50 17800 750
rect 17850 50 17950 750
rect 18000 50 18100 750
rect 18150 50 18250 750
rect 18300 50 18400 750
rect 18450 50 18550 750
rect 18600 50 18700 750
rect 18750 50 18850 750
rect 18900 50 19000 750
rect 19050 50 19150 750
rect 19200 50 19300 750
rect 19350 50 19450 750
rect 19500 50 19600 750
rect 19650 50 19750 750
rect 19800 50 19900 750
rect 19950 50 20050 750
rect 20100 50 20200 750
rect 20250 50 20350 750
rect 20400 50 20500 750
rect 20550 50 20650 750
rect 20700 50 20800 750
rect 20850 50 20950 750
rect 21000 50 21100 750
rect 21150 50 21250 750
rect 21300 50 21400 750
rect 21450 50 21550 750
rect 21600 50 21700 750
rect 21750 50 21850 750
rect 21900 50 22000 750
rect 22050 50 22150 750
rect 22200 50 22300 750
rect 22350 50 22450 750
rect 22500 50 22600 750
rect 22650 50 22750 750
rect 22800 50 22900 750
rect 22950 50 23050 750
rect 23100 50 23200 750
rect 23250 50 23350 750
rect 23400 50 23500 750
rect 23550 50 23650 750
rect 23700 50 23800 750
rect 23850 50 23950 750
rect 24000 50 24100 750
rect 24150 50 24250 750
rect 24300 50 24400 750
rect 24450 50 24550 750
rect 24600 50 24700 750
rect 24750 50 24850 750
rect 24900 50 25000 750
rect 25050 50 25150 750
rect 25200 50 25300 750
rect 25350 50 25450 750
rect 25500 50 25600 750
rect 25650 50 25750 750
rect 25800 50 25900 750
rect 25950 50 26050 750
rect 26100 50 26200 750
rect 26250 50 26350 750
rect 26400 50 26500 750
rect 26550 50 26650 750
rect 26700 50 26800 750
rect 26850 50 26950 750
rect 27000 50 27100 750
rect 27150 50 27250 750
rect 27300 50 27400 750
rect 27450 50 27550 750
rect 27600 50 27700 750
rect 27750 50 27850 750
rect 27900 50 28000 750
rect 28050 50 28150 750
rect 28200 50 28300 750
rect 28350 50 28450 750
rect 28500 50 28600 750
rect 28650 50 28750 750
rect -600 -800 -500 -100
rect -450 -800 -350 -100
rect -300 -800 -200 -100
rect -150 -800 -50 -100
rect 0 -800 100 -100
rect 150 -800 250 -100
rect 300 -800 400 -100
rect 450 -800 550 -100
rect 600 -800 700 -100
rect 750 -800 850 -100
rect 900 -800 1000 -100
rect 1050 -800 1150 -100
rect 1200 -800 1300 -100
rect 1350 -800 1450 -100
rect 1500 -800 1600 -100
rect 1650 -800 1750 -100
rect 1800 -800 1900 -100
rect 1950 -800 2050 -100
rect 2100 -800 2200 -100
rect 2250 -800 2350 -100
rect 2400 -800 2500 -100
rect 2550 -800 2650 -100
rect 2700 -800 2800 -100
rect 2850 -800 2950 -100
rect 3000 -800 3100 -100
rect 3150 -800 3250 -100
rect 3300 -800 3400 -100
rect 3450 -800 3550 -100
rect 3600 -800 3700 -100
rect 3750 -800 3850 -100
rect 3900 -800 4000 -100
rect 4050 -800 4150 -100
rect 4200 -800 4300 -100
rect 4350 -800 4450 -100
rect 4500 -800 4600 -100
rect 4650 -800 4750 -100
rect 4800 -800 4900 -100
rect 4950 -800 5050 -100
rect 5100 -800 5200 -100
rect 5250 -800 5350 -100
rect 5400 -800 5500 -100
rect 5550 -800 5650 -100
rect 5700 -800 5800 -100
rect 5850 -800 5950 -100
rect 6000 -800 6100 -100
rect 6150 -800 6250 -100
rect 6300 -800 6400 -100
rect 6450 -800 6550 -100
rect 6600 -800 6700 -100
rect 6750 -800 6850 -100
rect 6900 -800 7000 -100
rect 7050 -800 7150 -100
rect 7200 -800 7300 -100
rect 7350 -800 7450 -100
rect 7500 -800 7600 -100
rect 7650 -800 7750 -100
rect 7800 -800 7900 -100
rect 7950 -800 8050 -100
rect 8100 -800 8200 -100
rect 8250 -800 8350 -100
rect 8400 -800 8500 -100
rect 8550 -800 8650 -100
rect 8700 -800 8800 -100
rect 8850 -800 8950 -100
rect 9000 -800 9100 -100
rect 9150 -800 9250 -100
rect 9300 -800 9400 -100
rect 9450 -800 9550 -100
rect 9600 -800 9700 -100
rect 9750 -800 9850 -100
rect 9900 -800 10000 -100
rect 10050 -800 10150 -100
rect 10200 -800 10300 -100
rect 10350 -800 10450 -100
rect 10500 -800 10600 -100
rect 10650 -800 10750 -100
rect 10800 -800 10900 -100
rect 10950 -800 11050 -100
rect 11100 -800 11200 -100
rect 11250 -800 11350 -100
rect 11400 -800 11500 -100
rect 11550 -800 11650 -100
rect 11700 -800 11800 -100
rect 11850 -800 11950 -100
rect 12000 -800 12100 -100
rect 12150 -800 12250 -100
rect 12300 -800 12400 -100
rect 12450 -800 12550 -100
rect 12600 -800 12700 -100
rect 12750 -800 12850 -100
rect 12900 -800 13000 -100
rect 13050 -800 13150 -100
rect 13200 -800 13300 -100
rect 13350 -800 13450 -100
rect 13500 -800 13600 -100
rect 13650 -800 13750 -100
rect 13800 -800 13900 -100
rect 13950 -800 14050 -100
rect 14100 -800 14200 -100
rect 14250 -800 14350 -100
rect 14400 -800 14500 -100
rect 14550 -800 14650 -100
rect 14700 -800 14800 -100
rect 14850 -800 14950 -100
rect 15000 -800 15100 -100
rect 15150 -800 15250 -100
rect 15300 -800 15400 -100
rect 15450 -800 15550 -100
rect 15600 -800 15700 -100
rect 15750 -800 15850 -100
rect 15900 -800 16000 -100
rect 16050 -800 16150 -100
rect 16200 -800 16300 -100
rect 16350 -800 16450 -100
rect 16500 -800 16600 -100
rect 16650 -800 16750 -100
rect 16800 -800 16900 -100
rect 16950 -800 17050 -100
rect 17100 -800 17200 -100
rect 17250 -800 17350 -100
rect 17400 -800 17500 -100
rect 17550 -800 17650 -100
rect 17700 -800 17800 -100
rect 17850 -800 17950 -100
rect 18000 -800 18100 -100
rect 18150 -800 18250 -100
rect 18300 -800 18400 -100
rect 18450 -800 18550 -100
rect 18600 -800 18700 -100
rect 18750 -800 18850 -100
rect 18900 -800 19000 -100
rect 19050 -800 19150 -100
rect 19200 -800 19300 -100
rect 19350 -800 19450 -100
rect 19500 -800 19600 -100
rect 19650 -800 19750 -100
rect 19800 -800 19900 -100
rect 19950 -800 20050 -100
rect 20100 -800 20200 -100
rect 20250 -800 20350 -100
rect 20400 -800 20500 -100
rect 20550 -800 20650 -100
rect 20700 -800 20800 -100
rect 20850 -800 20950 -100
rect 21000 -800 21100 -100
rect 21150 -800 21250 -100
rect 21300 -800 21400 -100
rect 21450 -800 21550 -100
rect 21600 -800 21700 -100
rect 21750 -800 21850 -100
rect 21900 -800 22000 -100
rect 22050 -800 22150 -100
rect 22200 -800 22300 -100
rect 22350 -800 22450 -100
rect 22500 -800 22600 -100
rect 22650 -800 22750 -100
rect 22800 -800 22900 -100
rect 22950 -800 23050 -100
rect 23100 -800 23200 -100
rect 23250 -800 23350 -100
rect 23400 -800 23500 -100
rect 23550 -800 23650 -100
rect 23700 -800 23800 -100
rect 23850 -800 23950 -100
rect 24000 -800 24100 -100
rect 24150 -800 24250 -100
rect 24300 -800 24400 -100
rect 24450 -800 24550 -100
rect 24600 -800 24700 -100
rect 24750 -800 24850 -100
rect 24900 -800 25000 -100
rect 25050 -800 25150 -100
rect 25200 -800 25300 -100
rect 25350 -800 25450 -100
rect 25500 -800 25600 -100
rect 25650 -800 25750 -100
rect 25800 -800 25900 -100
rect 25950 -800 26050 -100
rect 26100 -800 26200 -100
rect 26250 -800 26350 -100
rect 26400 -800 26500 -100
rect 26550 -800 26650 -100
rect 26700 -800 26800 -100
rect 26850 -800 26950 -100
rect 27000 -800 27100 -100
rect 27150 -800 27250 -100
rect 27300 -800 27400 -100
rect 27450 -800 27550 -100
rect 27600 -800 27700 -100
rect 27750 -800 27850 -100
rect 27900 -800 28000 -100
rect 28050 -800 28150 -100
rect 28200 -800 28300 -100
rect 28350 -800 28450 -100
rect 28500 -800 28600 -100
rect 28650 -800 28750 -100
rect -600 -1650 -500 -950
rect -450 -1650 -350 -950
rect -300 -1650 -200 -950
rect -150 -1650 -50 -950
rect 0 -1650 100 -950
rect 150 -1650 250 -950
rect 300 -1650 400 -950
rect 450 -1650 550 -950
rect 600 -1650 700 -950
rect 750 -1650 850 -950
rect 900 -1650 1000 -950
rect 1050 -1650 1150 -950
rect 1200 -1650 1300 -950
rect 1350 -1650 1450 -950
rect 1500 -1650 1600 -950
rect 1650 -1650 1750 -950
rect 1800 -1650 1900 -950
rect 1950 -1650 2050 -950
rect 2100 -1650 2200 -950
rect 2250 -1650 2350 -950
rect 2400 -1650 2500 -950
rect 2550 -1650 2650 -950
rect 2700 -1650 2800 -950
rect 2850 -1650 2950 -950
rect 3000 -1650 3100 -950
rect 3150 -1650 3250 -950
rect 3300 -1650 3400 -950
rect 3450 -1650 3550 -950
rect 3600 -1650 3700 -950
rect 3750 -1650 3850 -950
rect 3900 -1650 4000 -950
rect 4050 -1650 4150 -950
rect 4200 -1650 4300 -950
rect 4350 -1650 4450 -950
rect 4500 -1650 4600 -950
rect 4650 -1650 4750 -950
rect 4800 -1650 4900 -950
rect 4950 -1650 5050 -950
rect 5100 -1650 5200 -950
rect 5250 -1650 5350 -950
rect 5400 -1650 5500 -950
rect 5550 -1650 5650 -950
rect 5700 -1650 5800 -950
rect 5850 -1650 5950 -950
rect 6000 -1650 6100 -950
rect 6150 -1650 6250 -950
rect 6300 -1650 6400 -950
rect 6450 -1650 6550 -950
rect 6600 -1650 6700 -950
rect 6750 -1650 6850 -950
rect 6900 -1650 7000 -950
rect 7050 -1650 7150 -950
rect 7200 -1650 7300 -950
rect 7350 -1650 7450 -950
rect 7500 -1650 7600 -950
rect 7650 -1650 7750 -950
rect 7800 -1650 7900 -950
rect 7950 -1650 8050 -950
rect 8100 -1650 8200 -950
rect 8250 -1650 8350 -950
rect 8400 -1650 8500 -950
rect 8550 -1650 8650 -950
rect 8700 -1650 8800 -950
rect 8850 -1650 8950 -950
rect 9000 -1650 9100 -950
rect 9150 -1650 9250 -950
rect 9300 -1650 9400 -950
rect 9450 -1650 9550 -950
rect 9600 -1650 9700 -950
rect 9750 -1650 9850 -950
rect 9900 -1650 10000 -950
rect 10050 -1650 10150 -950
rect 10200 -1650 10300 -950
rect 10350 -1650 10450 -950
rect 10500 -1650 10600 -950
rect 10650 -1650 10750 -950
rect 10800 -1650 10900 -950
rect 10950 -1650 11050 -950
rect 11100 -1650 11200 -950
rect 11250 -1650 11350 -950
rect 11400 -1650 11500 -950
rect 11550 -1650 11650 -950
rect 11700 -1650 11800 -950
rect 11850 -1650 11950 -950
rect 12000 -1650 12100 -950
rect 12150 -1650 12250 -950
rect 12300 -1650 12400 -950
rect 12450 -1650 12550 -950
rect 12600 -1650 12700 -950
rect 12750 -1650 12850 -950
rect 12900 -1650 13000 -950
rect 13050 -1650 13150 -950
rect 13200 -1650 13300 -950
rect 13350 -1650 13450 -950
rect 13500 -1650 13600 -950
rect 13650 -1650 13750 -950
rect 13800 -1650 13900 -950
rect 13950 -1650 14050 -950
rect 14100 -1650 14200 -950
rect 14250 -1650 14350 -950
rect 14400 -1650 14500 -950
rect 14550 -1650 14650 -950
rect 14700 -1650 14800 -950
rect 14850 -1650 14950 -950
rect 15000 -1650 15100 -950
rect 15150 -1650 15250 -950
rect 15300 -1650 15400 -950
rect 15450 -1650 15550 -950
rect 15600 -1650 15700 -950
rect 15750 -1650 15850 -950
rect 15900 -1650 16000 -950
rect 16050 -1650 16150 -950
rect 16200 -1650 16300 -950
rect 16350 -1650 16450 -950
rect 16500 -1650 16600 -950
rect 16650 -1650 16750 -950
rect 16800 -1650 16900 -950
rect 16950 -1650 17050 -950
rect 17100 -1650 17200 -950
rect 17250 -1650 17350 -950
rect 17400 -1650 17500 -950
rect 17550 -1650 17650 -950
rect 17700 -1650 17800 -950
rect 17850 -1650 17950 -950
rect 18000 -1650 18100 -950
rect 18150 -1650 18250 -950
rect 18300 -1650 18400 -950
rect 18450 -1650 18550 -950
rect 18600 -1650 18700 -950
rect 18750 -1650 18850 -950
rect 18900 -1650 19000 -950
rect 19050 -1650 19150 -950
rect 19200 -1650 19300 -950
rect 19350 -1650 19450 -950
rect 19500 -1650 19600 -950
rect 19650 -1650 19750 -950
rect 19800 -1650 19900 -950
rect 19950 -1650 20050 -950
rect 20100 -1650 20200 -950
rect 20250 -1650 20350 -950
rect 20400 -1650 20500 -950
rect 20550 -1650 20650 -950
rect 20700 -1650 20800 -950
rect 20850 -1650 20950 -950
rect 21000 -1650 21100 -950
rect 21150 -1650 21250 -950
rect 21300 -1650 21400 -950
rect 21450 -1650 21550 -950
rect 21600 -1650 21700 -950
rect 21750 -1650 21850 -950
rect 21900 -1650 22000 -950
rect 22050 -1650 22150 -950
rect 22200 -1650 22300 -950
rect 22350 -1650 22450 -950
rect 22500 -1650 22600 -950
rect 22650 -1650 22750 -950
rect 22800 -1650 22900 -950
rect 22950 -1650 23050 -950
rect 23100 -1650 23200 -950
rect 23250 -1650 23350 -950
rect 23400 -1650 23500 -950
rect 23550 -1650 23650 -950
rect 23700 -1650 23800 -950
rect 23850 -1650 23950 -950
rect 24000 -1650 24100 -950
rect 24150 -1650 24250 -950
rect 24300 -1650 24400 -950
rect 24450 -1650 24550 -950
rect 24600 -1650 24700 -950
rect 24750 -1650 24850 -950
rect 24900 -1650 25000 -950
rect 25050 -1650 25150 -950
rect 25200 -1650 25300 -950
rect 25350 -1650 25450 -950
rect 25500 -1650 25600 -950
rect 25650 -1650 25750 -950
rect 25800 -1650 25900 -950
rect 25950 -1650 26050 -950
rect 26100 -1650 26200 -950
rect 26250 -1650 26350 -950
rect 26400 -1650 26500 -950
rect 26550 -1650 26650 -950
rect 26700 -1650 26800 -950
rect 26850 -1650 26950 -950
rect 27000 -1650 27100 -950
rect 27150 -1650 27250 -950
rect 27300 -1650 27400 -950
rect 27450 -1650 27550 -950
rect 27600 -1650 27700 -950
rect 27750 -1650 27850 -950
rect 27900 -1650 28000 -950
rect 28050 -1650 28150 -950
rect 28200 -1650 28300 -950
rect 28350 -1650 28450 -950
rect 28500 -1650 28600 -950
rect 28650 -1650 28750 -950
<< mvpmos >>
rect -600 5000 -500 5500
rect -450 5000 -350 5500
rect -300 5000 -200 5500
rect -150 5000 -50 5500
rect 0 5000 100 5500
rect 150 5000 250 5500
rect 300 5000 400 5500
rect 450 5000 550 5500
rect 600 5000 700 5500
rect 750 5000 850 5500
rect 900 5000 1000 5500
rect 1050 5000 1150 5500
rect 1200 5000 1300 5500
rect 1350 5000 1450 5500
rect 1500 5000 1600 5500
rect 1650 5000 1750 5500
rect 1800 5000 1900 5500
rect 1950 5000 2050 5500
rect 2100 5000 2200 5500
rect 2250 5000 2350 5500
rect 2400 5000 2500 5500
rect 2550 5000 2650 5500
rect 2700 5000 2800 5500
rect 2850 5000 2950 5500
rect 3000 5000 3100 5500
rect 3150 5000 3250 5500
rect 3300 5000 3400 5500
rect 3450 5000 3550 5500
rect 3600 5000 3700 5500
rect 3750 5000 3850 5500
rect 3900 5000 4000 5500
rect 4050 5000 4150 5500
rect 4200 5000 4300 5500
rect 4350 5000 4450 5500
rect 4500 5000 4600 5500
rect 4650 5000 4750 5500
rect 4800 5000 4900 5500
rect 4950 5000 5050 5500
rect 5100 5000 5200 5500
rect 5250 5000 5350 5500
rect 5400 5000 5500 5500
rect 5550 5000 5650 5500
rect 5700 5000 5800 5500
rect 5850 5000 5950 5500
rect 6000 5000 6100 5500
rect 6150 5000 6250 5500
rect 6300 5000 6400 5500
rect 6450 5000 6550 5500
rect 6600 5000 6700 5500
rect 6750 5000 6850 5500
rect 6900 5000 7000 5500
rect 7050 5000 7150 5500
rect 7200 5000 7300 5500
rect 7350 5000 7450 5500
rect 7500 5000 7600 5500
rect 7650 5000 7750 5500
rect 7800 5000 7900 5500
rect 7950 5000 8050 5500
rect 8100 5000 8200 5500
rect 8250 5000 8350 5500
rect 8400 5000 8500 5500
rect 8550 5000 8650 5500
rect 8700 5000 8800 5500
rect 8850 5000 8950 5500
rect 9000 5000 9100 5500
rect 9150 5000 9250 5500
rect 9300 5000 9400 5500
rect 9450 5000 9550 5500
rect 9600 5000 9700 5500
rect 9750 5000 9850 5500
rect 9900 5000 10000 5500
rect 10050 5000 10150 5500
rect 10200 5000 10300 5500
rect 10350 5000 10450 5500
rect 10500 5000 10600 5500
rect 10650 5000 10750 5500
rect 10800 5000 10900 5500
rect 10950 5000 11050 5500
rect 11100 5000 11200 5500
rect 11250 5000 11350 5500
rect 11400 5000 11500 5500
rect 11550 5000 11650 5500
rect 11700 5000 11800 5500
rect 11850 5000 11950 5500
rect 12000 5000 12100 5500
rect 12150 5000 12250 5500
rect 12300 5000 12400 5500
rect 12450 5000 12550 5500
rect 12600 5000 12700 5500
rect 12750 5000 12850 5500
rect 12900 5000 13000 5500
rect 13050 5000 13150 5500
rect 13200 5000 13300 5500
rect 13350 5000 13450 5500
rect 13500 5000 13600 5500
rect 13650 5000 13750 5500
rect 13800 5000 13900 5500
rect 13950 5000 14050 5500
rect 14100 5000 14200 5500
rect 14250 5000 14350 5500
rect 14400 5000 14500 5500
rect 14550 5000 14650 5500
rect 14700 5000 14800 5500
rect 14850 5000 14950 5500
rect 15000 5000 15100 5500
rect 15150 5000 15250 5500
rect 15300 5000 15400 5500
rect 15450 5000 15550 5500
rect 15600 5000 15700 5500
rect 15750 5000 15850 5500
rect 15900 5000 16000 5500
rect 16050 5000 16150 5500
rect 16200 5000 16300 5500
rect 16350 5000 16450 5500
rect 16500 5000 16600 5500
rect 16650 5000 16750 5500
rect 16800 5000 16900 5500
rect 16950 5000 17050 5500
rect 17100 5000 17200 5500
rect 17250 5000 17350 5500
rect 17400 5000 17500 5500
rect 17550 5000 17650 5500
rect 17700 5000 17800 5500
rect 17850 5000 17950 5500
rect 18000 5000 18100 5500
rect 18150 5000 18250 5500
rect 18300 5000 18400 5500
rect 18450 5000 18550 5500
rect 18600 5000 18700 5500
rect 18750 5000 18850 5500
rect 18900 5000 19000 5500
rect 19050 5000 19150 5500
rect 19200 5000 19300 5500
rect 19350 5000 19450 5500
rect 19500 5000 19600 5500
rect 19650 5000 19750 5500
rect 19800 5000 19900 5500
rect 19950 5000 20050 5500
rect 20100 5000 20200 5500
rect 20250 5000 20350 5500
rect 20400 5000 20500 5500
rect 20550 5000 20650 5500
rect 20700 5000 20800 5500
rect 20850 5000 20950 5500
rect 21000 5000 21100 5500
rect 21150 5000 21250 5500
rect 21300 5000 21400 5500
rect 21450 5000 21550 5500
rect 21600 5000 21700 5500
rect 21750 5000 21850 5500
rect 21900 5000 22000 5500
rect 22050 5000 22150 5500
rect 22200 5000 22300 5500
rect 22350 5000 22450 5500
rect 22500 5000 22600 5500
rect 22650 5000 22750 5500
rect 22800 5000 22900 5500
rect 22950 5000 23050 5500
rect 23100 5000 23200 5500
rect 23250 5000 23350 5500
rect 23400 5000 23500 5500
rect 23550 5000 23650 5500
rect 23700 5000 23800 5500
rect 23850 5000 23950 5500
rect 24000 5000 24100 5500
rect 24150 5000 24250 5500
rect 24300 5000 24400 5500
rect 24450 5000 24550 5500
rect 24600 5000 24700 5500
rect 24750 5000 24850 5500
rect 24900 5000 25000 5500
rect 25050 5000 25150 5500
rect 25200 5000 25300 5500
rect 25350 5000 25450 5500
rect 25500 5000 25600 5500
rect 25650 5000 25750 5500
rect 25800 5000 25900 5500
rect 25950 5000 26050 5500
rect 26100 5000 26200 5500
rect 26250 5000 26350 5500
rect 26400 5000 26500 5500
rect 26550 5000 26650 5500
rect 26700 5000 26800 5500
rect 26850 5000 26950 5500
rect 27000 5000 27100 5500
rect 27150 5000 27250 5500
rect 27300 5000 27400 5500
rect 27450 5000 27550 5500
rect 27600 5000 27700 5500
rect 27750 5000 27850 5500
rect 27900 5000 28000 5500
rect 28050 5000 28150 5500
rect 28200 5000 28300 5500
rect 28350 5000 28450 5500
rect 28500 5000 28600 5500
rect 28650 5000 28750 5500
rect 28800 5000 28900 5500
rect 28950 5000 29050 5500
rect 29100 5000 29200 5500
rect 29250 5000 29350 5500
rect 29400 5000 29500 5500
rect 29550 5000 29650 5500
rect 29700 5000 29800 5500
rect 29850 5000 29950 5500
rect 30000 5000 30100 5500
rect 30150 5000 30250 5500
rect 30300 5000 30400 5500
rect 30450 5000 30550 5500
rect 30600 5000 30700 5500
rect 30750 5000 30850 5500
rect 30900 5000 31000 5500
rect 31050 5000 31150 5500
rect 31200 5000 31300 5500
rect 31350 5000 31450 5500
rect 31500 5000 31600 5500
rect 31650 5000 31750 5500
rect 31800 5000 31900 5500
rect 31950 5000 32050 5500
rect -600 4350 -500 4850
rect -450 4350 -350 4850
rect -300 4350 -200 4850
rect -150 4350 -50 4850
rect 0 4350 100 4850
rect 150 4350 250 4850
rect 300 4350 400 4850
rect 450 4350 550 4850
rect 600 4350 700 4850
rect 750 4350 850 4850
rect 900 4350 1000 4850
rect 1050 4350 1150 4850
rect 1200 4350 1300 4850
rect 1350 4350 1450 4850
rect 1500 4350 1600 4850
rect 1650 4350 1750 4850
rect 1800 4350 1900 4850
rect 1950 4350 2050 4850
rect 2100 4350 2200 4850
rect 2250 4350 2350 4850
rect 2400 4350 2500 4850
rect 2550 4350 2650 4850
rect 2700 4350 2800 4850
rect 2850 4350 2950 4850
rect 3000 4350 3100 4850
rect 3150 4350 3250 4850
rect 3300 4350 3400 4850
rect 3450 4350 3550 4850
rect 3600 4350 3700 4850
rect 3750 4350 3850 4850
rect 3900 4350 4000 4850
rect 4050 4350 4150 4850
rect 4200 4350 4300 4850
rect 4350 4350 4450 4850
rect 4500 4350 4600 4850
rect 4650 4350 4750 4850
rect 4800 4350 4900 4850
rect 4950 4350 5050 4850
rect 5100 4350 5200 4850
rect 5250 4350 5350 4850
rect 5400 4350 5500 4850
rect 5550 4350 5650 4850
rect 5700 4350 5800 4850
rect 5850 4350 5950 4850
rect 6000 4350 6100 4850
rect 6150 4350 6250 4850
rect 6300 4350 6400 4850
rect 6450 4350 6550 4850
rect 6600 4350 6700 4850
rect 6750 4350 6850 4850
rect 6900 4350 7000 4850
rect 7050 4350 7150 4850
rect 7200 4350 7300 4850
rect 7350 4350 7450 4850
rect 7500 4350 7600 4850
rect 7650 4350 7750 4850
rect 7800 4350 7900 4850
rect 7950 4350 8050 4850
rect 8100 4350 8200 4850
rect 8250 4350 8350 4850
rect 8400 4350 8500 4850
rect 8550 4350 8650 4850
rect 8700 4350 8800 4850
rect 8850 4350 8950 4850
rect 9000 4350 9100 4850
rect 9150 4350 9250 4850
rect 9300 4350 9400 4850
rect 9450 4350 9550 4850
rect 9600 4350 9700 4850
rect 9750 4350 9850 4850
rect 9900 4350 10000 4850
rect 10050 4350 10150 4850
rect 10200 4350 10300 4850
rect 10350 4350 10450 4850
rect 10500 4350 10600 4850
rect 10650 4350 10750 4850
rect 10800 4350 10900 4850
rect 10950 4350 11050 4850
rect 11100 4350 11200 4850
rect 11250 4350 11350 4850
rect 11400 4350 11500 4850
rect 11550 4350 11650 4850
rect 11700 4350 11800 4850
rect 11850 4350 11950 4850
rect 12000 4350 12100 4850
rect 12150 4350 12250 4850
rect 12300 4350 12400 4850
rect 12450 4350 12550 4850
rect 12600 4350 12700 4850
rect 12750 4350 12850 4850
rect 12900 4350 13000 4850
rect 13050 4350 13150 4850
rect 13200 4350 13300 4850
rect 13350 4350 13450 4850
rect 13500 4350 13600 4850
rect 13650 4350 13750 4850
rect 13800 4350 13900 4850
rect 13950 4350 14050 4850
rect 14100 4350 14200 4850
rect 14250 4350 14350 4850
rect 14400 4350 14500 4850
rect 14550 4350 14650 4850
rect 14700 4350 14800 4850
rect 14850 4350 14950 4850
rect 15000 4350 15100 4850
rect 15150 4350 15250 4850
rect 15300 4350 15400 4850
rect 15450 4350 15550 4850
rect 15600 4350 15700 4850
rect 15750 4350 15850 4850
rect 15900 4350 16000 4850
rect 16050 4350 16150 4850
rect 16200 4350 16300 4850
rect 16350 4350 16450 4850
rect 16500 4350 16600 4850
rect 16650 4350 16750 4850
rect 16800 4350 16900 4850
rect 16950 4350 17050 4850
rect 17100 4350 17200 4850
rect 17250 4350 17350 4850
rect 17400 4350 17500 4850
rect 17550 4350 17650 4850
rect 17700 4350 17800 4850
rect 17850 4350 17950 4850
rect 18000 4350 18100 4850
rect 18150 4350 18250 4850
rect 18300 4350 18400 4850
rect 18450 4350 18550 4850
rect 18600 4350 18700 4850
rect 18750 4350 18850 4850
rect 18900 4350 19000 4850
rect 19050 4350 19150 4850
rect 19200 4350 19300 4850
rect 19350 4350 19450 4850
rect 19500 4350 19600 4850
rect 19650 4350 19750 4850
rect 19800 4350 19900 4850
rect 19950 4350 20050 4850
rect 20100 4350 20200 4850
rect 20250 4350 20350 4850
rect 20400 4350 20500 4850
rect 20550 4350 20650 4850
rect 20700 4350 20800 4850
rect 20850 4350 20950 4850
rect 21000 4350 21100 4850
rect 21150 4350 21250 4850
rect 21300 4350 21400 4850
rect 21450 4350 21550 4850
rect 21600 4350 21700 4850
rect 21750 4350 21850 4850
rect 21900 4350 22000 4850
rect 22050 4350 22150 4850
rect 22200 4350 22300 4850
rect 22350 4350 22450 4850
rect 22500 4350 22600 4850
rect 22650 4350 22750 4850
rect 22800 4350 22900 4850
rect 22950 4350 23050 4850
rect 23100 4350 23200 4850
rect 23250 4350 23350 4850
rect 23400 4350 23500 4850
rect 23550 4350 23650 4850
rect 23700 4350 23800 4850
rect 23850 4350 23950 4850
rect 24000 4350 24100 4850
rect 24150 4350 24250 4850
rect 24300 4350 24400 4850
rect 24450 4350 24550 4850
rect 24600 4350 24700 4850
rect 24750 4350 24850 4850
rect 24900 4350 25000 4850
rect 25050 4350 25150 4850
rect 25200 4350 25300 4850
rect 25350 4350 25450 4850
rect 25500 4350 25600 4850
rect 25650 4350 25750 4850
rect 25800 4350 25900 4850
rect 25950 4350 26050 4850
rect 26100 4350 26200 4850
rect 26250 4350 26350 4850
rect 26400 4350 26500 4850
rect 26550 4350 26650 4850
rect 26700 4350 26800 4850
rect 26850 4350 26950 4850
rect 27000 4350 27100 4850
rect 27150 4350 27250 4850
rect 27300 4350 27400 4850
rect 27450 4350 27550 4850
rect 27600 4350 27700 4850
rect 27750 4350 27850 4850
rect 27900 4350 28000 4850
rect 28050 4350 28150 4850
rect 28200 4350 28300 4850
rect 28350 4350 28450 4850
rect 28500 4350 28600 4850
rect 28650 4350 28750 4850
rect 28800 4350 28900 4850
rect 28950 4350 29050 4850
rect 29100 4350 29200 4850
rect 29250 4350 29350 4850
rect 29400 4350 29500 4850
rect 29550 4350 29650 4850
rect 29700 4350 29800 4850
rect 29850 4350 29950 4850
rect 30000 4350 30100 4850
rect 30150 4350 30250 4850
rect 30300 4350 30400 4850
rect 30450 4350 30550 4850
rect 30600 4350 30700 4850
rect 30750 4350 30850 4850
rect 30900 4350 31000 4850
rect 31050 4350 31150 4850
rect 31200 4350 31300 4850
rect 31350 4350 31450 4850
rect 31500 4350 31600 4850
rect 31650 4350 31750 4850
rect 31800 4350 31900 4850
rect 31950 4350 32050 4850
rect -600 3700 -500 4200
rect -450 3700 -350 4200
rect -300 3700 -200 4200
rect -150 3700 -50 4200
rect 0 3700 100 4200
rect 150 3700 250 4200
rect 300 3700 400 4200
rect 450 3700 550 4200
rect 600 3700 700 4200
rect 750 3700 850 4200
rect 900 3700 1000 4200
rect 1050 3700 1150 4200
rect 1200 3700 1300 4200
rect 1350 3700 1450 4200
rect 1500 3700 1600 4200
rect 1650 3700 1750 4200
rect 1800 3700 1900 4200
rect 1950 3700 2050 4200
rect 2100 3700 2200 4200
rect 2250 3700 2350 4200
rect 2400 3700 2500 4200
rect 2550 3700 2650 4200
rect 2700 3700 2800 4200
rect 2850 3700 2950 4200
rect 3000 3700 3100 4200
rect 3150 3700 3250 4200
rect 3300 3700 3400 4200
rect 3450 3700 3550 4200
rect 3600 3700 3700 4200
rect 3750 3700 3850 4200
rect 3900 3700 4000 4200
rect 4050 3700 4150 4200
rect 4200 3700 4300 4200
rect 4350 3700 4450 4200
rect 4500 3700 4600 4200
rect 4650 3700 4750 4200
rect 4800 3700 4900 4200
rect 4950 3700 5050 4200
rect 5100 3700 5200 4200
rect 5250 3700 5350 4200
rect 5400 3700 5500 4200
rect 5550 3700 5650 4200
rect 5700 3700 5800 4200
rect 5850 3700 5950 4200
rect 6000 3700 6100 4200
rect 6150 3700 6250 4200
rect 6300 3700 6400 4200
rect 6450 3700 6550 4200
rect 6600 3700 6700 4200
rect 6750 3700 6850 4200
rect 6900 3700 7000 4200
rect 7050 3700 7150 4200
rect 7200 3700 7300 4200
rect 7350 3700 7450 4200
rect 7500 3700 7600 4200
rect 7650 3700 7750 4200
rect 7800 3700 7900 4200
rect 7950 3700 8050 4200
rect 8100 3700 8200 4200
rect 8250 3700 8350 4200
rect 8400 3700 8500 4200
rect 8550 3700 8650 4200
rect 8700 3700 8800 4200
rect 8850 3700 8950 4200
rect 9000 3700 9100 4200
rect 9150 3700 9250 4200
rect 9300 3700 9400 4200
rect 9450 3700 9550 4200
rect 9600 3700 9700 4200
rect 9750 3700 9850 4200
rect 9900 3700 10000 4200
rect 10050 3700 10150 4200
rect 10200 3700 10300 4200
rect 10350 3700 10450 4200
rect 10500 3700 10600 4200
rect 10650 3700 10750 4200
rect 10800 3700 10900 4200
rect 10950 3700 11050 4200
rect 11100 3700 11200 4200
rect 11250 3700 11350 4200
rect 11400 3700 11500 4200
rect 11550 3700 11650 4200
rect 11700 3700 11800 4200
rect 11850 3700 11950 4200
rect 12000 3700 12100 4200
rect 12150 3700 12250 4200
rect 12300 3700 12400 4200
rect 12450 3700 12550 4200
rect 12600 3700 12700 4200
rect 12750 3700 12850 4200
rect 12900 3700 13000 4200
rect 13050 3700 13150 4200
rect 13200 3700 13300 4200
rect 13350 3700 13450 4200
rect 13500 3700 13600 4200
rect 13650 3700 13750 4200
rect 13800 3700 13900 4200
rect 13950 3700 14050 4200
rect 14100 3700 14200 4200
rect 14250 3700 14350 4200
rect 14400 3700 14500 4200
rect 14550 3700 14650 4200
rect 14700 3700 14800 4200
rect 14850 3700 14950 4200
rect 15000 3700 15100 4200
rect 15150 3700 15250 4200
rect 15300 3700 15400 4200
rect 15450 3700 15550 4200
rect 15600 3700 15700 4200
rect 15750 3700 15850 4200
rect 15900 3700 16000 4200
rect 16050 3700 16150 4200
rect 16200 3700 16300 4200
rect 16350 3700 16450 4200
rect 16500 3700 16600 4200
rect 16650 3700 16750 4200
rect 16800 3700 16900 4200
rect 16950 3700 17050 4200
rect 17100 3700 17200 4200
rect 17250 3700 17350 4200
rect 17400 3700 17500 4200
rect 17550 3700 17650 4200
rect 17700 3700 17800 4200
rect 17850 3700 17950 4200
rect 18000 3700 18100 4200
rect 18150 3700 18250 4200
rect 18300 3700 18400 4200
rect 18450 3700 18550 4200
rect 18600 3700 18700 4200
rect 18750 3700 18850 4200
rect 18900 3700 19000 4200
rect 19050 3700 19150 4200
rect 19200 3700 19300 4200
rect 19350 3700 19450 4200
rect 19500 3700 19600 4200
rect 19650 3700 19750 4200
rect 19800 3700 19900 4200
rect 19950 3700 20050 4200
rect 20100 3700 20200 4200
rect 20250 3700 20350 4200
rect 20400 3700 20500 4200
rect 20550 3700 20650 4200
rect 20700 3700 20800 4200
rect 20850 3700 20950 4200
rect 21000 3700 21100 4200
rect 21150 3700 21250 4200
rect 21300 3700 21400 4200
rect 21450 3700 21550 4200
rect 21600 3700 21700 4200
rect 21750 3700 21850 4200
rect 21900 3700 22000 4200
rect 22050 3700 22150 4200
rect 22200 3700 22300 4200
rect 22350 3700 22450 4200
rect 22500 3700 22600 4200
rect 22650 3700 22750 4200
rect 22800 3700 22900 4200
rect 22950 3700 23050 4200
rect 23100 3700 23200 4200
rect 23250 3700 23350 4200
rect 23400 3700 23500 4200
rect 23550 3700 23650 4200
rect 23700 3700 23800 4200
rect 23850 3700 23950 4200
rect 24000 3700 24100 4200
rect 24150 3700 24250 4200
rect 24300 3700 24400 4200
rect 24450 3700 24550 4200
rect 24600 3700 24700 4200
rect 24750 3700 24850 4200
rect 24900 3700 25000 4200
rect 25050 3700 25150 4200
rect 25200 3700 25300 4200
rect 25350 3700 25450 4200
rect 25500 3700 25600 4200
rect 25650 3700 25750 4200
rect 25800 3700 25900 4200
rect 25950 3700 26050 4200
rect 26100 3700 26200 4200
rect 26250 3700 26350 4200
rect 26400 3700 26500 4200
rect 26550 3700 26650 4200
rect 26700 3700 26800 4200
rect 26850 3700 26950 4200
rect 27000 3700 27100 4200
rect 27150 3700 27250 4200
rect 27300 3700 27400 4200
rect 27450 3700 27550 4200
rect 27600 3700 27700 4200
rect 27750 3700 27850 4200
rect 27900 3700 28000 4200
rect 28050 3700 28150 4200
rect 28200 3700 28300 4200
rect 28350 3700 28450 4200
rect 28500 3700 28600 4200
rect 28650 3700 28750 4200
rect 28800 3700 28900 4200
rect 28950 3700 29050 4200
rect 29100 3700 29200 4200
rect 29250 3700 29350 4200
rect 29400 3700 29500 4200
rect 29550 3700 29650 4200
rect 29700 3700 29800 4200
rect 29850 3700 29950 4200
rect 30000 3700 30100 4200
rect 30150 3700 30250 4200
rect 30300 3700 30400 4200
rect 30450 3700 30550 4200
rect 30600 3700 30700 4200
rect 30750 3700 30850 4200
rect 30900 3700 31000 4200
rect 31050 3700 31150 4200
rect 31200 3700 31300 4200
rect 31350 3700 31450 4200
rect 31500 3700 31600 4200
rect 31650 3700 31750 4200
rect 31800 3700 31900 4200
rect 31950 3700 32050 4200
rect -600 3050 -500 3550
rect -450 3050 -350 3550
rect -300 3050 -200 3550
rect -150 3050 -50 3550
rect 0 3050 100 3550
rect 150 3050 250 3550
rect 300 3050 400 3550
rect 450 3050 550 3550
rect 600 3050 700 3550
rect 750 3050 850 3550
rect 900 3050 1000 3550
rect 1050 3050 1150 3550
rect 1200 3050 1300 3550
rect 1350 3050 1450 3550
rect 1500 3050 1600 3550
rect 1650 3050 1750 3550
rect 1800 3050 1900 3550
rect 1950 3050 2050 3550
rect 2100 3050 2200 3550
rect 2250 3050 2350 3550
rect 2400 3050 2500 3550
rect 2550 3050 2650 3550
rect 2700 3050 2800 3550
rect 2850 3050 2950 3550
rect 3000 3050 3100 3550
rect 3150 3050 3250 3550
rect 3300 3050 3400 3550
rect 3450 3050 3550 3550
rect 3600 3050 3700 3550
rect 3750 3050 3850 3550
rect 3900 3050 4000 3550
rect 4050 3050 4150 3550
rect 4200 3050 4300 3550
rect 4350 3050 4450 3550
rect 4500 3050 4600 3550
rect 4650 3050 4750 3550
rect 4800 3050 4900 3550
rect 4950 3050 5050 3550
rect 5100 3050 5200 3550
rect 5250 3050 5350 3550
rect 5400 3050 5500 3550
rect 5550 3050 5650 3550
rect 5700 3050 5800 3550
rect 5850 3050 5950 3550
rect 6000 3050 6100 3550
rect 6150 3050 6250 3550
rect 6300 3050 6400 3550
rect 6450 3050 6550 3550
rect 6600 3050 6700 3550
rect 6750 3050 6850 3550
rect 6900 3050 7000 3550
rect 7050 3050 7150 3550
rect 7200 3050 7300 3550
rect 7350 3050 7450 3550
rect 7500 3050 7600 3550
rect 7650 3050 7750 3550
rect 7800 3050 7900 3550
rect 7950 3050 8050 3550
rect 8100 3050 8200 3550
rect 8250 3050 8350 3550
rect 8400 3050 8500 3550
rect 8550 3050 8650 3550
rect 8700 3050 8800 3550
rect 8850 3050 8950 3550
rect 9000 3050 9100 3550
rect 9150 3050 9250 3550
rect 9300 3050 9400 3550
rect 9450 3050 9550 3550
rect 9600 3050 9700 3550
rect 9750 3050 9850 3550
rect 9900 3050 10000 3550
rect 10050 3050 10150 3550
rect 10200 3050 10300 3550
rect 10350 3050 10450 3550
rect 10500 3050 10600 3550
rect 10650 3050 10750 3550
rect 10800 3050 10900 3550
rect 10950 3050 11050 3550
rect 11100 3050 11200 3550
rect 11250 3050 11350 3550
rect 11400 3050 11500 3550
rect 11550 3050 11650 3550
rect 11700 3050 11800 3550
rect 11850 3050 11950 3550
rect 12000 3050 12100 3550
rect 12150 3050 12250 3550
rect 12300 3050 12400 3550
rect 12450 3050 12550 3550
rect 12600 3050 12700 3550
rect 12750 3050 12850 3550
rect 12900 3050 13000 3550
rect 13050 3050 13150 3550
rect 13200 3050 13300 3550
rect 13350 3050 13450 3550
rect 13500 3050 13600 3550
rect 13650 3050 13750 3550
rect 13800 3050 13900 3550
rect 13950 3050 14050 3550
rect 14100 3050 14200 3550
rect 14250 3050 14350 3550
rect 14400 3050 14500 3550
rect 14550 3050 14650 3550
rect 14700 3050 14800 3550
rect 14850 3050 14950 3550
rect 15000 3050 15100 3550
rect 15150 3050 15250 3550
rect 15300 3050 15400 3550
rect 15450 3050 15550 3550
rect 15600 3050 15700 3550
rect 15750 3050 15850 3550
rect 15900 3050 16000 3550
rect 16050 3050 16150 3550
rect 16200 3050 16300 3550
rect 16350 3050 16450 3550
rect 16500 3050 16600 3550
rect 16650 3050 16750 3550
rect 16800 3050 16900 3550
rect 16950 3050 17050 3550
rect 17100 3050 17200 3550
rect 17250 3050 17350 3550
rect 17400 3050 17500 3550
rect 17550 3050 17650 3550
rect 17700 3050 17800 3550
rect 17850 3050 17950 3550
rect 18000 3050 18100 3550
rect 18150 3050 18250 3550
rect 18300 3050 18400 3550
rect 18450 3050 18550 3550
rect 18600 3050 18700 3550
rect 18750 3050 18850 3550
rect 18900 3050 19000 3550
rect 19050 3050 19150 3550
rect 19200 3050 19300 3550
rect 19350 3050 19450 3550
rect 19500 3050 19600 3550
rect 19650 3050 19750 3550
rect 19800 3050 19900 3550
rect 19950 3050 20050 3550
rect 20100 3050 20200 3550
rect 20250 3050 20350 3550
rect 20400 3050 20500 3550
rect 20550 3050 20650 3550
rect 20700 3050 20800 3550
rect 20850 3050 20950 3550
rect 21000 3050 21100 3550
rect 21150 3050 21250 3550
rect 21300 3050 21400 3550
rect 21450 3050 21550 3550
rect 21600 3050 21700 3550
rect 21750 3050 21850 3550
rect 21900 3050 22000 3550
rect 22050 3050 22150 3550
rect 22200 3050 22300 3550
rect 22350 3050 22450 3550
rect 22500 3050 22600 3550
rect 22650 3050 22750 3550
rect 22800 3050 22900 3550
rect 22950 3050 23050 3550
rect 23100 3050 23200 3550
rect 23250 3050 23350 3550
rect 23400 3050 23500 3550
rect 23550 3050 23650 3550
rect 23700 3050 23800 3550
rect 23850 3050 23950 3550
rect 24000 3050 24100 3550
rect 24150 3050 24250 3550
rect 24300 3050 24400 3550
rect 24450 3050 24550 3550
rect 24600 3050 24700 3550
rect 24750 3050 24850 3550
rect 24900 3050 25000 3550
rect 25050 3050 25150 3550
rect 25200 3050 25300 3550
rect 25350 3050 25450 3550
rect 25500 3050 25600 3550
rect 25650 3050 25750 3550
rect 25800 3050 25900 3550
rect 25950 3050 26050 3550
rect 26100 3050 26200 3550
rect 26250 3050 26350 3550
rect 26400 3050 26500 3550
rect 26550 3050 26650 3550
rect 26700 3050 26800 3550
rect 26850 3050 26950 3550
rect 27000 3050 27100 3550
rect 27150 3050 27250 3550
rect 27300 3050 27400 3550
rect 27450 3050 27550 3550
rect 27600 3050 27700 3550
rect 27750 3050 27850 3550
rect 27900 3050 28000 3550
rect 28050 3050 28150 3550
rect 28200 3050 28300 3550
rect 28350 3050 28450 3550
rect 28500 3050 28600 3550
rect 28650 3050 28750 3550
rect 28800 3050 28900 3550
rect 28950 3050 29050 3550
rect 29100 3050 29200 3550
rect 29250 3050 29350 3550
rect 29400 3050 29500 3550
rect 29550 3050 29650 3550
rect 29700 3050 29800 3550
rect 29850 3050 29950 3550
rect 30000 3050 30100 3550
rect 30150 3050 30250 3550
rect 30300 3050 30400 3550
rect 30450 3050 30550 3550
rect 30600 3050 30700 3550
rect 30750 3050 30850 3550
rect 30900 3050 31000 3550
rect 31050 3050 31150 3550
rect 31200 3050 31300 3550
rect 31350 3050 31450 3550
rect 31500 3050 31600 3550
rect 31650 3050 31750 3550
rect 31800 3050 31900 3550
rect 31950 3050 32050 3550
<< mvndiff >>
rect -650 1585 -600 1600
rect -650 1565 -635 1585
rect -615 1565 -600 1585
rect -650 1535 -600 1565
rect -650 1515 -635 1535
rect -615 1515 -600 1535
rect -650 1485 -600 1515
rect -650 1465 -635 1485
rect -615 1465 -600 1485
rect -650 1435 -600 1465
rect -650 1415 -635 1435
rect -615 1415 -600 1435
rect -650 1385 -600 1415
rect -650 1365 -635 1385
rect -615 1365 -600 1385
rect -650 1335 -600 1365
rect -650 1315 -635 1335
rect -615 1315 -600 1335
rect -650 1285 -600 1315
rect -650 1265 -635 1285
rect -615 1265 -600 1285
rect -650 1235 -600 1265
rect -650 1215 -635 1235
rect -615 1215 -600 1235
rect -650 1185 -600 1215
rect -650 1165 -635 1185
rect -615 1165 -600 1185
rect -650 1135 -600 1165
rect -650 1115 -635 1135
rect -615 1115 -600 1135
rect -650 1085 -600 1115
rect -650 1065 -635 1085
rect -615 1065 -600 1085
rect -650 1035 -600 1065
rect -650 1015 -635 1035
rect -615 1015 -600 1035
rect -650 985 -600 1015
rect -650 965 -635 985
rect -615 965 -600 985
rect -650 935 -600 965
rect -650 915 -635 935
rect -615 915 -600 935
rect -650 900 -600 915
rect -500 1585 -450 1600
rect -500 1565 -485 1585
rect -465 1565 -450 1585
rect -500 1535 -450 1565
rect -500 1515 -485 1535
rect -465 1515 -450 1535
rect -500 1485 -450 1515
rect -500 1465 -485 1485
rect -465 1465 -450 1485
rect -500 1435 -450 1465
rect -500 1415 -485 1435
rect -465 1415 -450 1435
rect -500 1385 -450 1415
rect -500 1365 -485 1385
rect -465 1365 -450 1385
rect -500 1335 -450 1365
rect -500 1315 -485 1335
rect -465 1315 -450 1335
rect -500 1285 -450 1315
rect -500 1265 -485 1285
rect -465 1265 -450 1285
rect -500 1235 -450 1265
rect -500 1215 -485 1235
rect -465 1215 -450 1235
rect -500 1185 -450 1215
rect -500 1165 -485 1185
rect -465 1165 -450 1185
rect -500 1135 -450 1165
rect -500 1115 -485 1135
rect -465 1115 -450 1135
rect -500 1085 -450 1115
rect -500 1065 -485 1085
rect -465 1065 -450 1085
rect -500 1035 -450 1065
rect -500 1015 -485 1035
rect -465 1015 -450 1035
rect -500 985 -450 1015
rect -500 965 -485 985
rect -465 965 -450 985
rect -500 935 -450 965
rect -500 915 -485 935
rect -465 915 -450 935
rect -500 900 -450 915
rect -350 1585 -300 1600
rect -350 1565 -335 1585
rect -315 1565 -300 1585
rect -350 1535 -300 1565
rect -350 1515 -335 1535
rect -315 1515 -300 1535
rect -350 1485 -300 1515
rect -350 1465 -335 1485
rect -315 1465 -300 1485
rect -350 1435 -300 1465
rect -350 1415 -335 1435
rect -315 1415 -300 1435
rect -350 1385 -300 1415
rect -350 1365 -335 1385
rect -315 1365 -300 1385
rect -350 1335 -300 1365
rect -350 1315 -335 1335
rect -315 1315 -300 1335
rect -350 1285 -300 1315
rect -350 1265 -335 1285
rect -315 1265 -300 1285
rect -350 1235 -300 1265
rect -350 1215 -335 1235
rect -315 1215 -300 1235
rect -350 1185 -300 1215
rect -350 1165 -335 1185
rect -315 1165 -300 1185
rect -350 1135 -300 1165
rect -350 1115 -335 1135
rect -315 1115 -300 1135
rect -350 1085 -300 1115
rect -350 1065 -335 1085
rect -315 1065 -300 1085
rect -350 1035 -300 1065
rect -350 1015 -335 1035
rect -315 1015 -300 1035
rect -350 985 -300 1015
rect -350 965 -335 985
rect -315 965 -300 985
rect -350 935 -300 965
rect -350 915 -335 935
rect -315 915 -300 935
rect -350 900 -300 915
rect -200 1585 -150 1600
rect -200 1565 -185 1585
rect -165 1565 -150 1585
rect -200 1535 -150 1565
rect -200 1515 -185 1535
rect -165 1515 -150 1535
rect -200 1485 -150 1515
rect -200 1465 -185 1485
rect -165 1465 -150 1485
rect -200 1435 -150 1465
rect -200 1415 -185 1435
rect -165 1415 -150 1435
rect -200 1385 -150 1415
rect -200 1365 -185 1385
rect -165 1365 -150 1385
rect -200 1335 -150 1365
rect -200 1315 -185 1335
rect -165 1315 -150 1335
rect -200 1285 -150 1315
rect -200 1265 -185 1285
rect -165 1265 -150 1285
rect -200 1235 -150 1265
rect -200 1215 -185 1235
rect -165 1215 -150 1235
rect -200 1185 -150 1215
rect -200 1165 -185 1185
rect -165 1165 -150 1185
rect -200 1135 -150 1165
rect -200 1115 -185 1135
rect -165 1115 -150 1135
rect -200 1085 -150 1115
rect -200 1065 -185 1085
rect -165 1065 -150 1085
rect -200 1035 -150 1065
rect -200 1015 -185 1035
rect -165 1015 -150 1035
rect -200 985 -150 1015
rect -200 965 -185 985
rect -165 965 -150 985
rect -200 935 -150 965
rect -200 915 -185 935
rect -165 915 -150 935
rect -200 900 -150 915
rect -50 1585 0 1600
rect -50 1565 -35 1585
rect -15 1565 0 1585
rect -50 1535 0 1565
rect -50 1515 -35 1535
rect -15 1515 0 1535
rect -50 1485 0 1515
rect -50 1465 -35 1485
rect -15 1465 0 1485
rect -50 1435 0 1465
rect -50 1415 -35 1435
rect -15 1415 0 1435
rect -50 1385 0 1415
rect -50 1365 -35 1385
rect -15 1365 0 1385
rect -50 1335 0 1365
rect -50 1315 -35 1335
rect -15 1315 0 1335
rect -50 1285 0 1315
rect -50 1265 -35 1285
rect -15 1265 0 1285
rect -50 1235 0 1265
rect -50 1215 -35 1235
rect -15 1215 0 1235
rect -50 1185 0 1215
rect -50 1165 -35 1185
rect -15 1165 0 1185
rect -50 1135 0 1165
rect -50 1115 -35 1135
rect -15 1115 0 1135
rect -50 1085 0 1115
rect -50 1065 -35 1085
rect -15 1065 0 1085
rect -50 1035 0 1065
rect -50 1015 -35 1035
rect -15 1015 0 1035
rect -50 985 0 1015
rect -50 965 -35 985
rect -15 965 0 985
rect -50 935 0 965
rect -50 915 -35 935
rect -15 915 0 935
rect -50 900 0 915
rect 100 900 150 1600
rect 250 900 300 1600
rect 400 900 450 1600
rect 550 900 600 1600
rect 700 900 750 1600
rect 850 900 900 1600
rect 1000 900 1050 1600
rect 1150 1585 1200 1600
rect 1150 1565 1165 1585
rect 1185 1565 1200 1585
rect 1150 1535 1200 1565
rect 1150 1515 1165 1535
rect 1185 1515 1200 1535
rect 1150 1485 1200 1515
rect 1150 1465 1165 1485
rect 1185 1465 1200 1485
rect 1150 1435 1200 1465
rect 1150 1415 1165 1435
rect 1185 1415 1200 1435
rect 1150 1385 1200 1415
rect 1150 1365 1165 1385
rect 1185 1365 1200 1385
rect 1150 1335 1200 1365
rect 1150 1315 1165 1335
rect 1185 1315 1200 1335
rect 1150 1285 1200 1315
rect 1150 1265 1165 1285
rect 1185 1265 1200 1285
rect 1150 1235 1200 1265
rect 1150 1215 1165 1235
rect 1185 1215 1200 1235
rect 1150 1185 1200 1215
rect 1150 1165 1165 1185
rect 1185 1165 1200 1185
rect 1150 1135 1200 1165
rect 1150 1115 1165 1135
rect 1185 1115 1200 1135
rect 1150 1085 1200 1115
rect 1150 1065 1165 1085
rect 1185 1065 1200 1085
rect 1150 1035 1200 1065
rect 1150 1015 1165 1035
rect 1185 1015 1200 1035
rect 1150 985 1200 1015
rect 1150 965 1165 985
rect 1185 965 1200 985
rect 1150 935 1200 965
rect 1150 915 1165 935
rect 1185 915 1200 935
rect 1150 900 1200 915
rect 1300 900 1350 1600
rect 1450 1585 1500 1600
rect 1450 1565 1465 1585
rect 1485 1565 1500 1585
rect 1450 1535 1500 1565
rect 1450 1515 1465 1535
rect 1485 1515 1500 1535
rect 1450 1485 1500 1515
rect 1450 1465 1465 1485
rect 1485 1465 1500 1485
rect 1450 1435 1500 1465
rect 1450 1415 1465 1435
rect 1485 1415 1500 1435
rect 1450 1385 1500 1415
rect 1450 1365 1465 1385
rect 1485 1365 1500 1385
rect 1450 1335 1500 1365
rect 1450 1315 1465 1335
rect 1485 1315 1500 1335
rect 1450 1285 1500 1315
rect 1450 1265 1465 1285
rect 1485 1265 1500 1285
rect 1450 1235 1500 1265
rect 1450 1215 1465 1235
rect 1485 1215 1500 1235
rect 1450 1185 1500 1215
rect 1450 1165 1465 1185
rect 1485 1165 1500 1185
rect 1450 1135 1500 1165
rect 1450 1115 1465 1135
rect 1485 1115 1500 1135
rect 1450 1085 1500 1115
rect 1450 1065 1465 1085
rect 1485 1065 1500 1085
rect 1450 1035 1500 1065
rect 1450 1015 1465 1035
rect 1485 1015 1500 1035
rect 1450 985 1500 1015
rect 1450 965 1465 985
rect 1485 965 1500 985
rect 1450 935 1500 965
rect 1450 915 1465 935
rect 1485 915 1500 935
rect 1450 900 1500 915
rect 1600 900 1650 1600
rect 1750 1585 1800 1600
rect 1750 1565 1765 1585
rect 1785 1565 1800 1585
rect 1750 1535 1800 1565
rect 1750 1515 1765 1535
rect 1785 1515 1800 1535
rect 1750 1485 1800 1515
rect 1750 1465 1765 1485
rect 1785 1465 1800 1485
rect 1750 1435 1800 1465
rect 1750 1415 1765 1435
rect 1785 1415 1800 1435
rect 1750 1385 1800 1415
rect 1750 1365 1765 1385
rect 1785 1365 1800 1385
rect 1750 1335 1800 1365
rect 1750 1315 1765 1335
rect 1785 1315 1800 1335
rect 1750 1285 1800 1315
rect 1750 1265 1765 1285
rect 1785 1265 1800 1285
rect 1750 1235 1800 1265
rect 1750 1215 1765 1235
rect 1785 1215 1800 1235
rect 1750 1185 1800 1215
rect 1750 1165 1765 1185
rect 1785 1165 1800 1185
rect 1750 1135 1800 1165
rect 1750 1115 1765 1135
rect 1785 1115 1800 1135
rect 1750 1085 1800 1115
rect 1750 1065 1765 1085
rect 1785 1065 1800 1085
rect 1750 1035 1800 1065
rect 1750 1015 1765 1035
rect 1785 1015 1800 1035
rect 1750 985 1800 1015
rect 1750 965 1765 985
rect 1785 965 1800 985
rect 1750 935 1800 965
rect 1750 915 1765 935
rect 1785 915 1800 935
rect 1750 900 1800 915
rect 1900 900 1950 1600
rect 2050 1585 2100 1600
rect 2050 1565 2065 1585
rect 2085 1565 2100 1585
rect 2050 1535 2100 1565
rect 2050 1515 2065 1535
rect 2085 1515 2100 1535
rect 2050 1485 2100 1515
rect 2050 1465 2065 1485
rect 2085 1465 2100 1485
rect 2050 1435 2100 1465
rect 2050 1415 2065 1435
rect 2085 1415 2100 1435
rect 2050 1385 2100 1415
rect 2050 1365 2065 1385
rect 2085 1365 2100 1385
rect 2050 1335 2100 1365
rect 2050 1315 2065 1335
rect 2085 1315 2100 1335
rect 2050 1285 2100 1315
rect 2050 1265 2065 1285
rect 2085 1265 2100 1285
rect 2050 1235 2100 1265
rect 2050 1215 2065 1235
rect 2085 1215 2100 1235
rect 2050 1185 2100 1215
rect 2050 1165 2065 1185
rect 2085 1165 2100 1185
rect 2050 1135 2100 1165
rect 2050 1115 2065 1135
rect 2085 1115 2100 1135
rect 2050 1085 2100 1115
rect 2050 1065 2065 1085
rect 2085 1065 2100 1085
rect 2050 1035 2100 1065
rect 2050 1015 2065 1035
rect 2085 1015 2100 1035
rect 2050 985 2100 1015
rect 2050 965 2065 985
rect 2085 965 2100 985
rect 2050 935 2100 965
rect 2050 915 2065 935
rect 2085 915 2100 935
rect 2050 900 2100 915
rect 2200 900 2250 1600
rect 2350 1585 2400 1600
rect 2350 1565 2365 1585
rect 2385 1565 2400 1585
rect 2350 1535 2400 1565
rect 2350 1515 2365 1535
rect 2385 1515 2400 1535
rect 2350 1485 2400 1515
rect 2350 1465 2365 1485
rect 2385 1465 2400 1485
rect 2350 1435 2400 1465
rect 2350 1415 2365 1435
rect 2385 1415 2400 1435
rect 2350 1385 2400 1415
rect 2350 1365 2365 1385
rect 2385 1365 2400 1385
rect 2350 1335 2400 1365
rect 2350 1315 2365 1335
rect 2385 1315 2400 1335
rect 2350 1285 2400 1315
rect 2350 1265 2365 1285
rect 2385 1265 2400 1285
rect 2350 1235 2400 1265
rect 2350 1215 2365 1235
rect 2385 1215 2400 1235
rect 2350 1185 2400 1215
rect 2350 1165 2365 1185
rect 2385 1165 2400 1185
rect 2350 1135 2400 1165
rect 2350 1115 2365 1135
rect 2385 1115 2400 1135
rect 2350 1085 2400 1115
rect 2350 1065 2365 1085
rect 2385 1065 2400 1085
rect 2350 1035 2400 1065
rect 2350 1015 2365 1035
rect 2385 1015 2400 1035
rect 2350 985 2400 1015
rect 2350 965 2365 985
rect 2385 965 2400 985
rect 2350 935 2400 965
rect 2350 915 2365 935
rect 2385 915 2400 935
rect 2350 900 2400 915
rect 2500 900 2550 1600
rect 2650 1585 2700 1600
rect 2650 1565 2665 1585
rect 2685 1565 2700 1585
rect 2650 1535 2700 1565
rect 2650 1515 2665 1535
rect 2685 1515 2700 1535
rect 2650 1485 2700 1515
rect 2650 1465 2665 1485
rect 2685 1465 2700 1485
rect 2650 1435 2700 1465
rect 2650 1415 2665 1435
rect 2685 1415 2700 1435
rect 2650 1385 2700 1415
rect 2650 1365 2665 1385
rect 2685 1365 2700 1385
rect 2650 1335 2700 1365
rect 2650 1315 2665 1335
rect 2685 1315 2700 1335
rect 2650 1285 2700 1315
rect 2650 1265 2665 1285
rect 2685 1265 2700 1285
rect 2650 1235 2700 1265
rect 2650 1215 2665 1235
rect 2685 1215 2700 1235
rect 2650 1185 2700 1215
rect 2650 1165 2665 1185
rect 2685 1165 2700 1185
rect 2650 1135 2700 1165
rect 2650 1115 2665 1135
rect 2685 1115 2700 1135
rect 2650 1085 2700 1115
rect 2650 1065 2665 1085
rect 2685 1065 2700 1085
rect 2650 1035 2700 1065
rect 2650 1015 2665 1035
rect 2685 1015 2700 1035
rect 2650 985 2700 1015
rect 2650 965 2665 985
rect 2685 965 2700 985
rect 2650 935 2700 965
rect 2650 915 2665 935
rect 2685 915 2700 935
rect 2650 900 2700 915
rect 2800 900 2850 1600
rect 2950 1585 3000 1600
rect 2950 1565 2965 1585
rect 2985 1565 3000 1585
rect 2950 1535 3000 1565
rect 2950 1515 2965 1535
rect 2985 1515 3000 1535
rect 2950 1485 3000 1515
rect 2950 1465 2965 1485
rect 2985 1465 3000 1485
rect 2950 1435 3000 1465
rect 2950 1415 2965 1435
rect 2985 1415 3000 1435
rect 2950 1385 3000 1415
rect 2950 1365 2965 1385
rect 2985 1365 3000 1385
rect 2950 1335 3000 1365
rect 2950 1315 2965 1335
rect 2985 1315 3000 1335
rect 2950 1285 3000 1315
rect 2950 1265 2965 1285
rect 2985 1265 3000 1285
rect 2950 1235 3000 1265
rect 2950 1215 2965 1235
rect 2985 1215 3000 1235
rect 2950 1185 3000 1215
rect 2950 1165 2965 1185
rect 2985 1165 3000 1185
rect 2950 1135 3000 1165
rect 2950 1115 2965 1135
rect 2985 1115 3000 1135
rect 2950 1085 3000 1115
rect 2950 1065 2965 1085
rect 2985 1065 3000 1085
rect 2950 1035 3000 1065
rect 2950 1015 2965 1035
rect 2985 1015 3000 1035
rect 2950 985 3000 1015
rect 2950 965 2965 985
rect 2985 965 3000 985
rect 2950 935 3000 965
rect 2950 915 2965 935
rect 2985 915 3000 935
rect 2950 900 3000 915
rect 3100 900 3150 1600
rect 3250 1585 3300 1600
rect 3250 1565 3265 1585
rect 3285 1565 3300 1585
rect 3250 1535 3300 1565
rect 3250 1515 3265 1535
rect 3285 1515 3300 1535
rect 3250 1485 3300 1515
rect 3250 1465 3265 1485
rect 3285 1465 3300 1485
rect 3250 1435 3300 1465
rect 3250 1415 3265 1435
rect 3285 1415 3300 1435
rect 3250 1385 3300 1415
rect 3250 1365 3265 1385
rect 3285 1365 3300 1385
rect 3250 1335 3300 1365
rect 3250 1315 3265 1335
rect 3285 1315 3300 1335
rect 3250 1285 3300 1315
rect 3250 1265 3265 1285
rect 3285 1265 3300 1285
rect 3250 1235 3300 1265
rect 3250 1215 3265 1235
rect 3285 1215 3300 1235
rect 3250 1185 3300 1215
rect 3250 1165 3265 1185
rect 3285 1165 3300 1185
rect 3250 1135 3300 1165
rect 3250 1115 3265 1135
rect 3285 1115 3300 1135
rect 3250 1085 3300 1115
rect 3250 1065 3265 1085
rect 3285 1065 3300 1085
rect 3250 1035 3300 1065
rect 3250 1015 3265 1035
rect 3285 1015 3300 1035
rect 3250 985 3300 1015
rect 3250 965 3265 985
rect 3285 965 3300 985
rect 3250 935 3300 965
rect 3250 915 3265 935
rect 3285 915 3300 935
rect 3250 900 3300 915
rect 3400 900 3450 1600
rect 3550 1585 3600 1600
rect 3550 1565 3565 1585
rect 3585 1565 3600 1585
rect 3550 1535 3600 1565
rect 3550 1515 3565 1535
rect 3585 1515 3600 1535
rect 3550 1485 3600 1515
rect 3550 1465 3565 1485
rect 3585 1465 3600 1485
rect 3550 1435 3600 1465
rect 3550 1415 3565 1435
rect 3585 1415 3600 1435
rect 3550 1385 3600 1415
rect 3550 1365 3565 1385
rect 3585 1365 3600 1385
rect 3550 1335 3600 1365
rect 3550 1315 3565 1335
rect 3585 1315 3600 1335
rect 3550 1285 3600 1315
rect 3550 1265 3565 1285
rect 3585 1265 3600 1285
rect 3550 1235 3600 1265
rect 3550 1215 3565 1235
rect 3585 1215 3600 1235
rect 3550 1185 3600 1215
rect 3550 1165 3565 1185
rect 3585 1165 3600 1185
rect 3550 1135 3600 1165
rect 3550 1115 3565 1135
rect 3585 1115 3600 1135
rect 3550 1085 3600 1115
rect 3550 1065 3565 1085
rect 3585 1065 3600 1085
rect 3550 1035 3600 1065
rect 3550 1015 3565 1035
rect 3585 1015 3600 1035
rect 3550 985 3600 1015
rect 3550 965 3565 985
rect 3585 965 3600 985
rect 3550 935 3600 965
rect 3550 915 3565 935
rect 3585 915 3600 935
rect 3550 900 3600 915
rect 3700 1585 3750 1600
rect 3700 1565 3715 1585
rect 3735 1565 3750 1585
rect 3700 1535 3750 1565
rect 3700 1515 3715 1535
rect 3735 1515 3750 1535
rect 3700 1485 3750 1515
rect 3700 1465 3715 1485
rect 3735 1465 3750 1485
rect 3700 1435 3750 1465
rect 3700 1415 3715 1435
rect 3735 1415 3750 1435
rect 3700 1385 3750 1415
rect 3700 1365 3715 1385
rect 3735 1365 3750 1385
rect 3700 1335 3750 1365
rect 3700 1315 3715 1335
rect 3735 1315 3750 1335
rect 3700 1285 3750 1315
rect 3700 1265 3715 1285
rect 3735 1265 3750 1285
rect 3700 1235 3750 1265
rect 3700 1215 3715 1235
rect 3735 1215 3750 1235
rect 3700 1185 3750 1215
rect 3700 1165 3715 1185
rect 3735 1165 3750 1185
rect 3700 1135 3750 1165
rect 3700 1115 3715 1135
rect 3735 1115 3750 1135
rect 3700 1085 3750 1115
rect 3700 1065 3715 1085
rect 3735 1065 3750 1085
rect 3700 1035 3750 1065
rect 3700 1015 3715 1035
rect 3735 1015 3750 1035
rect 3700 985 3750 1015
rect 3700 965 3715 985
rect 3735 965 3750 985
rect 3700 935 3750 965
rect 3700 915 3715 935
rect 3735 915 3750 935
rect 3700 900 3750 915
rect 3850 1585 3900 1600
rect 3850 1565 3865 1585
rect 3885 1565 3900 1585
rect 3850 1535 3900 1565
rect 3850 1515 3865 1535
rect 3885 1515 3900 1535
rect 3850 1485 3900 1515
rect 3850 1465 3865 1485
rect 3885 1465 3900 1485
rect 3850 1435 3900 1465
rect 3850 1415 3865 1435
rect 3885 1415 3900 1435
rect 3850 1385 3900 1415
rect 3850 1365 3865 1385
rect 3885 1365 3900 1385
rect 3850 1335 3900 1365
rect 3850 1315 3865 1335
rect 3885 1315 3900 1335
rect 3850 1285 3900 1315
rect 3850 1265 3865 1285
rect 3885 1265 3900 1285
rect 3850 1235 3900 1265
rect 3850 1215 3865 1235
rect 3885 1215 3900 1235
rect 3850 1185 3900 1215
rect 3850 1165 3865 1185
rect 3885 1165 3900 1185
rect 3850 1135 3900 1165
rect 3850 1115 3865 1135
rect 3885 1115 3900 1135
rect 3850 1085 3900 1115
rect 3850 1065 3865 1085
rect 3885 1065 3900 1085
rect 3850 1035 3900 1065
rect 3850 1015 3865 1035
rect 3885 1015 3900 1035
rect 3850 985 3900 1015
rect 3850 965 3865 985
rect 3885 965 3900 985
rect 3850 935 3900 965
rect 3850 915 3865 935
rect 3885 915 3900 935
rect 3850 900 3900 915
rect 4000 1585 4050 1600
rect 4000 1565 4015 1585
rect 4035 1565 4050 1585
rect 4000 1535 4050 1565
rect 4000 1515 4015 1535
rect 4035 1515 4050 1535
rect 4000 1485 4050 1515
rect 4000 1465 4015 1485
rect 4035 1465 4050 1485
rect 4000 1435 4050 1465
rect 4000 1415 4015 1435
rect 4035 1415 4050 1435
rect 4000 1385 4050 1415
rect 4000 1365 4015 1385
rect 4035 1365 4050 1385
rect 4000 1335 4050 1365
rect 4000 1315 4015 1335
rect 4035 1315 4050 1335
rect 4000 1285 4050 1315
rect 4000 1265 4015 1285
rect 4035 1265 4050 1285
rect 4000 1235 4050 1265
rect 4000 1215 4015 1235
rect 4035 1215 4050 1235
rect 4000 1185 4050 1215
rect 4000 1165 4015 1185
rect 4035 1165 4050 1185
rect 4000 1135 4050 1165
rect 4000 1115 4015 1135
rect 4035 1115 4050 1135
rect 4000 1085 4050 1115
rect 4000 1065 4015 1085
rect 4035 1065 4050 1085
rect 4000 1035 4050 1065
rect 4000 1015 4015 1035
rect 4035 1015 4050 1035
rect 4000 985 4050 1015
rect 4000 965 4015 985
rect 4035 965 4050 985
rect 4000 935 4050 965
rect 4000 915 4015 935
rect 4035 915 4050 935
rect 4000 900 4050 915
rect 4150 1585 4200 1600
rect 4150 1565 4165 1585
rect 4185 1565 4200 1585
rect 4150 1535 4200 1565
rect 4150 1515 4165 1535
rect 4185 1515 4200 1535
rect 4150 1485 4200 1515
rect 4150 1465 4165 1485
rect 4185 1465 4200 1485
rect 4150 1435 4200 1465
rect 4150 1415 4165 1435
rect 4185 1415 4200 1435
rect 4150 1385 4200 1415
rect 4150 1365 4165 1385
rect 4185 1365 4200 1385
rect 4150 1335 4200 1365
rect 4150 1315 4165 1335
rect 4185 1315 4200 1335
rect 4150 1285 4200 1315
rect 4150 1265 4165 1285
rect 4185 1265 4200 1285
rect 4150 1235 4200 1265
rect 4150 1215 4165 1235
rect 4185 1215 4200 1235
rect 4150 1185 4200 1215
rect 4150 1165 4165 1185
rect 4185 1165 4200 1185
rect 4150 1135 4200 1165
rect 4150 1115 4165 1135
rect 4185 1115 4200 1135
rect 4150 1085 4200 1115
rect 4150 1065 4165 1085
rect 4185 1065 4200 1085
rect 4150 1035 4200 1065
rect 4150 1015 4165 1035
rect 4185 1015 4200 1035
rect 4150 985 4200 1015
rect 4150 965 4165 985
rect 4185 965 4200 985
rect 4150 935 4200 965
rect 4150 915 4165 935
rect 4185 915 4200 935
rect 4150 900 4200 915
rect 4300 1585 4350 1600
rect 4300 1565 4315 1585
rect 4335 1565 4350 1585
rect 4300 1535 4350 1565
rect 4300 1515 4315 1535
rect 4335 1515 4350 1535
rect 4300 1485 4350 1515
rect 4300 1465 4315 1485
rect 4335 1465 4350 1485
rect 4300 1435 4350 1465
rect 4300 1415 4315 1435
rect 4335 1415 4350 1435
rect 4300 1385 4350 1415
rect 4300 1365 4315 1385
rect 4335 1365 4350 1385
rect 4300 1335 4350 1365
rect 4300 1315 4315 1335
rect 4335 1315 4350 1335
rect 4300 1285 4350 1315
rect 4300 1265 4315 1285
rect 4335 1265 4350 1285
rect 4300 1235 4350 1265
rect 4300 1215 4315 1235
rect 4335 1215 4350 1235
rect 4300 1185 4350 1215
rect 4300 1165 4315 1185
rect 4335 1165 4350 1185
rect 4300 1135 4350 1165
rect 4300 1115 4315 1135
rect 4335 1115 4350 1135
rect 4300 1085 4350 1115
rect 4300 1065 4315 1085
rect 4335 1065 4350 1085
rect 4300 1035 4350 1065
rect 4300 1015 4315 1035
rect 4335 1015 4350 1035
rect 4300 985 4350 1015
rect 4300 965 4315 985
rect 4335 965 4350 985
rect 4300 935 4350 965
rect 4300 915 4315 935
rect 4335 915 4350 935
rect 4300 900 4350 915
rect 4450 1585 4500 1600
rect 4450 1565 4465 1585
rect 4485 1565 4500 1585
rect 4450 1535 4500 1565
rect 4450 1515 4465 1535
rect 4485 1515 4500 1535
rect 4450 1485 4500 1515
rect 4450 1465 4465 1485
rect 4485 1465 4500 1485
rect 4450 1435 4500 1465
rect 4450 1415 4465 1435
rect 4485 1415 4500 1435
rect 4450 1385 4500 1415
rect 4450 1365 4465 1385
rect 4485 1365 4500 1385
rect 4450 1335 4500 1365
rect 4450 1315 4465 1335
rect 4485 1315 4500 1335
rect 4450 1285 4500 1315
rect 4450 1265 4465 1285
rect 4485 1265 4500 1285
rect 4450 1235 4500 1265
rect 4450 1215 4465 1235
rect 4485 1215 4500 1235
rect 4450 1185 4500 1215
rect 4450 1165 4465 1185
rect 4485 1165 4500 1185
rect 4450 1135 4500 1165
rect 4450 1115 4465 1135
rect 4485 1115 4500 1135
rect 4450 1085 4500 1115
rect 4450 1065 4465 1085
rect 4485 1065 4500 1085
rect 4450 1035 4500 1065
rect 4450 1015 4465 1035
rect 4485 1015 4500 1035
rect 4450 985 4500 1015
rect 4450 965 4465 985
rect 4485 965 4500 985
rect 4450 935 4500 965
rect 4450 915 4465 935
rect 4485 915 4500 935
rect 4450 900 4500 915
rect 4600 1585 4650 1600
rect 4600 1565 4615 1585
rect 4635 1565 4650 1585
rect 4600 1535 4650 1565
rect 4600 1515 4615 1535
rect 4635 1515 4650 1535
rect 4600 1485 4650 1515
rect 4600 1465 4615 1485
rect 4635 1465 4650 1485
rect 4600 1435 4650 1465
rect 4600 1415 4615 1435
rect 4635 1415 4650 1435
rect 4600 1385 4650 1415
rect 4600 1365 4615 1385
rect 4635 1365 4650 1385
rect 4600 1335 4650 1365
rect 4600 1315 4615 1335
rect 4635 1315 4650 1335
rect 4600 1285 4650 1315
rect 4600 1265 4615 1285
rect 4635 1265 4650 1285
rect 4600 1235 4650 1265
rect 4600 1215 4615 1235
rect 4635 1215 4650 1235
rect 4600 1185 4650 1215
rect 4600 1165 4615 1185
rect 4635 1165 4650 1185
rect 4600 1135 4650 1165
rect 4600 1115 4615 1135
rect 4635 1115 4650 1135
rect 4600 1085 4650 1115
rect 4600 1065 4615 1085
rect 4635 1065 4650 1085
rect 4600 1035 4650 1065
rect 4600 1015 4615 1035
rect 4635 1015 4650 1035
rect 4600 985 4650 1015
rect 4600 965 4615 985
rect 4635 965 4650 985
rect 4600 935 4650 965
rect 4600 915 4615 935
rect 4635 915 4650 935
rect 4600 900 4650 915
rect 4750 1585 4800 1600
rect 4750 1565 4765 1585
rect 4785 1565 4800 1585
rect 4750 1535 4800 1565
rect 4750 1515 4765 1535
rect 4785 1515 4800 1535
rect 4750 1485 4800 1515
rect 4750 1465 4765 1485
rect 4785 1465 4800 1485
rect 4750 1435 4800 1465
rect 4750 1415 4765 1435
rect 4785 1415 4800 1435
rect 4750 1385 4800 1415
rect 4750 1365 4765 1385
rect 4785 1365 4800 1385
rect 4750 1335 4800 1365
rect 4750 1315 4765 1335
rect 4785 1315 4800 1335
rect 4750 1285 4800 1315
rect 4750 1265 4765 1285
rect 4785 1265 4800 1285
rect 4750 1235 4800 1265
rect 4750 1215 4765 1235
rect 4785 1215 4800 1235
rect 4750 1185 4800 1215
rect 4750 1165 4765 1185
rect 4785 1165 4800 1185
rect 4750 1135 4800 1165
rect 4750 1115 4765 1135
rect 4785 1115 4800 1135
rect 4750 1085 4800 1115
rect 4750 1065 4765 1085
rect 4785 1065 4800 1085
rect 4750 1035 4800 1065
rect 4750 1015 4765 1035
rect 4785 1015 4800 1035
rect 4750 985 4800 1015
rect 4750 965 4765 985
rect 4785 965 4800 985
rect 4750 935 4800 965
rect 4750 915 4765 935
rect 4785 915 4800 935
rect 4750 900 4800 915
rect 4900 900 4950 1600
rect 5050 1585 5100 1600
rect 5050 1565 5065 1585
rect 5085 1565 5100 1585
rect 5050 1535 5100 1565
rect 5050 1515 5065 1535
rect 5085 1515 5100 1535
rect 5050 1485 5100 1515
rect 5050 1465 5065 1485
rect 5085 1465 5100 1485
rect 5050 1435 5100 1465
rect 5050 1415 5065 1435
rect 5085 1415 5100 1435
rect 5050 1385 5100 1415
rect 5050 1365 5065 1385
rect 5085 1365 5100 1385
rect 5050 1335 5100 1365
rect 5050 1315 5065 1335
rect 5085 1315 5100 1335
rect 5050 1285 5100 1315
rect 5050 1265 5065 1285
rect 5085 1265 5100 1285
rect 5050 1235 5100 1265
rect 5050 1215 5065 1235
rect 5085 1215 5100 1235
rect 5050 1185 5100 1215
rect 5050 1165 5065 1185
rect 5085 1165 5100 1185
rect 5050 1135 5100 1165
rect 5050 1115 5065 1135
rect 5085 1115 5100 1135
rect 5050 1085 5100 1115
rect 5050 1065 5065 1085
rect 5085 1065 5100 1085
rect 5050 1035 5100 1065
rect 5050 1015 5065 1035
rect 5085 1015 5100 1035
rect 5050 985 5100 1015
rect 5050 965 5065 985
rect 5085 965 5100 985
rect 5050 935 5100 965
rect 5050 915 5065 935
rect 5085 915 5100 935
rect 5050 900 5100 915
rect 5200 900 5250 1600
rect 5350 1585 5400 1600
rect 5350 1565 5365 1585
rect 5385 1565 5400 1585
rect 5350 1535 5400 1565
rect 5350 1515 5365 1535
rect 5385 1515 5400 1535
rect 5350 1485 5400 1515
rect 5350 1465 5365 1485
rect 5385 1465 5400 1485
rect 5350 1435 5400 1465
rect 5350 1415 5365 1435
rect 5385 1415 5400 1435
rect 5350 1385 5400 1415
rect 5350 1365 5365 1385
rect 5385 1365 5400 1385
rect 5350 1335 5400 1365
rect 5350 1315 5365 1335
rect 5385 1315 5400 1335
rect 5350 1285 5400 1315
rect 5350 1265 5365 1285
rect 5385 1265 5400 1285
rect 5350 1235 5400 1265
rect 5350 1215 5365 1235
rect 5385 1215 5400 1235
rect 5350 1185 5400 1215
rect 5350 1165 5365 1185
rect 5385 1165 5400 1185
rect 5350 1135 5400 1165
rect 5350 1115 5365 1135
rect 5385 1115 5400 1135
rect 5350 1085 5400 1115
rect 5350 1065 5365 1085
rect 5385 1065 5400 1085
rect 5350 1035 5400 1065
rect 5350 1015 5365 1035
rect 5385 1015 5400 1035
rect 5350 985 5400 1015
rect 5350 965 5365 985
rect 5385 965 5400 985
rect 5350 935 5400 965
rect 5350 915 5365 935
rect 5385 915 5400 935
rect 5350 900 5400 915
rect 5500 900 5550 1600
rect 5650 1585 5700 1600
rect 5650 1565 5665 1585
rect 5685 1565 5700 1585
rect 5650 1535 5700 1565
rect 5650 1515 5665 1535
rect 5685 1515 5700 1535
rect 5650 1485 5700 1515
rect 5650 1465 5665 1485
rect 5685 1465 5700 1485
rect 5650 1435 5700 1465
rect 5650 1415 5665 1435
rect 5685 1415 5700 1435
rect 5650 1385 5700 1415
rect 5650 1365 5665 1385
rect 5685 1365 5700 1385
rect 5650 1335 5700 1365
rect 5650 1315 5665 1335
rect 5685 1315 5700 1335
rect 5650 1285 5700 1315
rect 5650 1265 5665 1285
rect 5685 1265 5700 1285
rect 5650 1235 5700 1265
rect 5650 1215 5665 1235
rect 5685 1215 5700 1235
rect 5650 1185 5700 1215
rect 5650 1165 5665 1185
rect 5685 1165 5700 1185
rect 5650 1135 5700 1165
rect 5650 1115 5665 1135
rect 5685 1115 5700 1135
rect 5650 1085 5700 1115
rect 5650 1065 5665 1085
rect 5685 1065 5700 1085
rect 5650 1035 5700 1065
rect 5650 1015 5665 1035
rect 5685 1015 5700 1035
rect 5650 985 5700 1015
rect 5650 965 5665 985
rect 5685 965 5700 985
rect 5650 935 5700 965
rect 5650 915 5665 935
rect 5685 915 5700 935
rect 5650 900 5700 915
rect 5800 900 5850 1600
rect 5950 1585 6000 1600
rect 5950 1565 5965 1585
rect 5985 1565 6000 1585
rect 5950 1535 6000 1565
rect 5950 1515 5965 1535
rect 5985 1515 6000 1535
rect 5950 1485 6000 1515
rect 5950 1465 5965 1485
rect 5985 1465 6000 1485
rect 5950 1435 6000 1465
rect 5950 1415 5965 1435
rect 5985 1415 6000 1435
rect 5950 1385 6000 1415
rect 5950 1365 5965 1385
rect 5985 1365 6000 1385
rect 5950 1335 6000 1365
rect 5950 1315 5965 1335
rect 5985 1315 6000 1335
rect 5950 1285 6000 1315
rect 5950 1265 5965 1285
rect 5985 1265 6000 1285
rect 5950 1235 6000 1265
rect 5950 1215 5965 1235
rect 5985 1215 6000 1235
rect 5950 1185 6000 1215
rect 5950 1165 5965 1185
rect 5985 1165 6000 1185
rect 5950 1135 6000 1165
rect 5950 1115 5965 1135
rect 5985 1115 6000 1135
rect 5950 1085 6000 1115
rect 5950 1065 5965 1085
rect 5985 1065 6000 1085
rect 5950 1035 6000 1065
rect 5950 1015 5965 1035
rect 5985 1015 6000 1035
rect 5950 985 6000 1015
rect 5950 965 5965 985
rect 5985 965 6000 985
rect 5950 935 6000 965
rect 5950 915 5965 935
rect 5985 915 6000 935
rect 5950 900 6000 915
rect 6100 900 6150 1600
rect 6250 1585 6300 1600
rect 6250 1565 6265 1585
rect 6285 1565 6300 1585
rect 6250 1535 6300 1565
rect 6250 1515 6265 1535
rect 6285 1515 6300 1535
rect 6250 1485 6300 1515
rect 6250 1465 6265 1485
rect 6285 1465 6300 1485
rect 6250 1435 6300 1465
rect 6250 1415 6265 1435
rect 6285 1415 6300 1435
rect 6250 1385 6300 1415
rect 6250 1365 6265 1385
rect 6285 1365 6300 1385
rect 6250 1335 6300 1365
rect 6250 1315 6265 1335
rect 6285 1315 6300 1335
rect 6250 1285 6300 1315
rect 6250 1265 6265 1285
rect 6285 1265 6300 1285
rect 6250 1235 6300 1265
rect 6250 1215 6265 1235
rect 6285 1215 6300 1235
rect 6250 1185 6300 1215
rect 6250 1165 6265 1185
rect 6285 1165 6300 1185
rect 6250 1135 6300 1165
rect 6250 1115 6265 1135
rect 6285 1115 6300 1135
rect 6250 1085 6300 1115
rect 6250 1065 6265 1085
rect 6285 1065 6300 1085
rect 6250 1035 6300 1065
rect 6250 1015 6265 1035
rect 6285 1015 6300 1035
rect 6250 985 6300 1015
rect 6250 965 6265 985
rect 6285 965 6300 985
rect 6250 935 6300 965
rect 6250 915 6265 935
rect 6285 915 6300 935
rect 6250 900 6300 915
rect 6400 900 6450 1600
rect 6550 1585 6600 1600
rect 6550 1565 6565 1585
rect 6585 1565 6600 1585
rect 6550 1535 6600 1565
rect 6550 1515 6565 1535
rect 6585 1515 6600 1535
rect 6550 1485 6600 1515
rect 6550 1465 6565 1485
rect 6585 1465 6600 1485
rect 6550 1435 6600 1465
rect 6550 1415 6565 1435
rect 6585 1415 6600 1435
rect 6550 1385 6600 1415
rect 6550 1365 6565 1385
rect 6585 1365 6600 1385
rect 6550 1335 6600 1365
rect 6550 1315 6565 1335
rect 6585 1315 6600 1335
rect 6550 1285 6600 1315
rect 6550 1265 6565 1285
rect 6585 1265 6600 1285
rect 6550 1235 6600 1265
rect 6550 1215 6565 1235
rect 6585 1215 6600 1235
rect 6550 1185 6600 1215
rect 6550 1165 6565 1185
rect 6585 1165 6600 1185
rect 6550 1135 6600 1165
rect 6550 1115 6565 1135
rect 6585 1115 6600 1135
rect 6550 1085 6600 1115
rect 6550 1065 6565 1085
rect 6585 1065 6600 1085
rect 6550 1035 6600 1065
rect 6550 1015 6565 1035
rect 6585 1015 6600 1035
rect 6550 985 6600 1015
rect 6550 965 6565 985
rect 6585 965 6600 985
rect 6550 935 6600 965
rect 6550 915 6565 935
rect 6585 915 6600 935
rect 6550 900 6600 915
rect 6700 900 6750 1600
rect 6850 1585 6900 1600
rect 6850 1565 6865 1585
rect 6885 1565 6900 1585
rect 6850 1535 6900 1565
rect 6850 1515 6865 1535
rect 6885 1515 6900 1535
rect 6850 1485 6900 1515
rect 6850 1465 6865 1485
rect 6885 1465 6900 1485
rect 6850 1435 6900 1465
rect 6850 1415 6865 1435
rect 6885 1415 6900 1435
rect 6850 1385 6900 1415
rect 6850 1365 6865 1385
rect 6885 1365 6900 1385
rect 6850 1335 6900 1365
rect 6850 1315 6865 1335
rect 6885 1315 6900 1335
rect 6850 1285 6900 1315
rect 6850 1265 6865 1285
rect 6885 1265 6900 1285
rect 6850 1235 6900 1265
rect 6850 1215 6865 1235
rect 6885 1215 6900 1235
rect 6850 1185 6900 1215
rect 6850 1165 6865 1185
rect 6885 1165 6900 1185
rect 6850 1135 6900 1165
rect 6850 1115 6865 1135
rect 6885 1115 6900 1135
rect 6850 1085 6900 1115
rect 6850 1065 6865 1085
rect 6885 1065 6900 1085
rect 6850 1035 6900 1065
rect 6850 1015 6865 1035
rect 6885 1015 6900 1035
rect 6850 985 6900 1015
rect 6850 965 6865 985
rect 6885 965 6900 985
rect 6850 935 6900 965
rect 6850 915 6865 935
rect 6885 915 6900 935
rect 6850 900 6900 915
rect 7000 900 7050 1600
rect 7150 1585 7200 1600
rect 7150 1565 7165 1585
rect 7185 1565 7200 1585
rect 7150 1535 7200 1565
rect 7150 1515 7165 1535
rect 7185 1515 7200 1535
rect 7150 1485 7200 1515
rect 7150 1465 7165 1485
rect 7185 1465 7200 1485
rect 7150 1435 7200 1465
rect 7150 1415 7165 1435
rect 7185 1415 7200 1435
rect 7150 1385 7200 1415
rect 7150 1365 7165 1385
rect 7185 1365 7200 1385
rect 7150 1335 7200 1365
rect 7150 1315 7165 1335
rect 7185 1315 7200 1335
rect 7150 1285 7200 1315
rect 7150 1265 7165 1285
rect 7185 1265 7200 1285
rect 7150 1235 7200 1265
rect 7150 1215 7165 1235
rect 7185 1215 7200 1235
rect 7150 1185 7200 1215
rect 7150 1165 7165 1185
rect 7185 1165 7200 1185
rect 7150 1135 7200 1165
rect 7150 1115 7165 1135
rect 7185 1115 7200 1135
rect 7150 1085 7200 1115
rect 7150 1065 7165 1085
rect 7185 1065 7200 1085
rect 7150 1035 7200 1065
rect 7150 1015 7165 1035
rect 7185 1015 7200 1035
rect 7150 985 7200 1015
rect 7150 965 7165 985
rect 7185 965 7200 985
rect 7150 935 7200 965
rect 7150 915 7165 935
rect 7185 915 7200 935
rect 7150 900 7200 915
rect 7300 900 7350 1600
rect 7450 900 7500 1600
rect 7600 900 7650 1600
rect 7750 900 7800 1600
rect 7900 900 7950 1600
rect 8050 900 8100 1600
rect 8200 900 8250 1600
rect 8350 1585 8400 1600
rect 8350 1565 8365 1585
rect 8385 1565 8400 1585
rect 8350 1535 8400 1565
rect 8350 1515 8365 1535
rect 8385 1515 8400 1535
rect 8350 1485 8400 1515
rect 8350 1465 8365 1485
rect 8385 1465 8400 1485
rect 8350 1435 8400 1465
rect 8350 1415 8365 1435
rect 8385 1415 8400 1435
rect 8350 1385 8400 1415
rect 8350 1365 8365 1385
rect 8385 1365 8400 1385
rect 8350 1335 8400 1365
rect 8350 1315 8365 1335
rect 8385 1315 8400 1335
rect 8350 1285 8400 1315
rect 8350 1265 8365 1285
rect 8385 1265 8400 1285
rect 8350 1235 8400 1265
rect 8350 1215 8365 1235
rect 8385 1215 8400 1235
rect 8350 1185 8400 1215
rect 8350 1165 8365 1185
rect 8385 1165 8400 1185
rect 8350 1135 8400 1165
rect 8350 1115 8365 1135
rect 8385 1115 8400 1135
rect 8350 1085 8400 1115
rect 8350 1065 8365 1085
rect 8385 1065 8400 1085
rect 8350 1035 8400 1065
rect 8350 1015 8365 1035
rect 8385 1015 8400 1035
rect 8350 985 8400 1015
rect 8350 965 8365 985
rect 8385 965 8400 985
rect 8350 935 8400 965
rect 8350 915 8365 935
rect 8385 915 8400 935
rect 8350 900 8400 915
rect 8500 900 8550 1600
rect 8650 900 8700 1600
rect 8800 900 8850 1600
rect 8950 900 9000 1600
rect 9100 900 9150 1600
rect 9250 900 9300 1600
rect 9400 900 9450 1600
rect 9550 1585 9600 1600
rect 9550 1565 9565 1585
rect 9585 1565 9600 1585
rect 9550 1535 9600 1565
rect 9550 1515 9565 1535
rect 9585 1515 9600 1535
rect 9550 1485 9600 1515
rect 9550 1465 9565 1485
rect 9585 1465 9600 1485
rect 9550 1435 9600 1465
rect 9550 1415 9565 1435
rect 9585 1415 9600 1435
rect 9550 1385 9600 1415
rect 9550 1365 9565 1385
rect 9585 1365 9600 1385
rect 9550 1335 9600 1365
rect 9550 1315 9565 1335
rect 9585 1315 9600 1335
rect 9550 1285 9600 1315
rect 9550 1265 9565 1285
rect 9585 1265 9600 1285
rect 9550 1235 9600 1265
rect 9550 1215 9565 1235
rect 9585 1215 9600 1235
rect 9550 1185 9600 1215
rect 9550 1165 9565 1185
rect 9585 1165 9600 1185
rect 9550 1135 9600 1165
rect 9550 1115 9565 1135
rect 9585 1115 9600 1135
rect 9550 1085 9600 1115
rect 9550 1065 9565 1085
rect 9585 1065 9600 1085
rect 9550 1035 9600 1065
rect 9550 1015 9565 1035
rect 9585 1015 9600 1035
rect 9550 985 9600 1015
rect 9550 965 9565 985
rect 9585 965 9600 985
rect 9550 935 9600 965
rect 9550 915 9565 935
rect 9585 915 9600 935
rect 9550 900 9600 915
rect 9700 900 9750 1600
rect 9850 900 9900 1600
rect 10000 900 10050 1600
rect 10150 900 10200 1600
rect 10300 900 10350 1600
rect 10450 900 10500 1600
rect 10600 900 10650 1600
rect 10750 1585 10800 1600
rect 10750 1565 10765 1585
rect 10785 1565 10800 1585
rect 10750 1535 10800 1565
rect 10750 1515 10765 1535
rect 10785 1515 10800 1535
rect 10750 1485 10800 1515
rect 10750 1465 10765 1485
rect 10785 1465 10800 1485
rect 10750 1435 10800 1465
rect 10750 1415 10765 1435
rect 10785 1415 10800 1435
rect 10750 1385 10800 1415
rect 10750 1365 10765 1385
rect 10785 1365 10800 1385
rect 10750 1335 10800 1365
rect 10750 1315 10765 1335
rect 10785 1315 10800 1335
rect 10750 1285 10800 1315
rect 10750 1265 10765 1285
rect 10785 1265 10800 1285
rect 10750 1235 10800 1265
rect 10750 1215 10765 1235
rect 10785 1215 10800 1235
rect 10750 1185 10800 1215
rect 10750 1165 10765 1185
rect 10785 1165 10800 1185
rect 10750 1135 10800 1165
rect 10750 1115 10765 1135
rect 10785 1115 10800 1135
rect 10750 1085 10800 1115
rect 10750 1065 10765 1085
rect 10785 1065 10800 1085
rect 10750 1035 10800 1065
rect 10750 1015 10765 1035
rect 10785 1015 10800 1035
rect 10750 985 10800 1015
rect 10750 965 10765 985
rect 10785 965 10800 985
rect 10750 935 10800 965
rect 10750 915 10765 935
rect 10785 915 10800 935
rect 10750 900 10800 915
rect 10900 900 10950 1600
rect 11050 900 11100 1600
rect 11200 900 11250 1600
rect 11350 900 11400 1600
rect 11500 900 11550 1600
rect 11650 900 11700 1600
rect 11800 900 11850 1600
rect 11950 1585 12000 1600
rect 11950 1565 11965 1585
rect 11985 1565 12000 1585
rect 11950 1535 12000 1565
rect 11950 1515 11965 1535
rect 11985 1515 12000 1535
rect 11950 1485 12000 1515
rect 11950 1465 11965 1485
rect 11985 1465 12000 1485
rect 11950 1435 12000 1465
rect 11950 1415 11965 1435
rect 11985 1415 12000 1435
rect 11950 1385 12000 1415
rect 11950 1365 11965 1385
rect 11985 1365 12000 1385
rect 11950 1335 12000 1365
rect 11950 1315 11965 1335
rect 11985 1315 12000 1335
rect 11950 1285 12000 1315
rect 11950 1265 11965 1285
rect 11985 1265 12000 1285
rect 11950 1235 12000 1265
rect 11950 1215 11965 1235
rect 11985 1215 12000 1235
rect 11950 1185 12000 1215
rect 11950 1165 11965 1185
rect 11985 1165 12000 1185
rect 11950 1135 12000 1165
rect 11950 1115 11965 1135
rect 11985 1115 12000 1135
rect 11950 1085 12000 1115
rect 11950 1065 11965 1085
rect 11985 1065 12000 1085
rect 11950 1035 12000 1065
rect 11950 1015 11965 1035
rect 11985 1015 12000 1035
rect 11950 985 12000 1015
rect 11950 965 11965 985
rect 11985 965 12000 985
rect 11950 935 12000 965
rect 11950 915 11965 935
rect 11985 915 12000 935
rect 11950 900 12000 915
rect 12100 900 12150 1600
rect 12250 1585 12300 1600
rect 12250 1565 12265 1585
rect 12285 1565 12300 1585
rect 12250 1535 12300 1565
rect 12250 1515 12265 1535
rect 12285 1515 12300 1535
rect 12250 1485 12300 1515
rect 12250 1465 12265 1485
rect 12285 1465 12300 1485
rect 12250 1435 12300 1465
rect 12250 1415 12265 1435
rect 12285 1415 12300 1435
rect 12250 1385 12300 1415
rect 12250 1365 12265 1385
rect 12285 1365 12300 1385
rect 12250 1335 12300 1365
rect 12250 1315 12265 1335
rect 12285 1315 12300 1335
rect 12250 1285 12300 1315
rect 12250 1265 12265 1285
rect 12285 1265 12300 1285
rect 12250 1235 12300 1265
rect 12250 1215 12265 1235
rect 12285 1215 12300 1235
rect 12250 1185 12300 1215
rect 12250 1165 12265 1185
rect 12285 1165 12300 1185
rect 12250 1135 12300 1165
rect 12250 1115 12265 1135
rect 12285 1115 12300 1135
rect 12250 1085 12300 1115
rect 12250 1065 12265 1085
rect 12285 1065 12300 1085
rect 12250 1035 12300 1065
rect 12250 1015 12265 1035
rect 12285 1015 12300 1035
rect 12250 985 12300 1015
rect 12250 965 12265 985
rect 12285 965 12300 985
rect 12250 935 12300 965
rect 12250 915 12265 935
rect 12285 915 12300 935
rect 12250 900 12300 915
rect 12400 900 12450 1600
rect 12550 1585 12600 1600
rect 12550 1565 12565 1585
rect 12585 1565 12600 1585
rect 12550 1535 12600 1565
rect 12550 1515 12565 1535
rect 12585 1515 12600 1535
rect 12550 1485 12600 1515
rect 12550 1465 12565 1485
rect 12585 1465 12600 1485
rect 12550 1435 12600 1465
rect 12550 1415 12565 1435
rect 12585 1415 12600 1435
rect 12550 1385 12600 1415
rect 12550 1365 12565 1385
rect 12585 1365 12600 1385
rect 12550 1335 12600 1365
rect 12550 1315 12565 1335
rect 12585 1315 12600 1335
rect 12550 1285 12600 1315
rect 12550 1265 12565 1285
rect 12585 1265 12600 1285
rect 12550 1235 12600 1265
rect 12550 1215 12565 1235
rect 12585 1215 12600 1235
rect 12550 1185 12600 1215
rect 12550 1165 12565 1185
rect 12585 1165 12600 1185
rect 12550 1135 12600 1165
rect 12550 1115 12565 1135
rect 12585 1115 12600 1135
rect 12550 1085 12600 1115
rect 12550 1065 12565 1085
rect 12585 1065 12600 1085
rect 12550 1035 12600 1065
rect 12550 1015 12565 1035
rect 12585 1015 12600 1035
rect 12550 985 12600 1015
rect 12550 965 12565 985
rect 12585 965 12600 985
rect 12550 935 12600 965
rect 12550 915 12565 935
rect 12585 915 12600 935
rect 12550 900 12600 915
rect 12700 900 12750 1600
rect 12850 1585 12900 1600
rect 12850 1565 12865 1585
rect 12885 1565 12900 1585
rect 12850 1535 12900 1565
rect 12850 1515 12865 1535
rect 12885 1515 12900 1535
rect 12850 1485 12900 1515
rect 12850 1465 12865 1485
rect 12885 1465 12900 1485
rect 12850 1435 12900 1465
rect 12850 1415 12865 1435
rect 12885 1415 12900 1435
rect 12850 1385 12900 1415
rect 12850 1365 12865 1385
rect 12885 1365 12900 1385
rect 12850 1335 12900 1365
rect 12850 1315 12865 1335
rect 12885 1315 12900 1335
rect 12850 1285 12900 1315
rect 12850 1265 12865 1285
rect 12885 1265 12900 1285
rect 12850 1235 12900 1265
rect 12850 1215 12865 1235
rect 12885 1215 12900 1235
rect 12850 1185 12900 1215
rect 12850 1165 12865 1185
rect 12885 1165 12900 1185
rect 12850 1135 12900 1165
rect 12850 1115 12865 1135
rect 12885 1115 12900 1135
rect 12850 1085 12900 1115
rect 12850 1065 12865 1085
rect 12885 1065 12900 1085
rect 12850 1035 12900 1065
rect 12850 1015 12865 1035
rect 12885 1015 12900 1035
rect 12850 985 12900 1015
rect 12850 965 12865 985
rect 12885 965 12900 985
rect 12850 935 12900 965
rect 12850 915 12865 935
rect 12885 915 12900 935
rect 12850 900 12900 915
rect 13000 900 13050 1600
rect 13150 1585 13200 1600
rect 13150 1565 13165 1585
rect 13185 1565 13200 1585
rect 13150 1535 13200 1565
rect 13150 1515 13165 1535
rect 13185 1515 13200 1535
rect 13150 1485 13200 1515
rect 13150 1465 13165 1485
rect 13185 1465 13200 1485
rect 13150 1435 13200 1465
rect 13150 1415 13165 1435
rect 13185 1415 13200 1435
rect 13150 1385 13200 1415
rect 13150 1365 13165 1385
rect 13185 1365 13200 1385
rect 13150 1335 13200 1365
rect 13150 1315 13165 1335
rect 13185 1315 13200 1335
rect 13150 1285 13200 1315
rect 13150 1265 13165 1285
rect 13185 1265 13200 1285
rect 13150 1235 13200 1265
rect 13150 1215 13165 1235
rect 13185 1215 13200 1235
rect 13150 1185 13200 1215
rect 13150 1165 13165 1185
rect 13185 1165 13200 1185
rect 13150 1135 13200 1165
rect 13150 1115 13165 1135
rect 13185 1115 13200 1135
rect 13150 1085 13200 1115
rect 13150 1065 13165 1085
rect 13185 1065 13200 1085
rect 13150 1035 13200 1065
rect 13150 1015 13165 1035
rect 13185 1015 13200 1035
rect 13150 985 13200 1015
rect 13150 965 13165 985
rect 13185 965 13200 985
rect 13150 935 13200 965
rect 13150 915 13165 935
rect 13185 915 13200 935
rect 13150 900 13200 915
rect 13300 900 13350 1600
rect 13450 1585 13500 1600
rect 13450 1565 13465 1585
rect 13485 1565 13500 1585
rect 13450 1535 13500 1565
rect 13450 1515 13465 1535
rect 13485 1515 13500 1535
rect 13450 1485 13500 1515
rect 13450 1465 13465 1485
rect 13485 1465 13500 1485
rect 13450 1435 13500 1465
rect 13450 1415 13465 1435
rect 13485 1415 13500 1435
rect 13450 1385 13500 1415
rect 13450 1365 13465 1385
rect 13485 1365 13500 1385
rect 13450 1335 13500 1365
rect 13450 1315 13465 1335
rect 13485 1315 13500 1335
rect 13450 1285 13500 1315
rect 13450 1265 13465 1285
rect 13485 1265 13500 1285
rect 13450 1235 13500 1265
rect 13450 1215 13465 1235
rect 13485 1215 13500 1235
rect 13450 1185 13500 1215
rect 13450 1165 13465 1185
rect 13485 1165 13500 1185
rect 13450 1135 13500 1165
rect 13450 1115 13465 1135
rect 13485 1115 13500 1135
rect 13450 1085 13500 1115
rect 13450 1065 13465 1085
rect 13485 1065 13500 1085
rect 13450 1035 13500 1065
rect 13450 1015 13465 1035
rect 13485 1015 13500 1035
rect 13450 985 13500 1015
rect 13450 965 13465 985
rect 13485 965 13500 985
rect 13450 935 13500 965
rect 13450 915 13465 935
rect 13485 915 13500 935
rect 13450 900 13500 915
rect 13600 900 13650 1600
rect 13750 1585 13800 1600
rect 13750 1565 13765 1585
rect 13785 1565 13800 1585
rect 13750 1535 13800 1565
rect 13750 1515 13765 1535
rect 13785 1515 13800 1535
rect 13750 1485 13800 1515
rect 13750 1465 13765 1485
rect 13785 1465 13800 1485
rect 13750 1435 13800 1465
rect 13750 1415 13765 1435
rect 13785 1415 13800 1435
rect 13750 1385 13800 1415
rect 13750 1365 13765 1385
rect 13785 1365 13800 1385
rect 13750 1335 13800 1365
rect 13750 1315 13765 1335
rect 13785 1315 13800 1335
rect 13750 1285 13800 1315
rect 13750 1265 13765 1285
rect 13785 1265 13800 1285
rect 13750 1235 13800 1265
rect 13750 1215 13765 1235
rect 13785 1215 13800 1235
rect 13750 1185 13800 1215
rect 13750 1165 13765 1185
rect 13785 1165 13800 1185
rect 13750 1135 13800 1165
rect 13750 1115 13765 1135
rect 13785 1115 13800 1135
rect 13750 1085 13800 1115
rect 13750 1065 13765 1085
rect 13785 1065 13800 1085
rect 13750 1035 13800 1065
rect 13750 1015 13765 1035
rect 13785 1015 13800 1035
rect 13750 985 13800 1015
rect 13750 965 13765 985
rect 13785 965 13800 985
rect 13750 935 13800 965
rect 13750 915 13765 935
rect 13785 915 13800 935
rect 13750 900 13800 915
rect 13900 900 13950 1600
rect 14050 1585 14100 1600
rect 14050 1565 14065 1585
rect 14085 1565 14100 1585
rect 14050 1535 14100 1565
rect 14050 1515 14065 1535
rect 14085 1515 14100 1535
rect 14050 1485 14100 1515
rect 14050 1465 14065 1485
rect 14085 1465 14100 1485
rect 14050 1435 14100 1465
rect 14050 1415 14065 1435
rect 14085 1415 14100 1435
rect 14050 1385 14100 1415
rect 14050 1365 14065 1385
rect 14085 1365 14100 1385
rect 14050 1335 14100 1365
rect 14050 1315 14065 1335
rect 14085 1315 14100 1335
rect 14050 1285 14100 1315
rect 14050 1265 14065 1285
rect 14085 1265 14100 1285
rect 14050 1235 14100 1265
rect 14050 1215 14065 1235
rect 14085 1215 14100 1235
rect 14050 1185 14100 1215
rect 14050 1165 14065 1185
rect 14085 1165 14100 1185
rect 14050 1135 14100 1165
rect 14050 1115 14065 1135
rect 14085 1115 14100 1135
rect 14050 1085 14100 1115
rect 14050 1065 14065 1085
rect 14085 1065 14100 1085
rect 14050 1035 14100 1065
rect 14050 1015 14065 1035
rect 14085 1015 14100 1035
rect 14050 985 14100 1015
rect 14050 965 14065 985
rect 14085 965 14100 985
rect 14050 935 14100 965
rect 14050 915 14065 935
rect 14085 915 14100 935
rect 14050 900 14100 915
rect 14200 900 14250 1600
rect 14350 1585 14400 1600
rect 14350 1565 14365 1585
rect 14385 1565 14400 1585
rect 14350 1535 14400 1565
rect 14350 1515 14365 1535
rect 14385 1515 14400 1535
rect 14350 1485 14400 1515
rect 14350 1465 14365 1485
rect 14385 1465 14400 1485
rect 14350 1435 14400 1465
rect 14350 1415 14365 1435
rect 14385 1415 14400 1435
rect 14350 1385 14400 1415
rect 14350 1365 14365 1385
rect 14385 1365 14400 1385
rect 14350 1335 14400 1365
rect 14350 1315 14365 1335
rect 14385 1315 14400 1335
rect 14350 1285 14400 1315
rect 14350 1265 14365 1285
rect 14385 1265 14400 1285
rect 14350 1235 14400 1265
rect 14350 1215 14365 1235
rect 14385 1215 14400 1235
rect 14350 1185 14400 1215
rect 14350 1165 14365 1185
rect 14385 1165 14400 1185
rect 14350 1135 14400 1165
rect 14350 1115 14365 1135
rect 14385 1115 14400 1135
rect 14350 1085 14400 1115
rect 14350 1065 14365 1085
rect 14385 1065 14400 1085
rect 14350 1035 14400 1065
rect 14350 1015 14365 1035
rect 14385 1015 14400 1035
rect 14350 985 14400 1015
rect 14350 965 14365 985
rect 14385 965 14400 985
rect 14350 935 14400 965
rect 14350 915 14365 935
rect 14385 915 14400 935
rect 14350 900 14400 915
rect 14500 900 14550 1600
rect 14650 900 14700 1600
rect 14800 900 14850 1600
rect 14950 900 15000 1600
rect 15100 900 15150 1600
rect 15250 900 15300 1600
rect 15400 900 15450 1600
rect 15550 1585 15600 1600
rect 15550 1565 15565 1585
rect 15585 1565 15600 1585
rect 15550 1535 15600 1565
rect 15550 1515 15565 1535
rect 15585 1515 15600 1535
rect 15550 1485 15600 1515
rect 15550 1465 15565 1485
rect 15585 1465 15600 1485
rect 15550 1435 15600 1465
rect 15550 1415 15565 1435
rect 15585 1415 15600 1435
rect 15550 1385 15600 1415
rect 15550 1365 15565 1385
rect 15585 1365 15600 1385
rect 15550 1335 15600 1365
rect 15550 1315 15565 1335
rect 15585 1315 15600 1335
rect 15550 1285 15600 1315
rect 15550 1265 15565 1285
rect 15585 1265 15600 1285
rect 15550 1235 15600 1265
rect 15550 1215 15565 1235
rect 15585 1215 15600 1235
rect 15550 1185 15600 1215
rect 15550 1165 15565 1185
rect 15585 1165 15600 1185
rect 15550 1135 15600 1165
rect 15550 1115 15565 1135
rect 15585 1115 15600 1135
rect 15550 1085 15600 1115
rect 15550 1065 15565 1085
rect 15585 1065 15600 1085
rect 15550 1035 15600 1065
rect 15550 1015 15565 1035
rect 15585 1015 15600 1035
rect 15550 985 15600 1015
rect 15550 965 15565 985
rect 15585 965 15600 985
rect 15550 935 15600 965
rect 15550 915 15565 935
rect 15585 915 15600 935
rect 15550 900 15600 915
rect 15700 900 15750 1600
rect 15850 900 15900 1600
rect 16000 900 16050 1600
rect 16150 900 16200 1600
rect 16300 900 16350 1600
rect 16450 900 16500 1600
rect 16600 900 16650 1600
rect 16750 1585 16800 1600
rect 16750 1565 16765 1585
rect 16785 1565 16800 1585
rect 16750 1535 16800 1565
rect 16750 1515 16765 1535
rect 16785 1515 16800 1535
rect 16750 1485 16800 1515
rect 16750 1465 16765 1485
rect 16785 1465 16800 1485
rect 16750 1435 16800 1465
rect 16750 1415 16765 1435
rect 16785 1415 16800 1435
rect 16750 1385 16800 1415
rect 16750 1365 16765 1385
rect 16785 1365 16800 1385
rect 16750 1335 16800 1365
rect 16750 1315 16765 1335
rect 16785 1315 16800 1335
rect 16750 1285 16800 1315
rect 16750 1265 16765 1285
rect 16785 1265 16800 1285
rect 16750 1235 16800 1265
rect 16750 1215 16765 1235
rect 16785 1215 16800 1235
rect 16750 1185 16800 1215
rect 16750 1165 16765 1185
rect 16785 1165 16800 1185
rect 16750 1135 16800 1165
rect 16750 1115 16765 1135
rect 16785 1115 16800 1135
rect 16750 1085 16800 1115
rect 16750 1065 16765 1085
rect 16785 1065 16800 1085
rect 16750 1035 16800 1065
rect 16750 1015 16765 1035
rect 16785 1015 16800 1035
rect 16750 985 16800 1015
rect 16750 965 16765 985
rect 16785 965 16800 985
rect 16750 935 16800 965
rect 16750 915 16765 935
rect 16785 915 16800 935
rect 16750 900 16800 915
rect 16900 900 16950 1600
rect 17050 900 17100 1600
rect 17200 900 17250 1600
rect 17350 900 17400 1600
rect 17500 900 17550 1600
rect 17650 900 17700 1600
rect 17800 900 17850 1600
rect 17950 1585 18000 1600
rect 17950 1565 17965 1585
rect 17985 1565 18000 1585
rect 17950 1535 18000 1565
rect 17950 1515 17965 1535
rect 17985 1515 18000 1535
rect 17950 1485 18000 1515
rect 17950 1465 17965 1485
rect 17985 1465 18000 1485
rect 17950 1435 18000 1465
rect 17950 1415 17965 1435
rect 17985 1415 18000 1435
rect 17950 1385 18000 1415
rect 17950 1365 17965 1385
rect 17985 1365 18000 1385
rect 17950 1335 18000 1365
rect 17950 1315 17965 1335
rect 17985 1315 18000 1335
rect 17950 1285 18000 1315
rect 17950 1265 17965 1285
rect 17985 1265 18000 1285
rect 17950 1235 18000 1265
rect 17950 1215 17965 1235
rect 17985 1215 18000 1235
rect 17950 1185 18000 1215
rect 17950 1165 17965 1185
rect 17985 1165 18000 1185
rect 17950 1135 18000 1165
rect 17950 1115 17965 1135
rect 17985 1115 18000 1135
rect 17950 1085 18000 1115
rect 17950 1065 17965 1085
rect 17985 1065 18000 1085
rect 17950 1035 18000 1065
rect 17950 1015 17965 1035
rect 17985 1015 18000 1035
rect 17950 985 18000 1015
rect 17950 965 17965 985
rect 17985 965 18000 985
rect 17950 935 18000 965
rect 17950 915 17965 935
rect 17985 915 18000 935
rect 17950 900 18000 915
rect 18100 900 18150 1600
rect 18250 900 18300 1600
rect 18400 900 18450 1600
rect 18550 900 18600 1600
rect 18700 900 18750 1600
rect 18850 900 18900 1600
rect 19000 900 19050 1600
rect 19150 1585 19200 1600
rect 19150 1565 19165 1585
rect 19185 1565 19200 1585
rect 19150 1535 19200 1565
rect 19150 1515 19165 1535
rect 19185 1515 19200 1535
rect 19150 1485 19200 1515
rect 19150 1465 19165 1485
rect 19185 1465 19200 1485
rect 19150 1435 19200 1465
rect 19150 1415 19165 1435
rect 19185 1415 19200 1435
rect 19150 1385 19200 1415
rect 19150 1365 19165 1385
rect 19185 1365 19200 1385
rect 19150 1335 19200 1365
rect 19150 1315 19165 1335
rect 19185 1315 19200 1335
rect 19150 1285 19200 1315
rect 19150 1265 19165 1285
rect 19185 1265 19200 1285
rect 19150 1235 19200 1265
rect 19150 1215 19165 1235
rect 19185 1215 19200 1235
rect 19150 1185 19200 1215
rect 19150 1165 19165 1185
rect 19185 1165 19200 1185
rect 19150 1135 19200 1165
rect 19150 1115 19165 1135
rect 19185 1115 19200 1135
rect 19150 1085 19200 1115
rect 19150 1065 19165 1085
rect 19185 1065 19200 1085
rect 19150 1035 19200 1065
rect 19150 1015 19165 1035
rect 19185 1015 19200 1035
rect 19150 985 19200 1015
rect 19150 965 19165 985
rect 19185 965 19200 985
rect 19150 935 19200 965
rect 19150 915 19165 935
rect 19185 915 19200 935
rect 19150 900 19200 915
rect 19300 900 19350 1600
rect 19450 900 19500 1600
rect 19600 900 19650 1600
rect 19750 900 19800 1600
rect 19900 900 19950 1600
rect 20050 900 20100 1600
rect 20200 900 20250 1600
rect 20350 1585 20400 1600
rect 20350 1565 20365 1585
rect 20385 1565 20400 1585
rect 20350 1535 20400 1565
rect 20350 1515 20365 1535
rect 20385 1515 20400 1535
rect 20350 1485 20400 1515
rect 20350 1465 20365 1485
rect 20385 1465 20400 1485
rect 20350 1435 20400 1465
rect 20350 1415 20365 1435
rect 20385 1415 20400 1435
rect 20350 1385 20400 1415
rect 20350 1365 20365 1385
rect 20385 1365 20400 1385
rect 20350 1335 20400 1365
rect 20350 1315 20365 1335
rect 20385 1315 20400 1335
rect 20350 1285 20400 1315
rect 20350 1265 20365 1285
rect 20385 1265 20400 1285
rect 20350 1235 20400 1265
rect 20350 1215 20365 1235
rect 20385 1215 20400 1235
rect 20350 1185 20400 1215
rect 20350 1165 20365 1185
rect 20385 1165 20400 1185
rect 20350 1135 20400 1165
rect 20350 1115 20365 1135
rect 20385 1115 20400 1135
rect 20350 1085 20400 1115
rect 20350 1065 20365 1085
rect 20385 1065 20400 1085
rect 20350 1035 20400 1065
rect 20350 1015 20365 1035
rect 20385 1015 20400 1035
rect 20350 985 20400 1015
rect 20350 965 20365 985
rect 20385 965 20400 985
rect 20350 935 20400 965
rect 20350 915 20365 935
rect 20385 915 20400 935
rect 20350 900 20400 915
rect 20500 900 20550 1600
rect 20650 900 20700 1600
rect 20800 900 20850 1600
rect 20950 900 21000 1600
rect 21100 900 21150 1600
rect 21250 900 21300 1600
rect 21400 900 21450 1600
rect 21550 1585 21600 1600
rect 21550 1565 21565 1585
rect 21585 1565 21600 1585
rect 21550 1535 21600 1565
rect 21550 1515 21565 1535
rect 21585 1515 21600 1535
rect 21550 1485 21600 1515
rect 21550 1465 21565 1485
rect 21585 1465 21600 1485
rect 21550 1435 21600 1465
rect 21550 1415 21565 1435
rect 21585 1415 21600 1435
rect 21550 1385 21600 1415
rect 21550 1365 21565 1385
rect 21585 1365 21600 1385
rect 21550 1335 21600 1365
rect 21550 1315 21565 1335
rect 21585 1315 21600 1335
rect 21550 1285 21600 1315
rect 21550 1265 21565 1285
rect 21585 1265 21600 1285
rect 21550 1235 21600 1265
rect 21550 1215 21565 1235
rect 21585 1215 21600 1235
rect 21550 1185 21600 1215
rect 21550 1165 21565 1185
rect 21585 1165 21600 1185
rect 21550 1135 21600 1165
rect 21550 1115 21565 1135
rect 21585 1115 21600 1135
rect 21550 1085 21600 1115
rect 21550 1065 21565 1085
rect 21585 1065 21600 1085
rect 21550 1035 21600 1065
rect 21550 1015 21565 1035
rect 21585 1015 21600 1035
rect 21550 985 21600 1015
rect 21550 965 21565 985
rect 21585 965 21600 985
rect 21550 935 21600 965
rect 21550 915 21565 935
rect 21585 915 21600 935
rect 21550 900 21600 915
rect 21700 900 21750 1600
rect 21850 900 21900 1600
rect 22000 900 22050 1600
rect 22150 900 22200 1600
rect 22300 900 22350 1600
rect 22450 1585 22500 1600
rect 22450 1565 22465 1585
rect 22485 1565 22500 1585
rect 22450 1535 22500 1565
rect 22450 1515 22465 1535
rect 22485 1515 22500 1535
rect 22450 1485 22500 1515
rect 22450 1465 22465 1485
rect 22485 1465 22500 1485
rect 22450 1435 22500 1465
rect 22450 1415 22465 1435
rect 22485 1415 22500 1435
rect 22450 1385 22500 1415
rect 22450 1365 22465 1385
rect 22485 1365 22500 1385
rect 22450 1335 22500 1365
rect 22450 1315 22465 1335
rect 22485 1315 22500 1335
rect 22450 1285 22500 1315
rect 22450 1265 22465 1285
rect 22485 1265 22500 1285
rect 22450 1235 22500 1265
rect 22450 1215 22465 1235
rect 22485 1215 22500 1235
rect 22450 1185 22500 1215
rect 22450 1165 22465 1185
rect 22485 1165 22500 1185
rect 22450 1135 22500 1165
rect 22450 1115 22465 1135
rect 22485 1115 22500 1135
rect 22450 1085 22500 1115
rect 22450 1065 22465 1085
rect 22485 1065 22500 1085
rect 22450 1035 22500 1065
rect 22450 1015 22465 1035
rect 22485 1015 22500 1035
rect 22450 985 22500 1015
rect 22450 965 22465 985
rect 22485 965 22500 985
rect 22450 935 22500 965
rect 22450 915 22465 935
rect 22485 915 22500 935
rect 22450 900 22500 915
rect 22600 900 22650 1600
rect 22750 900 22800 1600
rect 22900 900 22950 1600
rect 23050 900 23100 1600
rect 23200 900 23250 1600
rect 23350 1585 23400 1600
rect 23350 1565 23365 1585
rect 23385 1565 23400 1585
rect 23350 1535 23400 1565
rect 23350 1515 23365 1535
rect 23385 1515 23400 1535
rect 23350 1485 23400 1515
rect 23350 1465 23365 1485
rect 23385 1465 23400 1485
rect 23350 1435 23400 1465
rect 23350 1415 23365 1435
rect 23385 1415 23400 1435
rect 23350 1385 23400 1415
rect 23350 1365 23365 1385
rect 23385 1365 23400 1385
rect 23350 1335 23400 1365
rect 23350 1315 23365 1335
rect 23385 1315 23400 1335
rect 23350 1285 23400 1315
rect 23350 1265 23365 1285
rect 23385 1265 23400 1285
rect 23350 1235 23400 1265
rect 23350 1215 23365 1235
rect 23385 1215 23400 1235
rect 23350 1185 23400 1215
rect 23350 1165 23365 1185
rect 23385 1165 23400 1185
rect 23350 1135 23400 1165
rect 23350 1115 23365 1135
rect 23385 1115 23400 1135
rect 23350 1085 23400 1115
rect 23350 1065 23365 1085
rect 23385 1065 23400 1085
rect 23350 1035 23400 1065
rect 23350 1015 23365 1035
rect 23385 1015 23400 1035
rect 23350 985 23400 1015
rect 23350 965 23365 985
rect 23385 965 23400 985
rect 23350 935 23400 965
rect 23350 915 23365 935
rect 23385 915 23400 935
rect 23350 900 23400 915
rect 23500 900 23550 1600
rect 23650 900 23700 1600
rect 23800 900 23850 1600
rect 23950 900 24000 1600
rect 24100 900 24150 1600
rect 24250 900 24300 1600
rect 24400 900 24450 1600
rect 24550 1585 24600 1600
rect 24550 1565 24565 1585
rect 24585 1565 24600 1585
rect 24550 1535 24600 1565
rect 24550 1515 24565 1535
rect 24585 1515 24600 1535
rect 24550 1485 24600 1515
rect 24550 1465 24565 1485
rect 24585 1465 24600 1485
rect 24550 1435 24600 1465
rect 24550 1415 24565 1435
rect 24585 1415 24600 1435
rect 24550 1385 24600 1415
rect 24550 1365 24565 1385
rect 24585 1365 24600 1385
rect 24550 1335 24600 1365
rect 24550 1315 24565 1335
rect 24585 1315 24600 1335
rect 24550 1285 24600 1315
rect 24550 1265 24565 1285
rect 24585 1265 24600 1285
rect 24550 1235 24600 1265
rect 24550 1215 24565 1235
rect 24585 1215 24600 1235
rect 24550 1185 24600 1215
rect 24550 1165 24565 1185
rect 24585 1165 24600 1185
rect 24550 1135 24600 1165
rect 24550 1115 24565 1135
rect 24585 1115 24600 1135
rect 24550 1085 24600 1115
rect 24550 1065 24565 1085
rect 24585 1065 24600 1085
rect 24550 1035 24600 1065
rect 24550 1015 24565 1035
rect 24585 1015 24600 1035
rect 24550 985 24600 1015
rect 24550 965 24565 985
rect 24585 965 24600 985
rect 24550 935 24600 965
rect 24550 915 24565 935
rect 24585 915 24600 935
rect 24550 900 24600 915
rect 24700 900 24750 1600
rect 24850 900 24900 1600
rect 25000 900 25050 1600
rect 25150 900 25200 1600
rect 25300 900 25350 1600
rect 25450 900 25500 1600
rect 25600 900 25650 1600
rect 25750 1585 25800 1600
rect 25750 1565 25765 1585
rect 25785 1565 25800 1585
rect 25750 1535 25800 1565
rect 25750 1515 25765 1535
rect 25785 1515 25800 1535
rect 25750 1485 25800 1515
rect 25750 1465 25765 1485
rect 25785 1465 25800 1485
rect 25750 1435 25800 1465
rect 25750 1415 25765 1435
rect 25785 1415 25800 1435
rect 25750 1385 25800 1415
rect 25750 1365 25765 1385
rect 25785 1365 25800 1385
rect 25750 1335 25800 1365
rect 25750 1315 25765 1335
rect 25785 1315 25800 1335
rect 25750 1285 25800 1315
rect 25750 1265 25765 1285
rect 25785 1265 25800 1285
rect 25750 1235 25800 1265
rect 25750 1215 25765 1235
rect 25785 1215 25800 1235
rect 25750 1185 25800 1215
rect 25750 1165 25765 1185
rect 25785 1165 25800 1185
rect 25750 1135 25800 1165
rect 25750 1115 25765 1135
rect 25785 1115 25800 1135
rect 25750 1085 25800 1115
rect 25750 1065 25765 1085
rect 25785 1065 25800 1085
rect 25750 1035 25800 1065
rect 25750 1015 25765 1035
rect 25785 1015 25800 1035
rect 25750 985 25800 1015
rect 25750 965 25765 985
rect 25785 965 25800 985
rect 25750 935 25800 965
rect 25750 915 25765 935
rect 25785 915 25800 935
rect 25750 900 25800 915
rect 25900 900 25950 1600
rect 26050 900 26100 1600
rect 26200 900 26250 1600
rect 26350 900 26400 1600
rect 26500 900 26550 1600
rect 26650 1585 26700 1600
rect 26650 1565 26665 1585
rect 26685 1565 26700 1585
rect 26650 1535 26700 1565
rect 26650 1515 26665 1535
rect 26685 1515 26700 1535
rect 26650 1485 26700 1515
rect 26650 1465 26665 1485
rect 26685 1465 26700 1485
rect 26650 1435 26700 1465
rect 26650 1415 26665 1435
rect 26685 1415 26700 1435
rect 26650 1385 26700 1415
rect 26650 1365 26665 1385
rect 26685 1365 26700 1385
rect 26650 1335 26700 1365
rect 26650 1315 26665 1335
rect 26685 1315 26700 1335
rect 26650 1285 26700 1315
rect 26650 1265 26665 1285
rect 26685 1265 26700 1285
rect 26650 1235 26700 1265
rect 26650 1215 26665 1235
rect 26685 1215 26700 1235
rect 26650 1185 26700 1215
rect 26650 1165 26665 1185
rect 26685 1165 26700 1185
rect 26650 1135 26700 1165
rect 26650 1115 26665 1135
rect 26685 1115 26700 1135
rect 26650 1085 26700 1115
rect 26650 1065 26665 1085
rect 26685 1065 26700 1085
rect 26650 1035 26700 1065
rect 26650 1015 26665 1035
rect 26685 1015 26700 1035
rect 26650 985 26700 1015
rect 26650 965 26665 985
rect 26685 965 26700 985
rect 26650 935 26700 965
rect 26650 915 26665 935
rect 26685 915 26700 935
rect 26650 900 26700 915
rect 26800 900 26850 1600
rect 26950 900 27000 1600
rect 27100 900 27150 1600
rect 27250 900 27300 1600
rect 27400 900 27450 1600
rect 27550 1585 27600 1600
rect 27550 1565 27565 1585
rect 27585 1565 27600 1585
rect 27550 1535 27600 1565
rect 27550 1515 27565 1535
rect 27585 1515 27600 1535
rect 27550 1485 27600 1515
rect 27550 1465 27565 1485
rect 27585 1465 27600 1485
rect 27550 1435 27600 1465
rect 27550 1415 27565 1435
rect 27585 1415 27600 1435
rect 27550 1385 27600 1415
rect 27550 1365 27565 1385
rect 27585 1365 27600 1385
rect 27550 1335 27600 1365
rect 27550 1315 27565 1335
rect 27585 1315 27600 1335
rect 27550 1285 27600 1315
rect 27550 1265 27565 1285
rect 27585 1265 27600 1285
rect 27550 1235 27600 1265
rect 27550 1215 27565 1235
rect 27585 1215 27600 1235
rect 27550 1185 27600 1215
rect 27550 1165 27565 1185
rect 27585 1165 27600 1185
rect 27550 1135 27600 1165
rect 27550 1115 27565 1135
rect 27585 1115 27600 1135
rect 27550 1085 27600 1115
rect 27550 1065 27565 1085
rect 27585 1065 27600 1085
rect 27550 1035 27600 1065
rect 27550 1015 27565 1035
rect 27585 1015 27600 1035
rect 27550 985 27600 1015
rect 27550 965 27565 985
rect 27585 965 27600 985
rect 27550 935 27600 965
rect 27550 915 27565 935
rect 27585 915 27600 935
rect 27550 900 27600 915
rect 27700 900 27750 1600
rect 27850 900 27900 1600
rect 28000 900 28050 1600
rect 28150 900 28200 1600
rect 28300 900 28350 1600
rect 28450 900 28500 1600
rect 28600 900 28650 1600
rect 28750 1585 28800 1600
rect 28750 1565 28765 1585
rect 28785 1565 28800 1585
rect 28750 1535 28800 1565
rect 28750 1515 28765 1535
rect 28785 1515 28800 1535
rect 28750 1485 28800 1515
rect 28750 1465 28765 1485
rect 28785 1465 28800 1485
rect 28750 1435 28800 1465
rect 28750 1415 28765 1435
rect 28785 1415 28800 1435
rect 28750 1385 28800 1415
rect 28750 1365 28765 1385
rect 28785 1365 28800 1385
rect 28750 1335 28800 1365
rect 28750 1315 28765 1335
rect 28785 1315 28800 1335
rect 28750 1285 28800 1315
rect 28750 1265 28765 1285
rect 28785 1265 28800 1285
rect 28750 1235 28800 1265
rect 28750 1215 28765 1235
rect 28785 1215 28800 1235
rect 28750 1185 28800 1215
rect 28750 1165 28765 1185
rect 28785 1165 28800 1185
rect 28750 1135 28800 1165
rect 28750 1115 28765 1135
rect 28785 1115 28800 1135
rect 28750 1085 28800 1115
rect 28750 1065 28765 1085
rect 28785 1065 28800 1085
rect 28750 1035 28800 1065
rect 28750 1015 28765 1035
rect 28785 1015 28800 1035
rect 28750 985 28800 1015
rect 28750 965 28765 985
rect 28785 965 28800 985
rect 28750 935 28800 965
rect 28750 915 28765 935
rect 28785 915 28800 935
rect 28750 900 28800 915
rect -650 735 -600 750
rect -650 715 -635 735
rect -615 715 -600 735
rect -650 685 -600 715
rect -650 665 -635 685
rect -615 665 -600 685
rect -650 635 -600 665
rect -650 615 -635 635
rect -615 615 -600 635
rect -650 585 -600 615
rect -650 565 -635 585
rect -615 565 -600 585
rect -650 535 -600 565
rect -650 515 -635 535
rect -615 515 -600 535
rect -650 485 -600 515
rect -650 465 -635 485
rect -615 465 -600 485
rect -650 435 -600 465
rect -650 415 -635 435
rect -615 415 -600 435
rect -650 385 -600 415
rect -650 365 -635 385
rect -615 365 -600 385
rect -650 335 -600 365
rect -650 315 -635 335
rect -615 315 -600 335
rect -650 285 -600 315
rect -650 265 -635 285
rect -615 265 -600 285
rect -650 235 -600 265
rect -650 215 -635 235
rect -615 215 -600 235
rect -650 185 -600 215
rect -650 165 -635 185
rect -615 165 -600 185
rect -650 135 -600 165
rect -650 115 -635 135
rect -615 115 -600 135
rect -650 85 -600 115
rect -650 65 -635 85
rect -615 65 -600 85
rect -650 50 -600 65
rect -500 735 -450 750
rect -500 715 -485 735
rect -465 715 -450 735
rect -500 685 -450 715
rect -500 665 -485 685
rect -465 665 -450 685
rect -500 635 -450 665
rect -500 615 -485 635
rect -465 615 -450 635
rect -500 585 -450 615
rect -500 565 -485 585
rect -465 565 -450 585
rect -500 535 -450 565
rect -500 515 -485 535
rect -465 515 -450 535
rect -500 485 -450 515
rect -500 465 -485 485
rect -465 465 -450 485
rect -500 435 -450 465
rect -500 415 -485 435
rect -465 415 -450 435
rect -500 385 -450 415
rect -500 365 -485 385
rect -465 365 -450 385
rect -500 335 -450 365
rect -500 315 -485 335
rect -465 315 -450 335
rect -500 285 -450 315
rect -500 265 -485 285
rect -465 265 -450 285
rect -500 235 -450 265
rect -500 215 -485 235
rect -465 215 -450 235
rect -500 185 -450 215
rect -500 165 -485 185
rect -465 165 -450 185
rect -500 135 -450 165
rect -500 115 -485 135
rect -465 115 -450 135
rect -500 85 -450 115
rect -500 65 -485 85
rect -465 65 -450 85
rect -500 50 -450 65
rect -350 735 -300 750
rect -350 715 -335 735
rect -315 715 -300 735
rect -350 685 -300 715
rect -350 665 -335 685
rect -315 665 -300 685
rect -350 635 -300 665
rect -350 615 -335 635
rect -315 615 -300 635
rect -350 585 -300 615
rect -350 565 -335 585
rect -315 565 -300 585
rect -350 535 -300 565
rect -350 515 -335 535
rect -315 515 -300 535
rect -350 485 -300 515
rect -350 465 -335 485
rect -315 465 -300 485
rect -350 435 -300 465
rect -350 415 -335 435
rect -315 415 -300 435
rect -350 385 -300 415
rect -350 365 -335 385
rect -315 365 -300 385
rect -350 335 -300 365
rect -350 315 -335 335
rect -315 315 -300 335
rect -350 285 -300 315
rect -350 265 -335 285
rect -315 265 -300 285
rect -350 235 -300 265
rect -350 215 -335 235
rect -315 215 -300 235
rect -350 185 -300 215
rect -350 165 -335 185
rect -315 165 -300 185
rect -350 135 -300 165
rect -350 115 -335 135
rect -315 115 -300 135
rect -350 85 -300 115
rect -350 65 -335 85
rect -315 65 -300 85
rect -350 50 -300 65
rect -200 735 -150 750
rect -200 715 -185 735
rect -165 715 -150 735
rect -200 685 -150 715
rect -200 665 -185 685
rect -165 665 -150 685
rect -200 635 -150 665
rect -200 615 -185 635
rect -165 615 -150 635
rect -200 585 -150 615
rect -200 565 -185 585
rect -165 565 -150 585
rect -200 535 -150 565
rect -200 515 -185 535
rect -165 515 -150 535
rect -200 485 -150 515
rect -200 465 -185 485
rect -165 465 -150 485
rect -200 435 -150 465
rect -200 415 -185 435
rect -165 415 -150 435
rect -200 385 -150 415
rect -200 365 -185 385
rect -165 365 -150 385
rect -200 335 -150 365
rect -200 315 -185 335
rect -165 315 -150 335
rect -200 285 -150 315
rect -200 265 -185 285
rect -165 265 -150 285
rect -200 235 -150 265
rect -200 215 -185 235
rect -165 215 -150 235
rect -200 185 -150 215
rect -200 165 -185 185
rect -165 165 -150 185
rect -200 135 -150 165
rect -200 115 -185 135
rect -165 115 -150 135
rect -200 85 -150 115
rect -200 65 -185 85
rect -165 65 -150 85
rect -200 50 -150 65
rect -50 735 0 750
rect -50 715 -35 735
rect -15 715 0 735
rect -50 685 0 715
rect -50 665 -35 685
rect -15 665 0 685
rect -50 635 0 665
rect -50 615 -35 635
rect -15 615 0 635
rect -50 585 0 615
rect -50 565 -35 585
rect -15 565 0 585
rect -50 535 0 565
rect -50 515 -35 535
rect -15 515 0 535
rect -50 485 0 515
rect -50 465 -35 485
rect -15 465 0 485
rect -50 435 0 465
rect -50 415 -35 435
rect -15 415 0 435
rect -50 385 0 415
rect -50 365 -35 385
rect -15 365 0 385
rect -50 335 0 365
rect -50 315 -35 335
rect -15 315 0 335
rect -50 285 0 315
rect -50 265 -35 285
rect -15 265 0 285
rect -50 235 0 265
rect -50 215 -35 235
rect -15 215 0 235
rect -50 185 0 215
rect -50 165 -35 185
rect -15 165 0 185
rect -50 135 0 165
rect -50 115 -35 135
rect -15 115 0 135
rect -50 85 0 115
rect -50 65 -35 85
rect -15 65 0 85
rect -50 50 0 65
rect 100 50 150 750
rect 250 50 300 750
rect 400 50 450 750
rect 550 50 600 750
rect 700 50 750 750
rect 850 50 900 750
rect 1000 50 1050 750
rect 1150 735 1200 750
rect 1150 715 1165 735
rect 1185 715 1200 735
rect 1150 685 1200 715
rect 1150 665 1165 685
rect 1185 665 1200 685
rect 1150 635 1200 665
rect 1150 615 1165 635
rect 1185 615 1200 635
rect 1150 585 1200 615
rect 1150 565 1165 585
rect 1185 565 1200 585
rect 1150 535 1200 565
rect 1150 515 1165 535
rect 1185 515 1200 535
rect 1150 485 1200 515
rect 1150 465 1165 485
rect 1185 465 1200 485
rect 1150 435 1200 465
rect 1150 415 1165 435
rect 1185 415 1200 435
rect 1150 385 1200 415
rect 1150 365 1165 385
rect 1185 365 1200 385
rect 1150 335 1200 365
rect 1150 315 1165 335
rect 1185 315 1200 335
rect 1150 285 1200 315
rect 1150 265 1165 285
rect 1185 265 1200 285
rect 1150 235 1200 265
rect 1150 215 1165 235
rect 1185 215 1200 235
rect 1150 185 1200 215
rect 1150 165 1165 185
rect 1185 165 1200 185
rect 1150 135 1200 165
rect 1150 115 1165 135
rect 1185 115 1200 135
rect 1150 85 1200 115
rect 1150 65 1165 85
rect 1185 65 1200 85
rect 1150 50 1200 65
rect 1300 50 1350 750
rect 1450 735 1500 750
rect 1450 715 1465 735
rect 1485 715 1500 735
rect 1450 685 1500 715
rect 1450 665 1465 685
rect 1485 665 1500 685
rect 1450 635 1500 665
rect 1450 615 1465 635
rect 1485 615 1500 635
rect 1450 585 1500 615
rect 1450 565 1465 585
rect 1485 565 1500 585
rect 1450 535 1500 565
rect 1450 515 1465 535
rect 1485 515 1500 535
rect 1450 485 1500 515
rect 1450 465 1465 485
rect 1485 465 1500 485
rect 1450 435 1500 465
rect 1450 415 1465 435
rect 1485 415 1500 435
rect 1450 385 1500 415
rect 1450 365 1465 385
rect 1485 365 1500 385
rect 1450 335 1500 365
rect 1450 315 1465 335
rect 1485 315 1500 335
rect 1450 285 1500 315
rect 1450 265 1465 285
rect 1485 265 1500 285
rect 1450 235 1500 265
rect 1450 215 1465 235
rect 1485 215 1500 235
rect 1450 185 1500 215
rect 1450 165 1465 185
rect 1485 165 1500 185
rect 1450 135 1500 165
rect 1450 115 1465 135
rect 1485 115 1500 135
rect 1450 85 1500 115
rect 1450 65 1465 85
rect 1485 65 1500 85
rect 1450 50 1500 65
rect 1600 50 1650 750
rect 1750 735 1800 750
rect 1750 715 1765 735
rect 1785 715 1800 735
rect 1750 685 1800 715
rect 1750 665 1765 685
rect 1785 665 1800 685
rect 1750 635 1800 665
rect 1750 615 1765 635
rect 1785 615 1800 635
rect 1750 585 1800 615
rect 1750 565 1765 585
rect 1785 565 1800 585
rect 1750 535 1800 565
rect 1750 515 1765 535
rect 1785 515 1800 535
rect 1750 485 1800 515
rect 1750 465 1765 485
rect 1785 465 1800 485
rect 1750 435 1800 465
rect 1750 415 1765 435
rect 1785 415 1800 435
rect 1750 385 1800 415
rect 1750 365 1765 385
rect 1785 365 1800 385
rect 1750 335 1800 365
rect 1750 315 1765 335
rect 1785 315 1800 335
rect 1750 285 1800 315
rect 1750 265 1765 285
rect 1785 265 1800 285
rect 1750 235 1800 265
rect 1750 215 1765 235
rect 1785 215 1800 235
rect 1750 185 1800 215
rect 1750 165 1765 185
rect 1785 165 1800 185
rect 1750 135 1800 165
rect 1750 115 1765 135
rect 1785 115 1800 135
rect 1750 85 1800 115
rect 1750 65 1765 85
rect 1785 65 1800 85
rect 1750 50 1800 65
rect 1900 50 1950 750
rect 2050 735 2100 750
rect 2050 715 2065 735
rect 2085 715 2100 735
rect 2050 685 2100 715
rect 2050 665 2065 685
rect 2085 665 2100 685
rect 2050 635 2100 665
rect 2050 615 2065 635
rect 2085 615 2100 635
rect 2050 585 2100 615
rect 2050 565 2065 585
rect 2085 565 2100 585
rect 2050 535 2100 565
rect 2050 515 2065 535
rect 2085 515 2100 535
rect 2050 485 2100 515
rect 2050 465 2065 485
rect 2085 465 2100 485
rect 2050 435 2100 465
rect 2050 415 2065 435
rect 2085 415 2100 435
rect 2050 385 2100 415
rect 2050 365 2065 385
rect 2085 365 2100 385
rect 2050 335 2100 365
rect 2050 315 2065 335
rect 2085 315 2100 335
rect 2050 285 2100 315
rect 2050 265 2065 285
rect 2085 265 2100 285
rect 2050 235 2100 265
rect 2050 215 2065 235
rect 2085 215 2100 235
rect 2050 185 2100 215
rect 2050 165 2065 185
rect 2085 165 2100 185
rect 2050 135 2100 165
rect 2050 115 2065 135
rect 2085 115 2100 135
rect 2050 85 2100 115
rect 2050 65 2065 85
rect 2085 65 2100 85
rect 2050 50 2100 65
rect 2200 50 2250 750
rect 2350 735 2400 750
rect 2350 715 2365 735
rect 2385 715 2400 735
rect 2350 685 2400 715
rect 2350 665 2365 685
rect 2385 665 2400 685
rect 2350 635 2400 665
rect 2350 615 2365 635
rect 2385 615 2400 635
rect 2350 585 2400 615
rect 2350 565 2365 585
rect 2385 565 2400 585
rect 2350 535 2400 565
rect 2350 515 2365 535
rect 2385 515 2400 535
rect 2350 485 2400 515
rect 2350 465 2365 485
rect 2385 465 2400 485
rect 2350 435 2400 465
rect 2350 415 2365 435
rect 2385 415 2400 435
rect 2350 385 2400 415
rect 2350 365 2365 385
rect 2385 365 2400 385
rect 2350 335 2400 365
rect 2350 315 2365 335
rect 2385 315 2400 335
rect 2350 285 2400 315
rect 2350 265 2365 285
rect 2385 265 2400 285
rect 2350 235 2400 265
rect 2350 215 2365 235
rect 2385 215 2400 235
rect 2350 185 2400 215
rect 2350 165 2365 185
rect 2385 165 2400 185
rect 2350 135 2400 165
rect 2350 115 2365 135
rect 2385 115 2400 135
rect 2350 85 2400 115
rect 2350 65 2365 85
rect 2385 65 2400 85
rect 2350 50 2400 65
rect 2500 50 2550 750
rect 2650 735 2700 750
rect 2650 715 2665 735
rect 2685 715 2700 735
rect 2650 685 2700 715
rect 2650 665 2665 685
rect 2685 665 2700 685
rect 2650 635 2700 665
rect 2650 615 2665 635
rect 2685 615 2700 635
rect 2650 585 2700 615
rect 2650 565 2665 585
rect 2685 565 2700 585
rect 2650 535 2700 565
rect 2650 515 2665 535
rect 2685 515 2700 535
rect 2650 485 2700 515
rect 2650 465 2665 485
rect 2685 465 2700 485
rect 2650 435 2700 465
rect 2650 415 2665 435
rect 2685 415 2700 435
rect 2650 385 2700 415
rect 2650 365 2665 385
rect 2685 365 2700 385
rect 2650 335 2700 365
rect 2650 315 2665 335
rect 2685 315 2700 335
rect 2650 285 2700 315
rect 2650 265 2665 285
rect 2685 265 2700 285
rect 2650 235 2700 265
rect 2650 215 2665 235
rect 2685 215 2700 235
rect 2650 185 2700 215
rect 2650 165 2665 185
rect 2685 165 2700 185
rect 2650 135 2700 165
rect 2650 115 2665 135
rect 2685 115 2700 135
rect 2650 85 2700 115
rect 2650 65 2665 85
rect 2685 65 2700 85
rect 2650 50 2700 65
rect 2800 50 2850 750
rect 2950 735 3000 750
rect 2950 715 2965 735
rect 2985 715 3000 735
rect 2950 685 3000 715
rect 2950 665 2965 685
rect 2985 665 3000 685
rect 2950 635 3000 665
rect 2950 615 2965 635
rect 2985 615 3000 635
rect 2950 585 3000 615
rect 2950 565 2965 585
rect 2985 565 3000 585
rect 2950 535 3000 565
rect 2950 515 2965 535
rect 2985 515 3000 535
rect 2950 485 3000 515
rect 2950 465 2965 485
rect 2985 465 3000 485
rect 2950 435 3000 465
rect 2950 415 2965 435
rect 2985 415 3000 435
rect 2950 385 3000 415
rect 2950 365 2965 385
rect 2985 365 3000 385
rect 2950 335 3000 365
rect 2950 315 2965 335
rect 2985 315 3000 335
rect 2950 285 3000 315
rect 2950 265 2965 285
rect 2985 265 3000 285
rect 2950 235 3000 265
rect 2950 215 2965 235
rect 2985 215 3000 235
rect 2950 185 3000 215
rect 2950 165 2965 185
rect 2985 165 3000 185
rect 2950 135 3000 165
rect 2950 115 2965 135
rect 2985 115 3000 135
rect 2950 85 3000 115
rect 2950 65 2965 85
rect 2985 65 3000 85
rect 2950 50 3000 65
rect 3100 50 3150 750
rect 3250 735 3300 750
rect 3250 715 3265 735
rect 3285 715 3300 735
rect 3250 685 3300 715
rect 3250 665 3265 685
rect 3285 665 3300 685
rect 3250 635 3300 665
rect 3250 615 3265 635
rect 3285 615 3300 635
rect 3250 585 3300 615
rect 3250 565 3265 585
rect 3285 565 3300 585
rect 3250 535 3300 565
rect 3250 515 3265 535
rect 3285 515 3300 535
rect 3250 485 3300 515
rect 3250 465 3265 485
rect 3285 465 3300 485
rect 3250 435 3300 465
rect 3250 415 3265 435
rect 3285 415 3300 435
rect 3250 385 3300 415
rect 3250 365 3265 385
rect 3285 365 3300 385
rect 3250 335 3300 365
rect 3250 315 3265 335
rect 3285 315 3300 335
rect 3250 285 3300 315
rect 3250 265 3265 285
rect 3285 265 3300 285
rect 3250 235 3300 265
rect 3250 215 3265 235
rect 3285 215 3300 235
rect 3250 185 3300 215
rect 3250 165 3265 185
rect 3285 165 3300 185
rect 3250 135 3300 165
rect 3250 115 3265 135
rect 3285 115 3300 135
rect 3250 85 3300 115
rect 3250 65 3265 85
rect 3285 65 3300 85
rect 3250 50 3300 65
rect 3400 50 3450 750
rect 3550 735 3600 750
rect 3550 715 3565 735
rect 3585 715 3600 735
rect 3550 685 3600 715
rect 3550 665 3565 685
rect 3585 665 3600 685
rect 3550 635 3600 665
rect 3550 615 3565 635
rect 3585 615 3600 635
rect 3550 585 3600 615
rect 3550 565 3565 585
rect 3585 565 3600 585
rect 3550 535 3600 565
rect 3550 515 3565 535
rect 3585 515 3600 535
rect 3550 485 3600 515
rect 3550 465 3565 485
rect 3585 465 3600 485
rect 3550 435 3600 465
rect 3550 415 3565 435
rect 3585 415 3600 435
rect 3550 385 3600 415
rect 3550 365 3565 385
rect 3585 365 3600 385
rect 3550 335 3600 365
rect 3550 315 3565 335
rect 3585 315 3600 335
rect 3550 285 3600 315
rect 3550 265 3565 285
rect 3585 265 3600 285
rect 3550 235 3600 265
rect 3550 215 3565 235
rect 3585 215 3600 235
rect 3550 185 3600 215
rect 3550 165 3565 185
rect 3585 165 3600 185
rect 3550 135 3600 165
rect 3550 115 3565 135
rect 3585 115 3600 135
rect 3550 85 3600 115
rect 3550 65 3565 85
rect 3585 65 3600 85
rect 3550 50 3600 65
rect 3700 735 3750 750
rect 3700 715 3715 735
rect 3735 715 3750 735
rect 3700 685 3750 715
rect 3700 665 3715 685
rect 3735 665 3750 685
rect 3700 635 3750 665
rect 3700 615 3715 635
rect 3735 615 3750 635
rect 3700 585 3750 615
rect 3700 565 3715 585
rect 3735 565 3750 585
rect 3700 535 3750 565
rect 3700 515 3715 535
rect 3735 515 3750 535
rect 3700 485 3750 515
rect 3700 465 3715 485
rect 3735 465 3750 485
rect 3700 435 3750 465
rect 3700 415 3715 435
rect 3735 415 3750 435
rect 3700 385 3750 415
rect 3700 365 3715 385
rect 3735 365 3750 385
rect 3700 335 3750 365
rect 3700 315 3715 335
rect 3735 315 3750 335
rect 3700 285 3750 315
rect 3700 265 3715 285
rect 3735 265 3750 285
rect 3700 235 3750 265
rect 3700 215 3715 235
rect 3735 215 3750 235
rect 3700 185 3750 215
rect 3700 165 3715 185
rect 3735 165 3750 185
rect 3700 135 3750 165
rect 3700 115 3715 135
rect 3735 115 3750 135
rect 3700 85 3750 115
rect 3700 65 3715 85
rect 3735 65 3750 85
rect 3700 50 3750 65
rect 3850 735 3900 750
rect 3850 715 3865 735
rect 3885 715 3900 735
rect 3850 685 3900 715
rect 3850 665 3865 685
rect 3885 665 3900 685
rect 3850 635 3900 665
rect 3850 615 3865 635
rect 3885 615 3900 635
rect 3850 585 3900 615
rect 3850 565 3865 585
rect 3885 565 3900 585
rect 3850 535 3900 565
rect 3850 515 3865 535
rect 3885 515 3900 535
rect 3850 485 3900 515
rect 3850 465 3865 485
rect 3885 465 3900 485
rect 3850 435 3900 465
rect 3850 415 3865 435
rect 3885 415 3900 435
rect 3850 385 3900 415
rect 3850 365 3865 385
rect 3885 365 3900 385
rect 3850 335 3900 365
rect 3850 315 3865 335
rect 3885 315 3900 335
rect 3850 285 3900 315
rect 3850 265 3865 285
rect 3885 265 3900 285
rect 3850 235 3900 265
rect 3850 215 3865 235
rect 3885 215 3900 235
rect 3850 185 3900 215
rect 3850 165 3865 185
rect 3885 165 3900 185
rect 3850 135 3900 165
rect 3850 115 3865 135
rect 3885 115 3900 135
rect 3850 85 3900 115
rect 3850 65 3865 85
rect 3885 65 3900 85
rect 3850 50 3900 65
rect 4000 735 4050 750
rect 4000 715 4015 735
rect 4035 715 4050 735
rect 4000 685 4050 715
rect 4000 665 4015 685
rect 4035 665 4050 685
rect 4000 635 4050 665
rect 4000 615 4015 635
rect 4035 615 4050 635
rect 4000 585 4050 615
rect 4000 565 4015 585
rect 4035 565 4050 585
rect 4000 535 4050 565
rect 4000 515 4015 535
rect 4035 515 4050 535
rect 4000 485 4050 515
rect 4000 465 4015 485
rect 4035 465 4050 485
rect 4000 435 4050 465
rect 4000 415 4015 435
rect 4035 415 4050 435
rect 4000 385 4050 415
rect 4000 365 4015 385
rect 4035 365 4050 385
rect 4000 335 4050 365
rect 4000 315 4015 335
rect 4035 315 4050 335
rect 4000 285 4050 315
rect 4000 265 4015 285
rect 4035 265 4050 285
rect 4000 235 4050 265
rect 4000 215 4015 235
rect 4035 215 4050 235
rect 4000 185 4050 215
rect 4000 165 4015 185
rect 4035 165 4050 185
rect 4000 135 4050 165
rect 4000 115 4015 135
rect 4035 115 4050 135
rect 4000 85 4050 115
rect 4000 65 4015 85
rect 4035 65 4050 85
rect 4000 50 4050 65
rect 4150 735 4200 750
rect 4150 715 4165 735
rect 4185 715 4200 735
rect 4150 685 4200 715
rect 4150 665 4165 685
rect 4185 665 4200 685
rect 4150 635 4200 665
rect 4150 615 4165 635
rect 4185 615 4200 635
rect 4150 585 4200 615
rect 4150 565 4165 585
rect 4185 565 4200 585
rect 4150 535 4200 565
rect 4150 515 4165 535
rect 4185 515 4200 535
rect 4150 485 4200 515
rect 4150 465 4165 485
rect 4185 465 4200 485
rect 4150 435 4200 465
rect 4150 415 4165 435
rect 4185 415 4200 435
rect 4150 385 4200 415
rect 4150 365 4165 385
rect 4185 365 4200 385
rect 4150 335 4200 365
rect 4150 315 4165 335
rect 4185 315 4200 335
rect 4150 285 4200 315
rect 4150 265 4165 285
rect 4185 265 4200 285
rect 4150 235 4200 265
rect 4150 215 4165 235
rect 4185 215 4200 235
rect 4150 185 4200 215
rect 4150 165 4165 185
rect 4185 165 4200 185
rect 4150 135 4200 165
rect 4150 115 4165 135
rect 4185 115 4200 135
rect 4150 85 4200 115
rect 4150 65 4165 85
rect 4185 65 4200 85
rect 4150 50 4200 65
rect 4300 735 4350 750
rect 4300 715 4315 735
rect 4335 715 4350 735
rect 4300 685 4350 715
rect 4300 665 4315 685
rect 4335 665 4350 685
rect 4300 635 4350 665
rect 4300 615 4315 635
rect 4335 615 4350 635
rect 4300 585 4350 615
rect 4300 565 4315 585
rect 4335 565 4350 585
rect 4300 535 4350 565
rect 4300 515 4315 535
rect 4335 515 4350 535
rect 4300 485 4350 515
rect 4300 465 4315 485
rect 4335 465 4350 485
rect 4300 435 4350 465
rect 4300 415 4315 435
rect 4335 415 4350 435
rect 4300 385 4350 415
rect 4300 365 4315 385
rect 4335 365 4350 385
rect 4300 335 4350 365
rect 4300 315 4315 335
rect 4335 315 4350 335
rect 4300 285 4350 315
rect 4300 265 4315 285
rect 4335 265 4350 285
rect 4300 235 4350 265
rect 4300 215 4315 235
rect 4335 215 4350 235
rect 4300 185 4350 215
rect 4300 165 4315 185
rect 4335 165 4350 185
rect 4300 135 4350 165
rect 4300 115 4315 135
rect 4335 115 4350 135
rect 4300 85 4350 115
rect 4300 65 4315 85
rect 4335 65 4350 85
rect 4300 50 4350 65
rect 4450 735 4500 750
rect 4450 715 4465 735
rect 4485 715 4500 735
rect 4450 685 4500 715
rect 4450 665 4465 685
rect 4485 665 4500 685
rect 4450 635 4500 665
rect 4450 615 4465 635
rect 4485 615 4500 635
rect 4450 585 4500 615
rect 4450 565 4465 585
rect 4485 565 4500 585
rect 4450 535 4500 565
rect 4450 515 4465 535
rect 4485 515 4500 535
rect 4450 485 4500 515
rect 4450 465 4465 485
rect 4485 465 4500 485
rect 4450 435 4500 465
rect 4450 415 4465 435
rect 4485 415 4500 435
rect 4450 385 4500 415
rect 4450 365 4465 385
rect 4485 365 4500 385
rect 4450 335 4500 365
rect 4450 315 4465 335
rect 4485 315 4500 335
rect 4450 285 4500 315
rect 4450 265 4465 285
rect 4485 265 4500 285
rect 4450 235 4500 265
rect 4450 215 4465 235
rect 4485 215 4500 235
rect 4450 185 4500 215
rect 4450 165 4465 185
rect 4485 165 4500 185
rect 4450 135 4500 165
rect 4450 115 4465 135
rect 4485 115 4500 135
rect 4450 85 4500 115
rect 4450 65 4465 85
rect 4485 65 4500 85
rect 4450 50 4500 65
rect 4600 735 4650 750
rect 4600 715 4615 735
rect 4635 715 4650 735
rect 4600 685 4650 715
rect 4600 665 4615 685
rect 4635 665 4650 685
rect 4600 635 4650 665
rect 4600 615 4615 635
rect 4635 615 4650 635
rect 4600 585 4650 615
rect 4600 565 4615 585
rect 4635 565 4650 585
rect 4600 535 4650 565
rect 4600 515 4615 535
rect 4635 515 4650 535
rect 4600 485 4650 515
rect 4600 465 4615 485
rect 4635 465 4650 485
rect 4600 435 4650 465
rect 4600 415 4615 435
rect 4635 415 4650 435
rect 4600 385 4650 415
rect 4600 365 4615 385
rect 4635 365 4650 385
rect 4600 335 4650 365
rect 4600 315 4615 335
rect 4635 315 4650 335
rect 4600 285 4650 315
rect 4600 265 4615 285
rect 4635 265 4650 285
rect 4600 235 4650 265
rect 4600 215 4615 235
rect 4635 215 4650 235
rect 4600 185 4650 215
rect 4600 165 4615 185
rect 4635 165 4650 185
rect 4600 135 4650 165
rect 4600 115 4615 135
rect 4635 115 4650 135
rect 4600 85 4650 115
rect 4600 65 4615 85
rect 4635 65 4650 85
rect 4600 50 4650 65
rect 4750 735 4800 750
rect 4750 715 4765 735
rect 4785 715 4800 735
rect 4750 685 4800 715
rect 4750 665 4765 685
rect 4785 665 4800 685
rect 4750 635 4800 665
rect 4750 615 4765 635
rect 4785 615 4800 635
rect 4750 585 4800 615
rect 4750 565 4765 585
rect 4785 565 4800 585
rect 4750 535 4800 565
rect 4750 515 4765 535
rect 4785 515 4800 535
rect 4750 485 4800 515
rect 4750 465 4765 485
rect 4785 465 4800 485
rect 4750 435 4800 465
rect 4750 415 4765 435
rect 4785 415 4800 435
rect 4750 385 4800 415
rect 4750 365 4765 385
rect 4785 365 4800 385
rect 4750 335 4800 365
rect 4750 315 4765 335
rect 4785 315 4800 335
rect 4750 285 4800 315
rect 4750 265 4765 285
rect 4785 265 4800 285
rect 4750 235 4800 265
rect 4750 215 4765 235
rect 4785 215 4800 235
rect 4750 185 4800 215
rect 4750 165 4765 185
rect 4785 165 4800 185
rect 4750 135 4800 165
rect 4750 115 4765 135
rect 4785 115 4800 135
rect 4750 85 4800 115
rect 4750 65 4765 85
rect 4785 65 4800 85
rect 4750 50 4800 65
rect 4900 50 4950 750
rect 5050 735 5100 750
rect 5050 715 5065 735
rect 5085 715 5100 735
rect 5050 685 5100 715
rect 5050 665 5065 685
rect 5085 665 5100 685
rect 5050 635 5100 665
rect 5050 615 5065 635
rect 5085 615 5100 635
rect 5050 585 5100 615
rect 5050 565 5065 585
rect 5085 565 5100 585
rect 5050 535 5100 565
rect 5050 515 5065 535
rect 5085 515 5100 535
rect 5050 485 5100 515
rect 5050 465 5065 485
rect 5085 465 5100 485
rect 5050 435 5100 465
rect 5050 415 5065 435
rect 5085 415 5100 435
rect 5050 385 5100 415
rect 5050 365 5065 385
rect 5085 365 5100 385
rect 5050 335 5100 365
rect 5050 315 5065 335
rect 5085 315 5100 335
rect 5050 285 5100 315
rect 5050 265 5065 285
rect 5085 265 5100 285
rect 5050 235 5100 265
rect 5050 215 5065 235
rect 5085 215 5100 235
rect 5050 185 5100 215
rect 5050 165 5065 185
rect 5085 165 5100 185
rect 5050 135 5100 165
rect 5050 115 5065 135
rect 5085 115 5100 135
rect 5050 85 5100 115
rect 5050 65 5065 85
rect 5085 65 5100 85
rect 5050 50 5100 65
rect 5200 50 5250 750
rect 5350 735 5400 750
rect 5350 715 5365 735
rect 5385 715 5400 735
rect 5350 685 5400 715
rect 5350 665 5365 685
rect 5385 665 5400 685
rect 5350 635 5400 665
rect 5350 615 5365 635
rect 5385 615 5400 635
rect 5350 585 5400 615
rect 5350 565 5365 585
rect 5385 565 5400 585
rect 5350 535 5400 565
rect 5350 515 5365 535
rect 5385 515 5400 535
rect 5350 485 5400 515
rect 5350 465 5365 485
rect 5385 465 5400 485
rect 5350 435 5400 465
rect 5350 415 5365 435
rect 5385 415 5400 435
rect 5350 385 5400 415
rect 5350 365 5365 385
rect 5385 365 5400 385
rect 5350 335 5400 365
rect 5350 315 5365 335
rect 5385 315 5400 335
rect 5350 285 5400 315
rect 5350 265 5365 285
rect 5385 265 5400 285
rect 5350 235 5400 265
rect 5350 215 5365 235
rect 5385 215 5400 235
rect 5350 185 5400 215
rect 5350 165 5365 185
rect 5385 165 5400 185
rect 5350 135 5400 165
rect 5350 115 5365 135
rect 5385 115 5400 135
rect 5350 85 5400 115
rect 5350 65 5365 85
rect 5385 65 5400 85
rect 5350 50 5400 65
rect 5500 50 5550 750
rect 5650 735 5700 750
rect 5650 715 5665 735
rect 5685 715 5700 735
rect 5650 685 5700 715
rect 5650 665 5665 685
rect 5685 665 5700 685
rect 5650 635 5700 665
rect 5650 615 5665 635
rect 5685 615 5700 635
rect 5650 585 5700 615
rect 5650 565 5665 585
rect 5685 565 5700 585
rect 5650 535 5700 565
rect 5650 515 5665 535
rect 5685 515 5700 535
rect 5650 485 5700 515
rect 5650 465 5665 485
rect 5685 465 5700 485
rect 5650 435 5700 465
rect 5650 415 5665 435
rect 5685 415 5700 435
rect 5650 385 5700 415
rect 5650 365 5665 385
rect 5685 365 5700 385
rect 5650 335 5700 365
rect 5650 315 5665 335
rect 5685 315 5700 335
rect 5650 285 5700 315
rect 5650 265 5665 285
rect 5685 265 5700 285
rect 5650 235 5700 265
rect 5650 215 5665 235
rect 5685 215 5700 235
rect 5650 185 5700 215
rect 5650 165 5665 185
rect 5685 165 5700 185
rect 5650 135 5700 165
rect 5650 115 5665 135
rect 5685 115 5700 135
rect 5650 85 5700 115
rect 5650 65 5665 85
rect 5685 65 5700 85
rect 5650 50 5700 65
rect 5800 50 5850 750
rect 5950 735 6000 750
rect 5950 715 5965 735
rect 5985 715 6000 735
rect 5950 685 6000 715
rect 5950 665 5965 685
rect 5985 665 6000 685
rect 5950 635 6000 665
rect 5950 615 5965 635
rect 5985 615 6000 635
rect 5950 585 6000 615
rect 5950 565 5965 585
rect 5985 565 6000 585
rect 5950 535 6000 565
rect 5950 515 5965 535
rect 5985 515 6000 535
rect 5950 485 6000 515
rect 5950 465 5965 485
rect 5985 465 6000 485
rect 5950 435 6000 465
rect 5950 415 5965 435
rect 5985 415 6000 435
rect 5950 385 6000 415
rect 5950 365 5965 385
rect 5985 365 6000 385
rect 5950 335 6000 365
rect 5950 315 5965 335
rect 5985 315 6000 335
rect 5950 285 6000 315
rect 5950 265 5965 285
rect 5985 265 6000 285
rect 5950 235 6000 265
rect 5950 215 5965 235
rect 5985 215 6000 235
rect 5950 185 6000 215
rect 5950 165 5965 185
rect 5985 165 6000 185
rect 5950 135 6000 165
rect 5950 115 5965 135
rect 5985 115 6000 135
rect 5950 85 6000 115
rect 5950 65 5965 85
rect 5985 65 6000 85
rect 5950 50 6000 65
rect 6100 50 6150 750
rect 6250 735 6300 750
rect 6250 715 6265 735
rect 6285 715 6300 735
rect 6250 685 6300 715
rect 6250 665 6265 685
rect 6285 665 6300 685
rect 6250 635 6300 665
rect 6250 615 6265 635
rect 6285 615 6300 635
rect 6250 585 6300 615
rect 6250 565 6265 585
rect 6285 565 6300 585
rect 6250 535 6300 565
rect 6250 515 6265 535
rect 6285 515 6300 535
rect 6250 485 6300 515
rect 6250 465 6265 485
rect 6285 465 6300 485
rect 6250 435 6300 465
rect 6250 415 6265 435
rect 6285 415 6300 435
rect 6250 385 6300 415
rect 6250 365 6265 385
rect 6285 365 6300 385
rect 6250 335 6300 365
rect 6250 315 6265 335
rect 6285 315 6300 335
rect 6250 285 6300 315
rect 6250 265 6265 285
rect 6285 265 6300 285
rect 6250 235 6300 265
rect 6250 215 6265 235
rect 6285 215 6300 235
rect 6250 185 6300 215
rect 6250 165 6265 185
rect 6285 165 6300 185
rect 6250 135 6300 165
rect 6250 115 6265 135
rect 6285 115 6300 135
rect 6250 85 6300 115
rect 6250 65 6265 85
rect 6285 65 6300 85
rect 6250 50 6300 65
rect 6400 50 6450 750
rect 6550 735 6600 750
rect 6550 715 6565 735
rect 6585 715 6600 735
rect 6550 685 6600 715
rect 6550 665 6565 685
rect 6585 665 6600 685
rect 6550 635 6600 665
rect 6550 615 6565 635
rect 6585 615 6600 635
rect 6550 585 6600 615
rect 6550 565 6565 585
rect 6585 565 6600 585
rect 6550 535 6600 565
rect 6550 515 6565 535
rect 6585 515 6600 535
rect 6550 485 6600 515
rect 6550 465 6565 485
rect 6585 465 6600 485
rect 6550 435 6600 465
rect 6550 415 6565 435
rect 6585 415 6600 435
rect 6550 385 6600 415
rect 6550 365 6565 385
rect 6585 365 6600 385
rect 6550 335 6600 365
rect 6550 315 6565 335
rect 6585 315 6600 335
rect 6550 285 6600 315
rect 6550 265 6565 285
rect 6585 265 6600 285
rect 6550 235 6600 265
rect 6550 215 6565 235
rect 6585 215 6600 235
rect 6550 185 6600 215
rect 6550 165 6565 185
rect 6585 165 6600 185
rect 6550 135 6600 165
rect 6550 115 6565 135
rect 6585 115 6600 135
rect 6550 85 6600 115
rect 6550 65 6565 85
rect 6585 65 6600 85
rect 6550 50 6600 65
rect 6700 50 6750 750
rect 6850 735 6900 750
rect 6850 715 6865 735
rect 6885 715 6900 735
rect 6850 685 6900 715
rect 6850 665 6865 685
rect 6885 665 6900 685
rect 6850 635 6900 665
rect 6850 615 6865 635
rect 6885 615 6900 635
rect 6850 585 6900 615
rect 6850 565 6865 585
rect 6885 565 6900 585
rect 6850 535 6900 565
rect 6850 515 6865 535
rect 6885 515 6900 535
rect 6850 485 6900 515
rect 6850 465 6865 485
rect 6885 465 6900 485
rect 6850 435 6900 465
rect 6850 415 6865 435
rect 6885 415 6900 435
rect 6850 385 6900 415
rect 6850 365 6865 385
rect 6885 365 6900 385
rect 6850 335 6900 365
rect 6850 315 6865 335
rect 6885 315 6900 335
rect 6850 285 6900 315
rect 6850 265 6865 285
rect 6885 265 6900 285
rect 6850 235 6900 265
rect 6850 215 6865 235
rect 6885 215 6900 235
rect 6850 185 6900 215
rect 6850 165 6865 185
rect 6885 165 6900 185
rect 6850 135 6900 165
rect 6850 115 6865 135
rect 6885 115 6900 135
rect 6850 85 6900 115
rect 6850 65 6865 85
rect 6885 65 6900 85
rect 6850 50 6900 65
rect 7000 50 7050 750
rect 7150 735 7200 750
rect 7150 715 7165 735
rect 7185 715 7200 735
rect 7150 685 7200 715
rect 7150 665 7165 685
rect 7185 665 7200 685
rect 7150 635 7200 665
rect 7150 615 7165 635
rect 7185 615 7200 635
rect 7150 585 7200 615
rect 7150 565 7165 585
rect 7185 565 7200 585
rect 7150 535 7200 565
rect 7150 515 7165 535
rect 7185 515 7200 535
rect 7150 485 7200 515
rect 7150 465 7165 485
rect 7185 465 7200 485
rect 7150 435 7200 465
rect 7150 415 7165 435
rect 7185 415 7200 435
rect 7150 385 7200 415
rect 7150 365 7165 385
rect 7185 365 7200 385
rect 7150 335 7200 365
rect 7150 315 7165 335
rect 7185 315 7200 335
rect 7150 285 7200 315
rect 7150 265 7165 285
rect 7185 265 7200 285
rect 7150 235 7200 265
rect 7150 215 7165 235
rect 7185 215 7200 235
rect 7150 185 7200 215
rect 7150 165 7165 185
rect 7185 165 7200 185
rect 7150 135 7200 165
rect 7150 115 7165 135
rect 7185 115 7200 135
rect 7150 85 7200 115
rect 7150 65 7165 85
rect 7185 65 7200 85
rect 7150 50 7200 65
rect 7300 50 7350 750
rect 7450 50 7500 750
rect 7600 50 7650 750
rect 7750 50 7800 750
rect 7900 50 7950 750
rect 8050 50 8100 750
rect 8200 50 8250 750
rect 8350 735 8400 750
rect 8350 715 8365 735
rect 8385 715 8400 735
rect 8350 685 8400 715
rect 8350 665 8365 685
rect 8385 665 8400 685
rect 8350 635 8400 665
rect 8350 615 8365 635
rect 8385 615 8400 635
rect 8350 585 8400 615
rect 8350 565 8365 585
rect 8385 565 8400 585
rect 8350 535 8400 565
rect 8350 515 8365 535
rect 8385 515 8400 535
rect 8350 485 8400 515
rect 8350 465 8365 485
rect 8385 465 8400 485
rect 8350 435 8400 465
rect 8350 415 8365 435
rect 8385 415 8400 435
rect 8350 385 8400 415
rect 8350 365 8365 385
rect 8385 365 8400 385
rect 8350 335 8400 365
rect 8350 315 8365 335
rect 8385 315 8400 335
rect 8350 285 8400 315
rect 8350 265 8365 285
rect 8385 265 8400 285
rect 8350 235 8400 265
rect 8350 215 8365 235
rect 8385 215 8400 235
rect 8350 185 8400 215
rect 8350 165 8365 185
rect 8385 165 8400 185
rect 8350 135 8400 165
rect 8350 115 8365 135
rect 8385 115 8400 135
rect 8350 85 8400 115
rect 8350 65 8365 85
rect 8385 65 8400 85
rect 8350 50 8400 65
rect 8500 50 8550 750
rect 8650 50 8700 750
rect 8800 50 8850 750
rect 8950 50 9000 750
rect 9100 50 9150 750
rect 9250 50 9300 750
rect 9400 50 9450 750
rect 9550 735 9600 750
rect 9550 715 9565 735
rect 9585 715 9600 735
rect 9550 685 9600 715
rect 9550 665 9565 685
rect 9585 665 9600 685
rect 9550 635 9600 665
rect 9550 615 9565 635
rect 9585 615 9600 635
rect 9550 585 9600 615
rect 9550 565 9565 585
rect 9585 565 9600 585
rect 9550 535 9600 565
rect 9550 515 9565 535
rect 9585 515 9600 535
rect 9550 485 9600 515
rect 9550 465 9565 485
rect 9585 465 9600 485
rect 9550 435 9600 465
rect 9550 415 9565 435
rect 9585 415 9600 435
rect 9550 385 9600 415
rect 9550 365 9565 385
rect 9585 365 9600 385
rect 9550 335 9600 365
rect 9550 315 9565 335
rect 9585 315 9600 335
rect 9550 285 9600 315
rect 9550 265 9565 285
rect 9585 265 9600 285
rect 9550 235 9600 265
rect 9550 215 9565 235
rect 9585 215 9600 235
rect 9550 185 9600 215
rect 9550 165 9565 185
rect 9585 165 9600 185
rect 9550 135 9600 165
rect 9550 115 9565 135
rect 9585 115 9600 135
rect 9550 85 9600 115
rect 9550 65 9565 85
rect 9585 65 9600 85
rect 9550 50 9600 65
rect 9700 50 9750 750
rect 9850 50 9900 750
rect 10000 50 10050 750
rect 10150 50 10200 750
rect 10300 50 10350 750
rect 10450 50 10500 750
rect 10600 50 10650 750
rect 10750 735 10800 750
rect 10750 715 10765 735
rect 10785 715 10800 735
rect 10750 685 10800 715
rect 10750 665 10765 685
rect 10785 665 10800 685
rect 10750 635 10800 665
rect 10750 615 10765 635
rect 10785 615 10800 635
rect 10750 585 10800 615
rect 10750 565 10765 585
rect 10785 565 10800 585
rect 10750 535 10800 565
rect 10750 515 10765 535
rect 10785 515 10800 535
rect 10750 485 10800 515
rect 10750 465 10765 485
rect 10785 465 10800 485
rect 10750 435 10800 465
rect 10750 415 10765 435
rect 10785 415 10800 435
rect 10750 385 10800 415
rect 10750 365 10765 385
rect 10785 365 10800 385
rect 10750 335 10800 365
rect 10750 315 10765 335
rect 10785 315 10800 335
rect 10750 285 10800 315
rect 10750 265 10765 285
rect 10785 265 10800 285
rect 10750 235 10800 265
rect 10750 215 10765 235
rect 10785 215 10800 235
rect 10750 185 10800 215
rect 10750 165 10765 185
rect 10785 165 10800 185
rect 10750 135 10800 165
rect 10750 115 10765 135
rect 10785 115 10800 135
rect 10750 85 10800 115
rect 10750 65 10765 85
rect 10785 65 10800 85
rect 10750 50 10800 65
rect 10900 50 10950 750
rect 11050 50 11100 750
rect 11200 50 11250 750
rect 11350 50 11400 750
rect 11500 50 11550 750
rect 11650 50 11700 750
rect 11800 50 11850 750
rect 11950 735 12000 750
rect 11950 715 11965 735
rect 11985 715 12000 735
rect 11950 685 12000 715
rect 11950 665 11965 685
rect 11985 665 12000 685
rect 11950 635 12000 665
rect 11950 615 11965 635
rect 11985 615 12000 635
rect 11950 585 12000 615
rect 11950 565 11965 585
rect 11985 565 12000 585
rect 11950 535 12000 565
rect 11950 515 11965 535
rect 11985 515 12000 535
rect 11950 485 12000 515
rect 11950 465 11965 485
rect 11985 465 12000 485
rect 11950 435 12000 465
rect 11950 415 11965 435
rect 11985 415 12000 435
rect 11950 385 12000 415
rect 11950 365 11965 385
rect 11985 365 12000 385
rect 11950 335 12000 365
rect 11950 315 11965 335
rect 11985 315 12000 335
rect 11950 285 12000 315
rect 11950 265 11965 285
rect 11985 265 12000 285
rect 11950 235 12000 265
rect 11950 215 11965 235
rect 11985 215 12000 235
rect 11950 185 12000 215
rect 11950 165 11965 185
rect 11985 165 12000 185
rect 11950 135 12000 165
rect 11950 115 11965 135
rect 11985 115 12000 135
rect 11950 85 12000 115
rect 11950 65 11965 85
rect 11985 65 12000 85
rect 11950 50 12000 65
rect 12100 50 12150 750
rect 12250 735 12300 750
rect 12250 715 12265 735
rect 12285 715 12300 735
rect 12250 685 12300 715
rect 12250 665 12265 685
rect 12285 665 12300 685
rect 12250 635 12300 665
rect 12250 615 12265 635
rect 12285 615 12300 635
rect 12250 585 12300 615
rect 12250 565 12265 585
rect 12285 565 12300 585
rect 12250 535 12300 565
rect 12250 515 12265 535
rect 12285 515 12300 535
rect 12250 485 12300 515
rect 12250 465 12265 485
rect 12285 465 12300 485
rect 12250 435 12300 465
rect 12250 415 12265 435
rect 12285 415 12300 435
rect 12250 385 12300 415
rect 12250 365 12265 385
rect 12285 365 12300 385
rect 12250 335 12300 365
rect 12250 315 12265 335
rect 12285 315 12300 335
rect 12250 285 12300 315
rect 12250 265 12265 285
rect 12285 265 12300 285
rect 12250 235 12300 265
rect 12250 215 12265 235
rect 12285 215 12300 235
rect 12250 185 12300 215
rect 12250 165 12265 185
rect 12285 165 12300 185
rect 12250 135 12300 165
rect 12250 115 12265 135
rect 12285 115 12300 135
rect 12250 85 12300 115
rect 12250 65 12265 85
rect 12285 65 12300 85
rect 12250 50 12300 65
rect 12400 50 12450 750
rect 12550 735 12600 750
rect 12550 715 12565 735
rect 12585 715 12600 735
rect 12550 685 12600 715
rect 12550 665 12565 685
rect 12585 665 12600 685
rect 12550 635 12600 665
rect 12550 615 12565 635
rect 12585 615 12600 635
rect 12550 585 12600 615
rect 12550 565 12565 585
rect 12585 565 12600 585
rect 12550 535 12600 565
rect 12550 515 12565 535
rect 12585 515 12600 535
rect 12550 485 12600 515
rect 12550 465 12565 485
rect 12585 465 12600 485
rect 12550 435 12600 465
rect 12550 415 12565 435
rect 12585 415 12600 435
rect 12550 385 12600 415
rect 12550 365 12565 385
rect 12585 365 12600 385
rect 12550 335 12600 365
rect 12550 315 12565 335
rect 12585 315 12600 335
rect 12550 285 12600 315
rect 12550 265 12565 285
rect 12585 265 12600 285
rect 12550 235 12600 265
rect 12550 215 12565 235
rect 12585 215 12600 235
rect 12550 185 12600 215
rect 12550 165 12565 185
rect 12585 165 12600 185
rect 12550 135 12600 165
rect 12550 115 12565 135
rect 12585 115 12600 135
rect 12550 85 12600 115
rect 12550 65 12565 85
rect 12585 65 12600 85
rect 12550 50 12600 65
rect 12700 50 12750 750
rect 12850 735 12900 750
rect 12850 715 12865 735
rect 12885 715 12900 735
rect 12850 685 12900 715
rect 12850 665 12865 685
rect 12885 665 12900 685
rect 12850 635 12900 665
rect 12850 615 12865 635
rect 12885 615 12900 635
rect 12850 585 12900 615
rect 12850 565 12865 585
rect 12885 565 12900 585
rect 12850 535 12900 565
rect 12850 515 12865 535
rect 12885 515 12900 535
rect 12850 485 12900 515
rect 12850 465 12865 485
rect 12885 465 12900 485
rect 12850 435 12900 465
rect 12850 415 12865 435
rect 12885 415 12900 435
rect 12850 385 12900 415
rect 12850 365 12865 385
rect 12885 365 12900 385
rect 12850 335 12900 365
rect 12850 315 12865 335
rect 12885 315 12900 335
rect 12850 285 12900 315
rect 12850 265 12865 285
rect 12885 265 12900 285
rect 12850 235 12900 265
rect 12850 215 12865 235
rect 12885 215 12900 235
rect 12850 185 12900 215
rect 12850 165 12865 185
rect 12885 165 12900 185
rect 12850 135 12900 165
rect 12850 115 12865 135
rect 12885 115 12900 135
rect 12850 85 12900 115
rect 12850 65 12865 85
rect 12885 65 12900 85
rect 12850 50 12900 65
rect 13000 50 13050 750
rect 13150 735 13200 750
rect 13150 715 13165 735
rect 13185 715 13200 735
rect 13150 685 13200 715
rect 13150 665 13165 685
rect 13185 665 13200 685
rect 13150 635 13200 665
rect 13150 615 13165 635
rect 13185 615 13200 635
rect 13150 585 13200 615
rect 13150 565 13165 585
rect 13185 565 13200 585
rect 13150 535 13200 565
rect 13150 515 13165 535
rect 13185 515 13200 535
rect 13150 485 13200 515
rect 13150 465 13165 485
rect 13185 465 13200 485
rect 13150 435 13200 465
rect 13150 415 13165 435
rect 13185 415 13200 435
rect 13150 385 13200 415
rect 13150 365 13165 385
rect 13185 365 13200 385
rect 13150 335 13200 365
rect 13150 315 13165 335
rect 13185 315 13200 335
rect 13150 285 13200 315
rect 13150 265 13165 285
rect 13185 265 13200 285
rect 13150 235 13200 265
rect 13150 215 13165 235
rect 13185 215 13200 235
rect 13150 185 13200 215
rect 13150 165 13165 185
rect 13185 165 13200 185
rect 13150 135 13200 165
rect 13150 115 13165 135
rect 13185 115 13200 135
rect 13150 85 13200 115
rect 13150 65 13165 85
rect 13185 65 13200 85
rect 13150 50 13200 65
rect 13300 50 13350 750
rect 13450 735 13500 750
rect 13450 715 13465 735
rect 13485 715 13500 735
rect 13450 685 13500 715
rect 13450 665 13465 685
rect 13485 665 13500 685
rect 13450 635 13500 665
rect 13450 615 13465 635
rect 13485 615 13500 635
rect 13450 585 13500 615
rect 13450 565 13465 585
rect 13485 565 13500 585
rect 13450 535 13500 565
rect 13450 515 13465 535
rect 13485 515 13500 535
rect 13450 485 13500 515
rect 13450 465 13465 485
rect 13485 465 13500 485
rect 13450 435 13500 465
rect 13450 415 13465 435
rect 13485 415 13500 435
rect 13450 385 13500 415
rect 13450 365 13465 385
rect 13485 365 13500 385
rect 13450 335 13500 365
rect 13450 315 13465 335
rect 13485 315 13500 335
rect 13450 285 13500 315
rect 13450 265 13465 285
rect 13485 265 13500 285
rect 13450 235 13500 265
rect 13450 215 13465 235
rect 13485 215 13500 235
rect 13450 185 13500 215
rect 13450 165 13465 185
rect 13485 165 13500 185
rect 13450 135 13500 165
rect 13450 115 13465 135
rect 13485 115 13500 135
rect 13450 85 13500 115
rect 13450 65 13465 85
rect 13485 65 13500 85
rect 13450 50 13500 65
rect 13600 50 13650 750
rect 13750 735 13800 750
rect 13750 715 13765 735
rect 13785 715 13800 735
rect 13750 685 13800 715
rect 13750 665 13765 685
rect 13785 665 13800 685
rect 13750 635 13800 665
rect 13750 615 13765 635
rect 13785 615 13800 635
rect 13750 585 13800 615
rect 13750 565 13765 585
rect 13785 565 13800 585
rect 13750 535 13800 565
rect 13750 515 13765 535
rect 13785 515 13800 535
rect 13750 485 13800 515
rect 13750 465 13765 485
rect 13785 465 13800 485
rect 13750 435 13800 465
rect 13750 415 13765 435
rect 13785 415 13800 435
rect 13750 385 13800 415
rect 13750 365 13765 385
rect 13785 365 13800 385
rect 13750 335 13800 365
rect 13750 315 13765 335
rect 13785 315 13800 335
rect 13750 285 13800 315
rect 13750 265 13765 285
rect 13785 265 13800 285
rect 13750 235 13800 265
rect 13750 215 13765 235
rect 13785 215 13800 235
rect 13750 185 13800 215
rect 13750 165 13765 185
rect 13785 165 13800 185
rect 13750 135 13800 165
rect 13750 115 13765 135
rect 13785 115 13800 135
rect 13750 85 13800 115
rect 13750 65 13765 85
rect 13785 65 13800 85
rect 13750 50 13800 65
rect 13900 50 13950 750
rect 14050 735 14100 750
rect 14050 715 14065 735
rect 14085 715 14100 735
rect 14050 685 14100 715
rect 14050 665 14065 685
rect 14085 665 14100 685
rect 14050 635 14100 665
rect 14050 615 14065 635
rect 14085 615 14100 635
rect 14050 585 14100 615
rect 14050 565 14065 585
rect 14085 565 14100 585
rect 14050 535 14100 565
rect 14050 515 14065 535
rect 14085 515 14100 535
rect 14050 485 14100 515
rect 14050 465 14065 485
rect 14085 465 14100 485
rect 14050 435 14100 465
rect 14050 415 14065 435
rect 14085 415 14100 435
rect 14050 385 14100 415
rect 14050 365 14065 385
rect 14085 365 14100 385
rect 14050 335 14100 365
rect 14050 315 14065 335
rect 14085 315 14100 335
rect 14050 285 14100 315
rect 14050 265 14065 285
rect 14085 265 14100 285
rect 14050 235 14100 265
rect 14050 215 14065 235
rect 14085 215 14100 235
rect 14050 185 14100 215
rect 14050 165 14065 185
rect 14085 165 14100 185
rect 14050 135 14100 165
rect 14050 115 14065 135
rect 14085 115 14100 135
rect 14050 85 14100 115
rect 14050 65 14065 85
rect 14085 65 14100 85
rect 14050 50 14100 65
rect 14200 50 14250 750
rect 14350 735 14400 750
rect 14350 715 14365 735
rect 14385 715 14400 735
rect 14350 685 14400 715
rect 14350 665 14365 685
rect 14385 665 14400 685
rect 14350 635 14400 665
rect 14350 615 14365 635
rect 14385 615 14400 635
rect 14350 585 14400 615
rect 14350 565 14365 585
rect 14385 565 14400 585
rect 14350 535 14400 565
rect 14350 515 14365 535
rect 14385 515 14400 535
rect 14350 485 14400 515
rect 14350 465 14365 485
rect 14385 465 14400 485
rect 14350 435 14400 465
rect 14350 415 14365 435
rect 14385 415 14400 435
rect 14350 385 14400 415
rect 14350 365 14365 385
rect 14385 365 14400 385
rect 14350 335 14400 365
rect 14350 315 14365 335
rect 14385 315 14400 335
rect 14350 285 14400 315
rect 14350 265 14365 285
rect 14385 265 14400 285
rect 14350 235 14400 265
rect 14350 215 14365 235
rect 14385 215 14400 235
rect 14350 185 14400 215
rect 14350 165 14365 185
rect 14385 165 14400 185
rect 14350 135 14400 165
rect 14350 115 14365 135
rect 14385 115 14400 135
rect 14350 85 14400 115
rect 14350 65 14365 85
rect 14385 65 14400 85
rect 14350 50 14400 65
rect 14500 50 14550 750
rect 14650 50 14700 750
rect 14800 50 14850 750
rect 14950 50 15000 750
rect 15100 50 15150 750
rect 15250 50 15300 750
rect 15400 50 15450 750
rect 15550 735 15600 750
rect 15550 715 15565 735
rect 15585 715 15600 735
rect 15550 685 15600 715
rect 15550 665 15565 685
rect 15585 665 15600 685
rect 15550 635 15600 665
rect 15550 615 15565 635
rect 15585 615 15600 635
rect 15550 585 15600 615
rect 15550 565 15565 585
rect 15585 565 15600 585
rect 15550 535 15600 565
rect 15550 515 15565 535
rect 15585 515 15600 535
rect 15550 485 15600 515
rect 15550 465 15565 485
rect 15585 465 15600 485
rect 15550 435 15600 465
rect 15550 415 15565 435
rect 15585 415 15600 435
rect 15550 385 15600 415
rect 15550 365 15565 385
rect 15585 365 15600 385
rect 15550 335 15600 365
rect 15550 315 15565 335
rect 15585 315 15600 335
rect 15550 285 15600 315
rect 15550 265 15565 285
rect 15585 265 15600 285
rect 15550 235 15600 265
rect 15550 215 15565 235
rect 15585 215 15600 235
rect 15550 185 15600 215
rect 15550 165 15565 185
rect 15585 165 15600 185
rect 15550 135 15600 165
rect 15550 115 15565 135
rect 15585 115 15600 135
rect 15550 85 15600 115
rect 15550 65 15565 85
rect 15585 65 15600 85
rect 15550 50 15600 65
rect 15700 50 15750 750
rect 15850 50 15900 750
rect 16000 50 16050 750
rect 16150 50 16200 750
rect 16300 50 16350 750
rect 16450 50 16500 750
rect 16600 50 16650 750
rect 16750 735 16800 750
rect 16750 715 16765 735
rect 16785 715 16800 735
rect 16750 685 16800 715
rect 16750 665 16765 685
rect 16785 665 16800 685
rect 16750 635 16800 665
rect 16750 615 16765 635
rect 16785 615 16800 635
rect 16750 585 16800 615
rect 16750 565 16765 585
rect 16785 565 16800 585
rect 16750 535 16800 565
rect 16750 515 16765 535
rect 16785 515 16800 535
rect 16750 485 16800 515
rect 16750 465 16765 485
rect 16785 465 16800 485
rect 16750 435 16800 465
rect 16750 415 16765 435
rect 16785 415 16800 435
rect 16750 385 16800 415
rect 16750 365 16765 385
rect 16785 365 16800 385
rect 16750 335 16800 365
rect 16750 315 16765 335
rect 16785 315 16800 335
rect 16750 285 16800 315
rect 16750 265 16765 285
rect 16785 265 16800 285
rect 16750 235 16800 265
rect 16750 215 16765 235
rect 16785 215 16800 235
rect 16750 185 16800 215
rect 16750 165 16765 185
rect 16785 165 16800 185
rect 16750 135 16800 165
rect 16750 115 16765 135
rect 16785 115 16800 135
rect 16750 85 16800 115
rect 16750 65 16765 85
rect 16785 65 16800 85
rect 16750 50 16800 65
rect 16900 50 16950 750
rect 17050 50 17100 750
rect 17200 50 17250 750
rect 17350 50 17400 750
rect 17500 50 17550 750
rect 17650 50 17700 750
rect 17800 50 17850 750
rect 17950 735 18000 750
rect 17950 715 17965 735
rect 17985 715 18000 735
rect 17950 685 18000 715
rect 17950 665 17965 685
rect 17985 665 18000 685
rect 17950 635 18000 665
rect 17950 615 17965 635
rect 17985 615 18000 635
rect 17950 585 18000 615
rect 17950 565 17965 585
rect 17985 565 18000 585
rect 17950 535 18000 565
rect 17950 515 17965 535
rect 17985 515 18000 535
rect 17950 485 18000 515
rect 17950 465 17965 485
rect 17985 465 18000 485
rect 17950 435 18000 465
rect 17950 415 17965 435
rect 17985 415 18000 435
rect 17950 385 18000 415
rect 17950 365 17965 385
rect 17985 365 18000 385
rect 17950 335 18000 365
rect 17950 315 17965 335
rect 17985 315 18000 335
rect 17950 285 18000 315
rect 17950 265 17965 285
rect 17985 265 18000 285
rect 17950 235 18000 265
rect 17950 215 17965 235
rect 17985 215 18000 235
rect 17950 185 18000 215
rect 17950 165 17965 185
rect 17985 165 18000 185
rect 17950 135 18000 165
rect 17950 115 17965 135
rect 17985 115 18000 135
rect 17950 85 18000 115
rect 17950 65 17965 85
rect 17985 65 18000 85
rect 17950 50 18000 65
rect 18100 50 18150 750
rect 18250 50 18300 750
rect 18400 50 18450 750
rect 18550 50 18600 750
rect 18700 50 18750 750
rect 18850 50 18900 750
rect 19000 50 19050 750
rect 19150 735 19200 750
rect 19150 715 19165 735
rect 19185 715 19200 735
rect 19150 685 19200 715
rect 19150 665 19165 685
rect 19185 665 19200 685
rect 19150 635 19200 665
rect 19150 615 19165 635
rect 19185 615 19200 635
rect 19150 585 19200 615
rect 19150 565 19165 585
rect 19185 565 19200 585
rect 19150 535 19200 565
rect 19150 515 19165 535
rect 19185 515 19200 535
rect 19150 485 19200 515
rect 19150 465 19165 485
rect 19185 465 19200 485
rect 19150 435 19200 465
rect 19150 415 19165 435
rect 19185 415 19200 435
rect 19150 385 19200 415
rect 19150 365 19165 385
rect 19185 365 19200 385
rect 19150 335 19200 365
rect 19150 315 19165 335
rect 19185 315 19200 335
rect 19150 285 19200 315
rect 19150 265 19165 285
rect 19185 265 19200 285
rect 19150 235 19200 265
rect 19150 215 19165 235
rect 19185 215 19200 235
rect 19150 185 19200 215
rect 19150 165 19165 185
rect 19185 165 19200 185
rect 19150 135 19200 165
rect 19150 115 19165 135
rect 19185 115 19200 135
rect 19150 85 19200 115
rect 19150 65 19165 85
rect 19185 65 19200 85
rect 19150 50 19200 65
rect 19300 50 19350 750
rect 19450 50 19500 750
rect 19600 50 19650 750
rect 19750 50 19800 750
rect 19900 50 19950 750
rect 20050 50 20100 750
rect 20200 50 20250 750
rect 20350 735 20400 750
rect 20350 715 20365 735
rect 20385 715 20400 735
rect 20350 685 20400 715
rect 20350 665 20365 685
rect 20385 665 20400 685
rect 20350 635 20400 665
rect 20350 615 20365 635
rect 20385 615 20400 635
rect 20350 585 20400 615
rect 20350 565 20365 585
rect 20385 565 20400 585
rect 20350 535 20400 565
rect 20350 515 20365 535
rect 20385 515 20400 535
rect 20350 485 20400 515
rect 20350 465 20365 485
rect 20385 465 20400 485
rect 20350 435 20400 465
rect 20350 415 20365 435
rect 20385 415 20400 435
rect 20350 385 20400 415
rect 20350 365 20365 385
rect 20385 365 20400 385
rect 20350 335 20400 365
rect 20350 315 20365 335
rect 20385 315 20400 335
rect 20350 285 20400 315
rect 20350 265 20365 285
rect 20385 265 20400 285
rect 20350 235 20400 265
rect 20350 215 20365 235
rect 20385 215 20400 235
rect 20350 185 20400 215
rect 20350 165 20365 185
rect 20385 165 20400 185
rect 20350 135 20400 165
rect 20350 115 20365 135
rect 20385 115 20400 135
rect 20350 85 20400 115
rect 20350 65 20365 85
rect 20385 65 20400 85
rect 20350 50 20400 65
rect 20500 50 20550 750
rect 20650 50 20700 750
rect 20800 50 20850 750
rect 20950 50 21000 750
rect 21100 50 21150 750
rect 21250 50 21300 750
rect 21400 50 21450 750
rect 21550 735 21600 750
rect 21550 715 21565 735
rect 21585 715 21600 735
rect 21550 685 21600 715
rect 21550 665 21565 685
rect 21585 665 21600 685
rect 21550 635 21600 665
rect 21550 615 21565 635
rect 21585 615 21600 635
rect 21550 585 21600 615
rect 21550 565 21565 585
rect 21585 565 21600 585
rect 21550 535 21600 565
rect 21550 515 21565 535
rect 21585 515 21600 535
rect 21550 485 21600 515
rect 21550 465 21565 485
rect 21585 465 21600 485
rect 21550 435 21600 465
rect 21550 415 21565 435
rect 21585 415 21600 435
rect 21550 385 21600 415
rect 21550 365 21565 385
rect 21585 365 21600 385
rect 21550 335 21600 365
rect 21550 315 21565 335
rect 21585 315 21600 335
rect 21550 285 21600 315
rect 21550 265 21565 285
rect 21585 265 21600 285
rect 21550 235 21600 265
rect 21550 215 21565 235
rect 21585 215 21600 235
rect 21550 185 21600 215
rect 21550 165 21565 185
rect 21585 165 21600 185
rect 21550 135 21600 165
rect 21550 115 21565 135
rect 21585 115 21600 135
rect 21550 85 21600 115
rect 21550 65 21565 85
rect 21585 65 21600 85
rect 21550 50 21600 65
rect 21700 50 21750 750
rect 21850 50 21900 750
rect 22000 50 22050 750
rect 22150 50 22200 750
rect 22300 50 22350 750
rect 22450 735 22500 750
rect 22450 715 22465 735
rect 22485 715 22500 735
rect 22450 685 22500 715
rect 22450 665 22465 685
rect 22485 665 22500 685
rect 22450 635 22500 665
rect 22450 615 22465 635
rect 22485 615 22500 635
rect 22450 585 22500 615
rect 22450 565 22465 585
rect 22485 565 22500 585
rect 22450 535 22500 565
rect 22450 515 22465 535
rect 22485 515 22500 535
rect 22450 485 22500 515
rect 22450 465 22465 485
rect 22485 465 22500 485
rect 22450 435 22500 465
rect 22450 415 22465 435
rect 22485 415 22500 435
rect 22450 385 22500 415
rect 22450 365 22465 385
rect 22485 365 22500 385
rect 22450 335 22500 365
rect 22450 315 22465 335
rect 22485 315 22500 335
rect 22450 285 22500 315
rect 22450 265 22465 285
rect 22485 265 22500 285
rect 22450 235 22500 265
rect 22450 215 22465 235
rect 22485 215 22500 235
rect 22450 185 22500 215
rect 22450 165 22465 185
rect 22485 165 22500 185
rect 22450 135 22500 165
rect 22450 115 22465 135
rect 22485 115 22500 135
rect 22450 85 22500 115
rect 22450 65 22465 85
rect 22485 65 22500 85
rect 22450 50 22500 65
rect 22600 50 22650 750
rect 22750 50 22800 750
rect 22900 50 22950 750
rect 23050 50 23100 750
rect 23200 50 23250 750
rect 23350 735 23400 750
rect 23350 715 23365 735
rect 23385 715 23400 735
rect 23350 685 23400 715
rect 23350 665 23365 685
rect 23385 665 23400 685
rect 23350 635 23400 665
rect 23350 615 23365 635
rect 23385 615 23400 635
rect 23350 585 23400 615
rect 23350 565 23365 585
rect 23385 565 23400 585
rect 23350 535 23400 565
rect 23350 515 23365 535
rect 23385 515 23400 535
rect 23350 485 23400 515
rect 23350 465 23365 485
rect 23385 465 23400 485
rect 23350 435 23400 465
rect 23350 415 23365 435
rect 23385 415 23400 435
rect 23350 385 23400 415
rect 23350 365 23365 385
rect 23385 365 23400 385
rect 23350 335 23400 365
rect 23350 315 23365 335
rect 23385 315 23400 335
rect 23350 285 23400 315
rect 23350 265 23365 285
rect 23385 265 23400 285
rect 23350 235 23400 265
rect 23350 215 23365 235
rect 23385 215 23400 235
rect 23350 185 23400 215
rect 23350 165 23365 185
rect 23385 165 23400 185
rect 23350 135 23400 165
rect 23350 115 23365 135
rect 23385 115 23400 135
rect 23350 85 23400 115
rect 23350 65 23365 85
rect 23385 65 23400 85
rect 23350 50 23400 65
rect 23500 50 23550 750
rect 23650 50 23700 750
rect 23800 50 23850 750
rect 23950 50 24000 750
rect 24100 50 24150 750
rect 24250 50 24300 750
rect 24400 50 24450 750
rect 24550 735 24600 750
rect 24550 715 24565 735
rect 24585 715 24600 735
rect 24550 685 24600 715
rect 24550 665 24565 685
rect 24585 665 24600 685
rect 24550 635 24600 665
rect 24550 615 24565 635
rect 24585 615 24600 635
rect 24550 585 24600 615
rect 24550 565 24565 585
rect 24585 565 24600 585
rect 24550 535 24600 565
rect 24550 515 24565 535
rect 24585 515 24600 535
rect 24550 485 24600 515
rect 24550 465 24565 485
rect 24585 465 24600 485
rect 24550 435 24600 465
rect 24550 415 24565 435
rect 24585 415 24600 435
rect 24550 385 24600 415
rect 24550 365 24565 385
rect 24585 365 24600 385
rect 24550 335 24600 365
rect 24550 315 24565 335
rect 24585 315 24600 335
rect 24550 285 24600 315
rect 24550 265 24565 285
rect 24585 265 24600 285
rect 24550 235 24600 265
rect 24550 215 24565 235
rect 24585 215 24600 235
rect 24550 185 24600 215
rect 24550 165 24565 185
rect 24585 165 24600 185
rect 24550 135 24600 165
rect 24550 115 24565 135
rect 24585 115 24600 135
rect 24550 85 24600 115
rect 24550 65 24565 85
rect 24585 65 24600 85
rect 24550 50 24600 65
rect 24700 50 24750 750
rect 24850 50 24900 750
rect 25000 50 25050 750
rect 25150 50 25200 750
rect 25300 50 25350 750
rect 25450 50 25500 750
rect 25600 50 25650 750
rect 25750 735 25800 750
rect 25750 715 25765 735
rect 25785 715 25800 735
rect 25750 685 25800 715
rect 25750 665 25765 685
rect 25785 665 25800 685
rect 25750 635 25800 665
rect 25750 615 25765 635
rect 25785 615 25800 635
rect 25750 585 25800 615
rect 25750 565 25765 585
rect 25785 565 25800 585
rect 25750 535 25800 565
rect 25750 515 25765 535
rect 25785 515 25800 535
rect 25750 485 25800 515
rect 25750 465 25765 485
rect 25785 465 25800 485
rect 25750 435 25800 465
rect 25750 415 25765 435
rect 25785 415 25800 435
rect 25750 385 25800 415
rect 25750 365 25765 385
rect 25785 365 25800 385
rect 25750 335 25800 365
rect 25750 315 25765 335
rect 25785 315 25800 335
rect 25750 285 25800 315
rect 25750 265 25765 285
rect 25785 265 25800 285
rect 25750 235 25800 265
rect 25750 215 25765 235
rect 25785 215 25800 235
rect 25750 185 25800 215
rect 25750 165 25765 185
rect 25785 165 25800 185
rect 25750 135 25800 165
rect 25750 115 25765 135
rect 25785 115 25800 135
rect 25750 85 25800 115
rect 25750 65 25765 85
rect 25785 65 25800 85
rect 25750 50 25800 65
rect 25900 50 25950 750
rect 26050 50 26100 750
rect 26200 50 26250 750
rect 26350 50 26400 750
rect 26500 50 26550 750
rect 26650 735 26700 750
rect 26650 715 26665 735
rect 26685 715 26700 735
rect 26650 685 26700 715
rect 26650 665 26665 685
rect 26685 665 26700 685
rect 26650 635 26700 665
rect 26650 615 26665 635
rect 26685 615 26700 635
rect 26650 585 26700 615
rect 26650 565 26665 585
rect 26685 565 26700 585
rect 26650 535 26700 565
rect 26650 515 26665 535
rect 26685 515 26700 535
rect 26650 485 26700 515
rect 26650 465 26665 485
rect 26685 465 26700 485
rect 26650 435 26700 465
rect 26650 415 26665 435
rect 26685 415 26700 435
rect 26650 385 26700 415
rect 26650 365 26665 385
rect 26685 365 26700 385
rect 26650 335 26700 365
rect 26650 315 26665 335
rect 26685 315 26700 335
rect 26650 285 26700 315
rect 26650 265 26665 285
rect 26685 265 26700 285
rect 26650 235 26700 265
rect 26650 215 26665 235
rect 26685 215 26700 235
rect 26650 185 26700 215
rect 26650 165 26665 185
rect 26685 165 26700 185
rect 26650 135 26700 165
rect 26650 115 26665 135
rect 26685 115 26700 135
rect 26650 85 26700 115
rect 26650 65 26665 85
rect 26685 65 26700 85
rect 26650 50 26700 65
rect 26800 50 26850 750
rect 26950 50 27000 750
rect 27100 50 27150 750
rect 27250 50 27300 750
rect 27400 50 27450 750
rect 27550 735 27600 750
rect 27550 715 27565 735
rect 27585 715 27600 735
rect 27550 685 27600 715
rect 27550 665 27565 685
rect 27585 665 27600 685
rect 27550 635 27600 665
rect 27550 615 27565 635
rect 27585 615 27600 635
rect 27550 585 27600 615
rect 27550 565 27565 585
rect 27585 565 27600 585
rect 27550 535 27600 565
rect 27550 515 27565 535
rect 27585 515 27600 535
rect 27550 485 27600 515
rect 27550 465 27565 485
rect 27585 465 27600 485
rect 27550 435 27600 465
rect 27550 415 27565 435
rect 27585 415 27600 435
rect 27550 385 27600 415
rect 27550 365 27565 385
rect 27585 365 27600 385
rect 27550 335 27600 365
rect 27550 315 27565 335
rect 27585 315 27600 335
rect 27550 285 27600 315
rect 27550 265 27565 285
rect 27585 265 27600 285
rect 27550 235 27600 265
rect 27550 215 27565 235
rect 27585 215 27600 235
rect 27550 185 27600 215
rect 27550 165 27565 185
rect 27585 165 27600 185
rect 27550 135 27600 165
rect 27550 115 27565 135
rect 27585 115 27600 135
rect 27550 85 27600 115
rect 27550 65 27565 85
rect 27585 65 27600 85
rect 27550 50 27600 65
rect 27700 50 27750 750
rect 27850 50 27900 750
rect 28000 50 28050 750
rect 28150 50 28200 750
rect 28300 50 28350 750
rect 28450 50 28500 750
rect 28600 50 28650 750
rect 28750 735 28800 750
rect 28750 715 28765 735
rect 28785 715 28800 735
rect 28750 685 28800 715
rect 28750 665 28765 685
rect 28785 665 28800 685
rect 28750 635 28800 665
rect 28750 615 28765 635
rect 28785 615 28800 635
rect 28750 585 28800 615
rect 28750 565 28765 585
rect 28785 565 28800 585
rect 28750 535 28800 565
rect 28750 515 28765 535
rect 28785 515 28800 535
rect 28750 485 28800 515
rect 28750 465 28765 485
rect 28785 465 28800 485
rect 28750 435 28800 465
rect 28750 415 28765 435
rect 28785 415 28800 435
rect 28750 385 28800 415
rect 28750 365 28765 385
rect 28785 365 28800 385
rect 28750 335 28800 365
rect 28750 315 28765 335
rect 28785 315 28800 335
rect 28750 285 28800 315
rect 28750 265 28765 285
rect 28785 265 28800 285
rect 28750 235 28800 265
rect 28750 215 28765 235
rect 28785 215 28800 235
rect 28750 185 28800 215
rect 28750 165 28765 185
rect 28785 165 28800 185
rect 28750 135 28800 165
rect 28750 115 28765 135
rect 28785 115 28800 135
rect 28750 85 28800 115
rect 28750 65 28765 85
rect 28785 65 28800 85
rect 28750 50 28800 65
rect -650 -115 -600 -100
rect -650 -135 -635 -115
rect -615 -135 -600 -115
rect -650 -165 -600 -135
rect -650 -185 -635 -165
rect -615 -185 -600 -165
rect -650 -215 -600 -185
rect -650 -235 -635 -215
rect -615 -235 -600 -215
rect -650 -265 -600 -235
rect -650 -285 -635 -265
rect -615 -285 -600 -265
rect -650 -315 -600 -285
rect -650 -335 -635 -315
rect -615 -335 -600 -315
rect -650 -365 -600 -335
rect -650 -385 -635 -365
rect -615 -385 -600 -365
rect -650 -415 -600 -385
rect -650 -435 -635 -415
rect -615 -435 -600 -415
rect -650 -465 -600 -435
rect -650 -485 -635 -465
rect -615 -485 -600 -465
rect -650 -515 -600 -485
rect -650 -535 -635 -515
rect -615 -535 -600 -515
rect -650 -565 -600 -535
rect -650 -585 -635 -565
rect -615 -585 -600 -565
rect -650 -615 -600 -585
rect -650 -635 -635 -615
rect -615 -635 -600 -615
rect -650 -665 -600 -635
rect -650 -685 -635 -665
rect -615 -685 -600 -665
rect -650 -715 -600 -685
rect -650 -735 -635 -715
rect -615 -735 -600 -715
rect -650 -765 -600 -735
rect -650 -785 -635 -765
rect -615 -785 -600 -765
rect -650 -800 -600 -785
rect -500 -115 -450 -100
rect -500 -135 -485 -115
rect -465 -135 -450 -115
rect -500 -165 -450 -135
rect -500 -185 -485 -165
rect -465 -185 -450 -165
rect -500 -215 -450 -185
rect -500 -235 -485 -215
rect -465 -235 -450 -215
rect -500 -265 -450 -235
rect -500 -285 -485 -265
rect -465 -285 -450 -265
rect -500 -315 -450 -285
rect -500 -335 -485 -315
rect -465 -335 -450 -315
rect -500 -365 -450 -335
rect -500 -385 -485 -365
rect -465 -385 -450 -365
rect -500 -415 -450 -385
rect -500 -435 -485 -415
rect -465 -435 -450 -415
rect -500 -465 -450 -435
rect -500 -485 -485 -465
rect -465 -485 -450 -465
rect -500 -515 -450 -485
rect -500 -535 -485 -515
rect -465 -535 -450 -515
rect -500 -565 -450 -535
rect -500 -585 -485 -565
rect -465 -585 -450 -565
rect -500 -615 -450 -585
rect -500 -635 -485 -615
rect -465 -635 -450 -615
rect -500 -665 -450 -635
rect -500 -685 -485 -665
rect -465 -685 -450 -665
rect -500 -715 -450 -685
rect -500 -735 -485 -715
rect -465 -735 -450 -715
rect -500 -765 -450 -735
rect -500 -785 -485 -765
rect -465 -785 -450 -765
rect -500 -800 -450 -785
rect -350 -115 -300 -100
rect -350 -135 -335 -115
rect -315 -135 -300 -115
rect -350 -165 -300 -135
rect -350 -185 -335 -165
rect -315 -185 -300 -165
rect -350 -215 -300 -185
rect -350 -235 -335 -215
rect -315 -235 -300 -215
rect -350 -265 -300 -235
rect -350 -285 -335 -265
rect -315 -285 -300 -265
rect -350 -315 -300 -285
rect -350 -335 -335 -315
rect -315 -335 -300 -315
rect -350 -365 -300 -335
rect -350 -385 -335 -365
rect -315 -385 -300 -365
rect -350 -415 -300 -385
rect -350 -435 -335 -415
rect -315 -435 -300 -415
rect -350 -465 -300 -435
rect -350 -485 -335 -465
rect -315 -485 -300 -465
rect -350 -515 -300 -485
rect -350 -535 -335 -515
rect -315 -535 -300 -515
rect -350 -565 -300 -535
rect -350 -585 -335 -565
rect -315 -585 -300 -565
rect -350 -615 -300 -585
rect -350 -635 -335 -615
rect -315 -635 -300 -615
rect -350 -665 -300 -635
rect -350 -685 -335 -665
rect -315 -685 -300 -665
rect -350 -715 -300 -685
rect -350 -735 -335 -715
rect -315 -735 -300 -715
rect -350 -765 -300 -735
rect -350 -785 -335 -765
rect -315 -785 -300 -765
rect -350 -800 -300 -785
rect -200 -115 -150 -100
rect -200 -135 -185 -115
rect -165 -135 -150 -115
rect -200 -165 -150 -135
rect -200 -185 -185 -165
rect -165 -185 -150 -165
rect -200 -215 -150 -185
rect -200 -235 -185 -215
rect -165 -235 -150 -215
rect -200 -265 -150 -235
rect -200 -285 -185 -265
rect -165 -285 -150 -265
rect -200 -315 -150 -285
rect -200 -335 -185 -315
rect -165 -335 -150 -315
rect -200 -365 -150 -335
rect -200 -385 -185 -365
rect -165 -385 -150 -365
rect -200 -415 -150 -385
rect -200 -435 -185 -415
rect -165 -435 -150 -415
rect -200 -465 -150 -435
rect -200 -485 -185 -465
rect -165 -485 -150 -465
rect -200 -515 -150 -485
rect -200 -535 -185 -515
rect -165 -535 -150 -515
rect -200 -565 -150 -535
rect -200 -585 -185 -565
rect -165 -585 -150 -565
rect -200 -615 -150 -585
rect -200 -635 -185 -615
rect -165 -635 -150 -615
rect -200 -665 -150 -635
rect -200 -685 -185 -665
rect -165 -685 -150 -665
rect -200 -715 -150 -685
rect -200 -735 -185 -715
rect -165 -735 -150 -715
rect -200 -765 -150 -735
rect -200 -785 -185 -765
rect -165 -785 -150 -765
rect -200 -800 -150 -785
rect -50 -115 0 -100
rect -50 -135 -35 -115
rect -15 -135 0 -115
rect -50 -165 0 -135
rect -50 -185 -35 -165
rect -15 -185 0 -165
rect -50 -215 0 -185
rect -50 -235 -35 -215
rect -15 -235 0 -215
rect -50 -265 0 -235
rect -50 -285 -35 -265
rect -15 -285 0 -265
rect -50 -315 0 -285
rect -50 -335 -35 -315
rect -15 -335 0 -315
rect -50 -365 0 -335
rect -50 -385 -35 -365
rect -15 -385 0 -365
rect -50 -415 0 -385
rect -50 -435 -35 -415
rect -15 -435 0 -415
rect -50 -465 0 -435
rect -50 -485 -35 -465
rect -15 -485 0 -465
rect -50 -515 0 -485
rect -50 -535 -35 -515
rect -15 -535 0 -515
rect -50 -565 0 -535
rect -50 -585 -35 -565
rect -15 -585 0 -565
rect -50 -615 0 -585
rect -50 -635 -35 -615
rect -15 -635 0 -615
rect -50 -665 0 -635
rect -50 -685 -35 -665
rect -15 -685 0 -665
rect -50 -715 0 -685
rect -50 -735 -35 -715
rect -15 -735 0 -715
rect -50 -765 0 -735
rect -50 -785 -35 -765
rect -15 -785 0 -765
rect -50 -800 0 -785
rect 100 -800 150 -100
rect 250 -800 300 -100
rect 400 -800 450 -100
rect 550 -800 600 -100
rect 700 -800 750 -100
rect 850 -800 900 -100
rect 1000 -800 1050 -100
rect 1150 -115 1200 -100
rect 1150 -135 1165 -115
rect 1185 -135 1200 -115
rect 1150 -165 1200 -135
rect 1150 -185 1165 -165
rect 1185 -185 1200 -165
rect 1150 -215 1200 -185
rect 1150 -235 1165 -215
rect 1185 -235 1200 -215
rect 1150 -265 1200 -235
rect 1150 -285 1165 -265
rect 1185 -285 1200 -265
rect 1150 -315 1200 -285
rect 1150 -335 1165 -315
rect 1185 -335 1200 -315
rect 1150 -365 1200 -335
rect 1150 -385 1165 -365
rect 1185 -385 1200 -365
rect 1150 -415 1200 -385
rect 1150 -435 1165 -415
rect 1185 -435 1200 -415
rect 1150 -465 1200 -435
rect 1150 -485 1165 -465
rect 1185 -485 1200 -465
rect 1150 -515 1200 -485
rect 1150 -535 1165 -515
rect 1185 -535 1200 -515
rect 1150 -565 1200 -535
rect 1150 -585 1165 -565
rect 1185 -585 1200 -565
rect 1150 -615 1200 -585
rect 1150 -635 1165 -615
rect 1185 -635 1200 -615
rect 1150 -665 1200 -635
rect 1150 -685 1165 -665
rect 1185 -685 1200 -665
rect 1150 -715 1200 -685
rect 1150 -735 1165 -715
rect 1185 -735 1200 -715
rect 1150 -765 1200 -735
rect 1150 -785 1165 -765
rect 1185 -785 1200 -765
rect 1150 -800 1200 -785
rect 1300 -800 1350 -100
rect 1450 -115 1500 -100
rect 1450 -135 1465 -115
rect 1485 -135 1500 -115
rect 1450 -165 1500 -135
rect 1450 -185 1465 -165
rect 1485 -185 1500 -165
rect 1450 -215 1500 -185
rect 1450 -235 1465 -215
rect 1485 -235 1500 -215
rect 1450 -265 1500 -235
rect 1450 -285 1465 -265
rect 1485 -285 1500 -265
rect 1450 -315 1500 -285
rect 1450 -335 1465 -315
rect 1485 -335 1500 -315
rect 1450 -365 1500 -335
rect 1450 -385 1465 -365
rect 1485 -385 1500 -365
rect 1450 -415 1500 -385
rect 1450 -435 1465 -415
rect 1485 -435 1500 -415
rect 1450 -465 1500 -435
rect 1450 -485 1465 -465
rect 1485 -485 1500 -465
rect 1450 -515 1500 -485
rect 1450 -535 1465 -515
rect 1485 -535 1500 -515
rect 1450 -565 1500 -535
rect 1450 -585 1465 -565
rect 1485 -585 1500 -565
rect 1450 -615 1500 -585
rect 1450 -635 1465 -615
rect 1485 -635 1500 -615
rect 1450 -665 1500 -635
rect 1450 -685 1465 -665
rect 1485 -685 1500 -665
rect 1450 -715 1500 -685
rect 1450 -735 1465 -715
rect 1485 -735 1500 -715
rect 1450 -765 1500 -735
rect 1450 -785 1465 -765
rect 1485 -785 1500 -765
rect 1450 -800 1500 -785
rect 1600 -800 1650 -100
rect 1750 -115 1800 -100
rect 1750 -135 1765 -115
rect 1785 -135 1800 -115
rect 1750 -165 1800 -135
rect 1750 -185 1765 -165
rect 1785 -185 1800 -165
rect 1750 -215 1800 -185
rect 1750 -235 1765 -215
rect 1785 -235 1800 -215
rect 1750 -265 1800 -235
rect 1750 -285 1765 -265
rect 1785 -285 1800 -265
rect 1750 -315 1800 -285
rect 1750 -335 1765 -315
rect 1785 -335 1800 -315
rect 1750 -365 1800 -335
rect 1750 -385 1765 -365
rect 1785 -385 1800 -365
rect 1750 -415 1800 -385
rect 1750 -435 1765 -415
rect 1785 -435 1800 -415
rect 1750 -465 1800 -435
rect 1750 -485 1765 -465
rect 1785 -485 1800 -465
rect 1750 -515 1800 -485
rect 1750 -535 1765 -515
rect 1785 -535 1800 -515
rect 1750 -565 1800 -535
rect 1750 -585 1765 -565
rect 1785 -585 1800 -565
rect 1750 -615 1800 -585
rect 1750 -635 1765 -615
rect 1785 -635 1800 -615
rect 1750 -665 1800 -635
rect 1750 -685 1765 -665
rect 1785 -685 1800 -665
rect 1750 -715 1800 -685
rect 1750 -735 1765 -715
rect 1785 -735 1800 -715
rect 1750 -765 1800 -735
rect 1750 -785 1765 -765
rect 1785 -785 1800 -765
rect 1750 -800 1800 -785
rect 1900 -800 1950 -100
rect 2050 -115 2100 -100
rect 2050 -135 2065 -115
rect 2085 -135 2100 -115
rect 2050 -165 2100 -135
rect 2050 -185 2065 -165
rect 2085 -185 2100 -165
rect 2050 -215 2100 -185
rect 2050 -235 2065 -215
rect 2085 -235 2100 -215
rect 2050 -265 2100 -235
rect 2050 -285 2065 -265
rect 2085 -285 2100 -265
rect 2050 -315 2100 -285
rect 2050 -335 2065 -315
rect 2085 -335 2100 -315
rect 2050 -365 2100 -335
rect 2050 -385 2065 -365
rect 2085 -385 2100 -365
rect 2050 -415 2100 -385
rect 2050 -435 2065 -415
rect 2085 -435 2100 -415
rect 2050 -465 2100 -435
rect 2050 -485 2065 -465
rect 2085 -485 2100 -465
rect 2050 -515 2100 -485
rect 2050 -535 2065 -515
rect 2085 -535 2100 -515
rect 2050 -565 2100 -535
rect 2050 -585 2065 -565
rect 2085 -585 2100 -565
rect 2050 -615 2100 -585
rect 2050 -635 2065 -615
rect 2085 -635 2100 -615
rect 2050 -665 2100 -635
rect 2050 -685 2065 -665
rect 2085 -685 2100 -665
rect 2050 -715 2100 -685
rect 2050 -735 2065 -715
rect 2085 -735 2100 -715
rect 2050 -765 2100 -735
rect 2050 -785 2065 -765
rect 2085 -785 2100 -765
rect 2050 -800 2100 -785
rect 2200 -800 2250 -100
rect 2350 -115 2400 -100
rect 2350 -135 2365 -115
rect 2385 -135 2400 -115
rect 2350 -165 2400 -135
rect 2350 -185 2365 -165
rect 2385 -185 2400 -165
rect 2350 -215 2400 -185
rect 2350 -235 2365 -215
rect 2385 -235 2400 -215
rect 2350 -265 2400 -235
rect 2350 -285 2365 -265
rect 2385 -285 2400 -265
rect 2350 -315 2400 -285
rect 2350 -335 2365 -315
rect 2385 -335 2400 -315
rect 2350 -365 2400 -335
rect 2350 -385 2365 -365
rect 2385 -385 2400 -365
rect 2350 -415 2400 -385
rect 2350 -435 2365 -415
rect 2385 -435 2400 -415
rect 2350 -465 2400 -435
rect 2350 -485 2365 -465
rect 2385 -485 2400 -465
rect 2350 -515 2400 -485
rect 2350 -535 2365 -515
rect 2385 -535 2400 -515
rect 2350 -565 2400 -535
rect 2350 -585 2365 -565
rect 2385 -585 2400 -565
rect 2350 -615 2400 -585
rect 2350 -635 2365 -615
rect 2385 -635 2400 -615
rect 2350 -665 2400 -635
rect 2350 -685 2365 -665
rect 2385 -685 2400 -665
rect 2350 -715 2400 -685
rect 2350 -735 2365 -715
rect 2385 -735 2400 -715
rect 2350 -765 2400 -735
rect 2350 -785 2365 -765
rect 2385 -785 2400 -765
rect 2350 -800 2400 -785
rect 2500 -800 2550 -100
rect 2650 -115 2700 -100
rect 2650 -135 2665 -115
rect 2685 -135 2700 -115
rect 2650 -165 2700 -135
rect 2650 -185 2665 -165
rect 2685 -185 2700 -165
rect 2650 -215 2700 -185
rect 2650 -235 2665 -215
rect 2685 -235 2700 -215
rect 2650 -265 2700 -235
rect 2650 -285 2665 -265
rect 2685 -285 2700 -265
rect 2650 -315 2700 -285
rect 2650 -335 2665 -315
rect 2685 -335 2700 -315
rect 2650 -365 2700 -335
rect 2650 -385 2665 -365
rect 2685 -385 2700 -365
rect 2650 -415 2700 -385
rect 2650 -435 2665 -415
rect 2685 -435 2700 -415
rect 2650 -465 2700 -435
rect 2650 -485 2665 -465
rect 2685 -485 2700 -465
rect 2650 -515 2700 -485
rect 2650 -535 2665 -515
rect 2685 -535 2700 -515
rect 2650 -565 2700 -535
rect 2650 -585 2665 -565
rect 2685 -585 2700 -565
rect 2650 -615 2700 -585
rect 2650 -635 2665 -615
rect 2685 -635 2700 -615
rect 2650 -665 2700 -635
rect 2650 -685 2665 -665
rect 2685 -685 2700 -665
rect 2650 -715 2700 -685
rect 2650 -735 2665 -715
rect 2685 -735 2700 -715
rect 2650 -765 2700 -735
rect 2650 -785 2665 -765
rect 2685 -785 2700 -765
rect 2650 -800 2700 -785
rect 2800 -800 2850 -100
rect 2950 -115 3000 -100
rect 2950 -135 2965 -115
rect 2985 -135 3000 -115
rect 2950 -165 3000 -135
rect 2950 -185 2965 -165
rect 2985 -185 3000 -165
rect 2950 -215 3000 -185
rect 2950 -235 2965 -215
rect 2985 -235 3000 -215
rect 2950 -265 3000 -235
rect 2950 -285 2965 -265
rect 2985 -285 3000 -265
rect 2950 -315 3000 -285
rect 2950 -335 2965 -315
rect 2985 -335 3000 -315
rect 2950 -365 3000 -335
rect 2950 -385 2965 -365
rect 2985 -385 3000 -365
rect 2950 -415 3000 -385
rect 2950 -435 2965 -415
rect 2985 -435 3000 -415
rect 2950 -465 3000 -435
rect 2950 -485 2965 -465
rect 2985 -485 3000 -465
rect 2950 -515 3000 -485
rect 2950 -535 2965 -515
rect 2985 -535 3000 -515
rect 2950 -565 3000 -535
rect 2950 -585 2965 -565
rect 2985 -585 3000 -565
rect 2950 -615 3000 -585
rect 2950 -635 2965 -615
rect 2985 -635 3000 -615
rect 2950 -665 3000 -635
rect 2950 -685 2965 -665
rect 2985 -685 3000 -665
rect 2950 -715 3000 -685
rect 2950 -735 2965 -715
rect 2985 -735 3000 -715
rect 2950 -765 3000 -735
rect 2950 -785 2965 -765
rect 2985 -785 3000 -765
rect 2950 -800 3000 -785
rect 3100 -800 3150 -100
rect 3250 -115 3300 -100
rect 3250 -135 3265 -115
rect 3285 -135 3300 -115
rect 3250 -165 3300 -135
rect 3250 -185 3265 -165
rect 3285 -185 3300 -165
rect 3250 -215 3300 -185
rect 3250 -235 3265 -215
rect 3285 -235 3300 -215
rect 3250 -265 3300 -235
rect 3250 -285 3265 -265
rect 3285 -285 3300 -265
rect 3250 -315 3300 -285
rect 3250 -335 3265 -315
rect 3285 -335 3300 -315
rect 3250 -365 3300 -335
rect 3250 -385 3265 -365
rect 3285 -385 3300 -365
rect 3250 -415 3300 -385
rect 3250 -435 3265 -415
rect 3285 -435 3300 -415
rect 3250 -465 3300 -435
rect 3250 -485 3265 -465
rect 3285 -485 3300 -465
rect 3250 -515 3300 -485
rect 3250 -535 3265 -515
rect 3285 -535 3300 -515
rect 3250 -565 3300 -535
rect 3250 -585 3265 -565
rect 3285 -585 3300 -565
rect 3250 -615 3300 -585
rect 3250 -635 3265 -615
rect 3285 -635 3300 -615
rect 3250 -665 3300 -635
rect 3250 -685 3265 -665
rect 3285 -685 3300 -665
rect 3250 -715 3300 -685
rect 3250 -735 3265 -715
rect 3285 -735 3300 -715
rect 3250 -765 3300 -735
rect 3250 -785 3265 -765
rect 3285 -785 3300 -765
rect 3250 -800 3300 -785
rect 3400 -800 3450 -100
rect 3550 -115 3600 -100
rect 3550 -135 3565 -115
rect 3585 -135 3600 -115
rect 3550 -165 3600 -135
rect 3550 -185 3565 -165
rect 3585 -185 3600 -165
rect 3550 -215 3600 -185
rect 3550 -235 3565 -215
rect 3585 -235 3600 -215
rect 3550 -265 3600 -235
rect 3550 -285 3565 -265
rect 3585 -285 3600 -265
rect 3550 -315 3600 -285
rect 3550 -335 3565 -315
rect 3585 -335 3600 -315
rect 3550 -365 3600 -335
rect 3550 -385 3565 -365
rect 3585 -385 3600 -365
rect 3550 -415 3600 -385
rect 3550 -435 3565 -415
rect 3585 -435 3600 -415
rect 3550 -465 3600 -435
rect 3550 -485 3565 -465
rect 3585 -485 3600 -465
rect 3550 -515 3600 -485
rect 3550 -535 3565 -515
rect 3585 -535 3600 -515
rect 3550 -565 3600 -535
rect 3550 -585 3565 -565
rect 3585 -585 3600 -565
rect 3550 -615 3600 -585
rect 3550 -635 3565 -615
rect 3585 -635 3600 -615
rect 3550 -665 3600 -635
rect 3550 -685 3565 -665
rect 3585 -685 3600 -665
rect 3550 -715 3600 -685
rect 3550 -735 3565 -715
rect 3585 -735 3600 -715
rect 3550 -765 3600 -735
rect 3550 -785 3565 -765
rect 3585 -785 3600 -765
rect 3550 -800 3600 -785
rect 3700 -115 3750 -100
rect 3700 -135 3715 -115
rect 3735 -135 3750 -115
rect 3700 -165 3750 -135
rect 3700 -185 3715 -165
rect 3735 -185 3750 -165
rect 3700 -215 3750 -185
rect 3700 -235 3715 -215
rect 3735 -235 3750 -215
rect 3700 -265 3750 -235
rect 3700 -285 3715 -265
rect 3735 -285 3750 -265
rect 3700 -315 3750 -285
rect 3700 -335 3715 -315
rect 3735 -335 3750 -315
rect 3700 -365 3750 -335
rect 3700 -385 3715 -365
rect 3735 -385 3750 -365
rect 3700 -415 3750 -385
rect 3700 -435 3715 -415
rect 3735 -435 3750 -415
rect 3700 -465 3750 -435
rect 3700 -485 3715 -465
rect 3735 -485 3750 -465
rect 3700 -515 3750 -485
rect 3700 -535 3715 -515
rect 3735 -535 3750 -515
rect 3700 -565 3750 -535
rect 3700 -585 3715 -565
rect 3735 -585 3750 -565
rect 3700 -615 3750 -585
rect 3700 -635 3715 -615
rect 3735 -635 3750 -615
rect 3700 -665 3750 -635
rect 3700 -685 3715 -665
rect 3735 -685 3750 -665
rect 3700 -715 3750 -685
rect 3700 -735 3715 -715
rect 3735 -735 3750 -715
rect 3700 -765 3750 -735
rect 3700 -785 3715 -765
rect 3735 -785 3750 -765
rect 3700 -800 3750 -785
rect 3850 -115 3900 -100
rect 3850 -135 3865 -115
rect 3885 -135 3900 -115
rect 3850 -165 3900 -135
rect 3850 -185 3865 -165
rect 3885 -185 3900 -165
rect 3850 -215 3900 -185
rect 3850 -235 3865 -215
rect 3885 -235 3900 -215
rect 3850 -265 3900 -235
rect 3850 -285 3865 -265
rect 3885 -285 3900 -265
rect 3850 -315 3900 -285
rect 3850 -335 3865 -315
rect 3885 -335 3900 -315
rect 3850 -365 3900 -335
rect 3850 -385 3865 -365
rect 3885 -385 3900 -365
rect 3850 -415 3900 -385
rect 3850 -435 3865 -415
rect 3885 -435 3900 -415
rect 3850 -465 3900 -435
rect 3850 -485 3865 -465
rect 3885 -485 3900 -465
rect 3850 -515 3900 -485
rect 3850 -535 3865 -515
rect 3885 -535 3900 -515
rect 3850 -565 3900 -535
rect 3850 -585 3865 -565
rect 3885 -585 3900 -565
rect 3850 -615 3900 -585
rect 3850 -635 3865 -615
rect 3885 -635 3900 -615
rect 3850 -665 3900 -635
rect 3850 -685 3865 -665
rect 3885 -685 3900 -665
rect 3850 -715 3900 -685
rect 3850 -735 3865 -715
rect 3885 -735 3900 -715
rect 3850 -765 3900 -735
rect 3850 -785 3865 -765
rect 3885 -785 3900 -765
rect 3850 -800 3900 -785
rect 4000 -115 4050 -100
rect 4000 -135 4015 -115
rect 4035 -135 4050 -115
rect 4000 -165 4050 -135
rect 4000 -185 4015 -165
rect 4035 -185 4050 -165
rect 4000 -215 4050 -185
rect 4000 -235 4015 -215
rect 4035 -235 4050 -215
rect 4000 -265 4050 -235
rect 4000 -285 4015 -265
rect 4035 -285 4050 -265
rect 4000 -315 4050 -285
rect 4000 -335 4015 -315
rect 4035 -335 4050 -315
rect 4000 -365 4050 -335
rect 4000 -385 4015 -365
rect 4035 -385 4050 -365
rect 4000 -415 4050 -385
rect 4000 -435 4015 -415
rect 4035 -435 4050 -415
rect 4000 -465 4050 -435
rect 4000 -485 4015 -465
rect 4035 -485 4050 -465
rect 4000 -515 4050 -485
rect 4000 -535 4015 -515
rect 4035 -535 4050 -515
rect 4000 -565 4050 -535
rect 4000 -585 4015 -565
rect 4035 -585 4050 -565
rect 4000 -615 4050 -585
rect 4000 -635 4015 -615
rect 4035 -635 4050 -615
rect 4000 -665 4050 -635
rect 4000 -685 4015 -665
rect 4035 -685 4050 -665
rect 4000 -715 4050 -685
rect 4000 -735 4015 -715
rect 4035 -735 4050 -715
rect 4000 -765 4050 -735
rect 4000 -785 4015 -765
rect 4035 -785 4050 -765
rect 4000 -800 4050 -785
rect 4150 -115 4200 -100
rect 4150 -135 4165 -115
rect 4185 -135 4200 -115
rect 4150 -165 4200 -135
rect 4150 -185 4165 -165
rect 4185 -185 4200 -165
rect 4150 -215 4200 -185
rect 4150 -235 4165 -215
rect 4185 -235 4200 -215
rect 4150 -265 4200 -235
rect 4150 -285 4165 -265
rect 4185 -285 4200 -265
rect 4150 -315 4200 -285
rect 4150 -335 4165 -315
rect 4185 -335 4200 -315
rect 4150 -365 4200 -335
rect 4150 -385 4165 -365
rect 4185 -385 4200 -365
rect 4150 -415 4200 -385
rect 4150 -435 4165 -415
rect 4185 -435 4200 -415
rect 4150 -465 4200 -435
rect 4150 -485 4165 -465
rect 4185 -485 4200 -465
rect 4150 -515 4200 -485
rect 4150 -535 4165 -515
rect 4185 -535 4200 -515
rect 4150 -565 4200 -535
rect 4150 -585 4165 -565
rect 4185 -585 4200 -565
rect 4150 -615 4200 -585
rect 4150 -635 4165 -615
rect 4185 -635 4200 -615
rect 4150 -665 4200 -635
rect 4150 -685 4165 -665
rect 4185 -685 4200 -665
rect 4150 -715 4200 -685
rect 4150 -735 4165 -715
rect 4185 -735 4200 -715
rect 4150 -765 4200 -735
rect 4150 -785 4165 -765
rect 4185 -785 4200 -765
rect 4150 -800 4200 -785
rect 4300 -115 4350 -100
rect 4300 -135 4315 -115
rect 4335 -135 4350 -115
rect 4300 -165 4350 -135
rect 4300 -185 4315 -165
rect 4335 -185 4350 -165
rect 4300 -215 4350 -185
rect 4300 -235 4315 -215
rect 4335 -235 4350 -215
rect 4300 -265 4350 -235
rect 4300 -285 4315 -265
rect 4335 -285 4350 -265
rect 4300 -315 4350 -285
rect 4300 -335 4315 -315
rect 4335 -335 4350 -315
rect 4300 -365 4350 -335
rect 4300 -385 4315 -365
rect 4335 -385 4350 -365
rect 4300 -415 4350 -385
rect 4300 -435 4315 -415
rect 4335 -435 4350 -415
rect 4300 -465 4350 -435
rect 4300 -485 4315 -465
rect 4335 -485 4350 -465
rect 4300 -515 4350 -485
rect 4300 -535 4315 -515
rect 4335 -535 4350 -515
rect 4300 -565 4350 -535
rect 4300 -585 4315 -565
rect 4335 -585 4350 -565
rect 4300 -615 4350 -585
rect 4300 -635 4315 -615
rect 4335 -635 4350 -615
rect 4300 -665 4350 -635
rect 4300 -685 4315 -665
rect 4335 -685 4350 -665
rect 4300 -715 4350 -685
rect 4300 -735 4315 -715
rect 4335 -735 4350 -715
rect 4300 -765 4350 -735
rect 4300 -785 4315 -765
rect 4335 -785 4350 -765
rect 4300 -800 4350 -785
rect 4450 -115 4500 -100
rect 4450 -135 4465 -115
rect 4485 -135 4500 -115
rect 4450 -165 4500 -135
rect 4450 -185 4465 -165
rect 4485 -185 4500 -165
rect 4450 -215 4500 -185
rect 4450 -235 4465 -215
rect 4485 -235 4500 -215
rect 4450 -265 4500 -235
rect 4450 -285 4465 -265
rect 4485 -285 4500 -265
rect 4450 -315 4500 -285
rect 4450 -335 4465 -315
rect 4485 -335 4500 -315
rect 4450 -365 4500 -335
rect 4450 -385 4465 -365
rect 4485 -385 4500 -365
rect 4450 -415 4500 -385
rect 4450 -435 4465 -415
rect 4485 -435 4500 -415
rect 4450 -465 4500 -435
rect 4450 -485 4465 -465
rect 4485 -485 4500 -465
rect 4450 -515 4500 -485
rect 4450 -535 4465 -515
rect 4485 -535 4500 -515
rect 4450 -565 4500 -535
rect 4450 -585 4465 -565
rect 4485 -585 4500 -565
rect 4450 -615 4500 -585
rect 4450 -635 4465 -615
rect 4485 -635 4500 -615
rect 4450 -665 4500 -635
rect 4450 -685 4465 -665
rect 4485 -685 4500 -665
rect 4450 -715 4500 -685
rect 4450 -735 4465 -715
rect 4485 -735 4500 -715
rect 4450 -765 4500 -735
rect 4450 -785 4465 -765
rect 4485 -785 4500 -765
rect 4450 -800 4500 -785
rect 4600 -115 4650 -100
rect 4600 -135 4615 -115
rect 4635 -135 4650 -115
rect 4600 -165 4650 -135
rect 4600 -185 4615 -165
rect 4635 -185 4650 -165
rect 4600 -215 4650 -185
rect 4600 -235 4615 -215
rect 4635 -235 4650 -215
rect 4600 -265 4650 -235
rect 4600 -285 4615 -265
rect 4635 -285 4650 -265
rect 4600 -315 4650 -285
rect 4600 -335 4615 -315
rect 4635 -335 4650 -315
rect 4600 -365 4650 -335
rect 4600 -385 4615 -365
rect 4635 -385 4650 -365
rect 4600 -415 4650 -385
rect 4600 -435 4615 -415
rect 4635 -435 4650 -415
rect 4600 -465 4650 -435
rect 4600 -485 4615 -465
rect 4635 -485 4650 -465
rect 4600 -515 4650 -485
rect 4600 -535 4615 -515
rect 4635 -535 4650 -515
rect 4600 -565 4650 -535
rect 4600 -585 4615 -565
rect 4635 -585 4650 -565
rect 4600 -615 4650 -585
rect 4600 -635 4615 -615
rect 4635 -635 4650 -615
rect 4600 -665 4650 -635
rect 4600 -685 4615 -665
rect 4635 -685 4650 -665
rect 4600 -715 4650 -685
rect 4600 -735 4615 -715
rect 4635 -735 4650 -715
rect 4600 -765 4650 -735
rect 4600 -785 4615 -765
rect 4635 -785 4650 -765
rect 4600 -800 4650 -785
rect 4750 -115 4800 -100
rect 4750 -135 4765 -115
rect 4785 -135 4800 -115
rect 4750 -165 4800 -135
rect 4750 -185 4765 -165
rect 4785 -185 4800 -165
rect 4750 -215 4800 -185
rect 4750 -235 4765 -215
rect 4785 -235 4800 -215
rect 4750 -265 4800 -235
rect 4750 -285 4765 -265
rect 4785 -285 4800 -265
rect 4750 -315 4800 -285
rect 4750 -335 4765 -315
rect 4785 -335 4800 -315
rect 4750 -365 4800 -335
rect 4750 -385 4765 -365
rect 4785 -385 4800 -365
rect 4750 -415 4800 -385
rect 4750 -435 4765 -415
rect 4785 -435 4800 -415
rect 4750 -465 4800 -435
rect 4750 -485 4765 -465
rect 4785 -485 4800 -465
rect 4750 -515 4800 -485
rect 4750 -535 4765 -515
rect 4785 -535 4800 -515
rect 4750 -565 4800 -535
rect 4750 -585 4765 -565
rect 4785 -585 4800 -565
rect 4750 -615 4800 -585
rect 4750 -635 4765 -615
rect 4785 -635 4800 -615
rect 4750 -665 4800 -635
rect 4750 -685 4765 -665
rect 4785 -685 4800 -665
rect 4750 -715 4800 -685
rect 4750 -735 4765 -715
rect 4785 -735 4800 -715
rect 4750 -765 4800 -735
rect 4750 -785 4765 -765
rect 4785 -785 4800 -765
rect 4750 -800 4800 -785
rect 4900 -800 4950 -100
rect 5050 -115 5100 -100
rect 5050 -135 5065 -115
rect 5085 -135 5100 -115
rect 5050 -165 5100 -135
rect 5050 -185 5065 -165
rect 5085 -185 5100 -165
rect 5050 -215 5100 -185
rect 5050 -235 5065 -215
rect 5085 -235 5100 -215
rect 5050 -265 5100 -235
rect 5050 -285 5065 -265
rect 5085 -285 5100 -265
rect 5050 -315 5100 -285
rect 5050 -335 5065 -315
rect 5085 -335 5100 -315
rect 5050 -365 5100 -335
rect 5050 -385 5065 -365
rect 5085 -385 5100 -365
rect 5050 -415 5100 -385
rect 5050 -435 5065 -415
rect 5085 -435 5100 -415
rect 5050 -465 5100 -435
rect 5050 -485 5065 -465
rect 5085 -485 5100 -465
rect 5050 -515 5100 -485
rect 5050 -535 5065 -515
rect 5085 -535 5100 -515
rect 5050 -565 5100 -535
rect 5050 -585 5065 -565
rect 5085 -585 5100 -565
rect 5050 -615 5100 -585
rect 5050 -635 5065 -615
rect 5085 -635 5100 -615
rect 5050 -665 5100 -635
rect 5050 -685 5065 -665
rect 5085 -685 5100 -665
rect 5050 -715 5100 -685
rect 5050 -735 5065 -715
rect 5085 -735 5100 -715
rect 5050 -765 5100 -735
rect 5050 -785 5065 -765
rect 5085 -785 5100 -765
rect 5050 -800 5100 -785
rect 5200 -800 5250 -100
rect 5350 -115 5400 -100
rect 5350 -135 5365 -115
rect 5385 -135 5400 -115
rect 5350 -165 5400 -135
rect 5350 -185 5365 -165
rect 5385 -185 5400 -165
rect 5350 -215 5400 -185
rect 5350 -235 5365 -215
rect 5385 -235 5400 -215
rect 5350 -265 5400 -235
rect 5350 -285 5365 -265
rect 5385 -285 5400 -265
rect 5350 -315 5400 -285
rect 5350 -335 5365 -315
rect 5385 -335 5400 -315
rect 5350 -365 5400 -335
rect 5350 -385 5365 -365
rect 5385 -385 5400 -365
rect 5350 -415 5400 -385
rect 5350 -435 5365 -415
rect 5385 -435 5400 -415
rect 5350 -465 5400 -435
rect 5350 -485 5365 -465
rect 5385 -485 5400 -465
rect 5350 -515 5400 -485
rect 5350 -535 5365 -515
rect 5385 -535 5400 -515
rect 5350 -565 5400 -535
rect 5350 -585 5365 -565
rect 5385 -585 5400 -565
rect 5350 -615 5400 -585
rect 5350 -635 5365 -615
rect 5385 -635 5400 -615
rect 5350 -665 5400 -635
rect 5350 -685 5365 -665
rect 5385 -685 5400 -665
rect 5350 -715 5400 -685
rect 5350 -735 5365 -715
rect 5385 -735 5400 -715
rect 5350 -765 5400 -735
rect 5350 -785 5365 -765
rect 5385 -785 5400 -765
rect 5350 -800 5400 -785
rect 5500 -800 5550 -100
rect 5650 -115 5700 -100
rect 5650 -135 5665 -115
rect 5685 -135 5700 -115
rect 5650 -165 5700 -135
rect 5650 -185 5665 -165
rect 5685 -185 5700 -165
rect 5650 -215 5700 -185
rect 5650 -235 5665 -215
rect 5685 -235 5700 -215
rect 5650 -265 5700 -235
rect 5650 -285 5665 -265
rect 5685 -285 5700 -265
rect 5650 -315 5700 -285
rect 5650 -335 5665 -315
rect 5685 -335 5700 -315
rect 5650 -365 5700 -335
rect 5650 -385 5665 -365
rect 5685 -385 5700 -365
rect 5650 -415 5700 -385
rect 5650 -435 5665 -415
rect 5685 -435 5700 -415
rect 5650 -465 5700 -435
rect 5650 -485 5665 -465
rect 5685 -485 5700 -465
rect 5650 -515 5700 -485
rect 5650 -535 5665 -515
rect 5685 -535 5700 -515
rect 5650 -565 5700 -535
rect 5650 -585 5665 -565
rect 5685 -585 5700 -565
rect 5650 -615 5700 -585
rect 5650 -635 5665 -615
rect 5685 -635 5700 -615
rect 5650 -665 5700 -635
rect 5650 -685 5665 -665
rect 5685 -685 5700 -665
rect 5650 -715 5700 -685
rect 5650 -735 5665 -715
rect 5685 -735 5700 -715
rect 5650 -765 5700 -735
rect 5650 -785 5665 -765
rect 5685 -785 5700 -765
rect 5650 -800 5700 -785
rect 5800 -800 5850 -100
rect 5950 -115 6000 -100
rect 5950 -135 5965 -115
rect 5985 -135 6000 -115
rect 5950 -165 6000 -135
rect 5950 -185 5965 -165
rect 5985 -185 6000 -165
rect 5950 -215 6000 -185
rect 5950 -235 5965 -215
rect 5985 -235 6000 -215
rect 5950 -265 6000 -235
rect 5950 -285 5965 -265
rect 5985 -285 6000 -265
rect 5950 -315 6000 -285
rect 5950 -335 5965 -315
rect 5985 -335 6000 -315
rect 5950 -365 6000 -335
rect 5950 -385 5965 -365
rect 5985 -385 6000 -365
rect 5950 -415 6000 -385
rect 5950 -435 5965 -415
rect 5985 -435 6000 -415
rect 5950 -465 6000 -435
rect 5950 -485 5965 -465
rect 5985 -485 6000 -465
rect 5950 -515 6000 -485
rect 5950 -535 5965 -515
rect 5985 -535 6000 -515
rect 5950 -565 6000 -535
rect 5950 -585 5965 -565
rect 5985 -585 6000 -565
rect 5950 -615 6000 -585
rect 5950 -635 5965 -615
rect 5985 -635 6000 -615
rect 5950 -665 6000 -635
rect 5950 -685 5965 -665
rect 5985 -685 6000 -665
rect 5950 -715 6000 -685
rect 5950 -735 5965 -715
rect 5985 -735 6000 -715
rect 5950 -765 6000 -735
rect 5950 -785 5965 -765
rect 5985 -785 6000 -765
rect 5950 -800 6000 -785
rect 6100 -800 6150 -100
rect 6250 -115 6300 -100
rect 6250 -135 6265 -115
rect 6285 -135 6300 -115
rect 6250 -165 6300 -135
rect 6250 -185 6265 -165
rect 6285 -185 6300 -165
rect 6250 -215 6300 -185
rect 6250 -235 6265 -215
rect 6285 -235 6300 -215
rect 6250 -265 6300 -235
rect 6250 -285 6265 -265
rect 6285 -285 6300 -265
rect 6250 -315 6300 -285
rect 6250 -335 6265 -315
rect 6285 -335 6300 -315
rect 6250 -365 6300 -335
rect 6250 -385 6265 -365
rect 6285 -385 6300 -365
rect 6250 -415 6300 -385
rect 6250 -435 6265 -415
rect 6285 -435 6300 -415
rect 6250 -465 6300 -435
rect 6250 -485 6265 -465
rect 6285 -485 6300 -465
rect 6250 -515 6300 -485
rect 6250 -535 6265 -515
rect 6285 -535 6300 -515
rect 6250 -565 6300 -535
rect 6250 -585 6265 -565
rect 6285 -585 6300 -565
rect 6250 -615 6300 -585
rect 6250 -635 6265 -615
rect 6285 -635 6300 -615
rect 6250 -665 6300 -635
rect 6250 -685 6265 -665
rect 6285 -685 6300 -665
rect 6250 -715 6300 -685
rect 6250 -735 6265 -715
rect 6285 -735 6300 -715
rect 6250 -765 6300 -735
rect 6250 -785 6265 -765
rect 6285 -785 6300 -765
rect 6250 -800 6300 -785
rect 6400 -800 6450 -100
rect 6550 -115 6600 -100
rect 6550 -135 6565 -115
rect 6585 -135 6600 -115
rect 6550 -165 6600 -135
rect 6550 -185 6565 -165
rect 6585 -185 6600 -165
rect 6550 -215 6600 -185
rect 6550 -235 6565 -215
rect 6585 -235 6600 -215
rect 6550 -265 6600 -235
rect 6550 -285 6565 -265
rect 6585 -285 6600 -265
rect 6550 -315 6600 -285
rect 6550 -335 6565 -315
rect 6585 -335 6600 -315
rect 6550 -365 6600 -335
rect 6550 -385 6565 -365
rect 6585 -385 6600 -365
rect 6550 -415 6600 -385
rect 6550 -435 6565 -415
rect 6585 -435 6600 -415
rect 6550 -465 6600 -435
rect 6550 -485 6565 -465
rect 6585 -485 6600 -465
rect 6550 -515 6600 -485
rect 6550 -535 6565 -515
rect 6585 -535 6600 -515
rect 6550 -565 6600 -535
rect 6550 -585 6565 -565
rect 6585 -585 6600 -565
rect 6550 -615 6600 -585
rect 6550 -635 6565 -615
rect 6585 -635 6600 -615
rect 6550 -665 6600 -635
rect 6550 -685 6565 -665
rect 6585 -685 6600 -665
rect 6550 -715 6600 -685
rect 6550 -735 6565 -715
rect 6585 -735 6600 -715
rect 6550 -765 6600 -735
rect 6550 -785 6565 -765
rect 6585 -785 6600 -765
rect 6550 -800 6600 -785
rect 6700 -800 6750 -100
rect 6850 -115 6900 -100
rect 6850 -135 6865 -115
rect 6885 -135 6900 -115
rect 6850 -165 6900 -135
rect 6850 -185 6865 -165
rect 6885 -185 6900 -165
rect 6850 -215 6900 -185
rect 6850 -235 6865 -215
rect 6885 -235 6900 -215
rect 6850 -265 6900 -235
rect 6850 -285 6865 -265
rect 6885 -285 6900 -265
rect 6850 -315 6900 -285
rect 6850 -335 6865 -315
rect 6885 -335 6900 -315
rect 6850 -365 6900 -335
rect 6850 -385 6865 -365
rect 6885 -385 6900 -365
rect 6850 -415 6900 -385
rect 6850 -435 6865 -415
rect 6885 -435 6900 -415
rect 6850 -465 6900 -435
rect 6850 -485 6865 -465
rect 6885 -485 6900 -465
rect 6850 -515 6900 -485
rect 6850 -535 6865 -515
rect 6885 -535 6900 -515
rect 6850 -565 6900 -535
rect 6850 -585 6865 -565
rect 6885 -585 6900 -565
rect 6850 -615 6900 -585
rect 6850 -635 6865 -615
rect 6885 -635 6900 -615
rect 6850 -665 6900 -635
rect 6850 -685 6865 -665
rect 6885 -685 6900 -665
rect 6850 -715 6900 -685
rect 6850 -735 6865 -715
rect 6885 -735 6900 -715
rect 6850 -765 6900 -735
rect 6850 -785 6865 -765
rect 6885 -785 6900 -765
rect 6850 -800 6900 -785
rect 7000 -800 7050 -100
rect 7150 -115 7200 -100
rect 7150 -135 7165 -115
rect 7185 -135 7200 -115
rect 7150 -165 7200 -135
rect 7150 -185 7165 -165
rect 7185 -185 7200 -165
rect 7150 -215 7200 -185
rect 7150 -235 7165 -215
rect 7185 -235 7200 -215
rect 7150 -265 7200 -235
rect 7150 -285 7165 -265
rect 7185 -285 7200 -265
rect 7150 -315 7200 -285
rect 7150 -335 7165 -315
rect 7185 -335 7200 -315
rect 7150 -365 7200 -335
rect 7150 -385 7165 -365
rect 7185 -385 7200 -365
rect 7150 -415 7200 -385
rect 7150 -435 7165 -415
rect 7185 -435 7200 -415
rect 7150 -465 7200 -435
rect 7150 -485 7165 -465
rect 7185 -485 7200 -465
rect 7150 -515 7200 -485
rect 7150 -535 7165 -515
rect 7185 -535 7200 -515
rect 7150 -565 7200 -535
rect 7150 -585 7165 -565
rect 7185 -585 7200 -565
rect 7150 -615 7200 -585
rect 7150 -635 7165 -615
rect 7185 -635 7200 -615
rect 7150 -665 7200 -635
rect 7150 -685 7165 -665
rect 7185 -685 7200 -665
rect 7150 -715 7200 -685
rect 7150 -735 7165 -715
rect 7185 -735 7200 -715
rect 7150 -765 7200 -735
rect 7150 -785 7165 -765
rect 7185 -785 7200 -765
rect 7150 -800 7200 -785
rect 7300 -800 7350 -100
rect 7450 -800 7500 -100
rect 7600 -800 7650 -100
rect 7750 -800 7800 -100
rect 7900 -800 7950 -100
rect 8050 -800 8100 -100
rect 8200 -800 8250 -100
rect 8350 -115 8400 -100
rect 8350 -135 8365 -115
rect 8385 -135 8400 -115
rect 8350 -165 8400 -135
rect 8350 -185 8365 -165
rect 8385 -185 8400 -165
rect 8350 -215 8400 -185
rect 8350 -235 8365 -215
rect 8385 -235 8400 -215
rect 8350 -265 8400 -235
rect 8350 -285 8365 -265
rect 8385 -285 8400 -265
rect 8350 -315 8400 -285
rect 8350 -335 8365 -315
rect 8385 -335 8400 -315
rect 8350 -365 8400 -335
rect 8350 -385 8365 -365
rect 8385 -385 8400 -365
rect 8350 -415 8400 -385
rect 8350 -435 8365 -415
rect 8385 -435 8400 -415
rect 8350 -465 8400 -435
rect 8350 -485 8365 -465
rect 8385 -485 8400 -465
rect 8350 -515 8400 -485
rect 8350 -535 8365 -515
rect 8385 -535 8400 -515
rect 8350 -565 8400 -535
rect 8350 -585 8365 -565
rect 8385 -585 8400 -565
rect 8350 -615 8400 -585
rect 8350 -635 8365 -615
rect 8385 -635 8400 -615
rect 8350 -665 8400 -635
rect 8350 -685 8365 -665
rect 8385 -685 8400 -665
rect 8350 -715 8400 -685
rect 8350 -735 8365 -715
rect 8385 -735 8400 -715
rect 8350 -765 8400 -735
rect 8350 -785 8365 -765
rect 8385 -785 8400 -765
rect 8350 -800 8400 -785
rect 8500 -800 8550 -100
rect 8650 -800 8700 -100
rect 8800 -800 8850 -100
rect 8950 -800 9000 -100
rect 9100 -800 9150 -100
rect 9250 -800 9300 -100
rect 9400 -800 9450 -100
rect 9550 -115 9600 -100
rect 9550 -135 9565 -115
rect 9585 -135 9600 -115
rect 9550 -165 9600 -135
rect 9550 -185 9565 -165
rect 9585 -185 9600 -165
rect 9550 -215 9600 -185
rect 9550 -235 9565 -215
rect 9585 -235 9600 -215
rect 9550 -265 9600 -235
rect 9550 -285 9565 -265
rect 9585 -285 9600 -265
rect 9550 -315 9600 -285
rect 9550 -335 9565 -315
rect 9585 -335 9600 -315
rect 9550 -365 9600 -335
rect 9550 -385 9565 -365
rect 9585 -385 9600 -365
rect 9550 -415 9600 -385
rect 9550 -435 9565 -415
rect 9585 -435 9600 -415
rect 9550 -465 9600 -435
rect 9550 -485 9565 -465
rect 9585 -485 9600 -465
rect 9550 -515 9600 -485
rect 9550 -535 9565 -515
rect 9585 -535 9600 -515
rect 9550 -565 9600 -535
rect 9550 -585 9565 -565
rect 9585 -585 9600 -565
rect 9550 -615 9600 -585
rect 9550 -635 9565 -615
rect 9585 -635 9600 -615
rect 9550 -665 9600 -635
rect 9550 -685 9565 -665
rect 9585 -685 9600 -665
rect 9550 -715 9600 -685
rect 9550 -735 9565 -715
rect 9585 -735 9600 -715
rect 9550 -765 9600 -735
rect 9550 -785 9565 -765
rect 9585 -785 9600 -765
rect 9550 -800 9600 -785
rect 9700 -800 9750 -100
rect 9850 -800 9900 -100
rect 10000 -800 10050 -100
rect 10150 -800 10200 -100
rect 10300 -800 10350 -100
rect 10450 -800 10500 -100
rect 10600 -800 10650 -100
rect 10750 -115 10800 -100
rect 10750 -135 10765 -115
rect 10785 -135 10800 -115
rect 10750 -165 10800 -135
rect 10750 -185 10765 -165
rect 10785 -185 10800 -165
rect 10750 -215 10800 -185
rect 10750 -235 10765 -215
rect 10785 -235 10800 -215
rect 10750 -265 10800 -235
rect 10750 -285 10765 -265
rect 10785 -285 10800 -265
rect 10750 -315 10800 -285
rect 10750 -335 10765 -315
rect 10785 -335 10800 -315
rect 10750 -365 10800 -335
rect 10750 -385 10765 -365
rect 10785 -385 10800 -365
rect 10750 -415 10800 -385
rect 10750 -435 10765 -415
rect 10785 -435 10800 -415
rect 10750 -465 10800 -435
rect 10750 -485 10765 -465
rect 10785 -485 10800 -465
rect 10750 -515 10800 -485
rect 10750 -535 10765 -515
rect 10785 -535 10800 -515
rect 10750 -565 10800 -535
rect 10750 -585 10765 -565
rect 10785 -585 10800 -565
rect 10750 -615 10800 -585
rect 10750 -635 10765 -615
rect 10785 -635 10800 -615
rect 10750 -665 10800 -635
rect 10750 -685 10765 -665
rect 10785 -685 10800 -665
rect 10750 -715 10800 -685
rect 10750 -735 10765 -715
rect 10785 -735 10800 -715
rect 10750 -765 10800 -735
rect 10750 -785 10765 -765
rect 10785 -785 10800 -765
rect 10750 -800 10800 -785
rect 10900 -800 10950 -100
rect 11050 -800 11100 -100
rect 11200 -800 11250 -100
rect 11350 -800 11400 -100
rect 11500 -800 11550 -100
rect 11650 -800 11700 -100
rect 11800 -800 11850 -100
rect 11950 -115 12000 -100
rect 11950 -135 11965 -115
rect 11985 -135 12000 -115
rect 11950 -165 12000 -135
rect 11950 -185 11965 -165
rect 11985 -185 12000 -165
rect 11950 -215 12000 -185
rect 11950 -235 11965 -215
rect 11985 -235 12000 -215
rect 11950 -265 12000 -235
rect 11950 -285 11965 -265
rect 11985 -285 12000 -265
rect 11950 -315 12000 -285
rect 11950 -335 11965 -315
rect 11985 -335 12000 -315
rect 11950 -365 12000 -335
rect 11950 -385 11965 -365
rect 11985 -385 12000 -365
rect 11950 -415 12000 -385
rect 11950 -435 11965 -415
rect 11985 -435 12000 -415
rect 11950 -465 12000 -435
rect 11950 -485 11965 -465
rect 11985 -485 12000 -465
rect 11950 -515 12000 -485
rect 11950 -535 11965 -515
rect 11985 -535 12000 -515
rect 11950 -565 12000 -535
rect 11950 -585 11965 -565
rect 11985 -585 12000 -565
rect 11950 -615 12000 -585
rect 11950 -635 11965 -615
rect 11985 -635 12000 -615
rect 11950 -665 12000 -635
rect 11950 -685 11965 -665
rect 11985 -685 12000 -665
rect 11950 -715 12000 -685
rect 11950 -735 11965 -715
rect 11985 -735 12000 -715
rect 11950 -765 12000 -735
rect 11950 -785 11965 -765
rect 11985 -785 12000 -765
rect 11950 -800 12000 -785
rect 12100 -800 12150 -100
rect 12250 -115 12300 -100
rect 12250 -135 12265 -115
rect 12285 -135 12300 -115
rect 12250 -165 12300 -135
rect 12250 -185 12265 -165
rect 12285 -185 12300 -165
rect 12250 -215 12300 -185
rect 12250 -235 12265 -215
rect 12285 -235 12300 -215
rect 12250 -265 12300 -235
rect 12250 -285 12265 -265
rect 12285 -285 12300 -265
rect 12250 -315 12300 -285
rect 12250 -335 12265 -315
rect 12285 -335 12300 -315
rect 12250 -365 12300 -335
rect 12250 -385 12265 -365
rect 12285 -385 12300 -365
rect 12250 -415 12300 -385
rect 12250 -435 12265 -415
rect 12285 -435 12300 -415
rect 12250 -465 12300 -435
rect 12250 -485 12265 -465
rect 12285 -485 12300 -465
rect 12250 -515 12300 -485
rect 12250 -535 12265 -515
rect 12285 -535 12300 -515
rect 12250 -565 12300 -535
rect 12250 -585 12265 -565
rect 12285 -585 12300 -565
rect 12250 -615 12300 -585
rect 12250 -635 12265 -615
rect 12285 -635 12300 -615
rect 12250 -665 12300 -635
rect 12250 -685 12265 -665
rect 12285 -685 12300 -665
rect 12250 -715 12300 -685
rect 12250 -735 12265 -715
rect 12285 -735 12300 -715
rect 12250 -765 12300 -735
rect 12250 -785 12265 -765
rect 12285 -785 12300 -765
rect 12250 -800 12300 -785
rect 12400 -800 12450 -100
rect 12550 -115 12600 -100
rect 12550 -135 12565 -115
rect 12585 -135 12600 -115
rect 12550 -165 12600 -135
rect 12550 -185 12565 -165
rect 12585 -185 12600 -165
rect 12550 -215 12600 -185
rect 12550 -235 12565 -215
rect 12585 -235 12600 -215
rect 12550 -265 12600 -235
rect 12550 -285 12565 -265
rect 12585 -285 12600 -265
rect 12550 -315 12600 -285
rect 12550 -335 12565 -315
rect 12585 -335 12600 -315
rect 12550 -365 12600 -335
rect 12550 -385 12565 -365
rect 12585 -385 12600 -365
rect 12550 -415 12600 -385
rect 12550 -435 12565 -415
rect 12585 -435 12600 -415
rect 12550 -465 12600 -435
rect 12550 -485 12565 -465
rect 12585 -485 12600 -465
rect 12550 -515 12600 -485
rect 12550 -535 12565 -515
rect 12585 -535 12600 -515
rect 12550 -565 12600 -535
rect 12550 -585 12565 -565
rect 12585 -585 12600 -565
rect 12550 -615 12600 -585
rect 12550 -635 12565 -615
rect 12585 -635 12600 -615
rect 12550 -665 12600 -635
rect 12550 -685 12565 -665
rect 12585 -685 12600 -665
rect 12550 -715 12600 -685
rect 12550 -735 12565 -715
rect 12585 -735 12600 -715
rect 12550 -765 12600 -735
rect 12550 -785 12565 -765
rect 12585 -785 12600 -765
rect 12550 -800 12600 -785
rect 12700 -800 12750 -100
rect 12850 -115 12900 -100
rect 12850 -135 12865 -115
rect 12885 -135 12900 -115
rect 12850 -165 12900 -135
rect 12850 -185 12865 -165
rect 12885 -185 12900 -165
rect 12850 -215 12900 -185
rect 12850 -235 12865 -215
rect 12885 -235 12900 -215
rect 12850 -265 12900 -235
rect 12850 -285 12865 -265
rect 12885 -285 12900 -265
rect 12850 -315 12900 -285
rect 12850 -335 12865 -315
rect 12885 -335 12900 -315
rect 12850 -365 12900 -335
rect 12850 -385 12865 -365
rect 12885 -385 12900 -365
rect 12850 -415 12900 -385
rect 12850 -435 12865 -415
rect 12885 -435 12900 -415
rect 12850 -465 12900 -435
rect 12850 -485 12865 -465
rect 12885 -485 12900 -465
rect 12850 -515 12900 -485
rect 12850 -535 12865 -515
rect 12885 -535 12900 -515
rect 12850 -565 12900 -535
rect 12850 -585 12865 -565
rect 12885 -585 12900 -565
rect 12850 -615 12900 -585
rect 12850 -635 12865 -615
rect 12885 -635 12900 -615
rect 12850 -665 12900 -635
rect 12850 -685 12865 -665
rect 12885 -685 12900 -665
rect 12850 -715 12900 -685
rect 12850 -735 12865 -715
rect 12885 -735 12900 -715
rect 12850 -765 12900 -735
rect 12850 -785 12865 -765
rect 12885 -785 12900 -765
rect 12850 -800 12900 -785
rect 13000 -800 13050 -100
rect 13150 -115 13200 -100
rect 13150 -135 13165 -115
rect 13185 -135 13200 -115
rect 13150 -165 13200 -135
rect 13150 -185 13165 -165
rect 13185 -185 13200 -165
rect 13150 -215 13200 -185
rect 13150 -235 13165 -215
rect 13185 -235 13200 -215
rect 13150 -265 13200 -235
rect 13150 -285 13165 -265
rect 13185 -285 13200 -265
rect 13150 -315 13200 -285
rect 13150 -335 13165 -315
rect 13185 -335 13200 -315
rect 13150 -365 13200 -335
rect 13150 -385 13165 -365
rect 13185 -385 13200 -365
rect 13150 -415 13200 -385
rect 13150 -435 13165 -415
rect 13185 -435 13200 -415
rect 13150 -465 13200 -435
rect 13150 -485 13165 -465
rect 13185 -485 13200 -465
rect 13150 -515 13200 -485
rect 13150 -535 13165 -515
rect 13185 -535 13200 -515
rect 13150 -565 13200 -535
rect 13150 -585 13165 -565
rect 13185 -585 13200 -565
rect 13150 -615 13200 -585
rect 13150 -635 13165 -615
rect 13185 -635 13200 -615
rect 13150 -665 13200 -635
rect 13150 -685 13165 -665
rect 13185 -685 13200 -665
rect 13150 -715 13200 -685
rect 13150 -735 13165 -715
rect 13185 -735 13200 -715
rect 13150 -765 13200 -735
rect 13150 -785 13165 -765
rect 13185 -785 13200 -765
rect 13150 -800 13200 -785
rect 13300 -800 13350 -100
rect 13450 -115 13500 -100
rect 13450 -135 13465 -115
rect 13485 -135 13500 -115
rect 13450 -165 13500 -135
rect 13450 -185 13465 -165
rect 13485 -185 13500 -165
rect 13450 -215 13500 -185
rect 13450 -235 13465 -215
rect 13485 -235 13500 -215
rect 13450 -265 13500 -235
rect 13450 -285 13465 -265
rect 13485 -285 13500 -265
rect 13450 -315 13500 -285
rect 13450 -335 13465 -315
rect 13485 -335 13500 -315
rect 13450 -365 13500 -335
rect 13450 -385 13465 -365
rect 13485 -385 13500 -365
rect 13450 -415 13500 -385
rect 13450 -435 13465 -415
rect 13485 -435 13500 -415
rect 13450 -465 13500 -435
rect 13450 -485 13465 -465
rect 13485 -485 13500 -465
rect 13450 -515 13500 -485
rect 13450 -535 13465 -515
rect 13485 -535 13500 -515
rect 13450 -565 13500 -535
rect 13450 -585 13465 -565
rect 13485 -585 13500 -565
rect 13450 -615 13500 -585
rect 13450 -635 13465 -615
rect 13485 -635 13500 -615
rect 13450 -665 13500 -635
rect 13450 -685 13465 -665
rect 13485 -685 13500 -665
rect 13450 -715 13500 -685
rect 13450 -735 13465 -715
rect 13485 -735 13500 -715
rect 13450 -765 13500 -735
rect 13450 -785 13465 -765
rect 13485 -785 13500 -765
rect 13450 -800 13500 -785
rect 13600 -800 13650 -100
rect 13750 -115 13800 -100
rect 13750 -135 13765 -115
rect 13785 -135 13800 -115
rect 13750 -165 13800 -135
rect 13750 -185 13765 -165
rect 13785 -185 13800 -165
rect 13750 -215 13800 -185
rect 13750 -235 13765 -215
rect 13785 -235 13800 -215
rect 13750 -265 13800 -235
rect 13750 -285 13765 -265
rect 13785 -285 13800 -265
rect 13750 -315 13800 -285
rect 13750 -335 13765 -315
rect 13785 -335 13800 -315
rect 13750 -365 13800 -335
rect 13750 -385 13765 -365
rect 13785 -385 13800 -365
rect 13750 -415 13800 -385
rect 13750 -435 13765 -415
rect 13785 -435 13800 -415
rect 13750 -465 13800 -435
rect 13750 -485 13765 -465
rect 13785 -485 13800 -465
rect 13750 -515 13800 -485
rect 13750 -535 13765 -515
rect 13785 -535 13800 -515
rect 13750 -565 13800 -535
rect 13750 -585 13765 -565
rect 13785 -585 13800 -565
rect 13750 -615 13800 -585
rect 13750 -635 13765 -615
rect 13785 -635 13800 -615
rect 13750 -665 13800 -635
rect 13750 -685 13765 -665
rect 13785 -685 13800 -665
rect 13750 -715 13800 -685
rect 13750 -735 13765 -715
rect 13785 -735 13800 -715
rect 13750 -765 13800 -735
rect 13750 -785 13765 -765
rect 13785 -785 13800 -765
rect 13750 -800 13800 -785
rect 13900 -800 13950 -100
rect 14050 -115 14100 -100
rect 14050 -135 14065 -115
rect 14085 -135 14100 -115
rect 14050 -165 14100 -135
rect 14050 -185 14065 -165
rect 14085 -185 14100 -165
rect 14050 -215 14100 -185
rect 14050 -235 14065 -215
rect 14085 -235 14100 -215
rect 14050 -265 14100 -235
rect 14050 -285 14065 -265
rect 14085 -285 14100 -265
rect 14050 -315 14100 -285
rect 14050 -335 14065 -315
rect 14085 -335 14100 -315
rect 14050 -365 14100 -335
rect 14050 -385 14065 -365
rect 14085 -385 14100 -365
rect 14050 -415 14100 -385
rect 14050 -435 14065 -415
rect 14085 -435 14100 -415
rect 14050 -465 14100 -435
rect 14050 -485 14065 -465
rect 14085 -485 14100 -465
rect 14050 -515 14100 -485
rect 14050 -535 14065 -515
rect 14085 -535 14100 -515
rect 14050 -565 14100 -535
rect 14050 -585 14065 -565
rect 14085 -585 14100 -565
rect 14050 -615 14100 -585
rect 14050 -635 14065 -615
rect 14085 -635 14100 -615
rect 14050 -665 14100 -635
rect 14050 -685 14065 -665
rect 14085 -685 14100 -665
rect 14050 -715 14100 -685
rect 14050 -735 14065 -715
rect 14085 -735 14100 -715
rect 14050 -765 14100 -735
rect 14050 -785 14065 -765
rect 14085 -785 14100 -765
rect 14050 -800 14100 -785
rect 14200 -800 14250 -100
rect 14350 -115 14400 -100
rect 14350 -135 14365 -115
rect 14385 -135 14400 -115
rect 14350 -165 14400 -135
rect 14350 -185 14365 -165
rect 14385 -185 14400 -165
rect 14350 -215 14400 -185
rect 14350 -235 14365 -215
rect 14385 -235 14400 -215
rect 14350 -265 14400 -235
rect 14350 -285 14365 -265
rect 14385 -285 14400 -265
rect 14350 -315 14400 -285
rect 14350 -335 14365 -315
rect 14385 -335 14400 -315
rect 14350 -365 14400 -335
rect 14350 -385 14365 -365
rect 14385 -385 14400 -365
rect 14350 -415 14400 -385
rect 14350 -435 14365 -415
rect 14385 -435 14400 -415
rect 14350 -465 14400 -435
rect 14350 -485 14365 -465
rect 14385 -485 14400 -465
rect 14350 -515 14400 -485
rect 14350 -535 14365 -515
rect 14385 -535 14400 -515
rect 14350 -565 14400 -535
rect 14350 -585 14365 -565
rect 14385 -585 14400 -565
rect 14350 -615 14400 -585
rect 14350 -635 14365 -615
rect 14385 -635 14400 -615
rect 14350 -665 14400 -635
rect 14350 -685 14365 -665
rect 14385 -685 14400 -665
rect 14350 -715 14400 -685
rect 14350 -735 14365 -715
rect 14385 -735 14400 -715
rect 14350 -765 14400 -735
rect 14350 -785 14365 -765
rect 14385 -785 14400 -765
rect 14350 -800 14400 -785
rect 14500 -800 14550 -100
rect 14650 -800 14700 -100
rect 14800 -800 14850 -100
rect 14950 -800 15000 -100
rect 15100 -800 15150 -100
rect 15250 -800 15300 -100
rect 15400 -800 15450 -100
rect 15550 -115 15600 -100
rect 15550 -135 15565 -115
rect 15585 -135 15600 -115
rect 15550 -165 15600 -135
rect 15550 -185 15565 -165
rect 15585 -185 15600 -165
rect 15550 -215 15600 -185
rect 15550 -235 15565 -215
rect 15585 -235 15600 -215
rect 15550 -265 15600 -235
rect 15550 -285 15565 -265
rect 15585 -285 15600 -265
rect 15550 -315 15600 -285
rect 15550 -335 15565 -315
rect 15585 -335 15600 -315
rect 15550 -365 15600 -335
rect 15550 -385 15565 -365
rect 15585 -385 15600 -365
rect 15550 -415 15600 -385
rect 15550 -435 15565 -415
rect 15585 -435 15600 -415
rect 15550 -465 15600 -435
rect 15550 -485 15565 -465
rect 15585 -485 15600 -465
rect 15550 -515 15600 -485
rect 15550 -535 15565 -515
rect 15585 -535 15600 -515
rect 15550 -565 15600 -535
rect 15550 -585 15565 -565
rect 15585 -585 15600 -565
rect 15550 -615 15600 -585
rect 15550 -635 15565 -615
rect 15585 -635 15600 -615
rect 15550 -665 15600 -635
rect 15550 -685 15565 -665
rect 15585 -685 15600 -665
rect 15550 -715 15600 -685
rect 15550 -735 15565 -715
rect 15585 -735 15600 -715
rect 15550 -765 15600 -735
rect 15550 -785 15565 -765
rect 15585 -785 15600 -765
rect 15550 -800 15600 -785
rect 15700 -800 15750 -100
rect 15850 -800 15900 -100
rect 16000 -800 16050 -100
rect 16150 -800 16200 -100
rect 16300 -800 16350 -100
rect 16450 -800 16500 -100
rect 16600 -800 16650 -100
rect 16750 -115 16800 -100
rect 16750 -135 16765 -115
rect 16785 -135 16800 -115
rect 16750 -165 16800 -135
rect 16750 -185 16765 -165
rect 16785 -185 16800 -165
rect 16750 -215 16800 -185
rect 16750 -235 16765 -215
rect 16785 -235 16800 -215
rect 16750 -265 16800 -235
rect 16750 -285 16765 -265
rect 16785 -285 16800 -265
rect 16750 -315 16800 -285
rect 16750 -335 16765 -315
rect 16785 -335 16800 -315
rect 16750 -365 16800 -335
rect 16750 -385 16765 -365
rect 16785 -385 16800 -365
rect 16750 -415 16800 -385
rect 16750 -435 16765 -415
rect 16785 -435 16800 -415
rect 16750 -465 16800 -435
rect 16750 -485 16765 -465
rect 16785 -485 16800 -465
rect 16750 -515 16800 -485
rect 16750 -535 16765 -515
rect 16785 -535 16800 -515
rect 16750 -565 16800 -535
rect 16750 -585 16765 -565
rect 16785 -585 16800 -565
rect 16750 -615 16800 -585
rect 16750 -635 16765 -615
rect 16785 -635 16800 -615
rect 16750 -665 16800 -635
rect 16750 -685 16765 -665
rect 16785 -685 16800 -665
rect 16750 -715 16800 -685
rect 16750 -735 16765 -715
rect 16785 -735 16800 -715
rect 16750 -765 16800 -735
rect 16750 -785 16765 -765
rect 16785 -785 16800 -765
rect 16750 -800 16800 -785
rect 16900 -800 16950 -100
rect 17050 -800 17100 -100
rect 17200 -800 17250 -100
rect 17350 -800 17400 -100
rect 17500 -800 17550 -100
rect 17650 -800 17700 -100
rect 17800 -800 17850 -100
rect 17950 -115 18000 -100
rect 17950 -135 17965 -115
rect 17985 -135 18000 -115
rect 17950 -165 18000 -135
rect 17950 -185 17965 -165
rect 17985 -185 18000 -165
rect 17950 -215 18000 -185
rect 17950 -235 17965 -215
rect 17985 -235 18000 -215
rect 17950 -265 18000 -235
rect 17950 -285 17965 -265
rect 17985 -285 18000 -265
rect 17950 -315 18000 -285
rect 17950 -335 17965 -315
rect 17985 -335 18000 -315
rect 17950 -365 18000 -335
rect 17950 -385 17965 -365
rect 17985 -385 18000 -365
rect 17950 -415 18000 -385
rect 17950 -435 17965 -415
rect 17985 -435 18000 -415
rect 17950 -465 18000 -435
rect 17950 -485 17965 -465
rect 17985 -485 18000 -465
rect 17950 -515 18000 -485
rect 17950 -535 17965 -515
rect 17985 -535 18000 -515
rect 17950 -565 18000 -535
rect 17950 -585 17965 -565
rect 17985 -585 18000 -565
rect 17950 -615 18000 -585
rect 17950 -635 17965 -615
rect 17985 -635 18000 -615
rect 17950 -665 18000 -635
rect 17950 -685 17965 -665
rect 17985 -685 18000 -665
rect 17950 -715 18000 -685
rect 17950 -735 17965 -715
rect 17985 -735 18000 -715
rect 17950 -765 18000 -735
rect 17950 -785 17965 -765
rect 17985 -785 18000 -765
rect 17950 -800 18000 -785
rect 18100 -800 18150 -100
rect 18250 -800 18300 -100
rect 18400 -800 18450 -100
rect 18550 -800 18600 -100
rect 18700 -800 18750 -100
rect 18850 -800 18900 -100
rect 19000 -800 19050 -100
rect 19150 -115 19200 -100
rect 19150 -135 19165 -115
rect 19185 -135 19200 -115
rect 19150 -165 19200 -135
rect 19150 -185 19165 -165
rect 19185 -185 19200 -165
rect 19150 -215 19200 -185
rect 19150 -235 19165 -215
rect 19185 -235 19200 -215
rect 19150 -265 19200 -235
rect 19150 -285 19165 -265
rect 19185 -285 19200 -265
rect 19150 -315 19200 -285
rect 19150 -335 19165 -315
rect 19185 -335 19200 -315
rect 19150 -365 19200 -335
rect 19150 -385 19165 -365
rect 19185 -385 19200 -365
rect 19150 -415 19200 -385
rect 19150 -435 19165 -415
rect 19185 -435 19200 -415
rect 19150 -465 19200 -435
rect 19150 -485 19165 -465
rect 19185 -485 19200 -465
rect 19150 -515 19200 -485
rect 19150 -535 19165 -515
rect 19185 -535 19200 -515
rect 19150 -565 19200 -535
rect 19150 -585 19165 -565
rect 19185 -585 19200 -565
rect 19150 -615 19200 -585
rect 19150 -635 19165 -615
rect 19185 -635 19200 -615
rect 19150 -665 19200 -635
rect 19150 -685 19165 -665
rect 19185 -685 19200 -665
rect 19150 -715 19200 -685
rect 19150 -735 19165 -715
rect 19185 -735 19200 -715
rect 19150 -765 19200 -735
rect 19150 -785 19165 -765
rect 19185 -785 19200 -765
rect 19150 -800 19200 -785
rect 19300 -800 19350 -100
rect 19450 -800 19500 -100
rect 19600 -800 19650 -100
rect 19750 -800 19800 -100
rect 19900 -800 19950 -100
rect 20050 -800 20100 -100
rect 20200 -800 20250 -100
rect 20350 -115 20400 -100
rect 20350 -135 20365 -115
rect 20385 -135 20400 -115
rect 20350 -165 20400 -135
rect 20350 -185 20365 -165
rect 20385 -185 20400 -165
rect 20350 -215 20400 -185
rect 20350 -235 20365 -215
rect 20385 -235 20400 -215
rect 20350 -265 20400 -235
rect 20350 -285 20365 -265
rect 20385 -285 20400 -265
rect 20350 -315 20400 -285
rect 20350 -335 20365 -315
rect 20385 -335 20400 -315
rect 20350 -365 20400 -335
rect 20350 -385 20365 -365
rect 20385 -385 20400 -365
rect 20350 -415 20400 -385
rect 20350 -435 20365 -415
rect 20385 -435 20400 -415
rect 20350 -465 20400 -435
rect 20350 -485 20365 -465
rect 20385 -485 20400 -465
rect 20350 -515 20400 -485
rect 20350 -535 20365 -515
rect 20385 -535 20400 -515
rect 20350 -565 20400 -535
rect 20350 -585 20365 -565
rect 20385 -585 20400 -565
rect 20350 -615 20400 -585
rect 20350 -635 20365 -615
rect 20385 -635 20400 -615
rect 20350 -665 20400 -635
rect 20350 -685 20365 -665
rect 20385 -685 20400 -665
rect 20350 -715 20400 -685
rect 20350 -735 20365 -715
rect 20385 -735 20400 -715
rect 20350 -765 20400 -735
rect 20350 -785 20365 -765
rect 20385 -785 20400 -765
rect 20350 -800 20400 -785
rect 20500 -800 20550 -100
rect 20650 -800 20700 -100
rect 20800 -800 20850 -100
rect 20950 -800 21000 -100
rect 21100 -800 21150 -100
rect 21250 -800 21300 -100
rect 21400 -800 21450 -100
rect 21550 -115 21600 -100
rect 21550 -135 21565 -115
rect 21585 -135 21600 -115
rect 21550 -165 21600 -135
rect 21550 -185 21565 -165
rect 21585 -185 21600 -165
rect 21550 -215 21600 -185
rect 21550 -235 21565 -215
rect 21585 -235 21600 -215
rect 21550 -265 21600 -235
rect 21550 -285 21565 -265
rect 21585 -285 21600 -265
rect 21550 -315 21600 -285
rect 21550 -335 21565 -315
rect 21585 -335 21600 -315
rect 21550 -365 21600 -335
rect 21550 -385 21565 -365
rect 21585 -385 21600 -365
rect 21550 -415 21600 -385
rect 21550 -435 21565 -415
rect 21585 -435 21600 -415
rect 21550 -465 21600 -435
rect 21550 -485 21565 -465
rect 21585 -485 21600 -465
rect 21550 -515 21600 -485
rect 21550 -535 21565 -515
rect 21585 -535 21600 -515
rect 21550 -565 21600 -535
rect 21550 -585 21565 -565
rect 21585 -585 21600 -565
rect 21550 -615 21600 -585
rect 21550 -635 21565 -615
rect 21585 -635 21600 -615
rect 21550 -665 21600 -635
rect 21550 -685 21565 -665
rect 21585 -685 21600 -665
rect 21550 -715 21600 -685
rect 21550 -735 21565 -715
rect 21585 -735 21600 -715
rect 21550 -765 21600 -735
rect 21550 -785 21565 -765
rect 21585 -785 21600 -765
rect 21550 -800 21600 -785
rect 21700 -800 21750 -100
rect 21850 -800 21900 -100
rect 22000 -800 22050 -100
rect 22150 -800 22200 -100
rect 22300 -800 22350 -100
rect 22450 -115 22500 -100
rect 22450 -135 22465 -115
rect 22485 -135 22500 -115
rect 22450 -165 22500 -135
rect 22450 -185 22465 -165
rect 22485 -185 22500 -165
rect 22450 -215 22500 -185
rect 22450 -235 22465 -215
rect 22485 -235 22500 -215
rect 22450 -265 22500 -235
rect 22450 -285 22465 -265
rect 22485 -285 22500 -265
rect 22450 -315 22500 -285
rect 22450 -335 22465 -315
rect 22485 -335 22500 -315
rect 22450 -365 22500 -335
rect 22450 -385 22465 -365
rect 22485 -385 22500 -365
rect 22450 -415 22500 -385
rect 22450 -435 22465 -415
rect 22485 -435 22500 -415
rect 22450 -465 22500 -435
rect 22450 -485 22465 -465
rect 22485 -485 22500 -465
rect 22450 -515 22500 -485
rect 22450 -535 22465 -515
rect 22485 -535 22500 -515
rect 22450 -565 22500 -535
rect 22450 -585 22465 -565
rect 22485 -585 22500 -565
rect 22450 -615 22500 -585
rect 22450 -635 22465 -615
rect 22485 -635 22500 -615
rect 22450 -665 22500 -635
rect 22450 -685 22465 -665
rect 22485 -685 22500 -665
rect 22450 -715 22500 -685
rect 22450 -735 22465 -715
rect 22485 -735 22500 -715
rect 22450 -765 22500 -735
rect 22450 -785 22465 -765
rect 22485 -785 22500 -765
rect 22450 -800 22500 -785
rect 22600 -800 22650 -100
rect 22750 -800 22800 -100
rect 22900 -800 22950 -100
rect 23050 -800 23100 -100
rect 23200 -800 23250 -100
rect 23350 -115 23400 -100
rect 23350 -135 23365 -115
rect 23385 -135 23400 -115
rect 23350 -165 23400 -135
rect 23350 -185 23365 -165
rect 23385 -185 23400 -165
rect 23350 -215 23400 -185
rect 23350 -235 23365 -215
rect 23385 -235 23400 -215
rect 23350 -265 23400 -235
rect 23350 -285 23365 -265
rect 23385 -285 23400 -265
rect 23350 -315 23400 -285
rect 23350 -335 23365 -315
rect 23385 -335 23400 -315
rect 23350 -365 23400 -335
rect 23350 -385 23365 -365
rect 23385 -385 23400 -365
rect 23350 -415 23400 -385
rect 23350 -435 23365 -415
rect 23385 -435 23400 -415
rect 23350 -465 23400 -435
rect 23350 -485 23365 -465
rect 23385 -485 23400 -465
rect 23350 -515 23400 -485
rect 23350 -535 23365 -515
rect 23385 -535 23400 -515
rect 23350 -565 23400 -535
rect 23350 -585 23365 -565
rect 23385 -585 23400 -565
rect 23350 -615 23400 -585
rect 23350 -635 23365 -615
rect 23385 -635 23400 -615
rect 23350 -665 23400 -635
rect 23350 -685 23365 -665
rect 23385 -685 23400 -665
rect 23350 -715 23400 -685
rect 23350 -735 23365 -715
rect 23385 -735 23400 -715
rect 23350 -765 23400 -735
rect 23350 -785 23365 -765
rect 23385 -785 23400 -765
rect 23350 -800 23400 -785
rect 23500 -800 23550 -100
rect 23650 -800 23700 -100
rect 23800 -800 23850 -100
rect 23950 -800 24000 -100
rect 24100 -800 24150 -100
rect 24250 -800 24300 -100
rect 24400 -800 24450 -100
rect 24550 -115 24600 -100
rect 24550 -135 24565 -115
rect 24585 -135 24600 -115
rect 24550 -165 24600 -135
rect 24550 -185 24565 -165
rect 24585 -185 24600 -165
rect 24550 -215 24600 -185
rect 24550 -235 24565 -215
rect 24585 -235 24600 -215
rect 24550 -265 24600 -235
rect 24550 -285 24565 -265
rect 24585 -285 24600 -265
rect 24550 -315 24600 -285
rect 24550 -335 24565 -315
rect 24585 -335 24600 -315
rect 24550 -365 24600 -335
rect 24550 -385 24565 -365
rect 24585 -385 24600 -365
rect 24550 -415 24600 -385
rect 24550 -435 24565 -415
rect 24585 -435 24600 -415
rect 24550 -465 24600 -435
rect 24550 -485 24565 -465
rect 24585 -485 24600 -465
rect 24550 -515 24600 -485
rect 24550 -535 24565 -515
rect 24585 -535 24600 -515
rect 24550 -565 24600 -535
rect 24550 -585 24565 -565
rect 24585 -585 24600 -565
rect 24550 -615 24600 -585
rect 24550 -635 24565 -615
rect 24585 -635 24600 -615
rect 24550 -665 24600 -635
rect 24550 -685 24565 -665
rect 24585 -685 24600 -665
rect 24550 -715 24600 -685
rect 24550 -735 24565 -715
rect 24585 -735 24600 -715
rect 24550 -765 24600 -735
rect 24550 -785 24565 -765
rect 24585 -785 24600 -765
rect 24550 -800 24600 -785
rect 24700 -800 24750 -100
rect 24850 -800 24900 -100
rect 25000 -800 25050 -100
rect 25150 -800 25200 -100
rect 25300 -800 25350 -100
rect 25450 -800 25500 -100
rect 25600 -800 25650 -100
rect 25750 -115 25800 -100
rect 25750 -135 25765 -115
rect 25785 -135 25800 -115
rect 25750 -165 25800 -135
rect 25750 -185 25765 -165
rect 25785 -185 25800 -165
rect 25750 -215 25800 -185
rect 25750 -235 25765 -215
rect 25785 -235 25800 -215
rect 25750 -265 25800 -235
rect 25750 -285 25765 -265
rect 25785 -285 25800 -265
rect 25750 -315 25800 -285
rect 25750 -335 25765 -315
rect 25785 -335 25800 -315
rect 25750 -365 25800 -335
rect 25750 -385 25765 -365
rect 25785 -385 25800 -365
rect 25750 -415 25800 -385
rect 25750 -435 25765 -415
rect 25785 -435 25800 -415
rect 25750 -465 25800 -435
rect 25750 -485 25765 -465
rect 25785 -485 25800 -465
rect 25750 -515 25800 -485
rect 25750 -535 25765 -515
rect 25785 -535 25800 -515
rect 25750 -565 25800 -535
rect 25750 -585 25765 -565
rect 25785 -585 25800 -565
rect 25750 -615 25800 -585
rect 25750 -635 25765 -615
rect 25785 -635 25800 -615
rect 25750 -665 25800 -635
rect 25750 -685 25765 -665
rect 25785 -685 25800 -665
rect 25750 -715 25800 -685
rect 25750 -735 25765 -715
rect 25785 -735 25800 -715
rect 25750 -765 25800 -735
rect 25750 -785 25765 -765
rect 25785 -785 25800 -765
rect 25750 -800 25800 -785
rect 25900 -800 25950 -100
rect 26050 -800 26100 -100
rect 26200 -800 26250 -100
rect 26350 -800 26400 -100
rect 26500 -800 26550 -100
rect 26650 -115 26700 -100
rect 26650 -135 26665 -115
rect 26685 -135 26700 -115
rect 26650 -165 26700 -135
rect 26650 -185 26665 -165
rect 26685 -185 26700 -165
rect 26650 -215 26700 -185
rect 26650 -235 26665 -215
rect 26685 -235 26700 -215
rect 26650 -265 26700 -235
rect 26650 -285 26665 -265
rect 26685 -285 26700 -265
rect 26650 -315 26700 -285
rect 26650 -335 26665 -315
rect 26685 -335 26700 -315
rect 26650 -365 26700 -335
rect 26650 -385 26665 -365
rect 26685 -385 26700 -365
rect 26650 -415 26700 -385
rect 26650 -435 26665 -415
rect 26685 -435 26700 -415
rect 26650 -465 26700 -435
rect 26650 -485 26665 -465
rect 26685 -485 26700 -465
rect 26650 -515 26700 -485
rect 26650 -535 26665 -515
rect 26685 -535 26700 -515
rect 26650 -565 26700 -535
rect 26650 -585 26665 -565
rect 26685 -585 26700 -565
rect 26650 -615 26700 -585
rect 26650 -635 26665 -615
rect 26685 -635 26700 -615
rect 26650 -665 26700 -635
rect 26650 -685 26665 -665
rect 26685 -685 26700 -665
rect 26650 -715 26700 -685
rect 26650 -735 26665 -715
rect 26685 -735 26700 -715
rect 26650 -765 26700 -735
rect 26650 -785 26665 -765
rect 26685 -785 26700 -765
rect 26650 -800 26700 -785
rect 26800 -800 26850 -100
rect 26950 -800 27000 -100
rect 27100 -800 27150 -100
rect 27250 -800 27300 -100
rect 27400 -800 27450 -100
rect 27550 -115 27600 -100
rect 27550 -135 27565 -115
rect 27585 -135 27600 -115
rect 27550 -165 27600 -135
rect 27550 -185 27565 -165
rect 27585 -185 27600 -165
rect 27550 -215 27600 -185
rect 27550 -235 27565 -215
rect 27585 -235 27600 -215
rect 27550 -265 27600 -235
rect 27550 -285 27565 -265
rect 27585 -285 27600 -265
rect 27550 -315 27600 -285
rect 27550 -335 27565 -315
rect 27585 -335 27600 -315
rect 27550 -365 27600 -335
rect 27550 -385 27565 -365
rect 27585 -385 27600 -365
rect 27550 -415 27600 -385
rect 27550 -435 27565 -415
rect 27585 -435 27600 -415
rect 27550 -465 27600 -435
rect 27550 -485 27565 -465
rect 27585 -485 27600 -465
rect 27550 -515 27600 -485
rect 27550 -535 27565 -515
rect 27585 -535 27600 -515
rect 27550 -565 27600 -535
rect 27550 -585 27565 -565
rect 27585 -585 27600 -565
rect 27550 -615 27600 -585
rect 27550 -635 27565 -615
rect 27585 -635 27600 -615
rect 27550 -665 27600 -635
rect 27550 -685 27565 -665
rect 27585 -685 27600 -665
rect 27550 -715 27600 -685
rect 27550 -735 27565 -715
rect 27585 -735 27600 -715
rect 27550 -765 27600 -735
rect 27550 -785 27565 -765
rect 27585 -785 27600 -765
rect 27550 -800 27600 -785
rect 27700 -800 27750 -100
rect 27850 -800 27900 -100
rect 28000 -800 28050 -100
rect 28150 -800 28200 -100
rect 28300 -800 28350 -100
rect 28450 -800 28500 -100
rect 28600 -800 28650 -100
rect 28750 -115 28800 -100
rect 28750 -135 28765 -115
rect 28785 -135 28800 -115
rect 28750 -165 28800 -135
rect 28750 -185 28765 -165
rect 28785 -185 28800 -165
rect 28750 -215 28800 -185
rect 28750 -235 28765 -215
rect 28785 -235 28800 -215
rect 28750 -265 28800 -235
rect 28750 -285 28765 -265
rect 28785 -285 28800 -265
rect 28750 -315 28800 -285
rect 28750 -335 28765 -315
rect 28785 -335 28800 -315
rect 28750 -365 28800 -335
rect 28750 -385 28765 -365
rect 28785 -385 28800 -365
rect 28750 -415 28800 -385
rect 28750 -435 28765 -415
rect 28785 -435 28800 -415
rect 28750 -465 28800 -435
rect 28750 -485 28765 -465
rect 28785 -485 28800 -465
rect 28750 -515 28800 -485
rect 28750 -535 28765 -515
rect 28785 -535 28800 -515
rect 28750 -565 28800 -535
rect 28750 -585 28765 -565
rect 28785 -585 28800 -565
rect 28750 -615 28800 -585
rect 28750 -635 28765 -615
rect 28785 -635 28800 -615
rect 28750 -665 28800 -635
rect 28750 -685 28765 -665
rect 28785 -685 28800 -665
rect 28750 -715 28800 -685
rect 28750 -735 28765 -715
rect 28785 -735 28800 -715
rect 28750 -765 28800 -735
rect 28750 -785 28765 -765
rect 28785 -785 28800 -765
rect 28750 -800 28800 -785
rect -650 -965 -600 -950
rect -650 -985 -635 -965
rect -615 -985 -600 -965
rect -650 -1015 -600 -985
rect -650 -1035 -635 -1015
rect -615 -1035 -600 -1015
rect -650 -1065 -600 -1035
rect -650 -1085 -635 -1065
rect -615 -1085 -600 -1065
rect -650 -1115 -600 -1085
rect -650 -1135 -635 -1115
rect -615 -1135 -600 -1115
rect -650 -1165 -600 -1135
rect -650 -1185 -635 -1165
rect -615 -1185 -600 -1165
rect -650 -1215 -600 -1185
rect -650 -1235 -635 -1215
rect -615 -1235 -600 -1215
rect -650 -1265 -600 -1235
rect -650 -1285 -635 -1265
rect -615 -1285 -600 -1265
rect -650 -1315 -600 -1285
rect -650 -1335 -635 -1315
rect -615 -1335 -600 -1315
rect -650 -1365 -600 -1335
rect -650 -1385 -635 -1365
rect -615 -1385 -600 -1365
rect -650 -1415 -600 -1385
rect -650 -1435 -635 -1415
rect -615 -1435 -600 -1415
rect -650 -1465 -600 -1435
rect -650 -1485 -635 -1465
rect -615 -1485 -600 -1465
rect -650 -1515 -600 -1485
rect -650 -1535 -635 -1515
rect -615 -1535 -600 -1515
rect -650 -1565 -600 -1535
rect -650 -1585 -635 -1565
rect -615 -1585 -600 -1565
rect -650 -1615 -600 -1585
rect -650 -1635 -635 -1615
rect -615 -1635 -600 -1615
rect -650 -1650 -600 -1635
rect -500 -965 -450 -950
rect -500 -985 -485 -965
rect -465 -985 -450 -965
rect -500 -1015 -450 -985
rect -500 -1035 -485 -1015
rect -465 -1035 -450 -1015
rect -500 -1065 -450 -1035
rect -500 -1085 -485 -1065
rect -465 -1085 -450 -1065
rect -500 -1115 -450 -1085
rect -500 -1135 -485 -1115
rect -465 -1135 -450 -1115
rect -500 -1165 -450 -1135
rect -500 -1185 -485 -1165
rect -465 -1185 -450 -1165
rect -500 -1215 -450 -1185
rect -500 -1235 -485 -1215
rect -465 -1235 -450 -1215
rect -500 -1265 -450 -1235
rect -500 -1285 -485 -1265
rect -465 -1285 -450 -1265
rect -500 -1315 -450 -1285
rect -500 -1335 -485 -1315
rect -465 -1335 -450 -1315
rect -500 -1365 -450 -1335
rect -500 -1385 -485 -1365
rect -465 -1385 -450 -1365
rect -500 -1415 -450 -1385
rect -500 -1435 -485 -1415
rect -465 -1435 -450 -1415
rect -500 -1465 -450 -1435
rect -500 -1485 -485 -1465
rect -465 -1485 -450 -1465
rect -500 -1515 -450 -1485
rect -500 -1535 -485 -1515
rect -465 -1535 -450 -1515
rect -500 -1565 -450 -1535
rect -500 -1585 -485 -1565
rect -465 -1585 -450 -1565
rect -500 -1615 -450 -1585
rect -500 -1635 -485 -1615
rect -465 -1635 -450 -1615
rect -500 -1650 -450 -1635
rect -350 -965 -300 -950
rect -350 -985 -335 -965
rect -315 -985 -300 -965
rect -350 -1015 -300 -985
rect -350 -1035 -335 -1015
rect -315 -1035 -300 -1015
rect -350 -1065 -300 -1035
rect -350 -1085 -335 -1065
rect -315 -1085 -300 -1065
rect -350 -1115 -300 -1085
rect -350 -1135 -335 -1115
rect -315 -1135 -300 -1115
rect -350 -1165 -300 -1135
rect -350 -1185 -335 -1165
rect -315 -1185 -300 -1165
rect -350 -1215 -300 -1185
rect -350 -1235 -335 -1215
rect -315 -1235 -300 -1215
rect -350 -1265 -300 -1235
rect -350 -1285 -335 -1265
rect -315 -1285 -300 -1265
rect -350 -1315 -300 -1285
rect -350 -1335 -335 -1315
rect -315 -1335 -300 -1315
rect -350 -1365 -300 -1335
rect -350 -1385 -335 -1365
rect -315 -1385 -300 -1365
rect -350 -1415 -300 -1385
rect -350 -1435 -335 -1415
rect -315 -1435 -300 -1415
rect -350 -1465 -300 -1435
rect -350 -1485 -335 -1465
rect -315 -1485 -300 -1465
rect -350 -1515 -300 -1485
rect -350 -1535 -335 -1515
rect -315 -1535 -300 -1515
rect -350 -1565 -300 -1535
rect -350 -1585 -335 -1565
rect -315 -1585 -300 -1565
rect -350 -1615 -300 -1585
rect -350 -1635 -335 -1615
rect -315 -1635 -300 -1615
rect -350 -1650 -300 -1635
rect -200 -965 -150 -950
rect -200 -985 -185 -965
rect -165 -985 -150 -965
rect -200 -1015 -150 -985
rect -200 -1035 -185 -1015
rect -165 -1035 -150 -1015
rect -200 -1065 -150 -1035
rect -200 -1085 -185 -1065
rect -165 -1085 -150 -1065
rect -200 -1115 -150 -1085
rect -200 -1135 -185 -1115
rect -165 -1135 -150 -1115
rect -200 -1165 -150 -1135
rect -200 -1185 -185 -1165
rect -165 -1185 -150 -1165
rect -200 -1215 -150 -1185
rect -200 -1235 -185 -1215
rect -165 -1235 -150 -1215
rect -200 -1265 -150 -1235
rect -200 -1285 -185 -1265
rect -165 -1285 -150 -1265
rect -200 -1315 -150 -1285
rect -200 -1335 -185 -1315
rect -165 -1335 -150 -1315
rect -200 -1365 -150 -1335
rect -200 -1385 -185 -1365
rect -165 -1385 -150 -1365
rect -200 -1415 -150 -1385
rect -200 -1435 -185 -1415
rect -165 -1435 -150 -1415
rect -200 -1465 -150 -1435
rect -200 -1485 -185 -1465
rect -165 -1485 -150 -1465
rect -200 -1515 -150 -1485
rect -200 -1535 -185 -1515
rect -165 -1535 -150 -1515
rect -200 -1565 -150 -1535
rect -200 -1585 -185 -1565
rect -165 -1585 -150 -1565
rect -200 -1615 -150 -1585
rect -200 -1635 -185 -1615
rect -165 -1635 -150 -1615
rect -200 -1650 -150 -1635
rect -50 -965 0 -950
rect -50 -985 -35 -965
rect -15 -985 0 -965
rect -50 -1015 0 -985
rect -50 -1035 -35 -1015
rect -15 -1035 0 -1015
rect -50 -1065 0 -1035
rect -50 -1085 -35 -1065
rect -15 -1085 0 -1065
rect -50 -1115 0 -1085
rect -50 -1135 -35 -1115
rect -15 -1135 0 -1115
rect -50 -1165 0 -1135
rect -50 -1185 -35 -1165
rect -15 -1185 0 -1165
rect -50 -1215 0 -1185
rect -50 -1235 -35 -1215
rect -15 -1235 0 -1215
rect -50 -1265 0 -1235
rect -50 -1285 -35 -1265
rect -15 -1285 0 -1265
rect -50 -1315 0 -1285
rect -50 -1335 -35 -1315
rect -15 -1335 0 -1315
rect -50 -1365 0 -1335
rect -50 -1385 -35 -1365
rect -15 -1385 0 -1365
rect -50 -1415 0 -1385
rect -50 -1435 -35 -1415
rect -15 -1435 0 -1415
rect -50 -1465 0 -1435
rect -50 -1485 -35 -1465
rect -15 -1485 0 -1465
rect -50 -1515 0 -1485
rect -50 -1535 -35 -1515
rect -15 -1535 0 -1515
rect -50 -1565 0 -1535
rect -50 -1585 -35 -1565
rect -15 -1585 0 -1565
rect -50 -1615 0 -1585
rect -50 -1635 -35 -1615
rect -15 -1635 0 -1615
rect -50 -1650 0 -1635
rect 100 -1650 150 -950
rect 250 -1650 300 -950
rect 400 -1650 450 -950
rect 550 -1650 600 -950
rect 700 -1650 750 -950
rect 850 -1650 900 -950
rect 1000 -1650 1050 -950
rect 1150 -965 1200 -950
rect 1150 -985 1165 -965
rect 1185 -985 1200 -965
rect 1150 -1015 1200 -985
rect 1150 -1035 1165 -1015
rect 1185 -1035 1200 -1015
rect 1150 -1065 1200 -1035
rect 1150 -1085 1165 -1065
rect 1185 -1085 1200 -1065
rect 1150 -1115 1200 -1085
rect 1150 -1135 1165 -1115
rect 1185 -1135 1200 -1115
rect 1150 -1165 1200 -1135
rect 1150 -1185 1165 -1165
rect 1185 -1185 1200 -1165
rect 1150 -1215 1200 -1185
rect 1150 -1235 1165 -1215
rect 1185 -1235 1200 -1215
rect 1150 -1265 1200 -1235
rect 1150 -1285 1165 -1265
rect 1185 -1285 1200 -1265
rect 1150 -1315 1200 -1285
rect 1150 -1335 1165 -1315
rect 1185 -1335 1200 -1315
rect 1150 -1365 1200 -1335
rect 1150 -1385 1165 -1365
rect 1185 -1385 1200 -1365
rect 1150 -1415 1200 -1385
rect 1150 -1435 1165 -1415
rect 1185 -1435 1200 -1415
rect 1150 -1465 1200 -1435
rect 1150 -1485 1165 -1465
rect 1185 -1485 1200 -1465
rect 1150 -1515 1200 -1485
rect 1150 -1535 1165 -1515
rect 1185 -1535 1200 -1515
rect 1150 -1565 1200 -1535
rect 1150 -1585 1165 -1565
rect 1185 -1585 1200 -1565
rect 1150 -1615 1200 -1585
rect 1150 -1635 1165 -1615
rect 1185 -1635 1200 -1615
rect 1150 -1650 1200 -1635
rect 1300 -1650 1350 -950
rect 1450 -965 1500 -950
rect 1450 -985 1465 -965
rect 1485 -985 1500 -965
rect 1450 -1015 1500 -985
rect 1450 -1035 1465 -1015
rect 1485 -1035 1500 -1015
rect 1450 -1065 1500 -1035
rect 1450 -1085 1465 -1065
rect 1485 -1085 1500 -1065
rect 1450 -1115 1500 -1085
rect 1450 -1135 1465 -1115
rect 1485 -1135 1500 -1115
rect 1450 -1165 1500 -1135
rect 1450 -1185 1465 -1165
rect 1485 -1185 1500 -1165
rect 1450 -1215 1500 -1185
rect 1450 -1235 1465 -1215
rect 1485 -1235 1500 -1215
rect 1450 -1265 1500 -1235
rect 1450 -1285 1465 -1265
rect 1485 -1285 1500 -1265
rect 1450 -1315 1500 -1285
rect 1450 -1335 1465 -1315
rect 1485 -1335 1500 -1315
rect 1450 -1365 1500 -1335
rect 1450 -1385 1465 -1365
rect 1485 -1385 1500 -1365
rect 1450 -1415 1500 -1385
rect 1450 -1435 1465 -1415
rect 1485 -1435 1500 -1415
rect 1450 -1465 1500 -1435
rect 1450 -1485 1465 -1465
rect 1485 -1485 1500 -1465
rect 1450 -1515 1500 -1485
rect 1450 -1535 1465 -1515
rect 1485 -1535 1500 -1515
rect 1450 -1565 1500 -1535
rect 1450 -1585 1465 -1565
rect 1485 -1585 1500 -1565
rect 1450 -1615 1500 -1585
rect 1450 -1635 1465 -1615
rect 1485 -1635 1500 -1615
rect 1450 -1650 1500 -1635
rect 1600 -1650 1650 -950
rect 1750 -965 1800 -950
rect 1750 -985 1765 -965
rect 1785 -985 1800 -965
rect 1750 -1015 1800 -985
rect 1750 -1035 1765 -1015
rect 1785 -1035 1800 -1015
rect 1750 -1065 1800 -1035
rect 1750 -1085 1765 -1065
rect 1785 -1085 1800 -1065
rect 1750 -1115 1800 -1085
rect 1750 -1135 1765 -1115
rect 1785 -1135 1800 -1115
rect 1750 -1165 1800 -1135
rect 1750 -1185 1765 -1165
rect 1785 -1185 1800 -1165
rect 1750 -1215 1800 -1185
rect 1750 -1235 1765 -1215
rect 1785 -1235 1800 -1215
rect 1750 -1265 1800 -1235
rect 1750 -1285 1765 -1265
rect 1785 -1285 1800 -1265
rect 1750 -1315 1800 -1285
rect 1750 -1335 1765 -1315
rect 1785 -1335 1800 -1315
rect 1750 -1365 1800 -1335
rect 1750 -1385 1765 -1365
rect 1785 -1385 1800 -1365
rect 1750 -1415 1800 -1385
rect 1750 -1435 1765 -1415
rect 1785 -1435 1800 -1415
rect 1750 -1465 1800 -1435
rect 1750 -1485 1765 -1465
rect 1785 -1485 1800 -1465
rect 1750 -1515 1800 -1485
rect 1750 -1535 1765 -1515
rect 1785 -1535 1800 -1515
rect 1750 -1565 1800 -1535
rect 1750 -1585 1765 -1565
rect 1785 -1585 1800 -1565
rect 1750 -1615 1800 -1585
rect 1750 -1635 1765 -1615
rect 1785 -1635 1800 -1615
rect 1750 -1650 1800 -1635
rect 1900 -1650 1950 -950
rect 2050 -965 2100 -950
rect 2050 -985 2065 -965
rect 2085 -985 2100 -965
rect 2050 -1015 2100 -985
rect 2050 -1035 2065 -1015
rect 2085 -1035 2100 -1015
rect 2050 -1065 2100 -1035
rect 2050 -1085 2065 -1065
rect 2085 -1085 2100 -1065
rect 2050 -1115 2100 -1085
rect 2050 -1135 2065 -1115
rect 2085 -1135 2100 -1115
rect 2050 -1165 2100 -1135
rect 2050 -1185 2065 -1165
rect 2085 -1185 2100 -1165
rect 2050 -1215 2100 -1185
rect 2050 -1235 2065 -1215
rect 2085 -1235 2100 -1215
rect 2050 -1265 2100 -1235
rect 2050 -1285 2065 -1265
rect 2085 -1285 2100 -1265
rect 2050 -1315 2100 -1285
rect 2050 -1335 2065 -1315
rect 2085 -1335 2100 -1315
rect 2050 -1365 2100 -1335
rect 2050 -1385 2065 -1365
rect 2085 -1385 2100 -1365
rect 2050 -1415 2100 -1385
rect 2050 -1435 2065 -1415
rect 2085 -1435 2100 -1415
rect 2050 -1465 2100 -1435
rect 2050 -1485 2065 -1465
rect 2085 -1485 2100 -1465
rect 2050 -1515 2100 -1485
rect 2050 -1535 2065 -1515
rect 2085 -1535 2100 -1515
rect 2050 -1565 2100 -1535
rect 2050 -1585 2065 -1565
rect 2085 -1585 2100 -1565
rect 2050 -1615 2100 -1585
rect 2050 -1635 2065 -1615
rect 2085 -1635 2100 -1615
rect 2050 -1650 2100 -1635
rect 2200 -1650 2250 -950
rect 2350 -965 2400 -950
rect 2350 -985 2365 -965
rect 2385 -985 2400 -965
rect 2350 -1015 2400 -985
rect 2350 -1035 2365 -1015
rect 2385 -1035 2400 -1015
rect 2350 -1065 2400 -1035
rect 2350 -1085 2365 -1065
rect 2385 -1085 2400 -1065
rect 2350 -1115 2400 -1085
rect 2350 -1135 2365 -1115
rect 2385 -1135 2400 -1115
rect 2350 -1165 2400 -1135
rect 2350 -1185 2365 -1165
rect 2385 -1185 2400 -1165
rect 2350 -1215 2400 -1185
rect 2350 -1235 2365 -1215
rect 2385 -1235 2400 -1215
rect 2350 -1265 2400 -1235
rect 2350 -1285 2365 -1265
rect 2385 -1285 2400 -1265
rect 2350 -1315 2400 -1285
rect 2350 -1335 2365 -1315
rect 2385 -1335 2400 -1315
rect 2350 -1365 2400 -1335
rect 2350 -1385 2365 -1365
rect 2385 -1385 2400 -1365
rect 2350 -1415 2400 -1385
rect 2350 -1435 2365 -1415
rect 2385 -1435 2400 -1415
rect 2350 -1465 2400 -1435
rect 2350 -1485 2365 -1465
rect 2385 -1485 2400 -1465
rect 2350 -1515 2400 -1485
rect 2350 -1535 2365 -1515
rect 2385 -1535 2400 -1515
rect 2350 -1565 2400 -1535
rect 2350 -1585 2365 -1565
rect 2385 -1585 2400 -1565
rect 2350 -1615 2400 -1585
rect 2350 -1635 2365 -1615
rect 2385 -1635 2400 -1615
rect 2350 -1650 2400 -1635
rect 2500 -1650 2550 -950
rect 2650 -965 2700 -950
rect 2650 -985 2665 -965
rect 2685 -985 2700 -965
rect 2650 -1015 2700 -985
rect 2650 -1035 2665 -1015
rect 2685 -1035 2700 -1015
rect 2650 -1065 2700 -1035
rect 2650 -1085 2665 -1065
rect 2685 -1085 2700 -1065
rect 2650 -1115 2700 -1085
rect 2650 -1135 2665 -1115
rect 2685 -1135 2700 -1115
rect 2650 -1165 2700 -1135
rect 2650 -1185 2665 -1165
rect 2685 -1185 2700 -1165
rect 2650 -1215 2700 -1185
rect 2650 -1235 2665 -1215
rect 2685 -1235 2700 -1215
rect 2650 -1265 2700 -1235
rect 2650 -1285 2665 -1265
rect 2685 -1285 2700 -1265
rect 2650 -1315 2700 -1285
rect 2650 -1335 2665 -1315
rect 2685 -1335 2700 -1315
rect 2650 -1365 2700 -1335
rect 2650 -1385 2665 -1365
rect 2685 -1385 2700 -1365
rect 2650 -1415 2700 -1385
rect 2650 -1435 2665 -1415
rect 2685 -1435 2700 -1415
rect 2650 -1465 2700 -1435
rect 2650 -1485 2665 -1465
rect 2685 -1485 2700 -1465
rect 2650 -1515 2700 -1485
rect 2650 -1535 2665 -1515
rect 2685 -1535 2700 -1515
rect 2650 -1565 2700 -1535
rect 2650 -1585 2665 -1565
rect 2685 -1585 2700 -1565
rect 2650 -1615 2700 -1585
rect 2650 -1635 2665 -1615
rect 2685 -1635 2700 -1615
rect 2650 -1650 2700 -1635
rect 2800 -1650 2850 -950
rect 2950 -965 3000 -950
rect 2950 -985 2965 -965
rect 2985 -985 3000 -965
rect 2950 -1015 3000 -985
rect 2950 -1035 2965 -1015
rect 2985 -1035 3000 -1015
rect 2950 -1065 3000 -1035
rect 2950 -1085 2965 -1065
rect 2985 -1085 3000 -1065
rect 2950 -1115 3000 -1085
rect 2950 -1135 2965 -1115
rect 2985 -1135 3000 -1115
rect 2950 -1165 3000 -1135
rect 2950 -1185 2965 -1165
rect 2985 -1185 3000 -1165
rect 2950 -1215 3000 -1185
rect 2950 -1235 2965 -1215
rect 2985 -1235 3000 -1215
rect 2950 -1265 3000 -1235
rect 2950 -1285 2965 -1265
rect 2985 -1285 3000 -1265
rect 2950 -1315 3000 -1285
rect 2950 -1335 2965 -1315
rect 2985 -1335 3000 -1315
rect 2950 -1365 3000 -1335
rect 2950 -1385 2965 -1365
rect 2985 -1385 3000 -1365
rect 2950 -1415 3000 -1385
rect 2950 -1435 2965 -1415
rect 2985 -1435 3000 -1415
rect 2950 -1465 3000 -1435
rect 2950 -1485 2965 -1465
rect 2985 -1485 3000 -1465
rect 2950 -1515 3000 -1485
rect 2950 -1535 2965 -1515
rect 2985 -1535 3000 -1515
rect 2950 -1565 3000 -1535
rect 2950 -1585 2965 -1565
rect 2985 -1585 3000 -1565
rect 2950 -1615 3000 -1585
rect 2950 -1635 2965 -1615
rect 2985 -1635 3000 -1615
rect 2950 -1650 3000 -1635
rect 3100 -1650 3150 -950
rect 3250 -965 3300 -950
rect 3250 -985 3265 -965
rect 3285 -985 3300 -965
rect 3250 -1015 3300 -985
rect 3250 -1035 3265 -1015
rect 3285 -1035 3300 -1015
rect 3250 -1065 3300 -1035
rect 3250 -1085 3265 -1065
rect 3285 -1085 3300 -1065
rect 3250 -1115 3300 -1085
rect 3250 -1135 3265 -1115
rect 3285 -1135 3300 -1115
rect 3250 -1165 3300 -1135
rect 3250 -1185 3265 -1165
rect 3285 -1185 3300 -1165
rect 3250 -1215 3300 -1185
rect 3250 -1235 3265 -1215
rect 3285 -1235 3300 -1215
rect 3250 -1265 3300 -1235
rect 3250 -1285 3265 -1265
rect 3285 -1285 3300 -1265
rect 3250 -1315 3300 -1285
rect 3250 -1335 3265 -1315
rect 3285 -1335 3300 -1315
rect 3250 -1365 3300 -1335
rect 3250 -1385 3265 -1365
rect 3285 -1385 3300 -1365
rect 3250 -1415 3300 -1385
rect 3250 -1435 3265 -1415
rect 3285 -1435 3300 -1415
rect 3250 -1465 3300 -1435
rect 3250 -1485 3265 -1465
rect 3285 -1485 3300 -1465
rect 3250 -1515 3300 -1485
rect 3250 -1535 3265 -1515
rect 3285 -1535 3300 -1515
rect 3250 -1565 3300 -1535
rect 3250 -1585 3265 -1565
rect 3285 -1585 3300 -1565
rect 3250 -1615 3300 -1585
rect 3250 -1635 3265 -1615
rect 3285 -1635 3300 -1615
rect 3250 -1650 3300 -1635
rect 3400 -1650 3450 -950
rect 3550 -965 3600 -950
rect 3550 -985 3565 -965
rect 3585 -985 3600 -965
rect 3550 -1015 3600 -985
rect 3550 -1035 3565 -1015
rect 3585 -1035 3600 -1015
rect 3550 -1065 3600 -1035
rect 3550 -1085 3565 -1065
rect 3585 -1085 3600 -1065
rect 3550 -1115 3600 -1085
rect 3550 -1135 3565 -1115
rect 3585 -1135 3600 -1115
rect 3550 -1165 3600 -1135
rect 3550 -1185 3565 -1165
rect 3585 -1185 3600 -1165
rect 3550 -1215 3600 -1185
rect 3550 -1235 3565 -1215
rect 3585 -1235 3600 -1215
rect 3550 -1265 3600 -1235
rect 3550 -1285 3565 -1265
rect 3585 -1285 3600 -1265
rect 3550 -1315 3600 -1285
rect 3550 -1335 3565 -1315
rect 3585 -1335 3600 -1315
rect 3550 -1365 3600 -1335
rect 3550 -1385 3565 -1365
rect 3585 -1385 3600 -1365
rect 3550 -1415 3600 -1385
rect 3550 -1435 3565 -1415
rect 3585 -1435 3600 -1415
rect 3550 -1465 3600 -1435
rect 3550 -1485 3565 -1465
rect 3585 -1485 3600 -1465
rect 3550 -1515 3600 -1485
rect 3550 -1535 3565 -1515
rect 3585 -1535 3600 -1515
rect 3550 -1565 3600 -1535
rect 3550 -1585 3565 -1565
rect 3585 -1585 3600 -1565
rect 3550 -1615 3600 -1585
rect 3550 -1635 3565 -1615
rect 3585 -1635 3600 -1615
rect 3550 -1650 3600 -1635
rect 3700 -965 3750 -950
rect 3700 -985 3715 -965
rect 3735 -985 3750 -965
rect 3700 -1015 3750 -985
rect 3700 -1035 3715 -1015
rect 3735 -1035 3750 -1015
rect 3700 -1065 3750 -1035
rect 3700 -1085 3715 -1065
rect 3735 -1085 3750 -1065
rect 3700 -1115 3750 -1085
rect 3700 -1135 3715 -1115
rect 3735 -1135 3750 -1115
rect 3700 -1165 3750 -1135
rect 3700 -1185 3715 -1165
rect 3735 -1185 3750 -1165
rect 3700 -1215 3750 -1185
rect 3700 -1235 3715 -1215
rect 3735 -1235 3750 -1215
rect 3700 -1265 3750 -1235
rect 3700 -1285 3715 -1265
rect 3735 -1285 3750 -1265
rect 3700 -1315 3750 -1285
rect 3700 -1335 3715 -1315
rect 3735 -1335 3750 -1315
rect 3700 -1365 3750 -1335
rect 3700 -1385 3715 -1365
rect 3735 -1385 3750 -1365
rect 3700 -1415 3750 -1385
rect 3700 -1435 3715 -1415
rect 3735 -1435 3750 -1415
rect 3700 -1465 3750 -1435
rect 3700 -1485 3715 -1465
rect 3735 -1485 3750 -1465
rect 3700 -1515 3750 -1485
rect 3700 -1535 3715 -1515
rect 3735 -1535 3750 -1515
rect 3700 -1565 3750 -1535
rect 3700 -1585 3715 -1565
rect 3735 -1585 3750 -1565
rect 3700 -1615 3750 -1585
rect 3700 -1635 3715 -1615
rect 3735 -1635 3750 -1615
rect 3700 -1650 3750 -1635
rect 3850 -965 3900 -950
rect 3850 -985 3865 -965
rect 3885 -985 3900 -965
rect 3850 -1015 3900 -985
rect 3850 -1035 3865 -1015
rect 3885 -1035 3900 -1015
rect 3850 -1065 3900 -1035
rect 3850 -1085 3865 -1065
rect 3885 -1085 3900 -1065
rect 3850 -1115 3900 -1085
rect 3850 -1135 3865 -1115
rect 3885 -1135 3900 -1115
rect 3850 -1165 3900 -1135
rect 3850 -1185 3865 -1165
rect 3885 -1185 3900 -1165
rect 3850 -1215 3900 -1185
rect 3850 -1235 3865 -1215
rect 3885 -1235 3900 -1215
rect 3850 -1265 3900 -1235
rect 3850 -1285 3865 -1265
rect 3885 -1285 3900 -1265
rect 3850 -1315 3900 -1285
rect 3850 -1335 3865 -1315
rect 3885 -1335 3900 -1315
rect 3850 -1365 3900 -1335
rect 3850 -1385 3865 -1365
rect 3885 -1385 3900 -1365
rect 3850 -1415 3900 -1385
rect 3850 -1435 3865 -1415
rect 3885 -1435 3900 -1415
rect 3850 -1465 3900 -1435
rect 3850 -1485 3865 -1465
rect 3885 -1485 3900 -1465
rect 3850 -1515 3900 -1485
rect 3850 -1535 3865 -1515
rect 3885 -1535 3900 -1515
rect 3850 -1565 3900 -1535
rect 3850 -1585 3865 -1565
rect 3885 -1585 3900 -1565
rect 3850 -1615 3900 -1585
rect 3850 -1635 3865 -1615
rect 3885 -1635 3900 -1615
rect 3850 -1650 3900 -1635
rect 4000 -965 4050 -950
rect 4000 -985 4015 -965
rect 4035 -985 4050 -965
rect 4000 -1015 4050 -985
rect 4000 -1035 4015 -1015
rect 4035 -1035 4050 -1015
rect 4000 -1065 4050 -1035
rect 4000 -1085 4015 -1065
rect 4035 -1085 4050 -1065
rect 4000 -1115 4050 -1085
rect 4000 -1135 4015 -1115
rect 4035 -1135 4050 -1115
rect 4000 -1165 4050 -1135
rect 4000 -1185 4015 -1165
rect 4035 -1185 4050 -1165
rect 4000 -1215 4050 -1185
rect 4000 -1235 4015 -1215
rect 4035 -1235 4050 -1215
rect 4000 -1265 4050 -1235
rect 4000 -1285 4015 -1265
rect 4035 -1285 4050 -1265
rect 4000 -1315 4050 -1285
rect 4000 -1335 4015 -1315
rect 4035 -1335 4050 -1315
rect 4000 -1365 4050 -1335
rect 4000 -1385 4015 -1365
rect 4035 -1385 4050 -1365
rect 4000 -1415 4050 -1385
rect 4000 -1435 4015 -1415
rect 4035 -1435 4050 -1415
rect 4000 -1465 4050 -1435
rect 4000 -1485 4015 -1465
rect 4035 -1485 4050 -1465
rect 4000 -1515 4050 -1485
rect 4000 -1535 4015 -1515
rect 4035 -1535 4050 -1515
rect 4000 -1565 4050 -1535
rect 4000 -1585 4015 -1565
rect 4035 -1585 4050 -1565
rect 4000 -1615 4050 -1585
rect 4000 -1635 4015 -1615
rect 4035 -1635 4050 -1615
rect 4000 -1650 4050 -1635
rect 4150 -965 4200 -950
rect 4150 -985 4165 -965
rect 4185 -985 4200 -965
rect 4150 -1015 4200 -985
rect 4150 -1035 4165 -1015
rect 4185 -1035 4200 -1015
rect 4150 -1065 4200 -1035
rect 4150 -1085 4165 -1065
rect 4185 -1085 4200 -1065
rect 4150 -1115 4200 -1085
rect 4150 -1135 4165 -1115
rect 4185 -1135 4200 -1115
rect 4150 -1165 4200 -1135
rect 4150 -1185 4165 -1165
rect 4185 -1185 4200 -1165
rect 4150 -1215 4200 -1185
rect 4150 -1235 4165 -1215
rect 4185 -1235 4200 -1215
rect 4150 -1265 4200 -1235
rect 4150 -1285 4165 -1265
rect 4185 -1285 4200 -1265
rect 4150 -1315 4200 -1285
rect 4150 -1335 4165 -1315
rect 4185 -1335 4200 -1315
rect 4150 -1365 4200 -1335
rect 4150 -1385 4165 -1365
rect 4185 -1385 4200 -1365
rect 4150 -1415 4200 -1385
rect 4150 -1435 4165 -1415
rect 4185 -1435 4200 -1415
rect 4150 -1465 4200 -1435
rect 4150 -1485 4165 -1465
rect 4185 -1485 4200 -1465
rect 4150 -1515 4200 -1485
rect 4150 -1535 4165 -1515
rect 4185 -1535 4200 -1515
rect 4150 -1565 4200 -1535
rect 4150 -1585 4165 -1565
rect 4185 -1585 4200 -1565
rect 4150 -1615 4200 -1585
rect 4150 -1635 4165 -1615
rect 4185 -1635 4200 -1615
rect 4150 -1650 4200 -1635
rect 4300 -965 4350 -950
rect 4300 -985 4315 -965
rect 4335 -985 4350 -965
rect 4300 -1015 4350 -985
rect 4300 -1035 4315 -1015
rect 4335 -1035 4350 -1015
rect 4300 -1065 4350 -1035
rect 4300 -1085 4315 -1065
rect 4335 -1085 4350 -1065
rect 4300 -1115 4350 -1085
rect 4300 -1135 4315 -1115
rect 4335 -1135 4350 -1115
rect 4300 -1165 4350 -1135
rect 4300 -1185 4315 -1165
rect 4335 -1185 4350 -1165
rect 4300 -1215 4350 -1185
rect 4300 -1235 4315 -1215
rect 4335 -1235 4350 -1215
rect 4300 -1265 4350 -1235
rect 4300 -1285 4315 -1265
rect 4335 -1285 4350 -1265
rect 4300 -1315 4350 -1285
rect 4300 -1335 4315 -1315
rect 4335 -1335 4350 -1315
rect 4300 -1365 4350 -1335
rect 4300 -1385 4315 -1365
rect 4335 -1385 4350 -1365
rect 4300 -1415 4350 -1385
rect 4300 -1435 4315 -1415
rect 4335 -1435 4350 -1415
rect 4300 -1465 4350 -1435
rect 4300 -1485 4315 -1465
rect 4335 -1485 4350 -1465
rect 4300 -1515 4350 -1485
rect 4300 -1535 4315 -1515
rect 4335 -1535 4350 -1515
rect 4300 -1565 4350 -1535
rect 4300 -1585 4315 -1565
rect 4335 -1585 4350 -1565
rect 4300 -1615 4350 -1585
rect 4300 -1635 4315 -1615
rect 4335 -1635 4350 -1615
rect 4300 -1650 4350 -1635
rect 4450 -965 4500 -950
rect 4450 -985 4465 -965
rect 4485 -985 4500 -965
rect 4450 -1015 4500 -985
rect 4450 -1035 4465 -1015
rect 4485 -1035 4500 -1015
rect 4450 -1065 4500 -1035
rect 4450 -1085 4465 -1065
rect 4485 -1085 4500 -1065
rect 4450 -1115 4500 -1085
rect 4450 -1135 4465 -1115
rect 4485 -1135 4500 -1115
rect 4450 -1165 4500 -1135
rect 4450 -1185 4465 -1165
rect 4485 -1185 4500 -1165
rect 4450 -1215 4500 -1185
rect 4450 -1235 4465 -1215
rect 4485 -1235 4500 -1215
rect 4450 -1265 4500 -1235
rect 4450 -1285 4465 -1265
rect 4485 -1285 4500 -1265
rect 4450 -1315 4500 -1285
rect 4450 -1335 4465 -1315
rect 4485 -1335 4500 -1315
rect 4450 -1365 4500 -1335
rect 4450 -1385 4465 -1365
rect 4485 -1385 4500 -1365
rect 4450 -1415 4500 -1385
rect 4450 -1435 4465 -1415
rect 4485 -1435 4500 -1415
rect 4450 -1465 4500 -1435
rect 4450 -1485 4465 -1465
rect 4485 -1485 4500 -1465
rect 4450 -1515 4500 -1485
rect 4450 -1535 4465 -1515
rect 4485 -1535 4500 -1515
rect 4450 -1565 4500 -1535
rect 4450 -1585 4465 -1565
rect 4485 -1585 4500 -1565
rect 4450 -1615 4500 -1585
rect 4450 -1635 4465 -1615
rect 4485 -1635 4500 -1615
rect 4450 -1650 4500 -1635
rect 4600 -965 4650 -950
rect 4600 -985 4615 -965
rect 4635 -985 4650 -965
rect 4600 -1015 4650 -985
rect 4600 -1035 4615 -1015
rect 4635 -1035 4650 -1015
rect 4600 -1065 4650 -1035
rect 4600 -1085 4615 -1065
rect 4635 -1085 4650 -1065
rect 4600 -1115 4650 -1085
rect 4600 -1135 4615 -1115
rect 4635 -1135 4650 -1115
rect 4600 -1165 4650 -1135
rect 4600 -1185 4615 -1165
rect 4635 -1185 4650 -1165
rect 4600 -1215 4650 -1185
rect 4600 -1235 4615 -1215
rect 4635 -1235 4650 -1215
rect 4600 -1265 4650 -1235
rect 4600 -1285 4615 -1265
rect 4635 -1285 4650 -1265
rect 4600 -1315 4650 -1285
rect 4600 -1335 4615 -1315
rect 4635 -1335 4650 -1315
rect 4600 -1365 4650 -1335
rect 4600 -1385 4615 -1365
rect 4635 -1385 4650 -1365
rect 4600 -1415 4650 -1385
rect 4600 -1435 4615 -1415
rect 4635 -1435 4650 -1415
rect 4600 -1465 4650 -1435
rect 4600 -1485 4615 -1465
rect 4635 -1485 4650 -1465
rect 4600 -1515 4650 -1485
rect 4600 -1535 4615 -1515
rect 4635 -1535 4650 -1515
rect 4600 -1565 4650 -1535
rect 4600 -1585 4615 -1565
rect 4635 -1585 4650 -1565
rect 4600 -1615 4650 -1585
rect 4600 -1635 4615 -1615
rect 4635 -1635 4650 -1615
rect 4600 -1650 4650 -1635
rect 4750 -965 4800 -950
rect 4750 -985 4765 -965
rect 4785 -985 4800 -965
rect 4750 -1015 4800 -985
rect 4750 -1035 4765 -1015
rect 4785 -1035 4800 -1015
rect 4750 -1065 4800 -1035
rect 4750 -1085 4765 -1065
rect 4785 -1085 4800 -1065
rect 4750 -1115 4800 -1085
rect 4750 -1135 4765 -1115
rect 4785 -1135 4800 -1115
rect 4750 -1165 4800 -1135
rect 4750 -1185 4765 -1165
rect 4785 -1185 4800 -1165
rect 4750 -1215 4800 -1185
rect 4750 -1235 4765 -1215
rect 4785 -1235 4800 -1215
rect 4750 -1265 4800 -1235
rect 4750 -1285 4765 -1265
rect 4785 -1285 4800 -1265
rect 4750 -1315 4800 -1285
rect 4750 -1335 4765 -1315
rect 4785 -1335 4800 -1315
rect 4750 -1365 4800 -1335
rect 4750 -1385 4765 -1365
rect 4785 -1385 4800 -1365
rect 4750 -1415 4800 -1385
rect 4750 -1435 4765 -1415
rect 4785 -1435 4800 -1415
rect 4750 -1465 4800 -1435
rect 4750 -1485 4765 -1465
rect 4785 -1485 4800 -1465
rect 4750 -1515 4800 -1485
rect 4750 -1535 4765 -1515
rect 4785 -1535 4800 -1515
rect 4750 -1565 4800 -1535
rect 4750 -1585 4765 -1565
rect 4785 -1585 4800 -1565
rect 4750 -1615 4800 -1585
rect 4750 -1635 4765 -1615
rect 4785 -1635 4800 -1615
rect 4750 -1650 4800 -1635
rect 4900 -1650 4950 -950
rect 5050 -965 5100 -950
rect 5050 -985 5065 -965
rect 5085 -985 5100 -965
rect 5050 -1015 5100 -985
rect 5050 -1035 5065 -1015
rect 5085 -1035 5100 -1015
rect 5050 -1065 5100 -1035
rect 5050 -1085 5065 -1065
rect 5085 -1085 5100 -1065
rect 5050 -1115 5100 -1085
rect 5050 -1135 5065 -1115
rect 5085 -1135 5100 -1115
rect 5050 -1165 5100 -1135
rect 5050 -1185 5065 -1165
rect 5085 -1185 5100 -1165
rect 5050 -1215 5100 -1185
rect 5050 -1235 5065 -1215
rect 5085 -1235 5100 -1215
rect 5050 -1265 5100 -1235
rect 5050 -1285 5065 -1265
rect 5085 -1285 5100 -1265
rect 5050 -1315 5100 -1285
rect 5050 -1335 5065 -1315
rect 5085 -1335 5100 -1315
rect 5050 -1365 5100 -1335
rect 5050 -1385 5065 -1365
rect 5085 -1385 5100 -1365
rect 5050 -1415 5100 -1385
rect 5050 -1435 5065 -1415
rect 5085 -1435 5100 -1415
rect 5050 -1465 5100 -1435
rect 5050 -1485 5065 -1465
rect 5085 -1485 5100 -1465
rect 5050 -1515 5100 -1485
rect 5050 -1535 5065 -1515
rect 5085 -1535 5100 -1515
rect 5050 -1565 5100 -1535
rect 5050 -1585 5065 -1565
rect 5085 -1585 5100 -1565
rect 5050 -1615 5100 -1585
rect 5050 -1635 5065 -1615
rect 5085 -1635 5100 -1615
rect 5050 -1650 5100 -1635
rect 5200 -1650 5250 -950
rect 5350 -965 5400 -950
rect 5350 -985 5365 -965
rect 5385 -985 5400 -965
rect 5350 -1015 5400 -985
rect 5350 -1035 5365 -1015
rect 5385 -1035 5400 -1015
rect 5350 -1065 5400 -1035
rect 5350 -1085 5365 -1065
rect 5385 -1085 5400 -1065
rect 5350 -1115 5400 -1085
rect 5350 -1135 5365 -1115
rect 5385 -1135 5400 -1115
rect 5350 -1165 5400 -1135
rect 5350 -1185 5365 -1165
rect 5385 -1185 5400 -1165
rect 5350 -1215 5400 -1185
rect 5350 -1235 5365 -1215
rect 5385 -1235 5400 -1215
rect 5350 -1265 5400 -1235
rect 5350 -1285 5365 -1265
rect 5385 -1285 5400 -1265
rect 5350 -1315 5400 -1285
rect 5350 -1335 5365 -1315
rect 5385 -1335 5400 -1315
rect 5350 -1365 5400 -1335
rect 5350 -1385 5365 -1365
rect 5385 -1385 5400 -1365
rect 5350 -1415 5400 -1385
rect 5350 -1435 5365 -1415
rect 5385 -1435 5400 -1415
rect 5350 -1465 5400 -1435
rect 5350 -1485 5365 -1465
rect 5385 -1485 5400 -1465
rect 5350 -1515 5400 -1485
rect 5350 -1535 5365 -1515
rect 5385 -1535 5400 -1515
rect 5350 -1565 5400 -1535
rect 5350 -1585 5365 -1565
rect 5385 -1585 5400 -1565
rect 5350 -1615 5400 -1585
rect 5350 -1635 5365 -1615
rect 5385 -1635 5400 -1615
rect 5350 -1650 5400 -1635
rect 5500 -1650 5550 -950
rect 5650 -965 5700 -950
rect 5650 -985 5665 -965
rect 5685 -985 5700 -965
rect 5650 -1015 5700 -985
rect 5650 -1035 5665 -1015
rect 5685 -1035 5700 -1015
rect 5650 -1065 5700 -1035
rect 5650 -1085 5665 -1065
rect 5685 -1085 5700 -1065
rect 5650 -1115 5700 -1085
rect 5650 -1135 5665 -1115
rect 5685 -1135 5700 -1115
rect 5650 -1165 5700 -1135
rect 5650 -1185 5665 -1165
rect 5685 -1185 5700 -1165
rect 5650 -1215 5700 -1185
rect 5650 -1235 5665 -1215
rect 5685 -1235 5700 -1215
rect 5650 -1265 5700 -1235
rect 5650 -1285 5665 -1265
rect 5685 -1285 5700 -1265
rect 5650 -1315 5700 -1285
rect 5650 -1335 5665 -1315
rect 5685 -1335 5700 -1315
rect 5650 -1365 5700 -1335
rect 5650 -1385 5665 -1365
rect 5685 -1385 5700 -1365
rect 5650 -1415 5700 -1385
rect 5650 -1435 5665 -1415
rect 5685 -1435 5700 -1415
rect 5650 -1465 5700 -1435
rect 5650 -1485 5665 -1465
rect 5685 -1485 5700 -1465
rect 5650 -1515 5700 -1485
rect 5650 -1535 5665 -1515
rect 5685 -1535 5700 -1515
rect 5650 -1565 5700 -1535
rect 5650 -1585 5665 -1565
rect 5685 -1585 5700 -1565
rect 5650 -1615 5700 -1585
rect 5650 -1635 5665 -1615
rect 5685 -1635 5700 -1615
rect 5650 -1650 5700 -1635
rect 5800 -1650 5850 -950
rect 5950 -965 6000 -950
rect 5950 -985 5965 -965
rect 5985 -985 6000 -965
rect 5950 -1015 6000 -985
rect 5950 -1035 5965 -1015
rect 5985 -1035 6000 -1015
rect 5950 -1065 6000 -1035
rect 5950 -1085 5965 -1065
rect 5985 -1085 6000 -1065
rect 5950 -1115 6000 -1085
rect 5950 -1135 5965 -1115
rect 5985 -1135 6000 -1115
rect 5950 -1165 6000 -1135
rect 5950 -1185 5965 -1165
rect 5985 -1185 6000 -1165
rect 5950 -1215 6000 -1185
rect 5950 -1235 5965 -1215
rect 5985 -1235 6000 -1215
rect 5950 -1265 6000 -1235
rect 5950 -1285 5965 -1265
rect 5985 -1285 6000 -1265
rect 5950 -1315 6000 -1285
rect 5950 -1335 5965 -1315
rect 5985 -1335 6000 -1315
rect 5950 -1365 6000 -1335
rect 5950 -1385 5965 -1365
rect 5985 -1385 6000 -1365
rect 5950 -1415 6000 -1385
rect 5950 -1435 5965 -1415
rect 5985 -1435 6000 -1415
rect 5950 -1465 6000 -1435
rect 5950 -1485 5965 -1465
rect 5985 -1485 6000 -1465
rect 5950 -1515 6000 -1485
rect 5950 -1535 5965 -1515
rect 5985 -1535 6000 -1515
rect 5950 -1565 6000 -1535
rect 5950 -1585 5965 -1565
rect 5985 -1585 6000 -1565
rect 5950 -1615 6000 -1585
rect 5950 -1635 5965 -1615
rect 5985 -1635 6000 -1615
rect 5950 -1650 6000 -1635
rect 6100 -1650 6150 -950
rect 6250 -965 6300 -950
rect 6250 -985 6265 -965
rect 6285 -985 6300 -965
rect 6250 -1015 6300 -985
rect 6250 -1035 6265 -1015
rect 6285 -1035 6300 -1015
rect 6250 -1065 6300 -1035
rect 6250 -1085 6265 -1065
rect 6285 -1085 6300 -1065
rect 6250 -1115 6300 -1085
rect 6250 -1135 6265 -1115
rect 6285 -1135 6300 -1115
rect 6250 -1165 6300 -1135
rect 6250 -1185 6265 -1165
rect 6285 -1185 6300 -1165
rect 6250 -1215 6300 -1185
rect 6250 -1235 6265 -1215
rect 6285 -1235 6300 -1215
rect 6250 -1265 6300 -1235
rect 6250 -1285 6265 -1265
rect 6285 -1285 6300 -1265
rect 6250 -1315 6300 -1285
rect 6250 -1335 6265 -1315
rect 6285 -1335 6300 -1315
rect 6250 -1365 6300 -1335
rect 6250 -1385 6265 -1365
rect 6285 -1385 6300 -1365
rect 6250 -1415 6300 -1385
rect 6250 -1435 6265 -1415
rect 6285 -1435 6300 -1415
rect 6250 -1465 6300 -1435
rect 6250 -1485 6265 -1465
rect 6285 -1485 6300 -1465
rect 6250 -1515 6300 -1485
rect 6250 -1535 6265 -1515
rect 6285 -1535 6300 -1515
rect 6250 -1565 6300 -1535
rect 6250 -1585 6265 -1565
rect 6285 -1585 6300 -1565
rect 6250 -1615 6300 -1585
rect 6250 -1635 6265 -1615
rect 6285 -1635 6300 -1615
rect 6250 -1650 6300 -1635
rect 6400 -1650 6450 -950
rect 6550 -965 6600 -950
rect 6550 -985 6565 -965
rect 6585 -985 6600 -965
rect 6550 -1015 6600 -985
rect 6550 -1035 6565 -1015
rect 6585 -1035 6600 -1015
rect 6550 -1065 6600 -1035
rect 6550 -1085 6565 -1065
rect 6585 -1085 6600 -1065
rect 6550 -1115 6600 -1085
rect 6550 -1135 6565 -1115
rect 6585 -1135 6600 -1115
rect 6550 -1165 6600 -1135
rect 6550 -1185 6565 -1165
rect 6585 -1185 6600 -1165
rect 6550 -1215 6600 -1185
rect 6550 -1235 6565 -1215
rect 6585 -1235 6600 -1215
rect 6550 -1265 6600 -1235
rect 6550 -1285 6565 -1265
rect 6585 -1285 6600 -1265
rect 6550 -1315 6600 -1285
rect 6550 -1335 6565 -1315
rect 6585 -1335 6600 -1315
rect 6550 -1365 6600 -1335
rect 6550 -1385 6565 -1365
rect 6585 -1385 6600 -1365
rect 6550 -1415 6600 -1385
rect 6550 -1435 6565 -1415
rect 6585 -1435 6600 -1415
rect 6550 -1465 6600 -1435
rect 6550 -1485 6565 -1465
rect 6585 -1485 6600 -1465
rect 6550 -1515 6600 -1485
rect 6550 -1535 6565 -1515
rect 6585 -1535 6600 -1515
rect 6550 -1565 6600 -1535
rect 6550 -1585 6565 -1565
rect 6585 -1585 6600 -1565
rect 6550 -1615 6600 -1585
rect 6550 -1635 6565 -1615
rect 6585 -1635 6600 -1615
rect 6550 -1650 6600 -1635
rect 6700 -1650 6750 -950
rect 6850 -965 6900 -950
rect 6850 -985 6865 -965
rect 6885 -985 6900 -965
rect 6850 -1015 6900 -985
rect 6850 -1035 6865 -1015
rect 6885 -1035 6900 -1015
rect 6850 -1065 6900 -1035
rect 6850 -1085 6865 -1065
rect 6885 -1085 6900 -1065
rect 6850 -1115 6900 -1085
rect 6850 -1135 6865 -1115
rect 6885 -1135 6900 -1115
rect 6850 -1165 6900 -1135
rect 6850 -1185 6865 -1165
rect 6885 -1185 6900 -1165
rect 6850 -1215 6900 -1185
rect 6850 -1235 6865 -1215
rect 6885 -1235 6900 -1215
rect 6850 -1265 6900 -1235
rect 6850 -1285 6865 -1265
rect 6885 -1285 6900 -1265
rect 6850 -1315 6900 -1285
rect 6850 -1335 6865 -1315
rect 6885 -1335 6900 -1315
rect 6850 -1365 6900 -1335
rect 6850 -1385 6865 -1365
rect 6885 -1385 6900 -1365
rect 6850 -1415 6900 -1385
rect 6850 -1435 6865 -1415
rect 6885 -1435 6900 -1415
rect 6850 -1465 6900 -1435
rect 6850 -1485 6865 -1465
rect 6885 -1485 6900 -1465
rect 6850 -1515 6900 -1485
rect 6850 -1535 6865 -1515
rect 6885 -1535 6900 -1515
rect 6850 -1565 6900 -1535
rect 6850 -1585 6865 -1565
rect 6885 -1585 6900 -1565
rect 6850 -1615 6900 -1585
rect 6850 -1635 6865 -1615
rect 6885 -1635 6900 -1615
rect 6850 -1650 6900 -1635
rect 7000 -1650 7050 -950
rect 7150 -965 7200 -950
rect 7150 -985 7165 -965
rect 7185 -985 7200 -965
rect 7150 -1015 7200 -985
rect 7150 -1035 7165 -1015
rect 7185 -1035 7200 -1015
rect 7150 -1065 7200 -1035
rect 7150 -1085 7165 -1065
rect 7185 -1085 7200 -1065
rect 7150 -1115 7200 -1085
rect 7150 -1135 7165 -1115
rect 7185 -1135 7200 -1115
rect 7150 -1165 7200 -1135
rect 7150 -1185 7165 -1165
rect 7185 -1185 7200 -1165
rect 7150 -1215 7200 -1185
rect 7150 -1235 7165 -1215
rect 7185 -1235 7200 -1215
rect 7150 -1265 7200 -1235
rect 7150 -1285 7165 -1265
rect 7185 -1285 7200 -1265
rect 7150 -1315 7200 -1285
rect 7150 -1335 7165 -1315
rect 7185 -1335 7200 -1315
rect 7150 -1365 7200 -1335
rect 7150 -1385 7165 -1365
rect 7185 -1385 7200 -1365
rect 7150 -1415 7200 -1385
rect 7150 -1435 7165 -1415
rect 7185 -1435 7200 -1415
rect 7150 -1465 7200 -1435
rect 7150 -1485 7165 -1465
rect 7185 -1485 7200 -1465
rect 7150 -1515 7200 -1485
rect 7150 -1535 7165 -1515
rect 7185 -1535 7200 -1515
rect 7150 -1565 7200 -1535
rect 7150 -1585 7165 -1565
rect 7185 -1585 7200 -1565
rect 7150 -1615 7200 -1585
rect 7150 -1635 7165 -1615
rect 7185 -1635 7200 -1615
rect 7150 -1650 7200 -1635
rect 7300 -1650 7350 -950
rect 7450 -1650 7500 -950
rect 7600 -1650 7650 -950
rect 7750 -1650 7800 -950
rect 7900 -1650 7950 -950
rect 8050 -1650 8100 -950
rect 8200 -1650 8250 -950
rect 8350 -965 8400 -950
rect 8350 -985 8365 -965
rect 8385 -985 8400 -965
rect 8350 -1015 8400 -985
rect 8350 -1035 8365 -1015
rect 8385 -1035 8400 -1015
rect 8350 -1065 8400 -1035
rect 8350 -1085 8365 -1065
rect 8385 -1085 8400 -1065
rect 8350 -1115 8400 -1085
rect 8350 -1135 8365 -1115
rect 8385 -1135 8400 -1115
rect 8350 -1165 8400 -1135
rect 8350 -1185 8365 -1165
rect 8385 -1185 8400 -1165
rect 8350 -1215 8400 -1185
rect 8350 -1235 8365 -1215
rect 8385 -1235 8400 -1215
rect 8350 -1265 8400 -1235
rect 8350 -1285 8365 -1265
rect 8385 -1285 8400 -1265
rect 8350 -1315 8400 -1285
rect 8350 -1335 8365 -1315
rect 8385 -1335 8400 -1315
rect 8350 -1365 8400 -1335
rect 8350 -1385 8365 -1365
rect 8385 -1385 8400 -1365
rect 8350 -1415 8400 -1385
rect 8350 -1435 8365 -1415
rect 8385 -1435 8400 -1415
rect 8350 -1465 8400 -1435
rect 8350 -1485 8365 -1465
rect 8385 -1485 8400 -1465
rect 8350 -1515 8400 -1485
rect 8350 -1535 8365 -1515
rect 8385 -1535 8400 -1515
rect 8350 -1565 8400 -1535
rect 8350 -1585 8365 -1565
rect 8385 -1585 8400 -1565
rect 8350 -1615 8400 -1585
rect 8350 -1635 8365 -1615
rect 8385 -1635 8400 -1615
rect 8350 -1650 8400 -1635
rect 8500 -1650 8550 -950
rect 8650 -1650 8700 -950
rect 8800 -1650 8850 -950
rect 8950 -1650 9000 -950
rect 9100 -1650 9150 -950
rect 9250 -1650 9300 -950
rect 9400 -1650 9450 -950
rect 9550 -965 9600 -950
rect 9550 -985 9565 -965
rect 9585 -985 9600 -965
rect 9550 -1015 9600 -985
rect 9550 -1035 9565 -1015
rect 9585 -1035 9600 -1015
rect 9550 -1065 9600 -1035
rect 9550 -1085 9565 -1065
rect 9585 -1085 9600 -1065
rect 9550 -1115 9600 -1085
rect 9550 -1135 9565 -1115
rect 9585 -1135 9600 -1115
rect 9550 -1165 9600 -1135
rect 9550 -1185 9565 -1165
rect 9585 -1185 9600 -1165
rect 9550 -1215 9600 -1185
rect 9550 -1235 9565 -1215
rect 9585 -1235 9600 -1215
rect 9550 -1265 9600 -1235
rect 9550 -1285 9565 -1265
rect 9585 -1285 9600 -1265
rect 9550 -1315 9600 -1285
rect 9550 -1335 9565 -1315
rect 9585 -1335 9600 -1315
rect 9550 -1365 9600 -1335
rect 9550 -1385 9565 -1365
rect 9585 -1385 9600 -1365
rect 9550 -1415 9600 -1385
rect 9550 -1435 9565 -1415
rect 9585 -1435 9600 -1415
rect 9550 -1465 9600 -1435
rect 9550 -1485 9565 -1465
rect 9585 -1485 9600 -1465
rect 9550 -1515 9600 -1485
rect 9550 -1535 9565 -1515
rect 9585 -1535 9600 -1515
rect 9550 -1565 9600 -1535
rect 9550 -1585 9565 -1565
rect 9585 -1585 9600 -1565
rect 9550 -1615 9600 -1585
rect 9550 -1635 9565 -1615
rect 9585 -1635 9600 -1615
rect 9550 -1650 9600 -1635
rect 9700 -1650 9750 -950
rect 9850 -1650 9900 -950
rect 10000 -1650 10050 -950
rect 10150 -1650 10200 -950
rect 10300 -1650 10350 -950
rect 10450 -1650 10500 -950
rect 10600 -1650 10650 -950
rect 10750 -965 10800 -950
rect 10750 -985 10765 -965
rect 10785 -985 10800 -965
rect 10750 -1015 10800 -985
rect 10750 -1035 10765 -1015
rect 10785 -1035 10800 -1015
rect 10750 -1065 10800 -1035
rect 10750 -1085 10765 -1065
rect 10785 -1085 10800 -1065
rect 10750 -1115 10800 -1085
rect 10750 -1135 10765 -1115
rect 10785 -1135 10800 -1115
rect 10750 -1165 10800 -1135
rect 10750 -1185 10765 -1165
rect 10785 -1185 10800 -1165
rect 10750 -1215 10800 -1185
rect 10750 -1235 10765 -1215
rect 10785 -1235 10800 -1215
rect 10750 -1265 10800 -1235
rect 10750 -1285 10765 -1265
rect 10785 -1285 10800 -1265
rect 10750 -1315 10800 -1285
rect 10750 -1335 10765 -1315
rect 10785 -1335 10800 -1315
rect 10750 -1365 10800 -1335
rect 10750 -1385 10765 -1365
rect 10785 -1385 10800 -1365
rect 10750 -1415 10800 -1385
rect 10750 -1435 10765 -1415
rect 10785 -1435 10800 -1415
rect 10750 -1465 10800 -1435
rect 10750 -1485 10765 -1465
rect 10785 -1485 10800 -1465
rect 10750 -1515 10800 -1485
rect 10750 -1535 10765 -1515
rect 10785 -1535 10800 -1515
rect 10750 -1565 10800 -1535
rect 10750 -1585 10765 -1565
rect 10785 -1585 10800 -1565
rect 10750 -1615 10800 -1585
rect 10750 -1635 10765 -1615
rect 10785 -1635 10800 -1615
rect 10750 -1650 10800 -1635
rect 10900 -1650 10950 -950
rect 11050 -1650 11100 -950
rect 11200 -1650 11250 -950
rect 11350 -1650 11400 -950
rect 11500 -1650 11550 -950
rect 11650 -1650 11700 -950
rect 11800 -1650 11850 -950
rect 11950 -965 12000 -950
rect 11950 -985 11965 -965
rect 11985 -985 12000 -965
rect 11950 -1015 12000 -985
rect 11950 -1035 11965 -1015
rect 11985 -1035 12000 -1015
rect 11950 -1065 12000 -1035
rect 11950 -1085 11965 -1065
rect 11985 -1085 12000 -1065
rect 11950 -1115 12000 -1085
rect 11950 -1135 11965 -1115
rect 11985 -1135 12000 -1115
rect 11950 -1165 12000 -1135
rect 11950 -1185 11965 -1165
rect 11985 -1185 12000 -1165
rect 11950 -1215 12000 -1185
rect 11950 -1235 11965 -1215
rect 11985 -1235 12000 -1215
rect 11950 -1265 12000 -1235
rect 11950 -1285 11965 -1265
rect 11985 -1285 12000 -1265
rect 11950 -1315 12000 -1285
rect 11950 -1335 11965 -1315
rect 11985 -1335 12000 -1315
rect 11950 -1365 12000 -1335
rect 11950 -1385 11965 -1365
rect 11985 -1385 12000 -1365
rect 11950 -1415 12000 -1385
rect 11950 -1435 11965 -1415
rect 11985 -1435 12000 -1415
rect 11950 -1465 12000 -1435
rect 11950 -1485 11965 -1465
rect 11985 -1485 12000 -1465
rect 11950 -1515 12000 -1485
rect 11950 -1535 11965 -1515
rect 11985 -1535 12000 -1515
rect 11950 -1565 12000 -1535
rect 11950 -1585 11965 -1565
rect 11985 -1585 12000 -1565
rect 11950 -1615 12000 -1585
rect 11950 -1635 11965 -1615
rect 11985 -1635 12000 -1615
rect 11950 -1650 12000 -1635
rect 12100 -1650 12150 -950
rect 12250 -965 12300 -950
rect 12250 -985 12265 -965
rect 12285 -985 12300 -965
rect 12250 -1015 12300 -985
rect 12250 -1035 12265 -1015
rect 12285 -1035 12300 -1015
rect 12250 -1065 12300 -1035
rect 12250 -1085 12265 -1065
rect 12285 -1085 12300 -1065
rect 12250 -1115 12300 -1085
rect 12250 -1135 12265 -1115
rect 12285 -1135 12300 -1115
rect 12250 -1165 12300 -1135
rect 12250 -1185 12265 -1165
rect 12285 -1185 12300 -1165
rect 12250 -1215 12300 -1185
rect 12250 -1235 12265 -1215
rect 12285 -1235 12300 -1215
rect 12250 -1265 12300 -1235
rect 12250 -1285 12265 -1265
rect 12285 -1285 12300 -1265
rect 12250 -1315 12300 -1285
rect 12250 -1335 12265 -1315
rect 12285 -1335 12300 -1315
rect 12250 -1365 12300 -1335
rect 12250 -1385 12265 -1365
rect 12285 -1385 12300 -1365
rect 12250 -1415 12300 -1385
rect 12250 -1435 12265 -1415
rect 12285 -1435 12300 -1415
rect 12250 -1465 12300 -1435
rect 12250 -1485 12265 -1465
rect 12285 -1485 12300 -1465
rect 12250 -1515 12300 -1485
rect 12250 -1535 12265 -1515
rect 12285 -1535 12300 -1515
rect 12250 -1565 12300 -1535
rect 12250 -1585 12265 -1565
rect 12285 -1585 12300 -1565
rect 12250 -1615 12300 -1585
rect 12250 -1635 12265 -1615
rect 12285 -1635 12300 -1615
rect 12250 -1650 12300 -1635
rect 12400 -1650 12450 -950
rect 12550 -965 12600 -950
rect 12550 -985 12565 -965
rect 12585 -985 12600 -965
rect 12550 -1015 12600 -985
rect 12550 -1035 12565 -1015
rect 12585 -1035 12600 -1015
rect 12550 -1065 12600 -1035
rect 12550 -1085 12565 -1065
rect 12585 -1085 12600 -1065
rect 12550 -1115 12600 -1085
rect 12550 -1135 12565 -1115
rect 12585 -1135 12600 -1115
rect 12550 -1165 12600 -1135
rect 12550 -1185 12565 -1165
rect 12585 -1185 12600 -1165
rect 12550 -1215 12600 -1185
rect 12550 -1235 12565 -1215
rect 12585 -1235 12600 -1215
rect 12550 -1265 12600 -1235
rect 12550 -1285 12565 -1265
rect 12585 -1285 12600 -1265
rect 12550 -1315 12600 -1285
rect 12550 -1335 12565 -1315
rect 12585 -1335 12600 -1315
rect 12550 -1365 12600 -1335
rect 12550 -1385 12565 -1365
rect 12585 -1385 12600 -1365
rect 12550 -1415 12600 -1385
rect 12550 -1435 12565 -1415
rect 12585 -1435 12600 -1415
rect 12550 -1465 12600 -1435
rect 12550 -1485 12565 -1465
rect 12585 -1485 12600 -1465
rect 12550 -1515 12600 -1485
rect 12550 -1535 12565 -1515
rect 12585 -1535 12600 -1515
rect 12550 -1565 12600 -1535
rect 12550 -1585 12565 -1565
rect 12585 -1585 12600 -1565
rect 12550 -1615 12600 -1585
rect 12550 -1635 12565 -1615
rect 12585 -1635 12600 -1615
rect 12550 -1650 12600 -1635
rect 12700 -1650 12750 -950
rect 12850 -965 12900 -950
rect 12850 -985 12865 -965
rect 12885 -985 12900 -965
rect 12850 -1015 12900 -985
rect 12850 -1035 12865 -1015
rect 12885 -1035 12900 -1015
rect 12850 -1065 12900 -1035
rect 12850 -1085 12865 -1065
rect 12885 -1085 12900 -1065
rect 12850 -1115 12900 -1085
rect 12850 -1135 12865 -1115
rect 12885 -1135 12900 -1115
rect 12850 -1165 12900 -1135
rect 12850 -1185 12865 -1165
rect 12885 -1185 12900 -1165
rect 12850 -1215 12900 -1185
rect 12850 -1235 12865 -1215
rect 12885 -1235 12900 -1215
rect 12850 -1265 12900 -1235
rect 12850 -1285 12865 -1265
rect 12885 -1285 12900 -1265
rect 12850 -1315 12900 -1285
rect 12850 -1335 12865 -1315
rect 12885 -1335 12900 -1315
rect 12850 -1365 12900 -1335
rect 12850 -1385 12865 -1365
rect 12885 -1385 12900 -1365
rect 12850 -1415 12900 -1385
rect 12850 -1435 12865 -1415
rect 12885 -1435 12900 -1415
rect 12850 -1465 12900 -1435
rect 12850 -1485 12865 -1465
rect 12885 -1485 12900 -1465
rect 12850 -1515 12900 -1485
rect 12850 -1535 12865 -1515
rect 12885 -1535 12900 -1515
rect 12850 -1565 12900 -1535
rect 12850 -1585 12865 -1565
rect 12885 -1585 12900 -1565
rect 12850 -1615 12900 -1585
rect 12850 -1635 12865 -1615
rect 12885 -1635 12900 -1615
rect 12850 -1650 12900 -1635
rect 13000 -1650 13050 -950
rect 13150 -965 13200 -950
rect 13150 -985 13165 -965
rect 13185 -985 13200 -965
rect 13150 -1015 13200 -985
rect 13150 -1035 13165 -1015
rect 13185 -1035 13200 -1015
rect 13150 -1065 13200 -1035
rect 13150 -1085 13165 -1065
rect 13185 -1085 13200 -1065
rect 13150 -1115 13200 -1085
rect 13150 -1135 13165 -1115
rect 13185 -1135 13200 -1115
rect 13150 -1165 13200 -1135
rect 13150 -1185 13165 -1165
rect 13185 -1185 13200 -1165
rect 13150 -1215 13200 -1185
rect 13150 -1235 13165 -1215
rect 13185 -1235 13200 -1215
rect 13150 -1265 13200 -1235
rect 13150 -1285 13165 -1265
rect 13185 -1285 13200 -1265
rect 13150 -1315 13200 -1285
rect 13150 -1335 13165 -1315
rect 13185 -1335 13200 -1315
rect 13150 -1365 13200 -1335
rect 13150 -1385 13165 -1365
rect 13185 -1385 13200 -1365
rect 13150 -1415 13200 -1385
rect 13150 -1435 13165 -1415
rect 13185 -1435 13200 -1415
rect 13150 -1465 13200 -1435
rect 13150 -1485 13165 -1465
rect 13185 -1485 13200 -1465
rect 13150 -1515 13200 -1485
rect 13150 -1535 13165 -1515
rect 13185 -1535 13200 -1515
rect 13150 -1565 13200 -1535
rect 13150 -1585 13165 -1565
rect 13185 -1585 13200 -1565
rect 13150 -1615 13200 -1585
rect 13150 -1635 13165 -1615
rect 13185 -1635 13200 -1615
rect 13150 -1650 13200 -1635
rect 13300 -1650 13350 -950
rect 13450 -965 13500 -950
rect 13450 -985 13465 -965
rect 13485 -985 13500 -965
rect 13450 -1015 13500 -985
rect 13450 -1035 13465 -1015
rect 13485 -1035 13500 -1015
rect 13450 -1065 13500 -1035
rect 13450 -1085 13465 -1065
rect 13485 -1085 13500 -1065
rect 13450 -1115 13500 -1085
rect 13450 -1135 13465 -1115
rect 13485 -1135 13500 -1115
rect 13450 -1165 13500 -1135
rect 13450 -1185 13465 -1165
rect 13485 -1185 13500 -1165
rect 13450 -1215 13500 -1185
rect 13450 -1235 13465 -1215
rect 13485 -1235 13500 -1215
rect 13450 -1265 13500 -1235
rect 13450 -1285 13465 -1265
rect 13485 -1285 13500 -1265
rect 13450 -1315 13500 -1285
rect 13450 -1335 13465 -1315
rect 13485 -1335 13500 -1315
rect 13450 -1365 13500 -1335
rect 13450 -1385 13465 -1365
rect 13485 -1385 13500 -1365
rect 13450 -1415 13500 -1385
rect 13450 -1435 13465 -1415
rect 13485 -1435 13500 -1415
rect 13450 -1465 13500 -1435
rect 13450 -1485 13465 -1465
rect 13485 -1485 13500 -1465
rect 13450 -1515 13500 -1485
rect 13450 -1535 13465 -1515
rect 13485 -1535 13500 -1515
rect 13450 -1565 13500 -1535
rect 13450 -1585 13465 -1565
rect 13485 -1585 13500 -1565
rect 13450 -1615 13500 -1585
rect 13450 -1635 13465 -1615
rect 13485 -1635 13500 -1615
rect 13450 -1650 13500 -1635
rect 13600 -1650 13650 -950
rect 13750 -965 13800 -950
rect 13750 -985 13765 -965
rect 13785 -985 13800 -965
rect 13750 -1015 13800 -985
rect 13750 -1035 13765 -1015
rect 13785 -1035 13800 -1015
rect 13750 -1065 13800 -1035
rect 13750 -1085 13765 -1065
rect 13785 -1085 13800 -1065
rect 13750 -1115 13800 -1085
rect 13750 -1135 13765 -1115
rect 13785 -1135 13800 -1115
rect 13750 -1165 13800 -1135
rect 13750 -1185 13765 -1165
rect 13785 -1185 13800 -1165
rect 13750 -1215 13800 -1185
rect 13750 -1235 13765 -1215
rect 13785 -1235 13800 -1215
rect 13750 -1265 13800 -1235
rect 13750 -1285 13765 -1265
rect 13785 -1285 13800 -1265
rect 13750 -1315 13800 -1285
rect 13750 -1335 13765 -1315
rect 13785 -1335 13800 -1315
rect 13750 -1365 13800 -1335
rect 13750 -1385 13765 -1365
rect 13785 -1385 13800 -1365
rect 13750 -1415 13800 -1385
rect 13750 -1435 13765 -1415
rect 13785 -1435 13800 -1415
rect 13750 -1465 13800 -1435
rect 13750 -1485 13765 -1465
rect 13785 -1485 13800 -1465
rect 13750 -1515 13800 -1485
rect 13750 -1535 13765 -1515
rect 13785 -1535 13800 -1515
rect 13750 -1565 13800 -1535
rect 13750 -1585 13765 -1565
rect 13785 -1585 13800 -1565
rect 13750 -1615 13800 -1585
rect 13750 -1635 13765 -1615
rect 13785 -1635 13800 -1615
rect 13750 -1650 13800 -1635
rect 13900 -1650 13950 -950
rect 14050 -965 14100 -950
rect 14050 -985 14065 -965
rect 14085 -985 14100 -965
rect 14050 -1015 14100 -985
rect 14050 -1035 14065 -1015
rect 14085 -1035 14100 -1015
rect 14050 -1065 14100 -1035
rect 14050 -1085 14065 -1065
rect 14085 -1085 14100 -1065
rect 14050 -1115 14100 -1085
rect 14050 -1135 14065 -1115
rect 14085 -1135 14100 -1115
rect 14050 -1165 14100 -1135
rect 14050 -1185 14065 -1165
rect 14085 -1185 14100 -1165
rect 14050 -1215 14100 -1185
rect 14050 -1235 14065 -1215
rect 14085 -1235 14100 -1215
rect 14050 -1265 14100 -1235
rect 14050 -1285 14065 -1265
rect 14085 -1285 14100 -1265
rect 14050 -1315 14100 -1285
rect 14050 -1335 14065 -1315
rect 14085 -1335 14100 -1315
rect 14050 -1365 14100 -1335
rect 14050 -1385 14065 -1365
rect 14085 -1385 14100 -1365
rect 14050 -1415 14100 -1385
rect 14050 -1435 14065 -1415
rect 14085 -1435 14100 -1415
rect 14050 -1465 14100 -1435
rect 14050 -1485 14065 -1465
rect 14085 -1485 14100 -1465
rect 14050 -1515 14100 -1485
rect 14050 -1535 14065 -1515
rect 14085 -1535 14100 -1515
rect 14050 -1565 14100 -1535
rect 14050 -1585 14065 -1565
rect 14085 -1585 14100 -1565
rect 14050 -1615 14100 -1585
rect 14050 -1635 14065 -1615
rect 14085 -1635 14100 -1615
rect 14050 -1650 14100 -1635
rect 14200 -1650 14250 -950
rect 14350 -965 14400 -950
rect 14350 -985 14365 -965
rect 14385 -985 14400 -965
rect 14350 -1015 14400 -985
rect 14350 -1035 14365 -1015
rect 14385 -1035 14400 -1015
rect 14350 -1065 14400 -1035
rect 14350 -1085 14365 -1065
rect 14385 -1085 14400 -1065
rect 14350 -1115 14400 -1085
rect 14350 -1135 14365 -1115
rect 14385 -1135 14400 -1115
rect 14350 -1165 14400 -1135
rect 14350 -1185 14365 -1165
rect 14385 -1185 14400 -1165
rect 14350 -1215 14400 -1185
rect 14350 -1235 14365 -1215
rect 14385 -1235 14400 -1215
rect 14350 -1265 14400 -1235
rect 14350 -1285 14365 -1265
rect 14385 -1285 14400 -1265
rect 14350 -1315 14400 -1285
rect 14350 -1335 14365 -1315
rect 14385 -1335 14400 -1315
rect 14350 -1365 14400 -1335
rect 14350 -1385 14365 -1365
rect 14385 -1385 14400 -1365
rect 14350 -1415 14400 -1385
rect 14350 -1435 14365 -1415
rect 14385 -1435 14400 -1415
rect 14350 -1465 14400 -1435
rect 14350 -1485 14365 -1465
rect 14385 -1485 14400 -1465
rect 14350 -1515 14400 -1485
rect 14350 -1535 14365 -1515
rect 14385 -1535 14400 -1515
rect 14350 -1565 14400 -1535
rect 14350 -1585 14365 -1565
rect 14385 -1585 14400 -1565
rect 14350 -1615 14400 -1585
rect 14350 -1635 14365 -1615
rect 14385 -1635 14400 -1615
rect 14350 -1650 14400 -1635
rect 14500 -1650 14550 -950
rect 14650 -1650 14700 -950
rect 14800 -1650 14850 -950
rect 14950 -1650 15000 -950
rect 15100 -1650 15150 -950
rect 15250 -1650 15300 -950
rect 15400 -1650 15450 -950
rect 15550 -965 15600 -950
rect 15550 -985 15565 -965
rect 15585 -985 15600 -965
rect 15550 -1015 15600 -985
rect 15550 -1035 15565 -1015
rect 15585 -1035 15600 -1015
rect 15550 -1065 15600 -1035
rect 15550 -1085 15565 -1065
rect 15585 -1085 15600 -1065
rect 15550 -1115 15600 -1085
rect 15550 -1135 15565 -1115
rect 15585 -1135 15600 -1115
rect 15550 -1165 15600 -1135
rect 15550 -1185 15565 -1165
rect 15585 -1185 15600 -1165
rect 15550 -1215 15600 -1185
rect 15550 -1235 15565 -1215
rect 15585 -1235 15600 -1215
rect 15550 -1265 15600 -1235
rect 15550 -1285 15565 -1265
rect 15585 -1285 15600 -1265
rect 15550 -1315 15600 -1285
rect 15550 -1335 15565 -1315
rect 15585 -1335 15600 -1315
rect 15550 -1365 15600 -1335
rect 15550 -1385 15565 -1365
rect 15585 -1385 15600 -1365
rect 15550 -1415 15600 -1385
rect 15550 -1435 15565 -1415
rect 15585 -1435 15600 -1415
rect 15550 -1465 15600 -1435
rect 15550 -1485 15565 -1465
rect 15585 -1485 15600 -1465
rect 15550 -1515 15600 -1485
rect 15550 -1535 15565 -1515
rect 15585 -1535 15600 -1515
rect 15550 -1565 15600 -1535
rect 15550 -1585 15565 -1565
rect 15585 -1585 15600 -1565
rect 15550 -1615 15600 -1585
rect 15550 -1635 15565 -1615
rect 15585 -1635 15600 -1615
rect 15550 -1650 15600 -1635
rect 15700 -1650 15750 -950
rect 15850 -1650 15900 -950
rect 16000 -1650 16050 -950
rect 16150 -1650 16200 -950
rect 16300 -1650 16350 -950
rect 16450 -1650 16500 -950
rect 16600 -1650 16650 -950
rect 16750 -965 16800 -950
rect 16750 -985 16765 -965
rect 16785 -985 16800 -965
rect 16750 -1015 16800 -985
rect 16750 -1035 16765 -1015
rect 16785 -1035 16800 -1015
rect 16750 -1065 16800 -1035
rect 16750 -1085 16765 -1065
rect 16785 -1085 16800 -1065
rect 16750 -1115 16800 -1085
rect 16750 -1135 16765 -1115
rect 16785 -1135 16800 -1115
rect 16750 -1165 16800 -1135
rect 16750 -1185 16765 -1165
rect 16785 -1185 16800 -1165
rect 16750 -1215 16800 -1185
rect 16750 -1235 16765 -1215
rect 16785 -1235 16800 -1215
rect 16750 -1265 16800 -1235
rect 16750 -1285 16765 -1265
rect 16785 -1285 16800 -1265
rect 16750 -1315 16800 -1285
rect 16750 -1335 16765 -1315
rect 16785 -1335 16800 -1315
rect 16750 -1365 16800 -1335
rect 16750 -1385 16765 -1365
rect 16785 -1385 16800 -1365
rect 16750 -1415 16800 -1385
rect 16750 -1435 16765 -1415
rect 16785 -1435 16800 -1415
rect 16750 -1465 16800 -1435
rect 16750 -1485 16765 -1465
rect 16785 -1485 16800 -1465
rect 16750 -1515 16800 -1485
rect 16750 -1535 16765 -1515
rect 16785 -1535 16800 -1515
rect 16750 -1565 16800 -1535
rect 16750 -1585 16765 -1565
rect 16785 -1585 16800 -1565
rect 16750 -1615 16800 -1585
rect 16750 -1635 16765 -1615
rect 16785 -1635 16800 -1615
rect 16750 -1650 16800 -1635
rect 16900 -1650 16950 -950
rect 17050 -1650 17100 -950
rect 17200 -1650 17250 -950
rect 17350 -1650 17400 -950
rect 17500 -1650 17550 -950
rect 17650 -1650 17700 -950
rect 17800 -1650 17850 -950
rect 17950 -965 18000 -950
rect 17950 -985 17965 -965
rect 17985 -985 18000 -965
rect 17950 -1015 18000 -985
rect 17950 -1035 17965 -1015
rect 17985 -1035 18000 -1015
rect 17950 -1065 18000 -1035
rect 17950 -1085 17965 -1065
rect 17985 -1085 18000 -1065
rect 17950 -1115 18000 -1085
rect 17950 -1135 17965 -1115
rect 17985 -1135 18000 -1115
rect 17950 -1165 18000 -1135
rect 17950 -1185 17965 -1165
rect 17985 -1185 18000 -1165
rect 17950 -1215 18000 -1185
rect 17950 -1235 17965 -1215
rect 17985 -1235 18000 -1215
rect 17950 -1265 18000 -1235
rect 17950 -1285 17965 -1265
rect 17985 -1285 18000 -1265
rect 17950 -1315 18000 -1285
rect 17950 -1335 17965 -1315
rect 17985 -1335 18000 -1315
rect 17950 -1365 18000 -1335
rect 17950 -1385 17965 -1365
rect 17985 -1385 18000 -1365
rect 17950 -1415 18000 -1385
rect 17950 -1435 17965 -1415
rect 17985 -1435 18000 -1415
rect 17950 -1465 18000 -1435
rect 17950 -1485 17965 -1465
rect 17985 -1485 18000 -1465
rect 17950 -1515 18000 -1485
rect 17950 -1535 17965 -1515
rect 17985 -1535 18000 -1515
rect 17950 -1565 18000 -1535
rect 17950 -1585 17965 -1565
rect 17985 -1585 18000 -1565
rect 17950 -1615 18000 -1585
rect 17950 -1635 17965 -1615
rect 17985 -1635 18000 -1615
rect 17950 -1650 18000 -1635
rect 18100 -1650 18150 -950
rect 18250 -1650 18300 -950
rect 18400 -1650 18450 -950
rect 18550 -1650 18600 -950
rect 18700 -1650 18750 -950
rect 18850 -1650 18900 -950
rect 19000 -1650 19050 -950
rect 19150 -965 19200 -950
rect 19150 -985 19165 -965
rect 19185 -985 19200 -965
rect 19150 -1015 19200 -985
rect 19150 -1035 19165 -1015
rect 19185 -1035 19200 -1015
rect 19150 -1065 19200 -1035
rect 19150 -1085 19165 -1065
rect 19185 -1085 19200 -1065
rect 19150 -1115 19200 -1085
rect 19150 -1135 19165 -1115
rect 19185 -1135 19200 -1115
rect 19150 -1165 19200 -1135
rect 19150 -1185 19165 -1165
rect 19185 -1185 19200 -1165
rect 19150 -1215 19200 -1185
rect 19150 -1235 19165 -1215
rect 19185 -1235 19200 -1215
rect 19150 -1265 19200 -1235
rect 19150 -1285 19165 -1265
rect 19185 -1285 19200 -1265
rect 19150 -1315 19200 -1285
rect 19150 -1335 19165 -1315
rect 19185 -1335 19200 -1315
rect 19150 -1365 19200 -1335
rect 19150 -1385 19165 -1365
rect 19185 -1385 19200 -1365
rect 19150 -1415 19200 -1385
rect 19150 -1435 19165 -1415
rect 19185 -1435 19200 -1415
rect 19150 -1465 19200 -1435
rect 19150 -1485 19165 -1465
rect 19185 -1485 19200 -1465
rect 19150 -1515 19200 -1485
rect 19150 -1535 19165 -1515
rect 19185 -1535 19200 -1515
rect 19150 -1565 19200 -1535
rect 19150 -1585 19165 -1565
rect 19185 -1585 19200 -1565
rect 19150 -1615 19200 -1585
rect 19150 -1635 19165 -1615
rect 19185 -1635 19200 -1615
rect 19150 -1650 19200 -1635
rect 19300 -1650 19350 -950
rect 19450 -1650 19500 -950
rect 19600 -1650 19650 -950
rect 19750 -1650 19800 -950
rect 19900 -1650 19950 -950
rect 20050 -1650 20100 -950
rect 20200 -1650 20250 -950
rect 20350 -965 20400 -950
rect 20350 -985 20365 -965
rect 20385 -985 20400 -965
rect 20350 -1015 20400 -985
rect 20350 -1035 20365 -1015
rect 20385 -1035 20400 -1015
rect 20350 -1065 20400 -1035
rect 20350 -1085 20365 -1065
rect 20385 -1085 20400 -1065
rect 20350 -1115 20400 -1085
rect 20350 -1135 20365 -1115
rect 20385 -1135 20400 -1115
rect 20350 -1165 20400 -1135
rect 20350 -1185 20365 -1165
rect 20385 -1185 20400 -1165
rect 20350 -1215 20400 -1185
rect 20350 -1235 20365 -1215
rect 20385 -1235 20400 -1215
rect 20350 -1265 20400 -1235
rect 20350 -1285 20365 -1265
rect 20385 -1285 20400 -1265
rect 20350 -1315 20400 -1285
rect 20350 -1335 20365 -1315
rect 20385 -1335 20400 -1315
rect 20350 -1365 20400 -1335
rect 20350 -1385 20365 -1365
rect 20385 -1385 20400 -1365
rect 20350 -1415 20400 -1385
rect 20350 -1435 20365 -1415
rect 20385 -1435 20400 -1415
rect 20350 -1465 20400 -1435
rect 20350 -1485 20365 -1465
rect 20385 -1485 20400 -1465
rect 20350 -1515 20400 -1485
rect 20350 -1535 20365 -1515
rect 20385 -1535 20400 -1515
rect 20350 -1565 20400 -1535
rect 20350 -1585 20365 -1565
rect 20385 -1585 20400 -1565
rect 20350 -1615 20400 -1585
rect 20350 -1635 20365 -1615
rect 20385 -1635 20400 -1615
rect 20350 -1650 20400 -1635
rect 20500 -1650 20550 -950
rect 20650 -1650 20700 -950
rect 20800 -1650 20850 -950
rect 20950 -1650 21000 -950
rect 21100 -1650 21150 -950
rect 21250 -1650 21300 -950
rect 21400 -1650 21450 -950
rect 21550 -965 21600 -950
rect 21550 -985 21565 -965
rect 21585 -985 21600 -965
rect 21550 -1015 21600 -985
rect 21550 -1035 21565 -1015
rect 21585 -1035 21600 -1015
rect 21550 -1065 21600 -1035
rect 21550 -1085 21565 -1065
rect 21585 -1085 21600 -1065
rect 21550 -1115 21600 -1085
rect 21550 -1135 21565 -1115
rect 21585 -1135 21600 -1115
rect 21550 -1165 21600 -1135
rect 21550 -1185 21565 -1165
rect 21585 -1185 21600 -1165
rect 21550 -1215 21600 -1185
rect 21550 -1235 21565 -1215
rect 21585 -1235 21600 -1215
rect 21550 -1265 21600 -1235
rect 21550 -1285 21565 -1265
rect 21585 -1285 21600 -1265
rect 21550 -1315 21600 -1285
rect 21550 -1335 21565 -1315
rect 21585 -1335 21600 -1315
rect 21550 -1365 21600 -1335
rect 21550 -1385 21565 -1365
rect 21585 -1385 21600 -1365
rect 21550 -1415 21600 -1385
rect 21550 -1435 21565 -1415
rect 21585 -1435 21600 -1415
rect 21550 -1465 21600 -1435
rect 21550 -1485 21565 -1465
rect 21585 -1485 21600 -1465
rect 21550 -1515 21600 -1485
rect 21550 -1535 21565 -1515
rect 21585 -1535 21600 -1515
rect 21550 -1565 21600 -1535
rect 21550 -1585 21565 -1565
rect 21585 -1585 21600 -1565
rect 21550 -1615 21600 -1585
rect 21550 -1635 21565 -1615
rect 21585 -1635 21600 -1615
rect 21550 -1650 21600 -1635
rect 21700 -1650 21750 -950
rect 21850 -1650 21900 -950
rect 22000 -1650 22050 -950
rect 22150 -1650 22200 -950
rect 22300 -1650 22350 -950
rect 22450 -965 22500 -950
rect 22450 -985 22465 -965
rect 22485 -985 22500 -965
rect 22450 -1015 22500 -985
rect 22450 -1035 22465 -1015
rect 22485 -1035 22500 -1015
rect 22450 -1065 22500 -1035
rect 22450 -1085 22465 -1065
rect 22485 -1085 22500 -1065
rect 22450 -1115 22500 -1085
rect 22450 -1135 22465 -1115
rect 22485 -1135 22500 -1115
rect 22450 -1165 22500 -1135
rect 22450 -1185 22465 -1165
rect 22485 -1185 22500 -1165
rect 22450 -1215 22500 -1185
rect 22450 -1235 22465 -1215
rect 22485 -1235 22500 -1215
rect 22450 -1265 22500 -1235
rect 22450 -1285 22465 -1265
rect 22485 -1285 22500 -1265
rect 22450 -1315 22500 -1285
rect 22450 -1335 22465 -1315
rect 22485 -1335 22500 -1315
rect 22450 -1365 22500 -1335
rect 22450 -1385 22465 -1365
rect 22485 -1385 22500 -1365
rect 22450 -1415 22500 -1385
rect 22450 -1435 22465 -1415
rect 22485 -1435 22500 -1415
rect 22450 -1465 22500 -1435
rect 22450 -1485 22465 -1465
rect 22485 -1485 22500 -1465
rect 22450 -1515 22500 -1485
rect 22450 -1535 22465 -1515
rect 22485 -1535 22500 -1515
rect 22450 -1565 22500 -1535
rect 22450 -1585 22465 -1565
rect 22485 -1585 22500 -1565
rect 22450 -1615 22500 -1585
rect 22450 -1635 22465 -1615
rect 22485 -1635 22500 -1615
rect 22450 -1650 22500 -1635
rect 22600 -1650 22650 -950
rect 22750 -1650 22800 -950
rect 22900 -1650 22950 -950
rect 23050 -1650 23100 -950
rect 23200 -1650 23250 -950
rect 23350 -965 23400 -950
rect 23350 -985 23365 -965
rect 23385 -985 23400 -965
rect 23350 -1015 23400 -985
rect 23350 -1035 23365 -1015
rect 23385 -1035 23400 -1015
rect 23350 -1065 23400 -1035
rect 23350 -1085 23365 -1065
rect 23385 -1085 23400 -1065
rect 23350 -1115 23400 -1085
rect 23350 -1135 23365 -1115
rect 23385 -1135 23400 -1115
rect 23350 -1165 23400 -1135
rect 23350 -1185 23365 -1165
rect 23385 -1185 23400 -1165
rect 23350 -1215 23400 -1185
rect 23350 -1235 23365 -1215
rect 23385 -1235 23400 -1215
rect 23350 -1265 23400 -1235
rect 23350 -1285 23365 -1265
rect 23385 -1285 23400 -1265
rect 23350 -1315 23400 -1285
rect 23350 -1335 23365 -1315
rect 23385 -1335 23400 -1315
rect 23350 -1365 23400 -1335
rect 23350 -1385 23365 -1365
rect 23385 -1385 23400 -1365
rect 23350 -1415 23400 -1385
rect 23350 -1435 23365 -1415
rect 23385 -1435 23400 -1415
rect 23350 -1465 23400 -1435
rect 23350 -1485 23365 -1465
rect 23385 -1485 23400 -1465
rect 23350 -1515 23400 -1485
rect 23350 -1535 23365 -1515
rect 23385 -1535 23400 -1515
rect 23350 -1565 23400 -1535
rect 23350 -1585 23365 -1565
rect 23385 -1585 23400 -1565
rect 23350 -1615 23400 -1585
rect 23350 -1635 23365 -1615
rect 23385 -1635 23400 -1615
rect 23350 -1650 23400 -1635
rect 23500 -1650 23550 -950
rect 23650 -1650 23700 -950
rect 23800 -1650 23850 -950
rect 23950 -1650 24000 -950
rect 24100 -1650 24150 -950
rect 24250 -1650 24300 -950
rect 24400 -1650 24450 -950
rect 24550 -965 24600 -950
rect 24550 -985 24565 -965
rect 24585 -985 24600 -965
rect 24550 -1015 24600 -985
rect 24550 -1035 24565 -1015
rect 24585 -1035 24600 -1015
rect 24550 -1065 24600 -1035
rect 24550 -1085 24565 -1065
rect 24585 -1085 24600 -1065
rect 24550 -1115 24600 -1085
rect 24550 -1135 24565 -1115
rect 24585 -1135 24600 -1115
rect 24550 -1165 24600 -1135
rect 24550 -1185 24565 -1165
rect 24585 -1185 24600 -1165
rect 24550 -1215 24600 -1185
rect 24550 -1235 24565 -1215
rect 24585 -1235 24600 -1215
rect 24550 -1265 24600 -1235
rect 24550 -1285 24565 -1265
rect 24585 -1285 24600 -1265
rect 24550 -1315 24600 -1285
rect 24550 -1335 24565 -1315
rect 24585 -1335 24600 -1315
rect 24550 -1365 24600 -1335
rect 24550 -1385 24565 -1365
rect 24585 -1385 24600 -1365
rect 24550 -1415 24600 -1385
rect 24550 -1435 24565 -1415
rect 24585 -1435 24600 -1415
rect 24550 -1465 24600 -1435
rect 24550 -1485 24565 -1465
rect 24585 -1485 24600 -1465
rect 24550 -1515 24600 -1485
rect 24550 -1535 24565 -1515
rect 24585 -1535 24600 -1515
rect 24550 -1565 24600 -1535
rect 24550 -1585 24565 -1565
rect 24585 -1585 24600 -1565
rect 24550 -1615 24600 -1585
rect 24550 -1635 24565 -1615
rect 24585 -1635 24600 -1615
rect 24550 -1650 24600 -1635
rect 24700 -1650 24750 -950
rect 24850 -1650 24900 -950
rect 25000 -1650 25050 -950
rect 25150 -1650 25200 -950
rect 25300 -1650 25350 -950
rect 25450 -1650 25500 -950
rect 25600 -1650 25650 -950
rect 25750 -965 25800 -950
rect 25750 -985 25765 -965
rect 25785 -985 25800 -965
rect 25750 -1015 25800 -985
rect 25750 -1035 25765 -1015
rect 25785 -1035 25800 -1015
rect 25750 -1065 25800 -1035
rect 25750 -1085 25765 -1065
rect 25785 -1085 25800 -1065
rect 25750 -1115 25800 -1085
rect 25750 -1135 25765 -1115
rect 25785 -1135 25800 -1115
rect 25750 -1165 25800 -1135
rect 25750 -1185 25765 -1165
rect 25785 -1185 25800 -1165
rect 25750 -1215 25800 -1185
rect 25750 -1235 25765 -1215
rect 25785 -1235 25800 -1215
rect 25750 -1265 25800 -1235
rect 25750 -1285 25765 -1265
rect 25785 -1285 25800 -1265
rect 25750 -1315 25800 -1285
rect 25750 -1335 25765 -1315
rect 25785 -1335 25800 -1315
rect 25750 -1365 25800 -1335
rect 25750 -1385 25765 -1365
rect 25785 -1385 25800 -1365
rect 25750 -1415 25800 -1385
rect 25750 -1435 25765 -1415
rect 25785 -1435 25800 -1415
rect 25750 -1465 25800 -1435
rect 25750 -1485 25765 -1465
rect 25785 -1485 25800 -1465
rect 25750 -1515 25800 -1485
rect 25750 -1535 25765 -1515
rect 25785 -1535 25800 -1515
rect 25750 -1565 25800 -1535
rect 25750 -1585 25765 -1565
rect 25785 -1585 25800 -1565
rect 25750 -1615 25800 -1585
rect 25750 -1635 25765 -1615
rect 25785 -1635 25800 -1615
rect 25750 -1650 25800 -1635
rect 25900 -1650 25950 -950
rect 26050 -1650 26100 -950
rect 26200 -1650 26250 -950
rect 26350 -1650 26400 -950
rect 26500 -1650 26550 -950
rect 26650 -965 26700 -950
rect 26650 -985 26665 -965
rect 26685 -985 26700 -965
rect 26650 -1015 26700 -985
rect 26650 -1035 26665 -1015
rect 26685 -1035 26700 -1015
rect 26650 -1065 26700 -1035
rect 26650 -1085 26665 -1065
rect 26685 -1085 26700 -1065
rect 26650 -1115 26700 -1085
rect 26650 -1135 26665 -1115
rect 26685 -1135 26700 -1115
rect 26650 -1165 26700 -1135
rect 26650 -1185 26665 -1165
rect 26685 -1185 26700 -1165
rect 26650 -1215 26700 -1185
rect 26650 -1235 26665 -1215
rect 26685 -1235 26700 -1215
rect 26650 -1265 26700 -1235
rect 26650 -1285 26665 -1265
rect 26685 -1285 26700 -1265
rect 26650 -1315 26700 -1285
rect 26650 -1335 26665 -1315
rect 26685 -1335 26700 -1315
rect 26650 -1365 26700 -1335
rect 26650 -1385 26665 -1365
rect 26685 -1385 26700 -1365
rect 26650 -1415 26700 -1385
rect 26650 -1435 26665 -1415
rect 26685 -1435 26700 -1415
rect 26650 -1465 26700 -1435
rect 26650 -1485 26665 -1465
rect 26685 -1485 26700 -1465
rect 26650 -1515 26700 -1485
rect 26650 -1535 26665 -1515
rect 26685 -1535 26700 -1515
rect 26650 -1565 26700 -1535
rect 26650 -1585 26665 -1565
rect 26685 -1585 26700 -1565
rect 26650 -1615 26700 -1585
rect 26650 -1635 26665 -1615
rect 26685 -1635 26700 -1615
rect 26650 -1650 26700 -1635
rect 26800 -1650 26850 -950
rect 26950 -1650 27000 -950
rect 27100 -1650 27150 -950
rect 27250 -1650 27300 -950
rect 27400 -1650 27450 -950
rect 27550 -965 27600 -950
rect 27550 -985 27565 -965
rect 27585 -985 27600 -965
rect 27550 -1015 27600 -985
rect 27550 -1035 27565 -1015
rect 27585 -1035 27600 -1015
rect 27550 -1065 27600 -1035
rect 27550 -1085 27565 -1065
rect 27585 -1085 27600 -1065
rect 27550 -1115 27600 -1085
rect 27550 -1135 27565 -1115
rect 27585 -1135 27600 -1115
rect 27550 -1165 27600 -1135
rect 27550 -1185 27565 -1165
rect 27585 -1185 27600 -1165
rect 27550 -1215 27600 -1185
rect 27550 -1235 27565 -1215
rect 27585 -1235 27600 -1215
rect 27550 -1265 27600 -1235
rect 27550 -1285 27565 -1265
rect 27585 -1285 27600 -1265
rect 27550 -1315 27600 -1285
rect 27550 -1335 27565 -1315
rect 27585 -1335 27600 -1315
rect 27550 -1365 27600 -1335
rect 27550 -1385 27565 -1365
rect 27585 -1385 27600 -1365
rect 27550 -1415 27600 -1385
rect 27550 -1435 27565 -1415
rect 27585 -1435 27600 -1415
rect 27550 -1465 27600 -1435
rect 27550 -1485 27565 -1465
rect 27585 -1485 27600 -1465
rect 27550 -1515 27600 -1485
rect 27550 -1535 27565 -1515
rect 27585 -1535 27600 -1515
rect 27550 -1565 27600 -1535
rect 27550 -1585 27565 -1565
rect 27585 -1585 27600 -1565
rect 27550 -1615 27600 -1585
rect 27550 -1635 27565 -1615
rect 27585 -1635 27600 -1615
rect 27550 -1650 27600 -1635
rect 27700 -1650 27750 -950
rect 27850 -1650 27900 -950
rect 28000 -1650 28050 -950
rect 28150 -1650 28200 -950
rect 28300 -1650 28350 -950
rect 28450 -1650 28500 -950
rect 28600 -1650 28650 -950
rect 28750 -965 28800 -950
rect 28750 -985 28765 -965
rect 28785 -985 28800 -965
rect 28750 -1015 28800 -985
rect 28750 -1035 28765 -1015
rect 28785 -1035 28800 -1015
rect 28750 -1065 28800 -1035
rect 28750 -1085 28765 -1065
rect 28785 -1085 28800 -1065
rect 28750 -1115 28800 -1085
rect 28750 -1135 28765 -1115
rect 28785 -1135 28800 -1115
rect 28750 -1165 28800 -1135
rect 28750 -1185 28765 -1165
rect 28785 -1185 28800 -1165
rect 28750 -1215 28800 -1185
rect 28750 -1235 28765 -1215
rect 28785 -1235 28800 -1215
rect 28750 -1265 28800 -1235
rect 28750 -1285 28765 -1265
rect 28785 -1285 28800 -1265
rect 28750 -1315 28800 -1285
rect 28750 -1335 28765 -1315
rect 28785 -1335 28800 -1315
rect 28750 -1365 28800 -1335
rect 28750 -1385 28765 -1365
rect 28785 -1385 28800 -1365
rect 28750 -1415 28800 -1385
rect 28750 -1435 28765 -1415
rect 28785 -1435 28800 -1415
rect 28750 -1465 28800 -1435
rect 28750 -1485 28765 -1465
rect 28785 -1485 28800 -1465
rect 28750 -1515 28800 -1485
rect 28750 -1535 28765 -1515
rect 28785 -1535 28800 -1515
rect 28750 -1565 28800 -1535
rect 28750 -1585 28765 -1565
rect 28785 -1585 28800 -1565
rect 28750 -1615 28800 -1585
rect 28750 -1635 28765 -1615
rect 28785 -1635 28800 -1615
rect 28750 -1650 28800 -1635
<< mvpdiff >>
rect -650 5485 -600 5500
rect -650 5465 -635 5485
rect -615 5465 -600 5485
rect -650 5435 -600 5465
rect -650 5415 -635 5435
rect -615 5415 -600 5435
rect -650 5385 -600 5415
rect -650 5365 -635 5385
rect -615 5365 -600 5385
rect -650 5335 -600 5365
rect -650 5315 -635 5335
rect -615 5315 -600 5335
rect -650 5285 -600 5315
rect -650 5265 -635 5285
rect -615 5265 -600 5285
rect -650 5235 -600 5265
rect -650 5215 -635 5235
rect -615 5215 -600 5235
rect -650 5185 -600 5215
rect -650 5165 -635 5185
rect -615 5165 -600 5185
rect -650 5135 -600 5165
rect -650 5115 -635 5135
rect -615 5115 -600 5135
rect -650 5085 -600 5115
rect -650 5065 -635 5085
rect -615 5065 -600 5085
rect -650 5035 -600 5065
rect -650 5015 -635 5035
rect -615 5015 -600 5035
rect -650 5000 -600 5015
rect -500 5485 -450 5500
rect -500 5465 -485 5485
rect -465 5465 -450 5485
rect -500 5435 -450 5465
rect -500 5415 -485 5435
rect -465 5415 -450 5435
rect -500 5385 -450 5415
rect -500 5365 -485 5385
rect -465 5365 -450 5385
rect -500 5335 -450 5365
rect -500 5315 -485 5335
rect -465 5315 -450 5335
rect -500 5285 -450 5315
rect -500 5265 -485 5285
rect -465 5265 -450 5285
rect -500 5235 -450 5265
rect -500 5215 -485 5235
rect -465 5215 -450 5235
rect -500 5185 -450 5215
rect -500 5165 -485 5185
rect -465 5165 -450 5185
rect -500 5135 -450 5165
rect -500 5115 -485 5135
rect -465 5115 -450 5135
rect -500 5085 -450 5115
rect -500 5065 -485 5085
rect -465 5065 -450 5085
rect -500 5035 -450 5065
rect -500 5015 -485 5035
rect -465 5015 -450 5035
rect -500 5000 -450 5015
rect -350 5485 -300 5500
rect -350 5465 -335 5485
rect -315 5465 -300 5485
rect -350 5435 -300 5465
rect -350 5415 -335 5435
rect -315 5415 -300 5435
rect -350 5385 -300 5415
rect -350 5365 -335 5385
rect -315 5365 -300 5385
rect -350 5335 -300 5365
rect -350 5315 -335 5335
rect -315 5315 -300 5335
rect -350 5285 -300 5315
rect -350 5265 -335 5285
rect -315 5265 -300 5285
rect -350 5235 -300 5265
rect -350 5215 -335 5235
rect -315 5215 -300 5235
rect -350 5185 -300 5215
rect -350 5165 -335 5185
rect -315 5165 -300 5185
rect -350 5135 -300 5165
rect -350 5115 -335 5135
rect -315 5115 -300 5135
rect -350 5085 -300 5115
rect -350 5065 -335 5085
rect -315 5065 -300 5085
rect -350 5035 -300 5065
rect -350 5015 -335 5035
rect -315 5015 -300 5035
rect -350 5000 -300 5015
rect -200 5485 -150 5500
rect -200 5465 -185 5485
rect -165 5465 -150 5485
rect -200 5435 -150 5465
rect -200 5415 -185 5435
rect -165 5415 -150 5435
rect -200 5385 -150 5415
rect -200 5365 -185 5385
rect -165 5365 -150 5385
rect -200 5335 -150 5365
rect -200 5315 -185 5335
rect -165 5315 -150 5335
rect -200 5285 -150 5315
rect -200 5265 -185 5285
rect -165 5265 -150 5285
rect -200 5235 -150 5265
rect -200 5215 -185 5235
rect -165 5215 -150 5235
rect -200 5185 -150 5215
rect -200 5165 -185 5185
rect -165 5165 -150 5185
rect -200 5135 -150 5165
rect -200 5115 -185 5135
rect -165 5115 -150 5135
rect -200 5085 -150 5115
rect -200 5065 -185 5085
rect -165 5065 -150 5085
rect -200 5035 -150 5065
rect -200 5015 -185 5035
rect -165 5015 -150 5035
rect -200 5000 -150 5015
rect -50 5485 0 5500
rect -50 5465 -35 5485
rect -15 5465 0 5485
rect -50 5435 0 5465
rect -50 5415 -35 5435
rect -15 5415 0 5435
rect -50 5385 0 5415
rect -50 5365 -35 5385
rect -15 5365 0 5385
rect -50 5335 0 5365
rect -50 5315 -35 5335
rect -15 5315 0 5335
rect -50 5285 0 5315
rect -50 5265 -35 5285
rect -15 5265 0 5285
rect -50 5235 0 5265
rect -50 5215 -35 5235
rect -15 5215 0 5235
rect -50 5185 0 5215
rect -50 5165 -35 5185
rect -15 5165 0 5185
rect -50 5135 0 5165
rect -50 5115 -35 5135
rect -15 5115 0 5135
rect -50 5085 0 5115
rect -50 5065 -35 5085
rect -15 5065 0 5085
rect -50 5035 0 5065
rect -50 5015 -35 5035
rect -15 5015 0 5035
rect -50 5000 0 5015
rect 100 5000 150 5500
rect 250 5000 300 5500
rect 400 5000 450 5500
rect 550 5485 600 5500
rect 550 5465 565 5485
rect 585 5465 600 5485
rect 550 5435 600 5465
rect 550 5415 565 5435
rect 585 5415 600 5435
rect 550 5385 600 5415
rect 550 5365 565 5385
rect 585 5365 600 5385
rect 550 5335 600 5365
rect 550 5315 565 5335
rect 585 5315 600 5335
rect 550 5285 600 5315
rect 550 5265 565 5285
rect 585 5265 600 5285
rect 550 5235 600 5265
rect 550 5215 565 5235
rect 585 5215 600 5235
rect 550 5185 600 5215
rect 550 5165 565 5185
rect 585 5165 600 5185
rect 550 5135 600 5165
rect 550 5115 565 5135
rect 585 5115 600 5135
rect 550 5085 600 5115
rect 550 5065 565 5085
rect 585 5065 600 5085
rect 550 5035 600 5065
rect 550 5015 565 5035
rect 585 5015 600 5035
rect 550 5000 600 5015
rect 700 5485 750 5500
rect 700 5465 715 5485
rect 735 5465 750 5485
rect 700 5435 750 5465
rect 700 5415 715 5435
rect 735 5415 750 5435
rect 700 5385 750 5415
rect 700 5365 715 5385
rect 735 5365 750 5385
rect 700 5335 750 5365
rect 700 5315 715 5335
rect 735 5315 750 5335
rect 700 5285 750 5315
rect 700 5265 715 5285
rect 735 5265 750 5285
rect 700 5235 750 5265
rect 700 5215 715 5235
rect 735 5215 750 5235
rect 700 5185 750 5215
rect 700 5165 715 5185
rect 735 5165 750 5185
rect 700 5135 750 5165
rect 700 5115 715 5135
rect 735 5115 750 5135
rect 700 5085 750 5115
rect 700 5065 715 5085
rect 735 5065 750 5085
rect 700 5035 750 5065
rect 700 5015 715 5035
rect 735 5015 750 5035
rect 700 5000 750 5015
rect 850 5485 900 5500
rect 850 5465 865 5485
rect 885 5465 900 5485
rect 850 5435 900 5465
rect 850 5415 865 5435
rect 885 5415 900 5435
rect 850 5385 900 5415
rect 850 5365 865 5385
rect 885 5365 900 5385
rect 850 5335 900 5365
rect 850 5315 865 5335
rect 885 5315 900 5335
rect 850 5285 900 5315
rect 850 5265 865 5285
rect 885 5265 900 5285
rect 850 5235 900 5265
rect 850 5215 865 5235
rect 885 5215 900 5235
rect 850 5185 900 5215
rect 850 5165 865 5185
rect 885 5165 900 5185
rect 850 5135 900 5165
rect 850 5115 865 5135
rect 885 5115 900 5135
rect 850 5085 900 5115
rect 850 5065 865 5085
rect 885 5065 900 5085
rect 850 5035 900 5065
rect 850 5015 865 5035
rect 885 5015 900 5035
rect 850 5000 900 5015
rect 1000 5485 1050 5500
rect 1000 5465 1015 5485
rect 1035 5465 1050 5485
rect 1000 5435 1050 5465
rect 1000 5415 1015 5435
rect 1035 5415 1050 5435
rect 1000 5385 1050 5415
rect 1000 5365 1015 5385
rect 1035 5365 1050 5385
rect 1000 5335 1050 5365
rect 1000 5315 1015 5335
rect 1035 5315 1050 5335
rect 1000 5285 1050 5315
rect 1000 5265 1015 5285
rect 1035 5265 1050 5285
rect 1000 5235 1050 5265
rect 1000 5215 1015 5235
rect 1035 5215 1050 5235
rect 1000 5185 1050 5215
rect 1000 5165 1015 5185
rect 1035 5165 1050 5185
rect 1000 5135 1050 5165
rect 1000 5115 1015 5135
rect 1035 5115 1050 5135
rect 1000 5085 1050 5115
rect 1000 5065 1015 5085
rect 1035 5065 1050 5085
rect 1000 5035 1050 5065
rect 1000 5015 1015 5035
rect 1035 5015 1050 5035
rect 1000 5000 1050 5015
rect 1150 5485 1200 5500
rect 1150 5465 1165 5485
rect 1185 5465 1200 5485
rect 1150 5435 1200 5465
rect 1150 5415 1165 5435
rect 1185 5415 1200 5435
rect 1150 5385 1200 5415
rect 1150 5365 1165 5385
rect 1185 5365 1200 5385
rect 1150 5335 1200 5365
rect 1150 5315 1165 5335
rect 1185 5315 1200 5335
rect 1150 5285 1200 5315
rect 1150 5265 1165 5285
rect 1185 5265 1200 5285
rect 1150 5235 1200 5265
rect 1150 5215 1165 5235
rect 1185 5215 1200 5235
rect 1150 5185 1200 5215
rect 1150 5165 1165 5185
rect 1185 5165 1200 5185
rect 1150 5135 1200 5165
rect 1150 5115 1165 5135
rect 1185 5115 1200 5135
rect 1150 5085 1200 5115
rect 1150 5065 1165 5085
rect 1185 5065 1200 5085
rect 1150 5035 1200 5065
rect 1150 5015 1165 5035
rect 1185 5015 1200 5035
rect 1150 5000 1200 5015
rect 1300 5485 1350 5500
rect 1300 5465 1315 5485
rect 1335 5465 1350 5485
rect 1300 5435 1350 5465
rect 1300 5415 1315 5435
rect 1335 5415 1350 5435
rect 1300 5385 1350 5415
rect 1300 5365 1315 5385
rect 1335 5365 1350 5385
rect 1300 5335 1350 5365
rect 1300 5315 1315 5335
rect 1335 5315 1350 5335
rect 1300 5285 1350 5315
rect 1300 5265 1315 5285
rect 1335 5265 1350 5285
rect 1300 5235 1350 5265
rect 1300 5215 1315 5235
rect 1335 5215 1350 5235
rect 1300 5185 1350 5215
rect 1300 5165 1315 5185
rect 1335 5165 1350 5185
rect 1300 5135 1350 5165
rect 1300 5115 1315 5135
rect 1335 5115 1350 5135
rect 1300 5085 1350 5115
rect 1300 5065 1315 5085
rect 1335 5065 1350 5085
rect 1300 5035 1350 5065
rect 1300 5015 1315 5035
rect 1335 5015 1350 5035
rect 1300 5000 1350 5015
rect 1450 5485 1500 5500
rect 1450 5465 1465 5485
rect 1485 5465 1500 5485
rect 1450 5435 1500 5465
rect 1450 5415 1465 5435
rect 1485 5415 1500 5435
rect 1450 5385 1500 5415
rect 1450 5365 1465 5385
rect 1485 5365 1500 5385
rect 1450 5335 1500 5365
rect 1450 5315 1465 5335
rect 1485 5315 1500 5335
rect 1450 5285 1500 5315
rect 1450 5265 1465 5285
rect 1485 5265 1500 5285
rect 1450 5235 1500 5265
rect 1450 5215 1465 5235
rect 1485 5215 1500 5235
rect 1450 5185 1500 5215
rect 1450 5165 1465 5185
rect 1485 5165 1500 5185
rect 1450 5135 1500 5165
rect 1450 5115 1465 5135
rect 1485 5115 1500 5135
rect 1450 5085 1500 5115
rect 1450 5065 1465 5085
rect 1485 5065 1500 5085
rect 1450 5035 1500 5065
rect 1450 5015 1465 5035
rect 1485 5015 1500 5035
rect 1450 5000 1500 5015
rect 1600 5485 1650 5500
rect 1600 5465 1615 5485
rect 1635 5465 1650 5485
rect 1600 5435 1650 5465
rect 1600 5415 1615 5435
rect 1635 5415 1650 5435
rect 1600 5385 1650 5415
rect 1600 5365 1615 5385
rect 1635 5365 1650 5385
rect 1600 5335 1650 5365
rect 1600 5315 1615 5335
rect 1635 5315 1650 5335
rect 1600 5285 1650 5315
rect 1600 5265 1615 5285
rect 1635 5265 1650 5285
rect 1600 5235 1650 5265
rect 1600 5215 1615 5235
rect 1635 5215 1650 5235
rect 1600 5185 1650 5215
rect 1600 5165 1615 5185
rect 1635 5165 1650 5185
rect 1600 5135 1650 5165
rect 1600 5115 1615 5135
rect 1635 5115 1650 5135
rect 1600 5085 1650 5115
rect 1600 5065 1615 5085
rect 1635 5065 1650 5085
rect 1600 5035 1650 5065
rect 1600 5015 1615 5035
rect 1635 5015 1650 5035
rect 1600 5000 1650 5015
rect 1750 5485 1800 5500
rect 1750 5465 1765 5485
rect 1785 5465 1800 5485
rect 1750 5435 1800 5465
rect 1750 5415 1765 5435
rect 1785 5415 1800 5435
rect 1750 5385 1800 5415
rect 1750 5365 1765 5385
rect 1785 5365 1800 5385
rect 1750 5335 1800 5365
rect 1750 5315 1765 5335
rect 1785 5315 1800 5335
rect 1750 5285 1800 5315
rect 1750 5265 1765 5285
rect 1785 5265 1800 5285
rect 1750 5235 1800 5265
rect 1750 5215 1765 5235
rect 1785 5215 1800 5235
rect 1750 5185 1800 5215
rect 1750 5165 1765 5185
rect 1785 5165 1800 5185
rect 1750 5135 1800 5165
rect 1750 5115 1765 5135
rect 1785 5115 1800 5135
rect 1750 5085 1800 5115
rect 1750 5065 1765 5085
rect 1785 5065 1800 5085
rect 1750 5035 1800 5065
rect 1750 5015 1765 5035
rect 1785 5015 1800 5035
rect 1750 5000 1800 5015
rect 1900 5485 1950 5500
rect 1900 5465 1915 5485
rect 1935 5465 1950 5485
rect 1900 5435 1950 5465
rect 1900 5415 1915 5435
rect 1935 5415 1950 5435
rect 1900 5385 1950 5415
rect 1900 5365 1915 5385
rect 1935 5365 1950 5385
rect 1900 5335 1950 5365
rect 1900 5315 1915 5335
rect 1935 5315 1950 5335
rect 1900 5285 1950 5315
rect 1900 5265 1915 5285
rect 1935 5265 1950 5285
rect 1900 5235 1950 5265
rect 1900 5215 1915 5235
rect 1935 5215 1950 5235
rect 1900 5185 1950 5215
rect 1900 5165 1915 5185
rect 1935 5165 1950 5185
rect 1900 5135 1950 5165
rect 1900 5115 1915 5135
rect 1935 5115 1950 5135
rect 1900 5085 1950 5115
rect 1900 5065 1915 5085
rect 1935 5065 1950 5085
rect 1900 5035 1950 5065
rect 1900 5015 1915 5035
rect 1935 5015 1950 5035
rect 1900 5000 1950 5015
rect 2050 5485 2100 5500
rect 2050 5465 2065 5485
rect 2085 5465 2100 5485
rect 2050 5435 2100 5465
rect 2050 5415 2065 5435
rect 2085 5415 2100 5435
rect 2050 5385 2100 5415
rect 2050 5365 2065 5385
rect 2085 5365 2100 5385
rect 2050 5335 2100 5365
rect 2050 5315 2065 5335
rect 2085 5315 2100 5335
rect 2050 5285 2100 5315
rect 2050 5265 2065 5285
rect 2085 5265 2100 5285
rect 2050 5235 2100 5265
rect 2050 5215 2065 5235
rect 2085 5215 2100 5235
rect 2050 5185 2100 5215
rect 2050 5165 2065 5185
rect 2085 5165 2100 5185
rect 2050 5135 2100 5165
rect 2050 5115 2065 5135
rect 2085 5115 2100 5135
rect 2050 5085 2100 5115
rect 2050 5065 2065 5085
rect 2085 5065 2100 5085
rect 2050 5035 2100 5065
rect 2050 5015 2065 5035
rect 2085 5015 2100 5035
rect 2050 5000 2100 5015
rect 2200 5485 2250 5500
rect 2200 5465 2215 5485
rect 2235 5465 2250 5485
rect 2200 5435 2250 5465
rect 2200 5415 2215 5435
rect 2235 5415 2250 5435
rect 2200 5385 2250 5415
rect 2200 5365 2215 5385
rect 2235 5365 2250 5385
rect 2200 5335 2250 5365
rect 2200 5315 2215 5335
rect 2235 5315 2250 5335
rect 2200 5285 2250 5315
rect 2200 5265 2215 5285
rect 2235 5265 2250 5285
rect 2200 5235 2250 5265
rect 2200 5215 2215 5235
rect 2235 5215 2250 5235
rect 2200 5185 2250 5215
rect 2200 5165 2215 5185
rect 2235 5165 2250 5185
rect 2200 5135 2250 5165
rect 2200 5115 2215 5135
rect 2235 5115 2250 5135
rect 2200 5085 2250 5115
rect 2200 5065 2215 5085
rect 2235 5065 2250 5085
rect 2200 5035 2250 5065
rect 2200 5015 2215 5035
rect 2235 5015 2250 5035
rect 2200 5000 2250 5015
rect 2350 5485 2400 5500
rect 2350 5465 2365 5485
rect 2385 5465 2400 5485
rect 2350 5435 2400 5465
rect 2350 5415 2365 5435
rect 2385 5415 2400 5435
rect 2350 5385 2400 5415
rect 2350 5365 2365 5385
rect 2385 5365 2400 5385
rect 2350 5335 2400 5365
rect 2350 5315 2365 5335
rect 2385 5315 2400 5335
rect 2350 5285 2400 5315
rect 2350 5265 2365 5285
rect 2385 5265 2400 5285
rect 2350 5235 2400 5265
rect 2350 5215 2365 5235
rect 2385 5215 2400 5235
rect 2350 5185 2400 5215
rect 2350 5165 2365 5185
rect 2385 5165 2400 5185
rect 2350 5135 2400 5165
rect 2350 5115 2365 5135
rect 2385 5115 2400 5135
rect 2350 5085 2400 5115
rect 2350 5065 2365 5085
rect 2385 5065 2400 5085
rect 2350 5035 2400 5065
rect 2350 5015 2365 5035
rect 2385 5015 2400 5035
rect 2350 5000 2400 5015
rect 2500 5485 2550 5500
rect 2500 5465 2515 5485
rect 2535 5465 2550 5485
rect 2500 5435 2550 5465
rect 2500 5415 2515 5435
rect 2535 5415 2550 5435
rect 2500 5385 2550 5415
rect 2500 5365 2515 5385
rect 2535 5365 2550 5385
rect 2500 5335 2550 5365
rect 2500 5315 2515 5335
rect 2535 5315 2550 5335
rect 2500 5285 2550 5315
rect 2500 5265 2515 5285
rect 2535 5265 2550 5285
rect 2500 5235 2550 5265
rect 2500 5215 2515 5235
rect 2535 5215 2550 5235
rect 2500 5185 2550 5215
rect 2500 5165 2515 5185
rect 2535 5165 2550 5185
rect 2500 5135 2550 5165
rect 2500 5115 2515 5135
rect 2535 5115 2550 5135
rect 2500 5085 2550 5115
rect 2500 5065 2515 5085
rect 2535 5065 2550 5085
rect 2500 5035 2550 5065
rect 2500 5015 2515 5035
rect 2535 5015 2550 5035
rect 2500 5000 2550 5015
rect 2650 5485 2700 5500
rect 2650 5465 2665 5485
rect 2685 5465 2700 5485
rect 2650 5435 2700 5465
rect 2650 5415 2665 5435
rect 2685 5415 2700 5435
rect 2650 5385 2700 5415
rect 2650 5365 2665 5385
rect 2685 5365 2700 5385
rect 2650 5335 2700 5365
rect 2650 5315 2665 5335
rect 2685 5315 2700 5335
rect 2650 5285 2700 5315
rect 2650 5265 2665 5285
rect 2685 5265 2700 5285
rect 2650 5235 2700 5265
rect 2650 5215 2665 5235
rect 2685 5215 2700 5235
rect 2650 5185 2700 5215
rect 2650 5165 2665 5185
rect 2685 5165 2700 5185
rect 2650 5135 2700 5165
rect 2650 5115 2665 5135
rect 2685 5115 2700 5135
rect 2650 5085 2700 5115
rect 2650 5065 2665 5085
rect 2685 5065 2700 5085
rect 2650 5035 2700 5065
rect 2650 5015 2665 5035
rect 2685 5015 2700 5035
rect 2650 5000 2700 5015
rect 2800 5485 2850 5500
rect 2800 5465 2815 5485
rect 2835 5465 2850 5485
rect 2800 5435 2850 5465
rect 2800 5415 2815 5435
rect 2835 5415 2850 5435
rect 2800 5385 2850 5415
rect 2800 5365 2815 5385
rect 2835 5365 2850 5385
rect 2800 5335 2850 5365
rect 2800 5315 2815 5335
rect 2835 5315 2850 5335
rect 2800 5285 2850 5315
rect 2800 5265 2815 5285
rect 2835 5265 2850 5285
rect 2800 5235 2850 5265
rect 2800 5215 2815 5235
rect 2835 5215 2850 5235
rect 2800 5185 2850 5215
rect 2800 5165 2815 5185
rect 2835 5165 2850 5185
rect 2800 5135 2850 5165
rect 2800 5115 2815 5135
rect 2835 5115 2850 5135
rect 2800 5085 2850 5115
rect 2800 5065 2815 5085
rect 2835 5065 2850 5085
rect 2800 5035 2850 5065
rect 2800 5015 2815 5035
rect 2835 5015 2850 5035
rect 2800 5000 2850 5015
rect 2950 5485 3000 5500
rect 2950 5465 2965 5485
rect 2985 5465 3000 5485
rect 2950 5435 3000 5465
rect 2950 5415 2965 5435
rect 2985 5415 3000 5435
rect 2950 5385 3000 5415
rect 2950 5365 2965 5385
rect 2985 5365 3000 5385
rect 2950 5335 3000 5365
rect 2950 5315 2965 5335
rect 2985 5315 3000 5335
rect 2950 5285 3000 5315
rect 2950 5265 2965 5285
rect 2985 5265 3000 5285
rect 2950 5235 3000 5265
rect 2950 5215 2965 5235
rect 2985 5215 3000 5235
rect 2950 5185 3000 5215
rect 2950 5165 2965 5185
rect 2985 5165 3000 5185
rect 2950 5135 3000 5165
rect 2950 5115 2965 5135
rect 2985 5115 3000 5135
rect 2950 5085 3000 5115
rect 2950 5065 2965 5085
rect 2985 5065 3000 5085
rect 2950 5035 3000 5065
rect 2950 5015 2965 5035
rect 2985 5015 3000 5035
rect 2950 5000 3000 5015
rect 3100 5485 3150 5500
rect 3100 5465 3115 5485
rect 3135 5465 3150 5485
rect 3100 5435 3150 5465
rect 3100 5415 3115 5435
rect 3135 5415 3150 5435
rect 3100 5385 3150 5415
rect 3100 5365 3115 5385
rect 3135 5365 3150 5385
rect 3100 5335 3150 5365
rect 3100 5315 3115 5335
rect 3135 5315 3150 5335
rect 3100 5285 3150 5315
rect 3100 5265 3115 5285
rect 3135 5265 3150 5285
rect 3100 5235 3150 5265
rect 3100 5215 3115 5235
rect 3135 5215 3150 5235
rect 3100 5185 3150 5215
rect 3100 5165 3115 5185
rect 3135 5165 3150 5185
rect 3100 5135 3150 5165
rect 3100 5115 3115 5135
rect 3135 5115 3150 5135
rect 3100 5085 3150 5115
rect 3100 5065 3115 5085
rect 3135 5065 3150 5085
rect 3100 5035 3150 5065
rect 3100 5015 3115 5035
rect 3135 5015 3150 5035
rect 3100 5000 3150 5015
rect 3250 5485 3300 5500
rect 3250 5465 3265 5485
rect 3285 5465 3300 5485
rect 3250 5435 3300 5465
rect 3250 5415 3265 5435
rect 3285 5415 3300 5435
rect 3250 5385 3300 5415
rect 3250 5365 3265 5385
rect 3285 5365 3300 5385
rect 3250 5335 3300 5365
rect 3250 5315 3265 5335
rect 3285 5315 3300 5335
rect 3250 5285 3300 5315
rect 3250 5265 3265 5285
rect 3285 5265 3300 5285
rect 3250 5235 3300 5265
rect 3250 5215 3265 5235
rect 3285 5215 3300 5235
rect 3250 5185 3300 5215
rect 3250 5165 3265 5185
rect 3285 5165 3300 5185
rect 3250 5135 3300 5165
rect 3250 5115 3265 5135
rect 3285 5115 3300 5135
rect 3250 5085 3300 5115
rect 3250 5065 3265 5085
rect 3285 5065 3300 5085
rect 3250 5035 3300 5065
rect 3250 5015 3265 5035
rect 3285 5015 3300 5035
rect 3250 5000 3300 5015
rect 3400 5485 3450 5500
rect 3400 5465 3415 5485
rect 3435 5465 3450 5485
rect 3400 5435 3450 5465
rect 3400 5415 3415 5435
rect 3435 5415 3450 5435
rect 3400 5385 3450 5415
rect 3400 5365 3415 5385
rect 3435 5365 3450 5385
rect 3400 5335 3450 5365
rect 3400 5315 3415 5335
rect 3435 5315 3450 5335
rect 3400 5285 3450 5315
rect 3400 5265 3415 5285
rect 3435 5265 3450 5285
rect 3400 5235 3450 5265
rect 3400 5215 3415 5235
rect 3435 5215 3450 5235
rect 3400 5185 3450 5215
rect 3400 5165 3415 5185
rect 3435 5165 3450 5185
rect 3400 5135 3450 5165
rect 3400 5115 3415 5135
rect 3435 5115 3450 5135
rect 3400 5085 3450 5115
rect 3400 5065 3415 5085
rect 3435 5065 3450 5085
rect 3400 5035 3450 5065
rect 3400 5015 3415 5035
rect 3435 5015 3450 5035
rect 3400 5000 3450 5015
rect 3550 5485 3600 5500
rect 3550 5465 3565 5485
rect 3585 5465 3600 5485
rect 3550 5435 3600 5465
rect 3550 5415 3565 5435
rect 3585 5415 3600 5435
rect 3550 5385 3600 5415
rect 3550 5365 3565 5385
rect 3585 5365 3600 5385
rect 3550 5335 3600 5365
rect 3550 5315 3565 5335
rect 3585 5315 3600 5335
rect 3550 5285 3600 5315
rect 3550 5265 3565 5285
rect 3585 5265 3600 5285
rect 3550 5235 3600 5265
rect 3550 5215 3565 5235
rect 3585 5215 3600 5235
rect 3550 5185 3600 5215
rect 3550 5165 3565 5185
rect 3585 5165 3600 5185
rect 3550 5135 3600 5165
rect 3550 5115 3565 5135
rect 3585 5115 3600 5135
rect 3550 5085 3600 5115
rect 3550 5065 3565 5085
rect 3585 5065 3600 5085
rect 3550 5035 3600 5065
rect 3550 5015 3565 5035
rect 3585 5015 3600 5035
rect 3550 5000 3600 5015
rect 3700 5000 3750 5500
rect 3850 5000 3900 5500
rect 4000 5000 4050 5500
rect 4150 5485 4200 5500
rect 4150 5465 4165 5485
rect 4185 5465 4200 5485
rect 4150 5435 4200 5465
rect 4150 5415 4165 5435
rect 4185 5415 4200 5435
rect 4150 5385 4200 5415
rect 4150 5365 4165 5385
rect 4185 5365 4200 5385
rect 4150 5335 4200 5365
rect 4150 5315 4165 5335
rect 4185 5315 4200 5335
rect 4150 5285 4200 5315
rect 4150 5265 4165 5285
rect 4185 5265 4200 5285
rect 4150 5235 4200 5265
rect 4150 5215 4165 5235
rect 4185 5215 4200 5235
rect 4150 5185 4200 5215
rect 4150 5165 4165 5185
rect 4185 5165 4200 5185
rect 4150 5135 4200 5165
rect 4150 5115 4165 5135
rect 4185 5115 4200 5135
rect 4150 5085 4200 5115
rect 4150 5065 4165 5085
rect 4185 5065 4200 5085
rect 4150 5035 4200 5065
rect 4150 5015 4165 5035
rect 4185 5015 4200 5035
rect 4150 5000 4200 5015
rect 4300 5000 4350 5500
rect 4450 5000 4500 5500
rect 4600 5000 4650 5500
rect 4750 5485 4800 5500
rect 4750 5465 4765 5485
rect 4785 5465 4800 5485
rect 4750 5435 4800 5465
rect 4750 5415 4765 5435
rect 4785 5415 4800 5435
rect 4750 5385 4800 5415
rect 4750 5365 4765 5385
rect 4785 5365 4800 5385
rect 4750 5335 4800 5365
rect 4750 5315 4765 5335
rect 4785 5315 4800 5335
rect 4750 5285 4800 5315
rect 4750 5265 4765 5285
rect 4785 5265 4800 5285
rect 4750 5235 4800 5265
rect 4750 5215 4765 5235
rect 4785 5215 4800 5235
rect 4750 5185 4800 5215
rect 4750 5165 4765 5185
rect 4785 5165 4800 5185
rect 4750 5135 4800 5165
rect 4750 5115 4765 5135
rect 4785 5115 4800 5135
rect 4750 5085 4800 5115
rect 4750 5065 4765 5085
rect 4785 5065 4800 5085
rect 4750 5035 4800 5065
rect 4750 5015 4765 5035
rect 4785 5015 4800 5035
rect 4750 5000 4800 5015
rect 4900 5485 4950 5500
rect 4900 5465 4915 5485
rect 4935 5465 4950 5485
rect 4900 5435 4950 5465
rect 4900 5415 4915 5435
rect 4935 5415 4950 5435
rect 4900 5385 4950 5415
rect 4900 5365 4915 5385
rect 4935 5365 4950 5385
rect 4900 5335 4950 5365
rect 4900 5315 4915 5335
rect 4935 5315 4950 5335
rect 4900 5285 4950 5315
rect 4900 5265 4915 5285
rect 4935 5265 4950 5285
rect 4900 5235 4950 5265
rect 4900 5215 4915 5235
rect 4935 5215 4950 5235
rect 4900 5185 4950 5215
rect 4900 5165 4915 5185
rect 4935 5165 4950 5185
rect 4900 5135 4950 5165
rect 4900 5115 4915 5135
rect 4935 5115 4950 5135
rect 4900 5085 4950 5115
rect 4900 5065 4915 5085
rect 4935 5065 4950 5085
rect 4900 5035 4950 5065
rect 4900 5015 4915 5035
rect 4935 5015 4950 5035
rect 4900 5000 4950 5015
rect 5050 5485 5100 5500
rect 5050 5465 5065 5485
rect 5085 5465 5100 5485
rect 5050 5435 5100 5465
rect 5050 5415 5065 5435
rect 5085 5415 5100 5435
rect 5050 5385 5100 5415
rect 5050 5365 5065 5385
rect 5085 5365 5100 5385
rect 5050 5335 5100 5365
rect 5050 5315 5065 5335
rect 5085 5315 5100 5335
rect 5050 5285 5100 5315
rect 5050 5265 5065 5285
rect 5085 5265 5100 5285
rect 5050 5235 5100 5265
rect 5050 5215 5065 5235
rect 5085 5215 5100 5235
rect 5050 5185 5100 5215
rect 5050 5165 5065 5185
rect 5085 5165 5100 5185
rect 5050 5135 5100 5165
rect 5050 5115 5065 5135
rect 5085 5115 5100 5135
rect 5050 5085 5100 5115
rect 5050 5065 5065 5085
rect 5085 5065 5100 5085
rect 5050 5035 5100 5065
rect 5050 5015 5065 5035
rect 5085 5015 5100 5035
rect 5050 5000 5100 5015
rect 5200 5485 5250 5500
rect 5200 5465 5215 5485
rect 5235 5465 5250 5485
rect 5200 5435 5250 5465
rect 5200 5415 5215 5435
rect 5235 5415 5250 5435
rect 5200 5385 5250 5415
rect 5200 5365 5215 5385
rect 5235 5365 5250 5385
rect 5200 5335 5250 5365
rect 5200 5315 5215 5335
rect 5235 5315 5250 5335
rect 5200 5285 5250 5315
rect 5200 5265 5215 5285
rect 5235 5265 5250 5285
rect 5200 5235 5250 5265
rect 5200 5215 5215 5235
rect 5235 5215 5250 5235
rect 5200 5185 5250 5215
rect 5200 5165 5215 5185
rect 5235 5165 5250 5185
rect 5200 5135 5250 5165
rect 5200 5115 5215 5135
rect 5235 5115 5250 5135
rect 5200 5085 5250 5115
rect 5200 5065 5215 5085
rect 5235 5065 5250 5085
rect 5200 5035 5250 5065
rect 5200 5015 5215 5035
rect 5235 5015 5250 5035
rect 5200 5000 5250 5015
rect 5350 5485 5400 5500
rect 5350 5465 5365 5485
rect 5385 5465 5400 5485
rect 5350 5435 5400 5465
rect 5350 5415 5365 5435
rect 5385 5415 5400 5435
rect 5350 5385 5400 5415
rect 5350 5365 5365 5385
rect 5385 5365 5400 5385
rect 5350 5335 5400 5365
rect 5350 5315 5365 5335
rect 5385 5315 5400 5335
rect 5350 5285 5400 5315
rect 5350 5265 5365 5285
rect 5385 5265 5400 5285
rect 5350 5235 5400 5265
rect 5350 5215 5365 5235
rect 5385 5215 5400 5235
rect 5350 5185 5400 5215
rect 5350 5165 5365 5185
rect 5385 5165 5400 5185
rect 5350 5135 5400 5165
rect 5350 5115 5365 5135
rect 5385 5115 5400 5135
rect 5350 5085 5400 5115
rect 5350 5065 5365 5085
rect 5385 5065 5400 5085
rect 5350 5035 5400 5065
rect 5350 5015 5365 5035
rect 5385 5015 5400 5035
rect 5350 5000 5400 5015
rect 5500 5485 5550 5500
rect 5500 5465 5515 5485
rect 5535 5465 5550 5485
rect 5500 5435 5550 5465
rect 5500 5415 5515 5435
rect 5535 5415 5550 5435
rect 5500 5385 5550 5415
rect 5500 5365 5515 5385
rect 5535 5365 5550 5385
rect 5500 5335 5550 5365
rect 5500 5315 5515 5335
rect 5535 5315 5550 5335
rect 5500 5285 5550 5315
rect 5500 5265 5515 5285
rect 5535 5265 5550 5285
rect 5500 5235 5550 5265
rect 5500 5215 5515 5235
rect 5535 5215 5550 5235
rect 5500 5185 5550 5215
rect 5500 5165 5515 5185
rect 5535 5165 5550 5185
rect 5500 5135 5550 5165
rect 5500 5115 5515 5135
rect 5535 5115 5550 5135
rect 5500 5085 5550 5115
rect 5500 5065 5515 5085
rect 5535 5065 5550 5085
rect 5500 5035 5550 5065
rect 5500 5015 5515 5035
rect 5535 5015 5550 5035
rect 5500 5000 5550 5015
rect 5650 5485 5700 5500
rect 5650 5465 5665 5485
rect 5685 5465 5700 5485
rect 5650 5435 5700 5465
rect 5650 5415 5665 5435
rect 5685 5415 5700 5435
rect 5650 5385 5700 5415
rect 5650 5365 5665 5385
rect 5685 5365 5700 5385
rect 5650 5335 5700 5365
rect 5650 5315 5665 5335
rect 5685 5315 5700 5335
rect 5650 5285 5700 5315
rect 5650 5265 5665 5285
rect 5685 5265 5700 5285
rect 5650 5235 5700 5265
rect 5650 5215 5665 5235
rect 5685 5215 5700 5235
rect 5650 5185 5700 5215
rect 5650 5165 5665 5185
rect 5685 5165 5700 5185
rect 5650 5135 5700 5165
rect 5650 5115 5665 5135
rect 5685 5115 5700 5135
rect 5650 5085 5700 5115
rect 5650 5065 5665 5085
rect 5685 5065 5700 5085
rect 5650 5035 5700 5065
rect 5650 5015 5665 5035
rect 5685 5015 5700 5035
rect 5650 5000 5700 5015
rect 5800 5485 5850 5500
rect 5800 5465 5815 5485
rect 5835 5465 5850 5485
rect 5800 5435 5850 5465
rect 5800 5415 5815 5435
rect 5835 5415 5850 5435
rect 5800 5385 5850 5415
rect 5800 5365 5815 5385
rect 5835 5365 5850 5385
rect 5800 5335 5850 5365
rect 5800 5315 5815 5335
rect 5835 5315 5850 5335
rect 5800 5285 5850 5315
rect 5800 5265 5815 5285
rect 5835 5265 5850 5285
rect 5800 5235 5850 5265
rect 5800 5215 5815 5235
rect 5835 5215 5850 5235
rect 5800 5185 5850 5215
rect 5800 5165 5815 5185
rect 5835 5165 5850 5185
rect 5800 5135 5850 5165
rect 5800 5115 5815 5135
rect 5835 5115 5850 5135
rect 5800 5085 5850 5115
rect 5800 5065 5815 5085
rect 5835 5065 5850 5085
rect 5800 5035 5850 5065
rect 5800 5015 5815 5035
rect 5835 5015 5850 5035
rect 5800 5000 5850 5015
rect 5950 5485 6000 5500
rect 5950 5465 5965 5485
rect 5985 5465 6000 5485
rect 5950 5435 6000 5465
rect 5950 5415 5965 5435
rect 5985 5415 6000 5435
rect 5950 5385 6000 5415
rect 5950 5365 5965 5385
rect 5985 5365 6000 5385
rect 5950 5335 6000 5365
rect 5950 5315 5965 5335
rect 5985 5315 6000 5335
rect 5950 5285 6000 5315
rect 5950 5265 5965 5285
rect 5985 5265 6000 5285
rect 5950 5235 6000 5265
rect 5950 5215 5965 5235
rect 5985 5215 6000 5235
rect 5950 5185 6000 5215
rect 5950 5165 5965 5185
rect 5985 5165 6000 5185
rect 5950 5135 6000 5165
rect 5950 5115 5965 5135
rect 5985 5115 6000 5135
rect 5950 5085 6000 5115
rect 5950 5065 5965 5085
rect 5985 5065 6000 5085
rect 5950 5035 6000 5065
rect 5950 5015 5965 5035
rect 5985 5015 6000 5035
rect 5950 5000 6000 5015
rect 6100 5485 6150 5500
rect 6100 5465 6115 5485
rect 6135 5465 6150 5485
rect 6100 5435 6150 5465
rect 6100 5415 6115 5435
rect 6135 5415 6150 5435
rect 6100 5385 6150 5415
rect 6100 5365 6115 5385
rect 6135 5365 6150 5385
rect 6100 5335 6150 5365
rect 6100 5315 6115 5335
rect 6135 5315 6150 5335
rect 6100 5285 6150 5315
rect 6100 5265 6115 5285
rect 6135 5265 6150 5285
rect 6100 5235 6150 5265
rect 6100 5215 6115 5235
rect 6135 5215 6150 5235
rect 6100 5185 6150 5215
rect 6100 5165 6115 5185
rect 6135 5165 6150 5185
rect 6100 5135 6150 5165
rect 6100 5115 6115 5135
rect 6135 5115 6150 5135
rect 6100 5085 6150 5115
rect 6100 5065 6115 5085
rect 6135 5065 6150 5085
rect 6100 5035 6150 5065
rect 6100 5015 6115 5035
rect 6135 5015 6150 5035
rect 6100 5000 6150 5015
rect 6250 5485 6300 5500
rect 6250 5465 6265 5485
rect 6285 5465 6300 5485
rect 6250 5435 6300 5465
rect 6250 5415 6265 5435
rect 6285 5415 6300 5435
rect 6250 5385 6300 5415
rect 6250 5365 6265 5385
rect 6285 5365 6300 5385
rect 6250 5335 6300 5365
rect 6250 5315 6265 5335
rect 6285 5315 6300 5335
rect 6250 5285 6300 5315
rect 6250 5265 6265 5285
rect 6285 5265 6300 5285
rect 6250 5235 6300 5265
rect 6250 5215 6265 5235
rect 6285 5215 6300 5235
rect 6250 5185 6300 5215
rect 6250 5165 6265 5185
rect 6285 5165 6300 5185
rect 6250 5135 6300 5165
rect 6250 5115 6265 5135
rect 6285 5115 6300 5135
rect 6250 5085 6300 5115
rect 6250 5065 6265 5085
rect 6285 5065 6300 5085
rect 6250 5035 6300 5065
rect 6250 5015 6265 5035
rect 6285 5015 6300 5035
rect 6250 5000 6300 5015
rect 6400 5485 6450 5500
rect 6400 5465 6415 5485
rect 6435 5465 6450 5485
rect 6400 5435 6450 5465
rect 6400 5415 6415 5435
rect 6435 5415 6450 5435
rect 6400 5385 6450 5415
rect 6400 5365 6415 5385
rect 6435 5365 6450 5385
rect 6400 5335 6450 5365
rect 6400 5315 6415 5335
rect 6435 5315 6450 5335
rect 6400 5285 6450 5315
rect 6400 5265 6415 5285
rect 6435 5265 6450 5285
rect 6400 5235 6450 5265
rect 6400 5215 6415 5235
rect 6435 5215 6450 5235
rect 6400 5185 6450 5215
rect 6400 5165 6415 5185
rect 6435 5165 6450 5185
rect 6400 5135 6450 5165
rect 6400 5115 6415 5135
rect 6435 5115 6450 5135
rect 6400 5085 6450 5115
rect 6400 5065 6415 5085
rect 6435 5065 6450 5085
rect 6400 5035 6450 5065
rect 6400 5015 6415 5035
rect 6435 5015 6450 5035
rect 6400 5000 6450 5015
rect 6550 5485 6600 5500
rect 6550 5465 6565 5485
rect 6585 5465 6600 5485
rect 6550 5435 6600 5465
rect 6550 5415 6565 5435
rect 6585 5415 6600 5435
rect 6550 5385 6600 5415
rect 6550 5365 6565 5385
rect 6585 5365 6600 5385
rect 6550 5335 6600 5365
rect 6550 5315 6565 5335
rect 6585 5315 6600 5335
rect 6550 5285 6600 5315
rect 6550 5265 6565 5285
rect 6585 5265 6600 5285
rect 6550 5235 6600 5265
rect 6550 5215 6565 5235
rect 6585 5215 6600 5235
rect 6550 5185 6600 5215
rect 6550 5165 6565 5185
rect 6585 5165 6600 5185
rect 6550 5135 6600 5165
rect 6550 5115 6565 5135
rect 6585 5115 6600 5135
rect 6550 5085 6600 5115
rect 6550 5065 6565 5085
rect 6585 5065 6600 5085
rect 6550 5035 6600 5065
rect 6550 5015 6565 5035
rect 6585 5015 6600 5035
rect 6550 5000 6600 5015
rect 6700 5485 6750 5500
rect 6700 5465 6715 5485
rect 6735 5465 6750 5485
rect 6700 5435 6750 5465
rect 6700 5415 6715 5435
rect 6735 5415 6750 5435
rect 6700 5385 6750 5415
rect 6700 5365 6715 5385
rect 6735 5365 6750 5385
rect 6700 5335 6750 5365
rect 6700 5315 6715 5335
rect 6735 5315 6750 5335
rect 6700 5285 6750 5315
rect 6700 5265 6715 5285
rect 6735 5265 6750 5285
rect 6700 5235 6750 5265
rect 6700 5215 6715 5235
rect 6735 5215 6750 5235
rect 6700 5185 6750 5215
rect 6700 5165 6715 5185
rect 6735 5165 6750 5185
rect 6700 5135 6750 5165
rect 6700 5115 6715 5135
rect 6735 5115 6750 5135
rect 6700 5085 6750 5115
rect 6700 5065 6715 5085
rect 6735 5065 6750 5085
rect 6700 5035 6750 5065
rect 6700 5015 6715 5035
rect 6735 5015 6750 5035
rect 6700 5000 6750 5015
rect 6850 5485 6900 5500
rect 6850 5465 6865 5485
rect 6885 5465 6900 5485
rect 6850 5435 6900 5465
rect 6850 5415 6865 5435
rect 6885 5415 6900 5435
rect 6850 5385 6900 5415
rect 6850 5365 6865 5385
rect 6885 5365 6900 5385
rect 6850 5335 6900 5365
rect 6850 5315 6865 5335
rect 6885 5315 6900 5335
rect 6850 5285 6900 5315
rect 6850 5265 6865 5285
rect 6885 5265 6900 5285
rect 6850 5235 6900 5265
rect 6850 5215 6865 5235
rect 6885 5215 6900 5235
rect 6850 5185 6900 5215
rect 6850 5165 6865 5185
rect 6885 5165 6900 5185
rect 6850 5135 6900 5165
rect 6850 5115 6865 5135
rect 6885 5115 6900 5135
rect 6850 5085 6900 5115
rect 6850 5065 6865 5085
rect 6885 5065 6900 5085
rect 6850 5035 6900 5065
rect 6850 5015 6865 5035
rect 6885 5015 6900 5035
rect 6850 5000 6900 5015
rect 7000 5485 7050 5500
rect 7000 5465 7015 5485
rect 7035 5465 7050 5485
rect 7000 5435 7050 5465
rect 7000 5415 7015 5435
rect 7035 5415 7050 5435
rect 7000 5385 7050 5415
rect 7000 5365 7015 5385
rect 7035 5365 7050 5385
rect 7000 5335 7050 5365
rect 7000 5315 7015 5335
rect 7035 5315 7050 5335
rect 7000 5285 7050 5315
rect 7000 5265 7015 5285
rect 7035 5265 7050 5285
rect 7000 5235 7050 5265
rect 7000 5215 7015 5235
rect 7035 5215 7050 5235
rect 7000 5185 7050 5215
rect 7000 5165 7015 5185
rect 7035 5165 7050 5185
rect 7000 5135 7050 5165
rect 7000 5115 7015 5135
rect 7035 5115 7050 5135
rect 7000 5085 7050 5115
rect 7000 5065 7015 5085
rect 7035 5065 7050 5085
rect 7000 5035 7050 5065
rect 7000 5015 7015 5035
rect 7035 5015 7050 5035
rect 7000 5000 7050 5015
rect 7150 5485 7200 5500
rect 7150 5465 7165 5485
rect 7185 5465 7200 5485
rect 7150 5435 7200 5465
rect 7150 5415 7165 5435
rect 7185 5415 7200 5435
rect 7150 5385 7200 5415
rect 7150 5365 7165 5385
rect 7185 5365 7200 5385
rect 7150 5335 7200 5365
rect 7150 5315 7165 5335
rect 7185 5315 7200 5335
rect 7150 5285 7200 5315
rect 7150 5265 7165 5285
rect 7185 5265 7200 5285
rect 7150 5235 7200 5265
rect 7150 5215 7165 5235
rect 7185 5215 7200 5235
rect 7150 5185 7200 5215
rect 7150 5165 7165 5185
rect 7185 5165 7200 5185
rect 7150 5135 7200 5165
rect 7150 5115 7165 5135
rect 7185 5115 7200 5135
rect 7150 5085 7200 5115
rect 7150 5065 7165 5085
rect 7185 5065 7200 5085
rect 7150 5035 7200 5065
rect 7150 5015 7165 5035
rect 7185 5015 7200 5035
rect 7150 5000 7200 5015
rect 7300 5485 7350 5500
rect 7300 5465 7315 5485
rect 7335 5465 7350 5485
rect 7300 5435 7350 5465
rect 7300 5415 7315 5435
rect 7335 5415 7350 5435
rect 7300 5385 7350 5415
rect 7300 5365 7315 5385
rect 7335 5365 7350 5385
rect 7300 5335 7350 5365
rect 7300 5315 7315 5335
rect 7335 5315 7350 5335
rect 7300 5285 7350 5315
rect 7300 5265 7315 5285
rect 7335 5265 7350 5285
rect 7300 5235 7350 5265
rect 7300 5215 7315 5235
rect 7335 5215 7350 5235
rect 7300 5185 7350 5215
rect 7300 5165 7315 5185
rect 7335 5165 7350 5185
rect 7300 5135 7350 5165
rect 7300 5115 7315 5135
rect 7335 5115 7350 5135
rect 7300 5085 7350 5115
rect 7300 5065 7315 5085
rect 7335 5065 7350 5085
rect 7300 5035 7350 5065
rect 7300 5015 7315 5035
rect 7335 5015 7350 5035
rect 7300 5000 7350 5015
rect 7450 5485 7500 5500
rect 7450 5465 7465 5485
rect 7485 5465 7500 5485
rect 7450 5435 7500 5465
rect 7450 5415 7465 5435
rect 7485 5415 7500 5435
rect 7450 5385 7500 5415
rect 7450 5365 7465 5385
rect 7485 5365 7500 5385
rect 7450 5335 7500 5365
rect 7450 5315 7465 5335
rect 7485 5315 7500 5335
rect 7450 5285 7500 5315
rect 7450 5265 7465 5285
rect 7485 5265 7500 5285
rect 7450 5235 7500 5265
rect 7450 5215 7465 5235
rect 7485 5215 7500 5235
rect 7450 5185 7500 5215
rect 7450 5165 7465 5185
rect 7485 5165 7500 5185
rect 7450 5135 7500 5165
rect 7450 5115 7465 5135
rect 7485 5115 7500 5135
rect 7450 5085 7500 5115
rect 7450 5065 7465 5085
rect 7485 5065 7500 5085
rect 7450 5035 7500 5065
rect 7450 5015 7465 5035
rect 7485 5015 7500 5035
rect 7450 5000 7500 5015
rect 7600 5485 7650 5500
rect 7600 5465 7615 5485
rect 7635 5465 7650 5485
rect 7600 5435 7650 5465
rect 7600 5415 7615 5435
rect 7635 5415 7650 5435
rect 7600 5385 7650 5415
rect 7600 5365 7615 5385
rect 7635 5365 7650 5385
rect 7600 5335 7650 5365
rect 7600 5315 7615 5335
rect 7635 5315 7650 5335
rect 7600 5285 7650 5315
rect 7600 5265 7615 5285
rect 7635 5265 7650 5285
rect 7600 5235 7650 5265
rect 7600 5215 7615 5235
rect 7635 5215 7650 5235
rect 7600 5185 7650 5215
rect 7600 5165 7615 5185
rect 7635 5165 7650 5185
rect 7600 5135 7650 5165
rect 7600 5115 7615 5135
rect 7635 5115 7650 5135
rect 7600 5085 7650 5115
rect 7600 5065 7615 5085
rect 7635 5065 7650 5085
rect 7600 5035 7650 5065
rect 7600 5015 7615 5035
rect 7635 5015 7650 5035
rect 7600 5000 7650 5015
rect 7750 5485 7800 5500
rect 7750 5465 7765 5485
rect 7785 5465 7800 5485
rect 7750 5435 7800 5465
rect 7750 5415 7765 5435
rect 7785 5415 7800 5435
rect 7750 5385 7800 5415
rect 7750 5365 7765 5385
rect 7785 5365 7800 5385
rect 7750 5335 7800 5365
rect 7750 5315 7765 5335
rect 7785 5315 7800 5335
rect 7750 5285 7800 5315
rect 7750 5265 7765 5285
rect 7785 5265 7800 5285
rect 7750 5235 7800 5265
rect 7750 5215 7765 5235
rect 7785 5215 7800 5235
rect 7750 5185 7800 5215
rect 7750 5165 7765 5185
rect 7785 5165 7800 5185
rect 7750 5135 7800 5165
rect 7750 5115 7765 5135
rect 7785 5115 7800 5135
rect 7750 5085 7800 5115
rect 7750 5065 7765 5085
rect 7785 5065 7800 5085
rect 7750 5035 7800 5065
rect 7750 5015 7765 5035
rect 7785 5015 7800 5035
rect 7750 5000 7800 5015
rect 7900 5000 7950 5500
rect 8050 5000 8100 5500
rect 8200 5000 8250 5500
rect 8350 5485 8400 5500
rect 8350 5465 8365 5485
rect 8385 5465 8400 5485
rect 8350 5435 8400 5465
rect 8350 5415 8365 5435
rect 8385 5415 8400 5435
rect 8350 5385 8400 5415
rect 8350 5365 8365 5385
rect 8385 5365 8400 5385
rect 8350 5335 8400 5365
rect 8350 5315 8365 5335
rect 8385 5315 8400 5335
rect 8350 5285 8400 5315
rect 8350 5265 8365 5285
rect 8385 5265 8400 5285
rect 8350 5235 8400 5265
rect 8350 5215 8365 5235
rect 8385 5215 8400 5235
rect 8350 5185 8400 5215
rect 8350 5165 8365 5185
rect 8385 5165 8400 5185
rect 8350 5135 8400 5165
rect 8350 5115 8365 5135
rect 8385 5115 8400 5135
rect 8350 5085 8400 5115
rect 8350 5065 8365 5085
rect 8385 5065 8400 5085
rect 8350 5035 8400 5065
rect 8350 5015 8365 5035
rect 8385 5015 8400 5035
rect 8350 5000 8400 5015
rect 8500 5485 8550 5500
rect 8500 5465 8515 5485
rect 8535 5465 8550 5485
rect 8500 5435 8550 5465
rect 8500 5415 8515 5435
rect 8535 5415 8550 5435
rect 8500 5385 8550 5415
rect 8500 5365 8515 5385
rect 8535 5365 8550 5385
rect 8500 5335 8550 5365
rect 8500 5315 8515 5335
rect 8535 5315 8550 5335
rect 8500 5285 8550 5315
rect 8500 5265 8515 5285
rect 8535 5265 8550 5285
rect 8500 5235 8550 5265
rect 8500 5215 8515 5235
rect 8535 5215 8550 5235
rect 8500 5185 8550 5215
rect 8500 5165 8515 5185
rect 8535 5165 8550 5185
rect 8500 5135 8550 5165
rect 8500 5115 8515 5135
rect 8535 5115 8550 5135
rect 8500 5085 8550 5115
rect 8500 5065 8515 5085
rect 8535 5065 8550 5085
rect 8500 5035 8550 5065
rect 8500 5015 8515 5035
rect 8535 5015 8550 5035
rect 8500 5000 8550 5015
rect 8650 5485 8700 5500
rect 8650 5465 8665 5485
rect 8685 5465 8700 5485
rect 8650 5435 8700 5465
rect 8650 5415 8665 5435
rect 8685 5415 8700 5435
rect 8650 5385 8700 5415
rect 8650 5365 8665 5385
rect 8685 5365 8700 5385
rect 8650 5335 8700 5365
rect 8650 5315 8665 5335
rect 8685 5315 8700 5335
rect 8650 5285 8700 5315
rect 8650 5265 8665 5285
rect 8685 5265 8700 5285
rect 8650 5235 8700 5265
rect 8650 5215 8665 5235
rect 8685 5215 8700 5235
rect 8650 5185 8700 5215
rect 8650 5165 8665 5185
rect 8685 5165 8700 5185
rect 8650 5135 8700 5165
rect 8650 5115 8665 5135
rect 8685 5115 8700 5135
rect 8650 5085 8700 5115
rect 8650 5065 8665 5085
rect 8685 5065 8700 5085
rect 8650 5035 8700 5065
rect 8650 5015 8665 5035
rect 8685 5015 8700 5035
rect 8650 5000 8700 5015
rect 8800 5485 8850 5500
rect 8800 5465 8815 5485
rect 8835 5465 8850 5485
rect 8800 5435 8850 5465
rect 8800 5415 8815 5435
rect 8835 5415 8850 5435
rect 8800 5385 8850 5415
rect 8800 5365 8815 5385
rect 8835 5365 8850 5385
rect 8800 5335 8850 5365
rect 8800 5315 8815 5335
rect 8835 5315 8850 5335
rect 8800 5285 8850 5315
rect 8800 5265 8815 5285
rect 8835 5265 8850 5285
rect 8800 5235 8850 5265
rect 8800 5215 8815 5235
rect 8835 5215 8850 5235
rect 8800 5185 8850 5215
rect 8800 5165 8815 5185
rect 8835 5165 8850 5185
rect 8800 5135 8850 5165
rect 8800 5115 8815 5135
rect 8835 5115 8850 5135
rect 8800 5085 8850 5115
rect 8800 5065 8815 5085
rect 8835 5065 8850 5085
rect 8800 5035 8850 5065
rect 8800 5015 8815 5035
rect 8835 5015 8850 5035
rect 8800 5000 8850 5015
rect 8950 5485 9000 5500
rect 8950 5465 8965 5485
rect 8985 5465 9000 5485
rect 8950 5435 9000 5465
rect 8950 5415 8965 5435
rect 8985 5415 9000 5435
rect 8950 5385 9000 5415
rect 8950 5365 8965 5385
rect 8985 5365 9000 5385
rect 8950 5335 9000 5365
rect 8950 5315 8965 5335
rect 8985 5315 9000 5335
rect 8950 5285 9000 5315
rect 8950 5265 8965 5285
rect 8985 5265 9000 5285
rect 8950 5235 9000 5265
rect 8950 5215 8965 5235
rect 8985 5215 9000 5235
rect 8950 5185 9000 5215
rect 8950 5165 8965 5185
rect 8985 5165 9000 5185
rect 8950 5135 9000 5165
rect 8950 5115 8965 5135
rect 8985 5115 9000 5135
rect 8950 5085 9000 5115
rect 8950 5065 8965 5085
rect 8985 5065 9000 5085
rect 8950 5035 9000 5065
rect 8950 5015 8965 5035
rect 8985 5015 9000 5035
rect 8950 5000 9000 5015
rect 9100 5485 9150 5500
rect 9100 5465 9115 5485
rect 9135 5465 9150 5485
rect 9100 5435 9150 5465
rect 9100 5415 9115 5435
rect 9135 5415 9150 5435
rect 9100 5385 9150 5415
rect 9100 5365 9115 5385
rect 9135 5365 9150 5385
rect 9100 5335 9150 5365
rect 9100 5315 9115 5335
rect 9135 5315 9150 5335
rect 9100 5285 9150 5315
rect 9100 5265 9115 5285
rect 9135 5265 9150 5285
rect 9100 5235 9150 5265
rect 9100 5215 9115 5235
rect 9135 5215 9150 5235
rect 9100 5185 9150 5215
rect 9100 5165 9115 5185
rect 9135 5165 9150 5185
rect 9100 5135 9150 5165
rect 9100 5115 9115 5135
rect 9135 5115 9150 5135
rect 9100 5085 9150 5115
rect 9100 5065 9115 5085
rect 9135 5065 9150 5085
rect 9100 5035 9150 5065
rect 9100 5015 9115 5035
rect 9135 5015 9150 5035
rect 9100 5000 9150 5015
rect 9250 5485 9300 5500
rect 9250 5465 9265 5485
rect 9285 5465 9300 5485
rect 9250 5435 9300 5465
rect 9250 5415 9265 5435
rect 9285 5415 9300 5435
rect 9250 5385 9300 5415
rect 9250 5365 9265 5385
rect 9285 5365 9300 5385
rect 9250 5335 9300 5365
rect 9250 5315 9265 5335
rect 9285 5315 9300 5335
rect 9250 5285 9300 5315
rect 9250 5265 9265 5285
rect 9285 5265 9300 5285
rect 9250 5235 9300 5265
rect 9250 5215 9265 5235
rect 9285 5215 9300 5235
rect 9250 5185 9300 5215
rect 9250 5165 9265 5185
rect 9285 5165 9300 5185
rect 9250 5135 9300 5165
rect 9250 5115 9265 5135
rect 9285 5115 9300 5135
rect 9250 5085 9300 5115
rect 9250 5065 9265 5085
rect 9285 5065 9300 5085
rect 9250 5035 9300 5065
rect 9250 5015 9265 5035
rect 9285 5015 9300 5035
rect 9250 5000 9300 5015
rect 9400 5485 9450 5500
rect 9400 5465 9415 5485
rect 9435 5465 9450 5485
rect 9400 5435 9450 5465
rect 9400 5415 9415 5435
rect 9435 5415 9450 5435
rect 9400 5385 9450 5415
rect 9400 5365 9415 5385
rect 9435 5365 9450 5385
rect 9400 5335 9450 5365
rect 9400 5315 9415 5335
rect 9435 5315 9450 5335
rect 9400 5285 9450 5315
rect 9400 5265 9415 5285
rect 9435 5265 9450 5285
rect 9400 5235 9450 5265
rect 9400 5215 9415 5235
rect 9435 5215 9450 5235
rect 9400 5185 9450 5215
rect 9400 5165 9415 5185
rect 9435 5165 9450 5185
rect 9400 5135 9450 5165
rect 9400 5115 9415 5135
rect 9435 5115 9450 5135
rect 9400 5085 9450 5115
rect 9400 5065 9415 5085
rect 9435 5065 9450 5085
rect 9400 5035 9450 5065
rect 9400 5015 9415 5035
rect 9435 5015 9450 5035
rect 9400 5000 9450 5015
rect 9550 5485 9600 5500
rect 9550 5465 9565 5485
rect 9585 5465 9600 5485
rect 9550 5435 9600 5465
rect 9550 5415 9565 5435
rect 9585 5415 9600 5435
rect 9550 5385 9600 5415
rect 9550 5365 9565 5385
rect 9585 5365 9600 5385
rect 9550 5335 9600 5365
rect 9550 5315 9565 5335
rect 9585 5315 9600 5335
rect 9550 5285 9600 5315
rect 9550 5265 9565 5285
rect 9585 5265 9600 5285
rect 9550 5235 9600 5265
rect 9550 5215 9565 5235
rect 9585 5215 9600 5235
rect 9550 5185 9600 5215
rect 9550 5165 9565 5185
rect 9585 5165 9600 5185
rect 9550 5135 9600 5165
rect 9550 5115 9565 5135
rect 9585 5115 9600 5135
rect 9550 5085 9600 5115
rect 9550 5065 9565 5085
rect 9585 5065 9600 5085
rect 9550 5035 9600 5065
rect 9550 5015 9565 5035
rect 9585 5015 9600 5035
rect 9550 5000 9600 5015
rect 9700 5485 9750 5500
rect 9700 5465 9715 5485
rect 9735 5465 9750 5485
rect 9700 5435 9750 5465
rect 9700 5415 9715 5435
rect 9735 5415 9750 5435
rect 9700 5385 9750 5415
rect 9700 5365 9715 5385
rect 9735 5365 9750 5385
rect 9700 5335 9750 5365
rect 9700 5315 9715 5335
rect 9735 5315 9750 5335
rect 9700 5285 9750 5315
rect 9700 5265 9715 5285
rect 9735 5265 9750 5285
rect 9700 5235 9750 5265
rect 9700 5215 9715 5235
rect 9735 5215 9750 5235
rect 9700 5185 9750 5215
rect 9700 5165 9715 5185
rect 9735 5165 9750 5185
rect 9700 5135 9750 5165
rect 9700 5115 9715 5135
rect 9735 5115 9750 5135
rect 9700 5085 9750 5115
rect 9700 5065 9715 5085
rect 9735 5065 9750 5085
rect 9700 5035 9750 5065
rect 9700 5015 9715 5035
rect 9735 5015 9750 5035
rect 9700 5000 9750 5015
rect 9850 5485 9900 5500
rect 9850 5465 9865 5485
rect 9885 5465 9900 5485
rect 9850 5435 9900 5465
rect 9850 5415 9865 5435
rect 9885 5415 9900 5435
rect 9850 5385 9900 5415
rect 9850 5365 9865 5385
rect 9885 5365 9900 5385
rect 9850 5335 9900 5365
rect 9850 5315 9865 5335
rect 9885 5315 9900 5335
rect 9850 5285 9900 5315
rect 9850 5265 9865 5285
rect 9885 5265 9900 5285
rect 9850 5235 9900 5265
rect 9850 5215 9865 5235
rect 9885 5215 9900 5235
rect 9850 5185 9900 5215
rect 9850 5165 9865 5185
rect 9885 5165 9900 5185
rect 9850 5135 9900 5165
rect 9850 5115 9865 5135
rect 9885 5115 9900 5135
rect 9850 5085 9900 5115
rect 9850 5065 9865 5085
rect 9885 5065 9900 5085
rect 9850 5035 9900 5065
rect 9850 5015 9865 5035
rect 9885 5015 9900 5035
rect 9850 5000 9900 5015
rect 10000 5485 10050 5500
rect 10000 5465 10015 5485
rect 10035 5465 10050 5485
rect 10000 5435 10050 5465
rect 10000 5415 10015 5435
rect 10035 5415 10050 5435
rect 10000 5385 10050 5415
rect 10000 5365 10015 5385
rect 10035 5365 10050 5385
rect 10000 5335 10050 5365
rect 10000 5315 10015 5335
rect 10035 5315 10050 5335
rect 10000 5285 10050 5315
rect 10000 5265 10015 5285
rect 10035 5265 10050 5285
rect 10000 5235 10050 5265
rect 10000 5215 10015 5235
rect 10035 5215 10050 5235
rect 10000 5185 10050 5215
rect 10000 5165 10015 5185
rect 10035 5165 10050 5185
rect 10000 5135 10050 5165
rect 10000 5115 10015 5135
rect 10035 5115 10050 5135
rect 10000 5085 10050 5115
rect 10000 5065 10015 5085
rect 10035 5065 10050 5085
rect 10000 5035 10050 5065
rect 10000 5015 10015 5035
rect 10035 5015 10050 5035
rect 10000 5000 10050 5015
rect 10150 5485 10200 5500
rect 10150 5465 10165 5485
rect 10185 5465 10200 5485
rect 10150 5435 10200 5465
rect 10150 5415 10165 5435
rect 10185 5415 10200 5435
rect 10150 5385 10200 5415
rect 10150 5365 10165 5385
rect 10185 5365 10200 5385
rect 10150 5335 10200 5365
rect 10150 5315 10165 5335
rect 10185 5315 10200 5335
rect 10150 5285 10200 5315
rect 10150 5265 10165 5285
rect 10185 5265 10200 5285
rect 10150 5235 10200 5265
rect 10150 5215 10165 5235
rect 10185 5215 10200 5235
rect 10150 5185 10200 5215
rect 10150 5165 10165 5185
rect 10185 5165 10200 5185
rect 10150 5135 10200 5165
rect 10150 5115 10165 5135
rect 10185 5115 10200 5135
rect 10150 5085 10200 5115
rect 10150 5065 10165 5085
rect 10185 5065 10200 5085
rect 10150 5035 10200 5065
rect 10150 5015 10165 5035
rect 10185 5015 10200 5035
rect 10150 5000 10200 5015
rect 10300 5485 10350 5500
rect 10300 5465 10315 5485
rect 10335 5465 10350 5485
rect 10300 5435 10350 5465
rect 10300 5415 10315 5435
rect 10335 5415 10350 5435
rect 10300 5385 10350 5415
rect 10300 5365 10315 5385
rect 10335 5365 10350 5385
rect 10300 5335 10350 5365
rect 10300 5315 10315 5335
rect 10335 5315 10350 5335
rect 10300 5285 10350 5315
rect 10300 5265 10315 5285
rect 10335 5265 10350 5285
rect 10300 5235 10350 5265
rect 10300 5215 10315 5235
rect 10335 5215 10350 5235
rect 10300 5185 10350 5215
rect 10300 5165 10315 5185
rect 10335 5165 10350 5185
rect 10300 5135 10350 5165
rect 10300 5115 10315 5135
rect 10335 5115 10350 5135
rect 10300 5085 10350 5115
rect 10300 5065 10315 5085
rect 10335 5065 10350 5085
rect 10300 5035 10350 5065
rect 10300 5015 10315 5035
rect 10335 5015 10350 5035
rect 10300 5000 10350 5015
rect 10450 5485 10500 5500
rect 10450 5465 10465 5485
rect 10485 5465 10500 5485
rect 10450 5435 10500 5465
rect 10450 5415 10465 5435
rect 10485 5415 10500 5435
rect 10450 5385 10500 5415
rect 10450 5365 10465 5385
rect 10485 5365 10500 5385
rect 10450 5335 10500 5365
rect 10450 5315 10465 5335
rect 10485 5315 10500 5335
rect 10450 5285 10500 5315
rect 10450 5265 10465 5285
rect 10485 5265 10500 5285
rect 10450 5235 10500 5265
rect 10450 5215 10465 5235
rect 10485 5215 10500 5235
rect 10450 5185 10500 5215
rect 10450 5165 10465 5185
rect 10485 5165 10500 5185
rect 10450 5135 10500 5165
rect 10450 5115 10465 5135
rect 10485 5115 10500 5135
rect 10450 5085 10500 5115
rect 10450 5065 10465 5085
rect 10485 5065 10500 5085
rect 10450 5035 10500 5065
rect 10450 5015 10465 5035
rect 10485 5015 10500 5035
rect 10450 5000 10500 5015
rect 10600 5485 10650 5500
rect 10600 5465 10615 5485
rect 10635 5465 10650 5485
rect 10600 5435 10650 5465
rect 10600 5415 10615 5435
rect 10635 5415 10650 5435
rect 10600 5385 10650 5415
rect 10600 5365 10615 5385
rect 10635 5365 10650 5385
rect 10600 5335 10650 5365
rect 10600 5315 10615 5335
rect 10635 5315 10650 5335
rect 10600 5285 10650 5315
rect 10600 5265 10615 5285
rect 10635 5265 10650 5285
rect 10600 5235 10650 5265
rect 10600 5215 10615 5235
rect 10635 5215 10650 5235
rect 10600 5185 10650 5215
rect 10600 5165 10615 5185
rect 10635 5165 10650 5185
rect 10600 5135 10650 5165
rect 10600 5115 10615 5135
rect 10635 5115 10650 5135
rect 10600 5085 10650 5115
rect 10600 5065 10615 5085
rect 10635 5065 10650 5085
rect 10600 5035 10650 5065
rect 10600 5015 10615 5035
rect 10635 5015 10650 5035
rect 10600 5000 10650 5015
rect 10750 5485 10800 5500
rect 10750 5465 10765 5485
rect 10785 5465 10800 5485
rect 10750 5435 10800 5465
rect 10750 5415 10765 5435
rect 10785 5415 10800 5435
rect 10750 5385 10800 5415
rect 10750 5365 10765 5385
rect 10785 5365 10800 5385
rect 10750 5335 10800 5365
rect 10750 5315 10765 5335
rect 10785 5315 10800 5335
rect 10750 5285 10800 5315
rect 10750 5265 10765 5285
rect 10785 5265 10800 5285
rect 10750 5235 10800 5265
rect 10750 5215 10765 5235
rect 10785 5215 10800 5235
rect 10750 5185 10800 5215
rect 10750 5165 10765 5185
rect 10785 5165 10800 5185
rect 10750 5135 10800 5165
rect 10750 5115 10765 5135
rect 10785 5115 10800 5135
rect 10750 5085 10800 5115
rect 10750 5065 10765 5085
rect 10785 5065 10800 5085
rect 10750 5035 10800 5065
rect 10750 5015 10765 5035
rect 10785 5015 10800 5035
rect 10750 5000 10800 5015
rect 10900 5000 10950 5500
rect 11050 5000 11100 5500
rect 11200 5000 11250 5500
rect 11350 5485 11400 5500
rect 11350 5465 11365 5485
rect 11385 5465 11400 5485
rect 11350 5435 11400 5465
rect 11350 5415 11365 5435
rect 11385 5415 11400 5435
rect 11350 5385 11400 5415
rect 11350 5365 11365 5385
rect 11385 5365 11400 5385
rect 11350 5335 11400 5365
rect 11350 5315 11365 5335
rect 11385 5315 11400 5335
rect 11350 5285 11400 5315
rect 11350 5265 11365 5285
rect 11385 5265 11400 5285
rect 11350 5235 11400 5265
rect 11350 5215 11365 5235
rect 11385 5215 11400 5235
rect 11350 5185 11400 5215
rect 11350 5165 11365 5185
rect 11385 5165 11400 5185
rect 11350 5135 11400 5165
rect 11350 5115 11365 5135
rect 11385 5115 11400 5135
rect 11350 5085 11400 5115
rect 11350 5065 11365 5085
rect 11385 5065 11400 5085
rect 11350 5035 11400 5065
rect 11350 5015 11365 5035
rect 11385 5015 11400 5035
rect 11350 5000 11400 5015
rect 11500 5000 11550 5500
rect 11650 5000 11700 5500
rect 11800 5000 11850 5500
rect 11950 5485 12000 5500
rect 11950 5465 11965 5485
rect 11985 5465 12000 5485
rect 11950 5435 12000 5465
rect 11950 5415 11965 5435
rect 11985 5415 12000 5435
rect 11950 5385 12000 5415
rect 11950 5365 11965 5385
rect 11985 5365 12000 5385
rect 11950 5335 12000 5365
rect 11950 5315 11965 5335
rect 11985 5315 12000 5335
rect 11950 5285 12000 5315
rect 11950 5265 11965 5285
rect 11985 5265 12000 5285
rect 11950 5235 12000 5265
rect 11950 5215 11965 5235
rect 11985 5215 12000 5235
rect 11950 5185 12000 5215
rect 11950 5165 11965 5185
rect 11985 5165 12000 5185
rect 11950 5135 12000 5165
rect 11950 5115 11965 5135
rect 11985 5115 12000 5135
rect 11950 5085 12000 5115
rect 11950 5065 11965 5085
rect 11985 5065 12000 5085
rect 11950 5035 12000 5065
rect 11950 5015 11965 5035
rect 11985 5015 12000 5035
rect 11950 5000 12000 5015
rect 12100 5000 12150 5500
rect 12250 5000 12300 5500
rect 12400 5000 12450 5500
rect 12550 5485 12600 5500
rect 12550 5465 12565 5485
rect 12585 5465 12600 5485
rect 12550 5435 12600 5465
rect 12550 5415 12565 5435
rect 12585 5415 12600 5435
rect 12550 5385 12600 5415
rect 12550 5365 12565 5385
rect 12585 5365 12600 5385
rect 12550 5335 12600 5365
rect 12550 5315 12565 5335
rect 12585 5315 12600 5335
rect 12550 5285 12600 5315
rect 12550 5265 12565 5285
rect 12585 5265 12600 5285
rect 12550 5235 12600 5265
rect 12550 5215 12565 5235
rect 12585 5215 12600 5235
rect 12550 5185 12600 5215
rect 12550 5165 12565 5185
rect 12585 5165 12600 5185
rect 12550 5135 12600 5165
rect 12550 5115 12565 5135
rect 12585 5115 12600 5135
rect 12550 5085 12600 5115
rect 12550 5065 12565 5085
rect 12585 5065 12600 5085
rect 12550 5035 12600 5065
rect 12550 5015 12565 5035
rect 12585 5015 12600 5035
rect 12550 5000 12600 5015
rect 12700 5000 12750 5500
rect 12850 5000 12900 5500
rect 13000 5000 13050 5500
rect 13150 5485 13200 5500
rect 13150 5465 13165 5485
rect 13185 5465 13200 5485
rect 13150 5435 13200 5465
rect 13150 5415 13165 5435
rect 13185 5415 13200 5435
rect 13150 5385 13200 5415
rect 13150 5365 13165 5385
rect 13185 5365 13200 5385
rect 13150 5335 13200 5365
rect 13150 5315 13165 5335
rect 13185 5315 13200 5335
rect 13150 5285 13200 5315
rect 13150 5265 13165 5285
rect 13185 5265 13200 5285
rect 13150 5235 13200 5265
rect 13150 5215 13165 5235
rect 13185 5215 13200 5235
rect 13150 5185 13200 5215
rect 13150 5165 13165 5185
rect 13185 5165 13200 5185
rect 13150 5135 13200 5165
rect 13150 5115 13165 5135
rect 13185 5115 13200 5135
rect 13150 5085 13200 5115
rect 13150 5065 13165 5085
rect 13185 5065 13200 5085
rect 13150 5035 13200 5065
rect 13150 5015 13165 5035
rect 13185 5015 13200 5035
rect 13150 5000 13200 5015
rect 13300 5000 13350 5500
rect 13450 5000 13500 5500
rect 13600 5000 13650 5500
rect 13750 5485 13800 5500
rect 13750 5465 13765 5485
rect 13785 5465 13800 5485
rect 13750 5435 13800 5465
rect 13750 5415 13765 5435
rect 13785 5415 13800 5435
rect 13750 5385 13800 5415
rect 13750 5365 13765 5385
rect 13785 5365 13800 5385
rect 13750 5335 13800 5365
rect 13750 5315 13765 5335
rect 13785 5315 13800 5335
rect 13750 5285 13800 5315
rect 13750 5265 13765 5285
rect 13785 5265 13800 5285
rect 13750 5235 13800 5265
rect 13750 5215 13765 5235
rect 13785 5215 13800 5235
rect 13750 5185 13800 5215
rect 13750 5165 13765 5185
rect 13785 5165 13800 5185
rect 13750 5135 13800 5165
rect 13750 5115 13765 5135
rect 13785 5115 13800 5135
rect 13750 5085 13800 5115
rect 13750 5065 13765 5085
rect 13785 5065 13800 5085
rect 13750 5035 13800 5065
rect 13750 5015 13765 5035
rect 13785 5015 13800 5035
rect 13750 5000 13800 5015
rect 13900 5000 13950 5500
rect 14050 5000 14100 5500
rect 14200 5000 14250 5500
rect 14350 5485 14400 5500
rect 14350 5465 14365 5485
rect 14385 5465 14400 5485
rect 14350 5435 14400 5465
rect 14350 5415 14365 5435
rect 14385 5415 14400 5435
rect 14350 5385 14400 5415
rect 14350 5365 14365 5385
rect 14385 5365 14400 5385
rect 14350 5335 14400 5365
rect 14350 5315 14365 5335
rect 14385 5315 14400 5335
rect 14350 5285 14400 5315
rect 14350 5265 14365 5285
rect 14385 5265 14400 5285
rect 14350 5235 14400 5265
rect 14350 5215 14365 5235
rect 14385 5215 14400 5235
rect 14350 5185 14400 5215
rect 14350 5165 14365 5185
rect 14385 5165 14400 5185
rect 14350 5135 14400 5165
rect 14350 5115 14365 5135
rect 14385 5115 14400 5135
rect 14350 5085 14400 5115
rect 14350 5065 14365 5085
rect 14385 5065 14400 5085
rect 14350 5035 14400 5065
rect 14350 5015 14365 5035
rect 14385 5015 14400 5035
rect 14350 5000 14400 5015
rect 14500 5000 14550 5500
rect 14650 5000 14700 5500
rect 14800 5000 14850 5500
rect 14950 5485 15000 5500
rect 14950 5465 14965 5485
rect 14985 5465 15000 5485
rect 14950 5435 15000 5465
rect 14950 5415 14965 5435
rect 14985 5415 15000 5435
rect 14950 5385 15000 5415
rect 14950 5365 14965 5385
rect 14985 5365 15000 5385
rect 14950 5335 15000 5365
rect 14950 5315 14965 5335
rect 14985 5315 15000 5335
rect 14950 5285 15000 5315
rect 14950 5265 14965 5285
rect 14985 5265 15000 5285
rect 14950 5235 15000 5265
rect 14950 5215 14965 5235
rect 14985 5215 15000 5235
rect 14950 5185 15000 5215
rect 14950 5165 14965 5185
rect 14985 5165 15000 5185
rect 14950 5135 15000 5165
rect 14950 5115 14965 5135
rect 14985 5115 15000 5135
rect 14950 5085 15000 5115
rect 14950 5065 14965 5085
rect 14985 5065 15000 5085
rect 14950 5035 15000 5065
rect 14950 5015 14965 5035
rect 14985 5015 15000 5035
rect 14950 5000 15000 5015
rect 15100 5000 15150 5500
rect 15250 5000 15300 5500
rect 15400 5000 15450 5500
rect 15550 5485 15600 5500
rect 15550 5465 15565 5485
rect 15585 5465 15600 5485
rect 15550 5435 15600 5465
rect 15550 5415 15565 5435
rect 15585 5415 15600 5435
rect 15550 5385 15600 5415
rect 15550 5365 15565 5385
rect 15585 5365 15600 5385
rect 15550 5335 15600 5365
rect 15550 5315 15565 5335
rect 15585 5315 15600 5335
rect 15550 5285 15600 5315
rect 15550 5265 15565 5285
rect 15585 5265 15600 5285
rect 15550 5235 15600 5265
rect 15550 5215 15565 5235
rect 15585 5215 15600 5235
rect 15550 5185 15600 5215
rect 15550 5165 15565 5185
rect 15585 5165 15600 5185
rect 15550 5135 15600 5165
rect 15550 5115 15565 5135
rect 15585 5115 15600 5135
rect 15550 5085 15600 5115
rect 15550 5065 15565 5085
rect 15585 5065 15600 5085
rect 15550 5035 15600 5065
rect 15550 5015 15565 5035
rect 15585 5015 15600 5035
rect 15550 5000 15600 5015
rect 15700 5000 15750 5500
rect 15850 5000 15900 5500
rect 16000 5000 16050 5500
rect 16150 5485 16200 5500
rect 16150 5465 16165 5485
rect 16185 5465 16200 5485
rect 16150 5435 16200 5465
rect 16150 5415 16165 5435
rect 16185 5415 16200 5435
rect 16150 5385 16200 5415
rect 16150 5365 16165 5385
rect 16185 5365 16200 5385
rect 16150 5335 16200 5365
rect 16150 5315 16165 5335
rect 16185 5315 16200 5335
rect 16150 5285 16200 5315
rect 16150 5265 16165 5285
rect 16185 5265 16200 5285
rect 16150 5235 16200 5265
rect 16150 5215 16165 5235
rect 16185 5215 16200 5235
rect 16150 5185 16200 5215
rect 16150 5165 16165 5185
rect 16185 5165 16200 5185
rect 16150 5135 16200 5165
rect 16150 5115 16165 5135
rect 16185 5115 16200 5135
rect 16150 5085 16200 5115
rect 16150 5065 16165 5085
rect 16185 5065 16200 5085
rect 16150 5035 16200 5065
rect 16150 5015 16165 5035
rect 16185 5015 16200 5035
rect 16150 5000 16200 5015
rect 16300 5485 16350 5500
rect 16300 5465 16315 5485
rect 16335 5465 16350 5485
rect 16300 5435 16350 5465
rect 16300 5415 16315 5435
rect 16335 5415 16350 5435
rect 16300 5385 16350 5415
rect 16300 5365 16315 5385
rect 16335 5365 16350 5385
rect 16300 5335 16350 5365
rect 16300 5315 16315 5335
rect 16335 5315 16350 5335
rect 16300 5285 16350 5315
rect 16300 5265 16315 5285
rect 16335 5265 16350 5285
rect 16300 5235 16350 5265
rect 16300 5215 16315 5235
rect 16335 5215 16350 5235
rect 16300 5185 16350 5215
rect 16300 5165 16315 5185
rect 16335 5165 16350 5185
rect 16300 5135 16350 5165
rect 16300 5115 16315 5135
rect 16335 5115 16350 5135
rect 16300 5085 16350 5115
rect 16300 5065 16315 5085
rect 16335 5065 16350 5085
rect 16300 5035 16350 5065
rect 16300 5015 16315 5035
rect 16335 5015 16350 5035
rect 16300 5000 16350 5015
rect 16450 5485 16500 5500
rect 16450 5465 16465 5485
rect 16485 5465 16500 5485
rect 16450 5435 16500 5465
rect 16450 5415 16465 5435
rect 16485 5415 16500 5435
rect 16450 5385 16500 5415
rect 16450 5365 16465 5385
rect 16485 5365 16500 5385
rect 16450 5335 16500 5365
rect 16450 5315 16465 5335
rect 16485 5315 16500 5335
rect 16450 5285 16500 5315
rect 16450 5265 16465 5285
rect 16485 5265 16500 5285
rect 16450 5235 16500 5265
rect 16450 5215 16465 5235
rect 16485 5215 16500 5235
rect 16450 5185 16500 5215
rect 16450 5165 16465 5185
rect 16485 5165 16500 5185
rect 16450 5135 16500 5165
rect 16450 5115 16465 5135
rect 16485 5115 16500 5135
rect 16450 5085 16500 5115
rect 16450 5065 16465 5085
rect 16485 5065 16500 5085
rect 16450 5035 16500 5065
rect 16450 5015 16465 5035
rect 16485 5015 16500 5035
rect 16450 5000 16500 5015
rect 16600 5485 16650 5500
rect 16600 5465 16615 5485
rect 16635 5465 16650 5485
rect 16600 5435 16650 5465
rect 16600 5415 16615 5435
rect 16635 5415 16650 5435
rect 16600 5385 16650 5415
rect 16600 5365 16615 5385
rect 16635 5365 16650 5385
rect 16600 5335 16650 5365
rect 16600 5315 16615 5335
rect 16635 5315 16650 5335
rect 16600 5285 16650 5315
rect 16600 5265 16615 5285
rect 16635 5265 16650 5285
rect 16600 5235 16650 5265
rect 16600 5215 16615 5235
rect 16635 5215 16650 5235
rect 16600 5185 16650 5215
rect 16600 5165 16615 5185
rect 16635 5165 16650 5185
rect 16600 5135 16650 5165
rect 16600 5115 16615 5135
rect 16635 5115 16650 5135
rect 16600 5085 16650 5115
rect 16600 5065 16615 5085
rect 16635 5065 16650 5085
rect 16600 5035 16650 5065
rect 16600 5015 16615 5035
rect 16635 5015 16650 5035
rect 16600 5000 16650 5015
rect 16750 5485 16800 5500
rect 16750 5465 16765 5485
rect 16785 5465 16800 5485
rect 16750 5435 16800 5465
rect 16750 5415 16765 5435
rect 16785 5415 16800 5435
rect 16750 5385 16800 5415
rect 16750 5365 16765 5385
rect 16785 5365 16800 5385
rect 16750 5335 16800 5365
rect 16750 5315 16765 5335
rect 16785 5315 16800 5335
rect 16750 5285 16800 5315
rect 16750 5265 16765 5285
rect 16785 5265 16800 5285
rect 16750 5235 16800 5265
rect 16750 5215 16765 5235
rect 16785 5215 16800 5235
rect 16750 5185 16800 5215
rect 16750 5165 16765 5185
rect 16785 5165 16800 5185
rect 16750 5135 16800 5165
rect 16750 5115 16765 5135
rect 16785 5115 16800 5135
rect 16750 5085 16800 5115
rect 16750 5065 16765 5085
rect 16785 5065 16800 5085
rect 16750 5035 16800 5065
rect 16750 5015 16765 5035
rect 16785 5015 16800 5035
rect 16750 5000 16800 5015
rect 16900 5485 16950 5500
rect 16900 5465 16915 5485
rect 16935 5465 16950 5485
rect 16900 5435 16950 5465
rect 16900 5415 16915 5435
rect 16935 5415 16950 5435
rect 16900 5385 16950 5415
rect 16900 5365 16915 5385
rect 16935 5365 16950 5385
rect 16900 5335 16950 5365
rect 16900 5315 16915 5335
rect 16935 5315 16950 5335
rect 16900 5285 16950 5315
rect 16900 5265 16915 5285
rect 16935 5265 16950 5285
rect 16900 5235 16950 5265
rect 16900 5215 16915 5235
rect 16935 5215 16950 5235
rect 16900 5185 16950 5215
rect 16900 5165 16915 5185
rect 16935 5165 16950 5185
rect 16900 5135 16950 5165
rect 16900 5115 16915 5135
rect 16935 5115 16950 5135
rect 16900 5085 16950 5115
rect 16900 5065 16915 5085
rect 16935 5065 16950 5085
rect 16900 5035 16950 5065
rect 16900 5015 16915 5035
rect 16935 5015 16950 5035
rect 16900 5000 16950 5015
rect 17050 5485 17100 5500
rect 17050 5465 17065 5485
rect 17085 5465 17100 5485
rect 17050 5435 17100 5465
rect 17050 5415 17065 5435
rect 17085 5415 17100 5435
rect 17050 5385 17100 5415
rect 17050 5365 17065 5385
rect 17085 5365 17100 5385
rect 17050 5335 17100 5365
rect 17050 5315 17065 5335
rect 17085 5315 17100 5335
rect 17050 5285 17100 5315
rect 17050 5265 17065 5285
rect 17085 5265 17100 5285
rect 17050 5235 17100 5265
rect 17050 5215 17065 5235
rect 17085 5215 17100 5235
rect 17050 5185 17100 5215
rect 17050 5165 17065 5185
rect 17085 5165 17100 5185
rect 17050 5135 17100 5165
rect 17050 5115 17065 5135
rect 17085 5115 17100 5135
rect 17050 5085 17100 5115
rect 17050 5065 17065 5085
rect 17085 5065 17100 5085
rect 17050 5035 17100 5065
rect 17050 5015 17065 5035
rect 17085 5015 17100 5035
rect 17050 5000 17100 5015
rect 17200 5485 17250 5500
rect 17200 5465 17215 5485
rect 17235 5465 17250 5485
rect 17200 5435 17250 5465
rect 17200 5415 17215 5435
rect 17235 5415 17250 5435
rect 17200 5385 17250 5415
rect 17200 5365 17215 5385
rect 17235 5365 17250 5385
rect 17200 5335 17250 5365
rect 17200 5315 17215 5335
rect 17235 5315 17250 5335
rect 17200 5285 17250 5315
rect 17200 5265 17215 5285
rect 17235 5265 17250 5285
rect 17200 5235 17250 5265
rect 17200 5215 17215 5235
rect 17235 5215 17250 5235
rect 17200 5185 17250 5215
rect 17200 5165 17215 5185
rect 17235 5165 17250 5185
rect 17200 5135 17250 5165
rect 17200 5115 17215 5135
rect 17235 5115 17250 5135
rect 17200 5085 17250 5115
rect 17200 5065 17215 5085
rect 17235 5065 17250 5085
rect 17200 5035 17250 5065
rect 17200 5015 17215 5035
rect 17235 5015 17250 5035
rect 17200 5000 17250 5015
rect 17350 5485 17400 5500
rect 17350 5465 17365 5485
rect 17385 5465 17400 5485
rect 17350 5435 17400 5465
rect 17350 5415 17365 5435
rect 17385 5415 17400 5435
rect 17350 5385 17400 5415
rect 17350 5365 17365 5385
rect 17385 5365 17400 5385
rect 17350 5335 17400 5365
rect 17350 5315 17365 5335
rect 17385 5315 17400 5335
rect 17350 5285 17400 5315
rect 17350 5265 17365 5285
rect 17385 5265 17400 5285
rect 17350 5235 17400 5265
rect 17350 5215 17365 5235
rect 17385 5215 17400 5235
rect 17350 5185 17400 5215
rect 17350 5165 17365 5185
rect 17385 5165 17400 5185
rect 17350 5135 17400 5165
rect 17350 5115 17365 5135
rect 17385 5115 17400 5135
rect 17350 5085 17400 5115
rect 17350 5065 17365 5085
rect 17385 5065 17400 5085
rect 17350 5035 17400 5065
rect 17350 5015 17365 5035
rect 17385 5015 17400 5035
rect 17350 5000 17400 5015
rect 17500 5000 17550 5500
rect 17650 5000 17700 5500
rect 17800 5000 17850 5500
rect 17950 5485 18000 5500
rect 17950 5465 17965 5485
rect 17985 5465 18000 5485
rect 17950 5435 18000 5465
rect 17950 5415 17965 5435
rect 17985 5415 18000 5435
rect 17950 5385 18000 5415
rect 17950 5365 17965 5385
rect 17985 5365 18000 5385
rect 17950 5335 18000 5365
rect 17950 5315 17965 5335
rect 17985 5315 18000 5335
rect 17950 5285 18000 5315
rect 17950 5265 17965 5285
rect 17985 5265 18000 5285
rect 17950 5235 18000 5265
rect 17950 5215 17965 5235
rect 17985 5215 18000 5235
rect 17950 5185 18000 5215
rect 17950 5165 17965 5185
rect 17985 5165 18000 5185
rect 17950 5135 18000 5165
rect 17950 5115 17965 5135
rect 17985 5115 18000 5135
rect 17950 5085 18000 5115
rect 17950 5065 17965 5085
rect 17985 5065 18000 5085
rect 17950 5035 18000 5065
rect 17950 5015 17965 5035
rect 17985 5015 18000 5035
rect 17950 5000 18000 5015
rect 18100 5000 18150 5500
rect 18250 5000 18300 5500
rect 18400 5000 18450 5500
rect 18550 5485 18600 5500
rect 18550 5465 18565 5485
rect 18585 5465 18600 5485
rect 18550 5435 18600 5465
rect 18550 5415 18565 5435
rect 18585 5415 18600 5435
rect 18550 5385 18600 5415
rect 18550 5365 18565 5385
rect 18585 5365 18600 5385
rect 18550 5335 18600 5365
rect 18550 5315 18565 5335
rect 18585 5315 18600 5335
rect 18550 5285 18600 5315
rect 18550 5265 18565 5285
rect 18585 5265 18600 5285
rect 18550 5235 18600 5265
rect 18550 5215 18565 5235
rect 18585 5215 18600 5235
rect 18550 5185 18600 5215
rect 18550 5165 18565 5185
rect 18585 5165 18600 5185
rect 18550 5135 18600 5165
rect 18550 5115 18565 5135
rect 18585 5115 18600 5135
rect 18550 5085 18600 5115
rect 18550 5065 18565 5085
rect 18585 5065 18600 5085
rect 18550 5035 18600 5065
rect 18550 5015 18565 5035
rect 18585 5015 18600 5035
rect 18550 5000 18600 5015
rect 18700 5485 18750 5500
rect 18700 5465 18715 5485
rect 18735 5465 18750 5485
rect 18700 5435 18750 5465
rect 18700 5415 18715 5435
rect 18735 5415 18750 5435
rect 18700 5385 18750 5415
rect 18700 5365 18715 5385
rect 18735 5365 18750 5385
rect 18700 5335 18750 5365
rect 18700 5315 18715 5335
rect 18735 5315 18750 5335
rect 18700 5285 18750 5315
rect 18700 5265 18715 5285
rect 18735 5265 18750 5285
rect 18700 5235 18750 5265
rect 18700 5215 18715 5235
rect 18735 5215 18750 5235
rect 18700 5185 18750 5215
rect 18700 5165 18715 5185
rect 18735 5165 18750 5185
rect 18700 5135 18750 5165
rect 18700 5115 18715 5135
rect 18735 5115 18750 5135
rect 18700 5085 18750 5115
rect 18700 5065 18715 5085
rect 18735 5065 18750 5085
rect 18700 5035 18750 5065
rect 18700 5015 18715 5035
rect 18735 5015 18750 5035
rect 18700 5000 18750 5015
rect 18850 5485 18900 5500
rect 18850 5465 18865 5485
rect 18885 5465 18900 5485
rect 18850 5435 18900 5465
rect 18850 5415 18865 5435
rect 18885 5415 18900 5435
rect 18850 5385 18900 5415
rect 18850 5365 18865 5385
rect 18885 5365 18900 5385
rect 18850 5335 18900 5365
rect 18850 5315 18865 5335
rect 18885 5315 18900 5335
rect 18850 5285 18900 5315
rect 18850 5265 18865 5285
rect 18885 5265 18900 5285
rect 18850 5235 18900 5265
rect 18850 5215 18865 5235
rect 18885 5215 18900 5235
rect 18850 5185 18900 5215
rect 18850 5165 18865 5185
rect 18885 5165 18900 5185
rect 18850 5135 18900 5165
rect 18850 5115 18865 5135
rect 18885 5115 18900 5135
rect 18850 5085 18900 5115
rect 18850 5065 18865 5085
rect 18885 5065 18900 5085
rect 18850 5035 18900 5065
rect 18850 5015 18865 5035
rect 18885 5015 18900 5035
rect 18850 5000 18900 5015
rect 19000 5485 19050 5500
rect 19000 5465 19015 5485
rect 19035 5465 19050 5485
rect 19000 5435 19050 5465
rect 19000 5415 19015 5435
rect 19035 5415 19050 5435
rect 19000 5385 19050 5415
rect 19000 5365 19015 5385
rect 19035 5365 19050 5385
rect 19000 5335 19050 5365
rect 19000 5315 19015 5335
rect 19035 5315 19050 5335
rect 19000 5285 19050 5315
rect 19000 5265 19015 5285
rect 19035 5265 19050 5285
rect 19000 5235 19050 5265
rect 19000 5215 19015 5235
rect 19035 5215 19050 5235
rect 19000 5185 19050 5215
rect 19000 5165 19015 5185
rect 19035 5165 19050 5185
rect 19000 5135 19050 5165
rect 19000 5115 19015 5135
rect 19035 5115 19050 5135
rect 19000 5085 19050 5115
rect 19000 5065 19015 5085
rect 19035 5065 19050 5085
rect 19000 5035 19050 5065
rect 19000 5015 19015 5035
rect 19035 5015 19050 5035
rect 19000 5000 19050 5015
rect 19150 5485 19200 5500
rect 19150 5465 19165 5485
rect 19185 5465 19200 5485
rect 19150 5435 19200 5465
rect 19150 5415 19165 5435
rect 19185 5415 19200 5435
rect 19150 5385 19200 5415
rect 19150 5365 19165 5385
rect 19185 5365 19200 5385
rect 19150 5335 19200 5365
rect 19150 5315 19165 5335
rect 19185 5315 19200 5335
rect 19150 5285 19200 5315
rect 19150 5265 19165 5285
rect 19185 5265 19200 5285
rect 19150 5235 19200 5265
rect 19150 5215 19165 5235
rect 19185 5215 19200 5235
rect 19150 5185 19200 5215
rect 19150 5165 19165 5185
rect 19185 5165 19200 5185
rect 19150 5135 19200 5165
rect 19150 5115 19165 5135
rect 19185 5115 19200 5135
rect 19150 5085 19200 5115
rect 19150 5065 19165 5085
rect 19185 5065 19200 5085
rect 19150 5035 19200 5065
rect 19150 5015 19165 5035
rect 19185 5015 19200 5035
rect 19150 5000 19200 5015
rect 19300 5485 19350 5500
rect 19300 5465 19315 5485
rect 19335 5465 19350 5485
rect 19300 5435 19350 5465
rect 19300 5415 19315 5435
rect 19335 5415 19350 5435
rect 19300 5385 19350 5415
rect 19300 5365 19315 5385
rect 19335 5365 19350 5385
rect 19300 5335 19350 5365
rect 19300 5315 19315 5335
rect 19335 5315 19350 5335
rect 19300 5285 19350 5315
rect 19300 5265 19315 5285
rect 19335 5265 19350 5285
rect 19300 5235 19350 5265
rect 19300 5215 19315 5235
rect 19335 5215 19350 5235
rect 19300 5185 19350 5215
rect 19300 5165 19315 5185
rect 19335 5165 19350 5185
rect 19300 5135 19350 5165
rect 19300 5115 19315 5135
rect 19335 5115 19350 5135
rect 19300 5085 19350 5115
rect 19300 5065 19315 5085
rect 19335 5065 19350 5085
rect 19300 5035 19350 5065
rect 19300 5015 19315 5035
rect 19335 5015 19350 5035
rect 19300 5000 19350 5015
rect 19450 5485 19500 5500
rect 19450 5465 19465 5485
rect 19485 5465 19500 5485
rect 19450 5435 19500 5465
rect 19450 5415 19465 5435
rect 19485 5415 19500 5435
rect 19450 5385 19500 5415
rect 19450 5365 19465 5385
rect 19485 5365 19500 5385
rect 19450 5335 19500 5365
rect 19450 5315 19465 5335
rect 19485 5315 19500 5335
rect 19450 5285 19500 5315
rect 19450 5265 19465 5285
rect 19485 5265 19500 5285
rect 19450 5235 19500 5265
rect 19450 5215 19465 5235
rect 19485 5215 19500 5235
rect 19450 5185 19500 5215
rect 19450 5165 19465 5185
rect 19485 5165 19500 5185
rect 19450 5135 19500 5165
rect 19450 5115 19465 5135
rect 19485 5115 19500 5135
rect 19450 5085 19500 5115
rect 19450 5065 19465 5085
rect 19485 5065 19500 5085
rect 19450 5035 19500 5065
rect 19450 5015 19465 5035
rect 19485 5015 19500 5035
rect 19450 5000 19500 5015
rect 19600 5485 19650 5500
rect 19600 5465 19615 5485
rect 19635 5465 19650 5485
rect 19600 5435 19650 5465
rect 19600 5415 19615 5435
rect 19635 5415 19650 5435
rect 19600 5385 19650 5415
rect 19600 5365 19615 5385
rect 19635 5365 19650 5385
rect 19600 5335 19650 5365
rect 19600 5315 19615 5335
rect 19635 5315 19650 5335
rect 19600 5285 19650 5315
rect 19600 5265 19615 5285
rect 19635 5265 19650 5285
rect 19600 5235 19650 5265
rect 19600 5215 19615 5235
rect 19635 5215 19650 5235
rect 19600 5185 19650 5215
rect 19600 5165 19615 5185
rect 19635 5165 19650 5185
rect 19600 5135 19650 5165
rect 19600 5115 19615 5135
rect 19635 5115 19650 5135
rect 19600 5085 19650 5115
rect 19600 5065 19615 5085
rect 19635 5065 19650 5085
rect 19600 5035 19650 5065
rect 19600 5015 19615 5035
rect 19635 5015 19650 5035
rect 19600 5000 19650 5015
rect 19750 5485 19800 5500
rect 19750 5465 19765 5485
rect 19785 5465 19800 5485
rect 19750 5435 19800 5465
rect 19750 5415 19765 5435
rect 19785 5415 19800 5435
rect 19750 5385 19800 5415
rect 19750 5365 19765 5385
rect 19785 5365 19800 5385
rect 19750 5335 19800 5365
rect 19750 5315 19765 5335
rect 19785 5315 19800 5335
rect 19750 5285 19800 5315
rect 19750 5265 19765 5285
rect 19785 5265 19800 5285
rect 19750 5235 19800 5265
rect 19750 5215 19765 5235
rect 19785 5215 19800 5235
rect 19750 5185 19800 5215
rect 19750 5165 19765 5185
rect 19785 5165 19800 5185
rect 19750 5135 19800 5165
rect 19750 5115 19765 5135
rect 19785 5115 19800 5135
rect 19750 5085 19800 5115
rect 19750 5065 19765 5085
rect 19785 5065 19800 5085
rect 19750 5035 19800 5065
rect 19750 5015 19765 5035
rect 19785 5015 19800 5035
rect 19750 5000 19800 5015
rect 19900 5000 19950 5500
rect 20050 5000 20100 5500
rect 20200 5000 20250 5500
rect 20350 5485 20400 5500
rect 20350 5465 20365 5485
rect 20385 5465 20400 5485
rect 20350 5435 20400 5465
rect 20350 5415 20365 5435
rect 20385 5415 20400 5435
rect 20350 5385 20400 5415
rect 20350 5365 20365 5385
rect 20385 5365 20400 5385
rect 20350 5335 20400 5365
rect 20350 5315 20365 5335
rect 20385 5315 20400 5335
rect 20350 5285 20400 5315
rect 20350 5265 20365 5285
rect 20385 5265 20400 5285
rect 20350 5235 20400 5265
rect 20350 5215 20365 5235
rect 20385 5215 20400 5235
rect 20350 5185 20400 5215
rect 20350 5165 20365 5185
rect 20385 5165 20400 5185
rect 20350 5135 20400 5165
rect 20350 5115 20365 5135
rect 20385 5115 20400 5135
rect 20350 5085 20400 5115
rect 20350 5065 20365 5085
rect 20385 5065 20400 5085
rect 20350 5035 20400 5065
rect 20350 5015 20365 5035
rect 20385 5015 20400 5035
rect 20350 5000 20400 5015
rect 20500 5000 20550 5500
rect 20650 5000 20700 5500
rect 20800 5000 20850 5500
rect 20950 5485 21000 5500
rect 20950 5465 20965 5485
rect 20985 5465 21000 5485
rect 20950 5435 21000 5465
rect 20950 5415 20965 5435
rect 20985 5415 21000 5435
rect 20950 5385 21000 5415
rect 20950 5365 20965 5385
rect 20985 5365 21000 5385
rect 20950 5335 21000 5365
rect 20950 5315 20965 5335
rect 20985 5315 21000 5335
rect 20950 5285 21000 5315
rect 20950 5265 20965 5285
rect 20985 5265 21000 5285
rect 20950 5235 21000 5265
rect 20950 5215 20965 5235
rect 20985 5215 21000 5235
rect 20950 5185 21000 5215
rect 20950 5165 20965 5185
rect 20985 5165 21000 5185
rect 20950 5135 21000 5165
rect 20950 5115 20965 5135
rect 20985 5115 21000 5135
rect 20950 5085 21000 5115
rect 20950 5065 20965 5085
rect 20985 5065 21000 5085
rect 20950 5035 21000 5065
rect 20950 5015 20965 5035
rect 20985 5015 21000 5035
rect 20950 5000 21000 5015
rect 21100 5000 21150 5500
rect 21250 5000 21300 5500
rect 21400 5485 21450 5500
rect 21400 5465 21415 5485
rect 21435 5465 21450 5485
rect 21400 5435 21450 5465
rect 21400 5415 21415 5435
rect 21435 5415 21450 5435
rect 21400 5385 21450 5415
rect 21400 5365 21415 5385
rect 21435 5365 21450 5385
rect 21400 5335 21450 5365
rect 21400 5315 21415 5335
rect 21435 5315 21450 5335
rect 21400 5285 21450 5315
rect 21400 5265 21415 5285
rect 21435 5265 21450 5285
rect 21400 5235 21450 5265
rect 21400 5215 21415 5235
rect 21435 5215 21450 5235
rect 21400 5185 21450 5215
rect 21400 5165 21415 5185
rect 21435 5165 21450 5185
rect 21400 5135 21450 5165
rect 21400 5115 21415 5135
rect 21435 5115 21450 5135
rect 21400 5085 21450 5115
rect 21400 5065 21415 5085
rect 21435 5065 21450 5085
rect 21400 5035 21450 5065
rect 21400 5015 21415 5035
rect 21435 5015 21450 5035
rect 21400 5000 21450 5015
rect 21550 5000 21600 5500
rect 21700 5000 21750 5500
rect 21850 5485 21900 5500
rect 21850 5465 21865 5485
rect 21885 5465 21900 5485
rect 21850 5435 21900 5465
rect 21850 5415 21865 5435
rect 21885 5415 21900 5435
rect 21850 5385 21900 5415
rect 21850 5365 21865 5385
rect 21885 5365 21900 5385
rect 21850 5335 21900 5365
rect 21850 5315 21865 5335
rect 21885 5315 21900 5335
rect 21850 5285 21900 5315
rect 21850 5265 21865 5285
rect 21885 5265 21900 5285
rect 21850 5235 21900 5265
rect 21850 5215 21865 5235
rect 21885 5215 21900 5235
rect 21850 5185 21900 5215
rect 21850 5165 21865 5185
rect 21885 5165 21900 5185
rect 21850 5135 21900 5165
rect 21850 5115 21865 5135
rect 21885 5115 21900 5135
rect 21850 5085 21900 5115
rect 21850 5065 21865 5085
rect 21885 5065 21900 5085
rect 21850 5035 21900 5065
rect 21850 5015 21865 5035
rect 21885 5015 21900 5035
rect 21850 5000 21900 5015
rect 22000 5000 22050 5500
rect 22150 5000 22200 5500
rect 22300 5000 22350 5500
rect 22450 5485 22500 5500
rect 22450 5465 22465 5485
rect 22485 5465 22500 5485
rect 22450 5435 22500 5465
rect 22450 5415 22465 5435
rect 22485 5415 22500 5435
rect 22450 5385 22500 5415
rect 22450 5365 22465 5385
rect 22485 5365 22500 5385
rect 22450 5335 22500 5365
rect 22450 5315 22465 5335
rect 22485 5315 22500 5335
rect 22450 5285 22500 5315
rect 22450 5265 22465 5285
rect 22485 5265 22500 5285
rect 22450 5235 22500 5265
rect 22450 5215 22465 5235
rect 22485 5215 22500 5235
rect 22450 5185 22500 5215
rect 22450 5165 22465 5185
rect 22485 5165 22500 5185
rect 22450 5135 22500 5165
rect 22450 5115 22465 5135
rect 22485 5115 22500 5135
rect 22450 5085 22500 5115
rect 22450 5065 22465 5085
rect 22485 5065 22500 5085
rect 22450 5035 22500 5065
rect 22450 5015 22465 5035
rect 22485 5015 22500 5035
rect 22450 5000 22500 5015
rect 22600 5000 22650 5500
rect 22750 5000 22800 5500
rect 22900 5000 22950 5500
rect 23050 5485 23100 5500
rect 23050 5465 23065 5485
rect 23085 5465 23100 5485
rect 23050 5435 23100 5465
rect 23050 5415 23065 5435
rect 23085 5415 23100 5435
rect 23050 5385 23100 5415
rect 23050 5365 23065 5385
rect 23085 5365 23100 5385
rect 23050 5335 23100 5365
rect 23050 5315 23065 5335
rect 23085 5315 23100 5335
rect 23050 5285 23100 5315
rect 23050 5265 23065 5285
rect 23085 5265 23100 5285
rect 23050 5235 23100 5265
rect 23050 5215 23065 5235
rect 23085 5215 23100 5235
rect 23050 5185 23100 5215
rect 23050 5165 23065 5185
rect 23085 5165 23100 5185
rect 23050 5135 23100 5165
rect 23050 5115 23065 5135
rect 23085 5115 23100 5135
rect 23050 5085 23100 5115
rect 23050 5065 23065 5085
rect 23085 5065 23100 5085
rect 23050 5035 23100 5065
rect 23050 5015 23065 5035
rect 23085 5015 23100 5035
rect 23050 5000 23100 5015
rect 23200 5000 23250 5500
rect 23350 5000 23400 5500
rect 23500 5485 23550 5500
rect 23500 5465 23515 5485
rect 23535 5465 23550 5485
rect 23500 5435 23550 5465
rect 23500 5415 23515 5435
rect 23535 5415 23550 5435
rect 23500 5385 23550 5415
rect 23500 5365 23515 5385
rect 23535 5365 23550 5385
rect 23500 5335 23550 5365
rect 23500 5315 23515 5335
rect 23535 5315 23550 5335
rect 23500 5285 23550 5315
rect 23500 5265 23515 5285
rect 23535 5265 23550 5285
rect 23500 5235 23550 5265
rect 23500 5215 23515 5235
rect 23535 5215 23550 5235
rect 23500 5185 23550 5215
rect 23500 5165 23515 5185
rect 23535 5165 23550 5185
rect 23500 5135 23550 5165
rect 23500 5115 23515 5135
rect 23535 5115 23550 5135
rect 23500 5085 23550 5115
rect 23500 5065 23515 5085
rect 23535 5065 23550 5085
rect 23500 5035 23550 5065
rect 23500 5015 23515 5035
rect 23535 5015 23550 5035
rect 23500 5000 23550 5015
rect 23650 5000 23700 5500
rect 23800 5000 23850 5500
rect 23950 5485 24000 5500
rect 23950 5465 23965 5485
rect 23985 5465 24000 5485
rect 23950 5435 24000 5465
rect 23950 5415 23965 5435
rect 23985 5415 24000 5435
rect 23950 5385 24000 5415
rect 23950 5365 23965 5385
rect 23985 5365 24000 5385
rect 23950 5335 24000 5365
rect 23950 5315 23965 5335
rect 23985 5315 24000 5335
rect 23950 5285 24000 5315
rect 23950 5265 23965 5285
rect 23985 5265 24000 5285
rect 23950 5235 24000 5265
rect 23950 5215 23965 5235
rect 23985 5215 24000 5235
rect 23950 5185 24000 5215
rect 23950 5165 23965 5185
rect 23985 5165 24000 5185
rect 23950 5135 24000 5165
rect 23950 5115 23965 5135
rect 23985 5115 24000 5135
rect 23950 5085 24000 5115
rect 23950 5065 23965 5085
rect 23985 5065 24000 5085
rect 23950 5035 24000 5065
rect 23950 5015 23965 5035
rect 23985 5015 24000 5035
rect 23950 5000 24000 5015
rect 24100 5000 24150 5500
rect 24250 5000 24300 5500
rect 24400 5000 24450 5500
rect 24550 5485 24600 5500
rect 24550 5465 24565 5485
rect 24585 5465 24600 5485
rect 24550 5435 24600 5465
rect 24550 5415 24565 5435
rect 24585 5415 24600 5435
rect 24550 5385 24600 5415
rect 24550 5365 24565 5385
rect 24585 5365 24600 5385
rect 24550 5335 24600 5365
rect 24550 5315 24565 5335
rect 24585 5315 24600 5335
rect 24550 5285 24600 5315
rect 24550 5265 24565 5285
rect 24585 5265 24600 5285
rect 24550 5235 24600 5265
rect 24550 5215 24565 5235
rect 24585 5215 24600 5235
rect 24550 5185 24600 5215
rect 24550 5165 24565 5185
rect 24585 5165 24600 5185
rect 24550 5135 24600 5165
rect 24550 5115 24565 5135
rect 24585 5115 24600 5135
rect 24550 5085 24600 5115
rect 24550 5065 24565 5085
rect 24585 5065 24600 5085
rect 24550 5035 24600 5065
rect 24550 5015 24565 5035
rect 24585 5015 24600 5035
rect 24550 5000 24600 5015
rect 24700 5000 24750 5500
rect 24850 5000 24900 5500
rect 25000 5000 25050 5500
rect 25150 5485 25200 5500
rect 25150 5465 25165 5485
rect 25185 5465 25200 5485
rect 25150 5435 25200 5465
rect 25150 5415 25165 5435
rect 25185 5415 25200 5435
rect 25150 5385 25200 5415
rect 25150 5365 25165 5385
rect 25185 5365 25200 5385
rect 25150 5335 25200 5365
rect 25150 5315 25165 5335
rect 25185 5315 25200 5335
rect 25150 5285 25200 5315
rect 25150 5265 25165 5285
rect 25185 5265 25200 5285
rect 25150 5235 25200 5265
rect 25150 5215 25165 5235
rect 25185 5215 25200 5235
rect 25150 5185 25200 5215
rect 25150 5165 25165 5185
rect 25185 5165 25200 5185
rect 25150 5135 25200 5165
rect 25150 5115 25165 5135
rect 25185 5115 25200 5135
rect 25150 5085 25200 5115
rect 25150 5065 25165 5085
rect 25185 5065 25200 5085
rect 25150 5035 25200 5065
rect 25150 5015 25165 5035
rect 25185 5015 25200 5035
rect 25150 5000 25200 5015
rect 25300 5000 25350 5500
rect 25450 5000 25500 5500
rect 25600 5485 25650 5500
rect 25600 5465 25615 5485
rect 25635 5465 25650 5485
rect 25600 5435 25650 5465
rect 25600 5415 25615 5435
rect 25635 5415 25650 5435
rect 25600 5385 25650 5415
rect 25600 5365 25615 5385
rect 25635 5365 25650 5385
rect 25600 5335 25650 5365
rect 25600 5315 25615 5335
rect 25635 5315 25650 5335
rect 25600 5285 25650 5315
rect 25600 5265 25615 5285
rect 25635 5265 25650 5285
rect 25600 5235 25650 5265
rect 25600 5215 25615 5235
rect 25635 5215 25650 5235
rect 25600 5185 25650 5215
rect 25600 5165 25615 5185
rect 25635 5165 25650 5185
rect 25600 5135 25650 5165
rect 25600 5115 25615 5135
rect 25635 5115 25650 5135
rect 25600 5085 25650 5115
rect 25600 5065 25615 5085
rect 25635 5065 25650 5085
rect 25600 5035 25650 5065
rect 25600 5015 25615 5035
rect 25635 5015 25650 5035
rect 25600 5000 25650 5015
rect 25750 5000 25800 5500
rect 25900 5000 25950 5500
rect 26050 5485 26100 5500
rect 26050 5465 26065 5485
rect 26085 5465 26100 5485
rect 26050 5435 26100 5465
rect 26050 5415 26065 5435
rect 26085 5415 26100 5435
rect 26050 5385 26100 5415
rect 26050 5365 26065 5385
rect 26085 5365 26100 5385
rect 26050 5335 26100 5365
rect 26050 5315 26065 5335
rect 26085 5315 26100 5335
rect 26050 5285 26100 5315
rect 26050 5265 26065 5285
rect 26085 5265 26100 5285
rect 26050 5235 26100 5265
rect 26050 5215 26065 5235
rect 26085 5215 26100 5235
rect 26050 5185 26100 5215
rect 26050 5165 26065 5185
rect 26085 5165 26100 5185
rect 26050 5135 26100 5165
rect 26050 5115 26065 5135
rect 26085 5115 26100 5135
rect 26050 5085 26100 5115
rect 26050 5065 26065 5085
rect 26085 5065 26100 5085
rect 26050 5035 26100 5065
rect 26050 5015 26065 5035
rect 26085 5015 26100 5035
rect 26050 5000 26100 5015
rect 26200 5000 26250 5500
rect 26350 5000 26400 5500
rect 26500 5000 26550 5500
rect 26650 5485 26700 5500
rect 26650 5465 26665 5485
rect 26685 5465 26700 5485
rect 26650 5435 26700 5465
rect 26650 5415 26665 5435
rect 26685 5415 26700 5435
rect 26650 5385 26700 5415
rect 26650 5365 26665 5385
rect 26685 5365 26700 5385
rect 26650 5335 26700 5365
rect 26650 5315 26665 5335
rect 26685 5315 26700 5335
rect 26650 5285 26700 5315
rect 26650 5265 26665 5285
rect 26685 5265 26700 5285
rect 26650 5235 26700 5265
rect 26650 5215 26665 5235
rect 26685 5215 26700 5235
rect 26650 5185 26700 5215
rect 26650 5165 26665 5185
rect 26685 5165 26700 5185
rect 26650 5135 26700 5165
rect 26650 5115 26665 5135
rect 26685 5115 26700 5135
rect 26650 5085 26700 5115
rect 26650 5065 26665 5085
rect 26685 5065 26700 5085
rect 26650 5035 26700 5065
rect 26650 5015 26665 5035
rect 26685 5015 26700 5035
rect 26650 5000 26700 5015
rect 26800 5000 26850 5500
rect 26950 5000 27000 5500
rect 27100 5000 27150 5500
rect 27250 5485 27300 5500
rect 27250 5465 27265 5485
rect 27285 5465 27300 5485
rect 27250 5435 27300 5465
rect 27250 5415 27265 5435
rect 27285 5415 27300 5435
rect 27250 5385 27300 5415
rect 27250 5365 27265 5385
rect 27285 5365 27300 5385
rect 27250 5335 27300 5365
rect 27250 5315 27265 5335
rect 27285 5315 27300 5335
rect 27250 5285 27300 5315
rect 27250 5265 27265 5285
rect 27285 5265 27300 5285
rect 27250 5235 27300 5265
rect 27250 5215 27265 5235
rect 27285 5215 27300 5235
rect 27250 5185 27300 5215
rect 27250 5165 27265 5185
rect 27285 5165 27300 5185
rect 27250 5135 27300 5165
rect 27250 5115 27265 5135
rect 27285 5115 27300 5135
rect 27250 5085 27300 5115
rect 27250 5065 27265 5085
rect 27285 5065 27300 5085
rect 27250 5035 27300 5065
rect 27250 5015 27265 5035
rect 27285 5015 27300 5035
rect 27250 5000 27300 5015
rect 27400 5000 27450 5500
rect 27550 5000 27600 5500
rect 27700 5485 27750 5500
rect 27700 5465 27715 5485
rect 27735 5465 27750 5485
rect 27700 5435 27750 5465
rect 27700 5415 27715 5435
rect 27735 5415 27750 5435
rect 27700 5385 27750 5415
rect 27700 5365 27715 5385
rect 27735 5365 27750 5385
rect 27700 5335 27750 5365
rect 27700 5315 27715 5335
rect 27735 5315 27750 5335
rect 27700 5285 27750 5315
rect 27700 5265 27715 5285
rect 27735 5265 27750 5285
rect 27700 5235 27750 5265
rect 27700 5215 27715 5235
rect 27735 5215 27750 5235
rect 27700 5185 27750 5215
rect 27700 5165 27715 5185
rect 27735 5165 27750 5185
rect 27700 5135 27750 5165
rect 27700 5115 27715 5135
rect 27735 5115 27750 5135
rect 27700 5085 27750 5115
rect 27700 5065 27715 5085
rect 27735 5065 27750 5085
rect 27700 5035 27750 5065
rect 27700 5015 27715 5035
rect 27735 5015 27750 5035
rect 27700 5000 27750 5015
rect 27850 5000 27900 5500
rect 28000 5000 28050 5500
rect 28150 5485 28200 5500
rect 28150 5465 28165 5485
rect 28185 5465 28200 5485
rect 28150 5435 28200 5465
rect 28150 5415 28165 5435
rect 28185 5415 28200 5435
rect 28150 5385 28200 5415
rect 28150 5365 28165 5385
rect 28185 5365 28200 5385
rect 28150 5335 28200 5365
rect 28150 5315 28165 5335
rect 28185 5315 28200 5335
rect 28150 5285 28200 5315
rect 28150 5265 28165 5285
rect 28185 5265 28200 5285
rect 28150 5235 28200 5265
rect 28150 5215 28165 5235
rect 28185 5215 28200 5235
rect 28150 5185 28200 5215
rect 28150 5165 28165 5185
rect 28185 5165 28200 5185
rect 28150 5135 28200 5165
rect 28150 5115 28165 5135
rect 28185 5115 28200 5135
rect 28150 5085 28200 5115
rect 28150 5065 28165 5085
rect 28185 5065 28200 5085
rect 28150 5035 28200 5065
rect 28150 5015 28165 5035
rect 28185 5015 28200 5035
rect 28150 5000 28200 5015
rect 28300 5000 28350 5500
rect 28450 5000 28500 5500
rect 28600 5000 28650 5500
rect 28750 5485 28800 5500
rect 28750 5465 28765 5485
rect 28785 5465 28800 5485
rect 28750 5435 28800 5465
rect 28750 5415 28765 5435
rect 28785 5415 28800 5435
rect 28750 5385 28800 5415
rect 28750 5365 28765 5385
rect 28785 5365 28800 5385
rect 28750 5335 28800 5365
rect 28750 5315 28765 5335
rect 28785 5315 28800 5335
rect 28750 5285 28800 5315
rect 28750 5265 28765 5285
rect 28785 5265 28800 5285
rect 28750 5235 28800 5265
rect 28750 5215 28765 5235
rect 28785 5215 28800 5235
rect 28750 5185 28800 5215
rect 28750 5165 28765 5185
rect 28785 5165 28800 5185
rect 28750 5135 28800 5165
rect 28750 5115 28765 5135
rect 28785 5115 28800 5135
rect 28750 5085 28800 5115
rect 28750 5065 28765 5085
rect 28785 5065 28800 5085
rect 28750 5035 28800 5065
rect 28750 5015 28765 5035
rect 28785 5015 28800 5035
rect 28750 5000 28800 5015
rect 28900 5000 28950 5500
rect 29050 5000 29100 5500
rect 29200 5000 29250 5500
rect 29350 5485 29400 5500
rect 29350 5465 29365 5485
rect 29385 5465 29400 5485
rect 29350 5435 29400 5465
rect 29350 5415 29365 5435
rect 29385 5415 29400 5435
rect 29350 5385 29400 5415
rect 29350 5365 29365 5385
rect 29385 5365 29400 5385
rect 29350 5335 29400 5365
rect 29350 5315 29365 5335
rect 29385 5315 29400 5335
rect 29350 5285 29400 5315
rect 29350 5265 29365 5285
rect 29385 5265 29400 5285
rect 29350 5235 29400 5265
rect 29350 5215 29365 5235
rect 29385 5215 29400 5235
rect 29350 5185 29400 5215
rect 29350 5165 29365 5185
rect 29385 5165 29400 5185
rect 29350 5135 29400 5165
rect 29350 5115 29365 5135
rect 29385 5115 29400 5135
rect 29350 5085 29400 5115
rect 29350 5065 29365 5085
rect 29385 5065 29400 5085
rect 29350 5035 29400 5065
rect 29350 5015 29365 5035
rect 29385 5015 29400 5035
rect 29350 5000 29400 5015
rect 29500 5485 29550 5500
rect 29500 5465 29515 5485
rect 29535 5465 29550 5485
rect 29500 5435 29550 5465
rect 29500 5415 29515 5435
rect 29535 5415 29550 5435
rect 29500 5385 29550 5415
rect 29500 5365 29515 5385
rect 29535 5365 29550 5385
rect 29500 5335 29550 5365
rect 29500 5315 29515 5335
rect 29535 5315 29550 5335
rect 29500 5285 29550 5315
rect 29500 5265 29515 5285
rect 29535 5265 29550 5285
rect 29500 5235 29550 5265
rect 29500 5215 29515 5235
rect 29535 5215 29550 5235
rect 29500 5185 29550 5215
rect 29500 5165 29515 5185
rect 29535 5165 29550 5185
rect 29500 5135 29550 5165
rect 29500 5115 29515 5135
rect 29535 5115 29550 5135
rect 29500 5085 29550 5115
rect 29500 5065 29515 5085
rect 29535 5065 29550 5085
rect 29500 5035 29550 5065
rect 29500 5015 29515 5035
rect 29535 5015 29550 5035
rect 29500 5000 29550 5015
rect 29650 5485 29700 5500
rect 29650 5465 29665 5485
rect 29685 5465 29700 5485
rect 29650 5435 29700 5465
rect 29650 5415 29665 5435
rect 29685 5415 29700 5435
rect 29650 5385 29700 5415
rect 29650 5365 29665 5385
rect 29685 5365 29700 5385
rect 29650 5335 29700 5365
rect 29650 5315 29665 5335
rect 29685 5315 29700 5335
rect 29650 5285 29700 5315
rect 29650 5265 29665 5285
rect 29685 5265 29700 5285
rect 29650 5235 29700 5265
rect 29650 5215 29665 5235
rect 29685 5215 29700 5235
rect 29650 5185 29700 5215
rect 29650 5165 29665 5185
rect 29685 5165 29700 5185
rect 29650 5135 29700 5165
rect 29650 5115 29665 5135
rect 29685 5115 29700 5135
rect 29650 5085 29700 5115
rect 29650 5065 29665 5085
rect 29685 5065 29700 5085
rect 29650 5035 29700 5065
rect 29650 5015 29665 5035
rect 29685 5015 29700 5035
rect 29650 5000 29700 5015
rect 29800 5485 29850 5500
rect 29800 5465 29815 5485
rect 29835 5465 29850 5485
rect 29800 5435 29850 5465
rect 29800 5415 29815 5435
rect 29835 5415 29850 5435
rect 29800 5385 29850 5415
rect 29800 5365 29815 5385
rect 29835 5365 29850 5385
rect 29800 5335 29850 5365
rect 29800 5315 29815 5335
rect 29835 5315 29850 5335
rect 29800 5285 29850 5315
rect 29800 5265 29815 5285
rect 29835 5265 29850 5285
rect 29800 5235 29850 5265
rect 29800 5215 29815 5235
rect 29835 5215 29850 5235
rect 29800 5185 29850 5215
rect 29800 5165 29815 5185
rect 29835 5165 29850 5185
rect 29800 5135 29850 5165
rect 29800 5115 29815 5135
rect 29835 5115 29850 5135
rect 29800 5085 29850 5115
rect 29800 5065 29815 5085
rect 29835 5065 29850 5085
rect 29800 5035 29850 5065
rect 29800 5015 29815 5035
rect 29835 5015 29850 5035
rect 29800 5000 29850 5015
rect 29950 5485 30000 5500
rect 29950 5465 29965 5485
rect 29985 5465 30000 5485
rect 29950 5435 30000 5465
rect 29950 5415 29965 5435
rect 29985 5415 30000 5435
rect 29950 5385 30000 5415
rect 29950 5365 29965 5385
rect 29985 5365 30000 5385
rect 29950 5335 30000 5365
rect 29950 5315 29965 5335
rect 29985 5315 30000 5335
rect 29950 5285 30000 5315
rect 29950 5265 29965 5285
rect 29985 5265 30000 5285
rect 29950 5235 30000 5265
rect 29950 5215 29965 5235
rect 29985 5215 30000 5235
rect 29950 5185 30000 5215
rect 29950 5165 29965 5185
rect 29985 5165 30000 5185
rect 29950 5135 30000 5165
rect 29950 5115 29965 5135
rect 29985 5115 30000 5135
rect 29950 5085 30000 5115
rect 29950 5065 29965 5085
rect 29985 5065 30000 5085
rect 29950 5035 30000 5065
rect 29950 5015 29965 5035
rect 29985 5015 30000 5035
rect 29950 5000 30000 5015
rect 30100 5485 30150 5500
rect 30100 5465 30115 5485
rect 30135 5465 30150 5485
rect 30100 5435 30150 5465
rect 30100 5415 30115 5435
rect 30135 5415 30150 5435
rect 30100 5385 30150 5415
rect 30100 5365 30115 5385
rect 30135 5365 30150 5385
rect 30100 5335 30150 5365
rect 30100 5315 30115 5335
rect 30135 5315 30150 5335
rect 30100 5285 30150 5315
rect 30100 5265 30115 5285
rect 30135 5265 30150 5285
rect 30100 5235 30150 5265
rect 30100 5215 30115 5235
rect 30135 5215 30150 5235
rect 30100 5185 30150 5215
rect 30100 5165 30115 5185
rect 30135 5165 30150 5185
rect 30100 5135 30150 5165
rect 30100 5115 30115 5135
rect 30135 5115 30150 5135
rect 30100 5085 30150 5115
rect 30100 5065 30115 5085
rect 30135 5065 30150 5085
rect 30100 5035 30150 5065
rect 30100 5015 30115 5035
rect 30135 5015 30150 5035
rect 30100 5000 30150 5015
rect 30250 5485 30300 5500
rect 30250 5465 30265 5485
rect 30285 5465 30300 5485
rect 30250 5435 30300 5465
rect 30250 5415 30265 5435
rect 30285 5415 30300 5435
rect 30250 5385 30300 5415
rect 30250 5365 30265 5385
rect 30285 5365 30300 5385
rect 30250 5335 30300 5365
rect 30250 5315 30265 5335
rect 30285 5315 30300 5335
rect 30250 5285 30300 5315
rect 30250 5265 30265 5285
rect 30285 5265 30300 5285
rect 30250 5235 30300 5265
rect 30250 5215 30265 5235
rect 30285 5215 30300 5235
rect 30250 5185 30300 5215
rect 30250 5165 30265 5185
rect 30285 5165 30300 5185
rect 30250 5135 30300 5165
rect 30250 5115 30265 5135
rect 30285 5115 30300 5135
rect 30250 5085 30300 5115
rect 30250 5065 30265 5085
rect 30285 5065 30300 5085
rect 30250 5035 30300 5065
rect 30250 5015 30265 5035
rect 30285 5015 30300 5035
rect 30250 5000 30300 5015
rect 30400 5485 30450 5500
rect 30400 5465 30415 5485
rect 30435 5465 30450 5485
rect 30400 5435 30450 5465
rect 30400 5415 30415 5435
rect 30435 5415 30450 5435
rect 30400 5385 30450 5415
rect 30400 5365 30415 5385
rect 30435 5365 30450 5385
rect 30400 5335 30450 5365
rect 30400 5315 30415 5335
rect 30435 5315 30450 5335
rect 30400 5285 30450 5315
rect 30400 5265 30415 5285
rect 30435 5265 30450 5285
rect 30400 5235 30450 5265
rect 30400 5215 30415 5235
rect 30435 5215 30450 5235
rect 30400 5185 30450 5215
rect 30400 5165 30415 5185
rect 30435 5165 30450 5185
rect 30400 5135 30450 5165
rect 30400 5115 30415 5135
rect 30435 5115 30450 5135
rect 30400 5085 30450 5115
rect 30400 5065 30415 5085
rect 30435 5065 30450 5085
rect 30400 5035 30450 5065
rect 30400 5015 30415 5035
rect 30435 5015 30450 5035
rect 30400 5000 30450 5015
rect 30550 5485 30600 5500
rect 30550 5465 30565 5485
rect 30585 5465 30600 5485
rect 30550 5435 30600 5465
rect 30550 5415 30565 5435
rect 30585 5415 30600 5435
rect 30550 5385 30600 5415
rect 30550 5365 30565 5385
rect 30585 5365 30600 5385
rect 30550 5335 30600 5365
rect 30550 5315 30565 5335
rect 30585 5315 30600 5335
rect 30550 5285 30600 5315
rect 30550 5265 30565 5285
rect 30585 5265 30600 5285
rect 30550 5235 30600 5265
rect 30550 5215 30565 5235
rect 30585 5215 30600 5235
rect 30550 5185 30600 5215
rect 30550 5165 30565 5185
rect 30585 5165 30600 5185
rect 30550 5135 30600 5165
rect 30550 5115 30565 5135
rect 30585 5115 30600 5135
rect 30550 5085 30600 5115
rect 30550 5065 30565 5085
rect 30585 5065 30600 5085
rect 30550 5035 30600 5065
rect 30550 5015 30565 5035
rect 30585 5015 30600 5035
rect 30550 5000 30600 5015
rect 30700 5485 30750 5500
rect 30700 5465 30715 5485
rect 30735 5465 30750 5485
rect 30700 5435 30750 5465
rect 30700 5415 30715 5435
rect 30735 5415 30750 5435
rect 30700 5385 30750 5415
rect 30700 5365 30715 5385
rect 30735 5365 30750 5385
rect 30700 5335 30750 5365
rect 30700 5315 30715 5335
rect 30735 5315 30750 5335
rect 30700 5285 30750 5315
rect 30700 5265 30715 5285
rect 30735 5265 30750 5285
rect 30700 5235 30750 5265
rect 30700 5215 30715 5235
rect 30735 5215 30750 5235
rect 30700 5185 30750 5215
rect 30700 5165 30715 5185
rect 30735 5165 30750 5185
rect 30700 5135 30750 5165
rect 30700 5115 30715 5135
rect 30735 5115 30750 5135
rect 30700 5085 30750 5115
rect 30700 5065 30715 5085
rect 30735 5065 30750 5085
rect 30700 5035 30750 5065
rect 30700 5015 30715 5035
rect 30735 5015 30750 5035
rect 30700 5000 30750 5015
rect 30850 5485 30900 5500
rect 30850 5465 30865 5485
rect 30885 5465 30900 5485
rect 30850 5435 30900 5465
rect 30850 5415 30865 5435
rect 30885 5415 30900 5435
rect 30850 5385 30900 5415
rect 30850 5365 30865 5385
rect 30885 5365 30900 5385
rect 30850 5335 30900 5365
rect 30850 5315 30865 5335
rect 30885 5315 30900 5335
rect 30850 5285 30900 5315
rect 30850 5265 30865 5285
rect 30885 5265 30900 5285
rect 30850 5235 30900 5265
rect 30850 5215 30865 5235
rect 30885 5215 30900 5235
rect 30850 5185 30900 5215
rect 30850 5165 30865 5185
rect 30885 5165 30900 5185
rect 30850 5135 30900 5165
rect 30850 5115 30865 5135
rect 30885 5115 30900 5135
rect 30850 5085 30900 5115
rect 30850 5065 30865 5085
rect 30885 5065 30900 5085
rect 30850 5035 30900 5065
rect 30850 5015 30865 5035
rect 30885 5015 30900 5035
rect 30850 5000 30900 5015
rect 31000 5485 31050 5500
rect 31000 5465 31015 5485
rect 31035 5465 31050 5485
rect 31000 5435 31050 5465
rect 31000 5415 31015 5435
rect 31035 5415 31050 5435
rect 31000 5385 31050 5415
rect 31000 5365 31015 5385
rect 31035 5365 31050 5385
rect 31000 5335 31050 5365
rect 31000 5315 31015 5335
rect 31035 5315 31050 5335
rect 31000 5285 31050 5315
rect 31000 5265 31015 5285
rect 31035 5265 31050 5285
rect 31000 5235 31050 5265
rect 31000 5215 31015 5235
rect 31035 5215 31050 5235
rect 31000 5185 31050 5215
rect 31000 5165 31015 5185
rect 31035 5165 31050 5185
rect 31000 5135 31050 5165
rect 31000 5115 31015 5135
rect 31035 5115 31050 5135
rect 31000 5085 31050 5115
rect 31000 5065 31015 5085
rect 31035 5065 31050 5085
rect 31000 5035 31050 5065
rect 31000 5015 31015 5035
rect 31035 5015 31050 5035
rect 31000 5000 31050 5015
rect 31150 5485 31200 5500
rect 31150 5465 31165 5485
rect 31185 5465 31200 5485
rect 31150 5435 31200 5465
rect 31150 5415 31165 5435
rect 31185 5415 31200 5435
rect 31150 5385 31200 5415
rect 31150 5365 31165 5385
rect 31185 5365 31200 5385
rect 31150 5335 31200 5365
rect 31150 5315 31165 5335
rect 31185 5315 31200 5335
rect 31150 5285 31200 5315
rect 31150 5265 31165 5285
rect 31185 5265 31200 5285
rect 31150 5235 31200 5265
rect 31150 5215 31165 5235
rect 31185 5215 31200 5235
rect 31150 5185 31200 5215
rect 31150 5165 31165 5185
rect 31185 5165 31200 5185
rect 31150 5135 31200 5165
rect 31150 5115 31165 5135
rect 31185 5115 31200 5135
rect 31150 5085 31200 5115
rect 31150 5065 31165 5085
rect 31185 5065 31200 5085
rect 31150 5035 31200 5065
rect 31150 5015 31165 5035
rect 31185 5015 31200 5035
rect 31150 5000 31200 5015
rect 31300 5485 31350 5500
rect 31300 5465 31315 5485
rect 31335 5465 31350 5485
rect 31300 5435 31350 5465
rect 31300 5415 31315 5435
rect 31335 5415 31350 5435
rect 31300 5385 31350 5415
rect 31300 5365 31315 5385
rect 31335 5365 31350 5385
rect 31300 5335 31350 5365
rect 31300 5315 31315 5335
rect 31335 5315 31350 5335
rect 31300 5285 31350 5315
rect 31300 5265 31315 5285
rect 31335 5265 31350 5285
rect 31300 5235 31350 5265
rect 31300 5215 31315 5235
rect 31335 5215 31350 5235
rect 31300 5185 31350 5215
rect 31300 5165 31315 5185
rect 31335 5165 31350 5185
rect 31300 5135 31350 5165
rect 31300 5115 31315 5135
rect 31335 5115 31350 5135
rect 31300 5085 31350 5115
rect 31300 5065 31315 5085
rect 31335 5065 31350 5085
rect 31300 5035 31350 5065
rect 31300 5015 31315 5035
rect 31335 5015 31350 5035
rect 31300 5000 31350 5015
rect 31450 5485 31500 5500
rect 31450 5465 31465 5485
rect 31485 5465 31500 5485
rect 31450 5435 31500 5465
rect 31450 5415 31465 5435
rect 31485 5415 31500 5435
rect 31450 5385 31500 5415
rect 31450 5365 31465 5385
rect 31485 5365 31500 5385
rect 31450 5335 31500 5365
rect 31450 5315 31465 5335
rect 31485 5315 31500 5335
rect 31450 5285 31500 5315
rect 31450 5265 31465 5285
rect 31485 5265 31500 5285
rect 31450 5235 31500 5265
rect 31450 5215 31465 5235
rect 31485 5215 31500 5235
rect 31450 5185 31500 5215
rect 31450 5165 31465 5185
rect 31485 5165 31500 5185
rect 31450 5135 31500 5165
rect 31450 5115 31465 5135
rect 31485 5115 31500 5135
rect 31450 5085 31500 5115
rect 31450 5065 31465 5085
rect 31485 5065 31500 5085
rect 31450 5035 31500 5065
rect 31450 5015 31465 5035
rect 31485 5015 31500 5035
rect 31450 5000 31500 5015
rect 31600 5000 31650 5500
rect 31750 5000 31800 5500
rect 31900 5000 31950 5500
rect 32050 5485 32100 5500
rect 32050 5465 32065 5485
rect 32085 5465 32100 5485
rect 32050 5435 32100 5465
rect 32050 5415 32065 5435
rect 32085 5415 32100 5435
rect 32050 5385 32100 5415
rect 32050 5365 32065 5385
rect 32085 5365 32100 5385
rect 32050 5335 32100 5365
rect 32050 5315 32065 5335
rect 32085 5315 32100 5335
rect 32050 5285 32100 5315
rect 32050 5265 32065 5285
rect 32085 5265 32100 5285
rect 32050 5235 32100 5265
rect 32050 5215 32065 5235
rect 32085 5215 32100 5235
rect 32050 5185 32100 5215
rect 32050 5165 32065 5185
rect 32085 5165 32100 5185
rect 32050 5135 32100 5165
rect 32050 5115 32065 5135
rect 32085 5115 32100 5135
rect 32050 5085 32100 5115
rect 32050 5065 32065 5085
rect 32085 5065 32100 5085
rect 32050 5035 32100 5065
rect 32050 5015 32065 5035
rect 32085 5015 32100 5035
rect 32050 5000 32100 5015
rect -650 4835 -600 4850
rect -650 4815 -635 4835
rect -615 4815 -600 4835
rect -650 4785 -600 4815
rect -650 4765 -635 4785
rect -615 4765 -600 4785
rect -650 4735 -600 4765
rect -650 4715 -635 4735
rect -615 4715 -600 4735
rect -650 4685 -600 4715
rect -650 4665 -635 4685
rect -615 4665 -600 4685
rect -650 4635 -600 4665
rect -650 4615 -635 4635
rect -615 4615 -600 4635
rect -650 4585 -600 4615
rect -650 4565 -635 4585
rect -615 4565 -600 4585
rect -650 4535 -600 4565
rect -650 4515 -635 4535
rect -615 4515 -600 4535
rect -650 4485 -600 4515
rect -650 4465 -635 4485
rect -615 4465 -600 4485
rect -650 4435 -600 4465
rect -650 4415 -635 4435
rect -615 4415 -600 4435
rect -650 4385 -600 4415
rect -650 4365 -635 4385
rect -615 4365 -600 4385
rect -650 4350 -600 4365
rect -500 4835 -450 4850
rect -500 4815 -485 4835
rect -465 4815 -450 4835
rect -500 4785 -450 4815
rect -500 4765 -485 4785
rect -465 4765 -450 4785
rect -500 4735 -450 4765
rect -500 4715 -485 4735
rect -465 4715 -450 4735
rect -500 4685 -450 4715
rect -500 4665 -485 4685
rect -465 4665 -450 4685
rect -500 4635 -450 4665
rect -500 4615 -485 4635
rect -465 4615 -450 4635
rect -500 4585 -450 4615
rect -500 4565 -485 4585
rect -465 4565 -450 4585
rect -500 4535 -450 4565
rect -500 4515 -485 4535
rect -465 4515 -450 4535
rect -500 4485 -450 4515
rect -500 4465 -485 4485
rect -465 4465 -450 4485
rect -500 4435 -450 4465
rect -500 4415 -485 4435
rect -465 4415 -450 4435
rect -500 4385 -450 4415
rect -500 4365 -485 4385
rect -465 4365 -450 4385
rect -500 4350 -450 4365
rect -350 4835 -300 4850
rect -350 4815 -335 4835
rect -315 4815 -300 4835
rect -350 4785 -300 4815
rect -350 4765 -335 4785
rect -315 4765 -300 4785
rect -350 4735 -300 4765
rect -350 4715 -335 4735
rect -315 4715 -300 4735
rect -350 4685 -300 4715
rect -350 4665 -335 4685
rect -315 4665 -300 4685
rect -350 4635 -300 4665
rect -350 4615 -335 4635
rect -315 4615 -300 4635
rect -350 4585 -300 4615
rect -350 4565 -335 4585
rect -315 4565 -300 4585
rect -350 4535 -300 4565
rect -350 4515 -335 4535
rect -315 4515 -300 4535
rect -350 4485 -300 4515
rect -350 4465 -335 4485
rect -315 4465 -300 4485
rect -350 4435 -300 4465
rect -350 4415 -335 4435
rect -315 4415 -300 4435
rect -350 4385 -300 4415
rect -350 4365 -335 4385
rect -315 4365 -300 4385
rect -350 4350 -300 4365
rect -200 4835 -150 4850
rect -200 4815 -185 4835
rect -165 4815 -150 4835
rect -200 4785 -150 4815
rect -200 4765 -185 4785
rect -165 4765 -150 4785
rect -200 4735 -150 4765
rect -200 4715 -185 4735
rect -165 4715 -150 4735
rect -200 4685 -150 4715
rect -200 4665 -185 4685
rect -165 4665 -150 4685
rect -200 4635 -150 4665
rect -200 4615 -185 4635
rect -165 4615 -150 4635
rect -200 4585 -150 4615
rect -200 4565 -185 4585
rect -165 4565 -150 4585
rect -200 4535 -150 4565
rect -200 4515 -185 4535
rect -165 4515 -150 4535
rect -200 4485 -150 4515
rect -200 4465 -185 4485
rect -165 4465 -150 4485
rect -200 4435 -150 4465
rect -200 4415 -185 4435
rect -165 4415 -150 4435
rect -200 4385 -150 4415
rect -200 4365 -185 4385
rect -165 4365 -150 4385
rect -200 4350 -150 4365
rect -50 4835 0 4850
rect -50 4815 -35 4835
rect -15 4815 0 4835
rect -50 4785 0 4815
rect -50 4765 -35 4785
rect -15 4765 0 4785
rect -50 4735 0 4765
rect -50 4715 -35 4735
rect -15 4715 0 4735
rect -50 4685 0 4715
rect -50 4665 -35 4685
rect -15 4665 0 4685
rect -50 4635 0 4665
rect -50 4615 -35 4635
rect -15 4615 0 4635
rect -50 4585 0 4615
rect -50 4565 -35 4585
rect -15 4565 0 4585
rect -50 4535 0 4565
rect -50 4515 -35 4535
rect -15 4515 0 4535
rect -50 4485 0 4515
rect -50 4465 -35 4485
rect -15 4465 0 4485
rect -50 4435 0 4465
rect -50 4415 -35 4435
rect -15 4415 0 4435
rect -50 4385 0 4415
rect -50 4365 -35 4385
rect -15 4365 0 4385
rect -50 4350 0 4365
rect 100 4350 150 4850
rect 250 4350 300 4850
rect 400 4350 450 4850
rect 550 4835 600 4850
rect 550 4815 565 4835
rect 585 4815 600 4835
rect 550 4785 600 4815
rect 550 4765 565 4785
rect 585 4765 600 4785
rect 550 4735 600 4765
rect 550 4715 565 4735
rect 585 4715 600 4735
rect 550 4685 600 4715
rect 550 4665 565 4685
rect 585 4665 600 4685
rect 550 4635 600 4665
rect 550 4615 565 4635
rect 585 4615 600 4635
rect 550 4585 600 4615
rect 550 4565 565 4585
rect 585 4565 600 4585
rect 550 4535 600 4565
rect 550 4515 565 4535
rect 585 4515 600 4535
rect 550 4485 600 4515
rect 550 4465 565 4485
rect 585 4465 600 4485
rect 550 4435 600 4465
rect 550 4415 565 4435
rect 585 4415 600 4435
rect 550 4385 600 4415
rect 550 4365 565 4385
rect 585 4365 600 4385
rect 550 4350 600 4365
rect 700 4835 750 4850
rect 700 4815 715 4835
rect 735 4815 750 4835
rect 700 4785 750 4815
rect 700 4765 715 4785
rect 735 4765 750 4785
rect 700 4735 750 4765
rect 700 4715 715 4735
rect 735 4715 750 4735
rect 700 4685 750 4715
rect 700 4665 715 4685
rect 735 4665 750 4685
rect 700 4635 750 4665
rect 700 4615 715 4635
rect 735 4615 750 4635
rect 700 4585 750 4615
rect 700 4565 715 4585
rect 735 4565 750 4585
rect 700 4535 750 4565
rect 700 4515 715 4535
rect 735 4515 750 4535
rect 700 4485 750 4515
rect 700 4465 715 4485
rect 735 4465 750 4485
rect 700 4435 750 4465
rect 700 4415 715 4435
rect 735 4415 750 4435
rect 700 4385 750 4415
rect 700 4365 715 4385
rect 735 4365 750 4385
rect 700 4350 750 4365
rect 850 4835 900 4850
rect 850 4815 865 4835
rect 885 4815 900 4835
rect 850 4785 900 4815
rect 850 4765 865 4785
rect 885 4765 900 4785
rect 850 4735 900 4765
rect 850 4715 865 4735
rect 885 4715 900 4735
rect 850 4685 900 4715
rect 850 4665 865 4685
rect 885 4665 900 4685
rect 850 4635 900 4665
rect 850 4615 865 4635
rect 885 4615 900 4635
rect 850 4585 900 4615
rect 850 4565 865 4585
rect 885 4565 900 4585
rect 850 4535 900 4565
rect 850 4515 865 4535
rect 885 4515 900 4535
rect 850 4485 900 4515
rect 850 4465 865 4485
rect 885 4465 900 4485
rect 850 4435 900 4465
rect 850 4415 865 4435
rect 885 4415 900 4435
rect 850 4385 900 4415
rect 850 4365 865 4385
rect 885 4365 900 4385
rect 850 4350 900 4365
rect 1000 4835 1050 4850
rect 1000 4815 1015 4835
rect 1035 4815 1050 4835
rect 1000 4785 1050 4815
rect 1000 4765 1015 4785
rect 1035 4765 1050 4785
rect 1000 4735 1050 4765
rect 1000 4715 1015 4735
rect 1035 4715 1050 4735
rect 1000 4685 1050 4715
rect 1000 4665 1015 4685
rect 1035 4665 1050 4685
rect 1000 4635 1050 4665
rect 1000 4615 1015 4635
rect 1035 4615 1050 4635
rect 1000 4585 1050 4615
rect 1000 4565 1015 4585
rect 1035 4565 1050 4585
rect 1000 4535 1050 4565
rect 1000 4515 1015 4535
rect 1035 4515 1050 4535
rect 1000 4485 1050 4515
rect 1000 4465 1015 4485
rect 1035 4465 1050 4485
rect 1000 4435 1050 4465
rect 1000 4415 1015 4435
rect 1035 4415 1050 4435
rect 1000 4385 1050 4415
rect 1000 4365 1015 4385
rect 1035 4365 1050 4385
rect 1000 4350 1050 4365
rect 1150 4835 1200 4850
rect 1150 4815 1165 4835
rect 1185 4815 1200 4835
rect 1150 4785 1200 4815
rect 1150 4765 1165 4785
rect 1185 4765 1200 4785
rect 1150 4735 1200 4765
rect 1150 4715 1165 4735
rect 1185 4715 1200 4735
rect 1150 4685 1200 4715
rect 1150 4665 1165 4685
rect 1185 4665 1200 4685
rect 1150 4635 1200 4665
rect 1150 4615 1165 4635
rect 1185 4615 1200 4635
rect 1150 4585 1200 4615
rect 1150 4565 1165 4585
rect 1185 4565 1200 4585
rect 1150 4535 1200 4565
rect 1150 4515 1165 4535
rect 1185 4515 1200 4535
rect 1150 4485 1200 4515
rect 1150 4465 1165 4485
rect 1185 4465 1200 4485
rect 1150 4435 1200 4465
rect 1150 4415 1165 4435
rect 1185 4415 1200 4435
rect 1150 4385 1200 4415
rect 1150 4365 1165 4385
rect 1185 4365 1200 4385
rect 1150 4350 1200 4365
rect 1300 4835 1350 4850
rect 1300 4815 1315 4835
rect 1335 4815 1350 4835
rect 1300 4785 1350 4815
rect 1300 4765 1315 4785
rect 1335 4765 1350 4785
rect 1300 4735 1350 4765
rect 1300 4715 1315 4735
rect 1335 4715 1350 4735
rect 1300 4685 1350 4715
rect 1300 4665 1315 4685
rect 1335 4665 1350 4685
rect 1300 4635 1350 4665
rect 1300 4615 1315 4635
rect 1335 4615 1350 4635
rect 1300 4585 1350 4615
rect 1300 4565 1315 4585
rect 1335 4565 1350 4585
rect 1300 4535 1350 4565
rect 1300 4515 1315 4535
rect 1335 4515 1350 4535
rect 1300 4485 1350 4515
rect 1300 4465 1315 4485
rect 1335 4465 1350 4485
rect 1300 4435 1350 4465
rect 1300 4415 1315 4435
rect 1335 4415 1350 4435
rect 1300 4385 1350 4415
rect 1300 4365 1315 4385
rect 1335 4365 1350 4385
rect 1300 4350 1350 4365
rect 1450 4835 1500 4850
rect 1450 4815 1465 4835
rect 1485 4815 1500 4835
rect 1450 4785 1500 4815
rect 1450 4765 1465 4785
rect 1485 4765 1500 4785
rect 1450 4735 1500 4765
rect 1450 4715 1465 4735
rect 1485 4715 1500 4735
rect 1450 4685 1500 4715
rect 1450 4665 1465 4685
rect 1485 4665 1500 4685
rect 1450 4635 1500 4665
rect 1450 4615 1465 4635
rect 1485 4615 1500 4635
rect 1450 4585 1500 4615
rect 1450 4565 1465 4585
rect 1485 4565 1500 4585
rect 1450 4535 1500 4565
rect 1450 4515 1465 4535
rect 1485 4515 1500 4535
rect 1450 4485 1500 4515
rect 1450 4465 1465 4485
rect 1485 4465 1500 4485
rect 1450 4435 1500 4465
rect 1450 4415 1465 4435
rect 1485 4415 1500 4435
rect 1450 4385 1500 4415
rect 1450 4365 1465 4385
rect 1485 4365 1500 4385
rect 1450 4350 1500 4365
rect 1600 4835 1650 4850
rect 1600 4815 1615 4835
rect 1635 4815 1650 4835
rect 1600 4785 1650 4815
rect 1600 4765 1615 4785
rect 1635 4765 1650 4785
rect 1600 4735 1650 4765
rect 1600 4715 1615 4735
rect 1635 4715 1650 4735
rect 1600 4685 1650 4715
rect 1600 4665 1615 4685
rect 1635 4665 1650 4685
rect 1600 4635 1650 4665
rect 1600 4615 1615 4635
rect 1635 4615 1650 4635
rect 1600 4585 1650 4615
rect 1600 4565 1615 4585
rect 1635 4565 1650 4585
rect 1600 4535 1650 4565
rect 1600 4515 1615 4535
rect 1635 4515 1650 4535
rect 1600 4485 1650 4515
rect 1600 4465 1615 4485
rect 1635 4465 1650 4485
rect 1600 4435 1650 4465
rect 1600 4415 1615 4435
rect 1635 4415 1650 4435
rect 1600 4385 1650 4415
rect 1600 4365 1615 4385
rect 1635 4365 1650 4385
rect 1600 4350 1650 4365
rect 1750 4835 1800 4850
rect 1750 4815 1765 4835
rect 1785 4815 1800 4835
rect 1750 4785 1800 4815
rect 1750 4765 1765 4785
rect 1785 4765 1800 4785
rect 1750 4735 1800 4765
rect 1750 4715 1765 4735
rect 1785 4715 1800 4735
rect 1750 4685 1800 4715
rect 1750 4665 1765 4685
rect 1785 4665 1800 4685
rect 1750 4635 1800 4665
rect 1750 4615 1765 4635
rect 1785 4615 1800 4635
rect 1750 4585 1800 4615
rect 1750 4565 1765 4585
rect 1785 4565 1800 4585
rect 1750 4535 1800 4565
rect 1750 4515 1765 4535
rect 1785 4515 1800 4535
rect 1750 4485 1800 4515
rect 1750 4465 1765 4485
rect 1785 4465 1800 4485
rect 1750 4435 1800 4465
rect 1750 4415 1765 4435
rect 1785 4415 1800 4435
rect 1750 4385 1800 4415
rect 1750 4365 1765 4385
rect 1785 4365 1800 4385
rect 1750 4350 1800 4365
rect 1900 4835 1950 4850
rect 1900 4815 1915 4835
rect 1935 4815 1950 4835
rect 1900 4785 1950 4815
rect 1900 4765 1915 4785
rect 1935 4765 1950 4785
rect 1900 4735 1950 4765
rect 1900 4715 1915 4735
rect 1935 4715 1950 4735
rect 1900 4685 1950 4715
rect 1900 4665 1915 4685
rect 1935 4665 1950 4685
rect 1900 4635 1950 4665
rect 1900 4615 1915 4635
rect 1935 4615 1950 4635
rect 1900 4585 1950 4615
rect 1900 4565 1915 4585
rect 1935 4565 1950 4585
rect 1900 4535 1950 4565
rect 1900 4515 1915 4535
rect 1935 4515 1950 4535
rect 1900 4485 1950 4515
rect 1900 4465 1915 4485
rect 1935 4465 1950 4485
rect 1900 4435 1950 4465
rect 1900 4415 1915 4435
rect 1935 4415 1950 4435
rect 1900 4385 1950 4415
rect 1900 4365 1915 4385
rect 1935 4365 1950 4385
rect 1900 4350 1950 4365
rect 2050 4835 2100 4850
rect 2050 4815 2065 4835
rect 2085 4815 2100 4835
rect 2050 4785 2100 4815
rect 2050 4765 2065 4785
rect 2085 4765 2100 4785
rect 2050 4735 2100 4765
rect 2050 4715 2065 4735
rect 2085 4715 2100 4735
rect 2050 4685 2100 4715
rect 2050 4665 2065 4685
rect 2085 4665 2100 4685
rect 2050 4635 2100 4665
rect 2050 4615 2065 4635
rect 2085 4615 2100 4635
rect 2050 4585 2100 4615
rect 2050 4565 2065 4585
rect 2085 4565 2100 4585
rect 2050 4535 2100 4565
rect 2050 4515 2065 4535
rect 2085 4515 2100 4535
rect 2050 4485 2100 4515
rect 2050 4465 2065 4485
rect 2085 4465 2100 4485
rect 2050 4435 2100 4465
rect 2050 4415 2065 4435
rect 2085 4415 2100 4435
rect 2050 4385 2100 4415
rect 2050 4365 2065 4385
rect 2085 4365 2100 4385
rect 2050 4350 2100 4365
rect 2200 4835 2250 4850
rect 2200 4815 2215 4835
rect 2235 4815 2250 4835
rect 2200 4785 2250 4815
rect 2200 4765 2215 4785
rect 2235 4765 2250 4785
rect 2200 4735 2250 4765
rect 2200 4715 2215 4735
rect 2235 4715 2250 4735
rect 2200 4685 2250 4715
rect 2200 4665 2215 4685
rect 2235 4665 2250 4685
rect 2200 4635 2250 4665
rect 2200 4615 2215 4635
rect 2235 4615 2250 4635
rect 2200 4585 2250 4615
rect 2200 4565 2215 4585
rect 2235 4565 2250 4585
rect 2200 4535 2250 4565
rect 2200 4515 2215 4535
rect 2235 4515 2250 4535
rect 2200 4485 2250 4515
rect 2200 4465 2215 4485
rect 2235 4465 2250 4485
rect 2200 4435 2250 4465
rect 2200 4415 2215 4435
rect 2235 4415 2250 4435
rect 2200 4385 2250 4415
rect 2200 4365 2215 4385
rect 2235 4365 2250 4385
rect 2200 4350 2250 4365
rect 2350 4835 2400 4850
rect 2350 4815 2365 4835
rect 2385 4815 2400 4835
rect 2350 4785 2400 4815
rect 2350 4765 2365 4785
rect 2385 4765 2400 4785
rect 2350 4735 2400 4765
rect 2350 4715 2365 4735
rect 2385 4715 2400 4735
rect 2350 4685 2400 4715
rect 2350 4665 2365 4685
rect 2385 4665 2400 4685
rect 2350 4635 2400 4665
rect 2350 4615 2365 4635
rect 2385 4615 2400 4635
rect 2350 4585 2400 4615
rect 2350 4565 2365 4585
rect 2385 4565 2400 4585
rect 2350 4535 2400 4565
rect 2350 4515 2365 4535
rect 2385 4515 2400 4535
rect 2350 4485 2400 4515
rect 2350 4465 2365 4485
rect 2385 4465 2400 4485
rect 2350 4435 2400 4465
rect 2350 4415 2365 4435
rect 2385 4415 2400 4435
rect 2350 4385 2400 4415
rect 2350 4365 2365 4385
rect 2385 4365 2400 4385
rect 2350 4350 2400 4365
rect 2500 4835 2550 4850
rect 2500 4815 2515 4835
rect 2535 4815 2550 4835
rect 2500 4785 2550 4815
rect 2500 4765 2515 4785
rect 2535 4765 2550 4785
rect 2500 4735 2550 4765
rect 2500 4715 2515 4735
rect 2535 4715 2550 4735
rect 2500 4685 2550 4715
rect 2500 4665 2515 4685
rect 2535 4665 2550 4685
rect 2500 4635 2550 4665
rect 2500 4615 2515 4635
rect 2535 4615 2550 4635
rect 2500 4585 2550 4615
rect 2500 4565 2515 4585
rect 2535 4565 2550 4585
rect 2500 4535 2550 4565
rect 2500 4515 2515 4535
rect 2535 4515 2550 4535
rect 2500 4485 2550 4515
rect 2500 4465 2515 4485
rect 2535 4465 2550 4485
rect 2500 4435 2550 4465
rect 2500 4415 2515 4435
rect 2535 4415 2550 4435
rect 2500 4385 2550 4415
rect 2500 4365 2515 4385
rect 2535 4365 2550 4385
rect 2500 4350 2550 4365
rect 2650 4835 2700 4850
rect 2650 4815 2665 4835
rect 2685 4815 2700 4835
rect 2650 4785 2700 4815
rect 2650 4765 2665 4785
rect 2685 4765 2700 4785
rect 2650 4735 2700 4765
rect 2650 4715 2665 4735
rect 2685 4715 2700 4735
rect 2650 4685 2700 4715
rect 2650 4665 2665 4685
rect 2685 4665 2700 4685
rect 2650 4635 2700 4665
rect 2650 4615 2665 4635
rect 2685 4615 2700 4635
rect 2650 4585 2700 4615
rect 2650 4565 2665 4585
rect 2685 4565 2700 4585
rect 2650 4535 2700 4565
rect 2650 4515 2665 4535
rect 2685 4515 2700 4535
rect 2650 4485 2700 4515
rect 2650 4465 2665 4485
rect 2685 4465 2700 4485
rect 2650 4435 2700 4465
rect 2650 4415 2665 4435
rect 2685 4415 2700 4435
rect 2650 4385 2700 4415
rect 2650 4365 2665 4385
rect 2685 4365 2700 4385
rect 2650 4350 2700 4365
rect 2800 4835 2850 4850
rect 2800 4815 2815 4835
rect 2835 4815 2850 4835
rect 2800 4785 2850 4815
rect 2800 4765 2815 4785
rect 2835 4765 2850 4785
rect 2800 4735 2850 4765
rect 2800 4715 2815 4735
rect 2835 4715 2850 4735
rect 2800 4685 2850 4715
rect 2800 4665 2815 4685
rect 2835 4665 2850 4685
rect 2800 4635 2850 4665
rect 2800 4615 2815 4635
rect 2835 4615 2850 4635
rect 2800 4585 2850 4615
rect 2800 4565 2815 4585
rect 2835 4565 2850 4585
rect 2800 4535 2850 4565
rect 2800 4515 2815 4535
rect 2835 4515 2850 4535
rect 2800 4485 2850 4515
rect 2800 4465 2815 4485
rect 2835 4465 2850 4485
rect 2800 4435 2850 4465
rect 2800 4415 2815 4435
rect 2835 4415 2850 4435
rect 2800 4385 2850 4415
rect 2800 4365 2815 4385
rect 2835 4365 2850 4385
rect 2800 4350 2850 4365
rect 2950 4835 3000 4850
rect 2950 4815 2965 4835
rect 2985 4815 3000 4835
rect 2950 4785 3000 4815
rect 2950 4765 2965 4785
rect 2985 4765 3000 4785
rect 2950 4735 3000 4765
rect 2950 4715 2965 4735
rect 2985 4715 3000 4735
rect 2950 4685 3000 4715
rect 2950 4665 2965 4685
rect 2985 4665 3000 4685
rect 2950 4635 3000 4665
rect 2950 4615 2965 4635
rect 2985 4615 3000 4635
rect 2950 4585 3000 4615
rect 2950 4565 2965 4585
rect 2985 4565 3000 4585
rect 2950 4535 3000 4565
rect 2950 4515 2965 4535
rect 2985 4515 3000 4535
rect 2950 4485 3000 4515
rect 2950 4465 2965 4485
rect 2985 4465 3000 4485
rect 2950 4435 3000 4465
rect 2950 4415 2965 4435
rect 2985 4415 3000 4435
rect 2950 4385 3000 4415
rect 2950 4365 2965 4385
rect 2985 4365 3000 4385
rect 2950 4350 3000 4365
rect 3100 4835 3150 4850
rect 3100 4815 3115 4835
rect 3135 4815 3150 4835
rect 3100 4785 3150 4815
rect 3100 4765 3115 4785
rect 3135 4765 3150 4785
rect 3100 4735 3150 4765
rect 3100 4715 3115 4735
rect 3135 4715 3150 4735
rect 3100 4685 3150 4715
rect 3100 4665 3115 4685
rect 3135 4665 3150 4685
rect 3100 4635 3150 4665
rect 3100 4615 3115 4635
rect 3135 4615 3150 4635
rect 3100 4585 3150 4615
rect 3100 4565 3115 4585
rect 3135 4565 3150 4585
rect 3100 4535 3150 4565
rect 3100 4515 3115 4535
rect 3135 4515 3150 4535
rect 3100 4485 3150 4515
rect 3100 4465 3115 4485
rect 3135 4465 3150 4485
rect 3100 4435 3150 4465
rect 3100 4415 3115 4435
rect 3135 4415 3150 4435
rect 3100 4385 3150 4415
rect 3100 4365 3115 4385
rect 3135 4365 3150 4385
rect 3100 4350 3150 4365
rect 3250 4835 3300 4850
rect 3250 4815 3265 4835
rect 3285 4815 3300 4835
rect 3250 4785 3300 4815
rect 3250 4765 3265 4785
rect 3285 4765 3300 4785
rect 3250 4735 3300 4765
rect 3250 4715 3265 4735
rect 3285 4715 3300 4735
rect 3250 4685 3300 4715
rect 3250 4665 3265 4685
rect 3285 4665 3300 4685
rect 3250 4635 3300 4665
rect 3250 4615 3265 4635
rect 3285 4615 3300 4635
rect 3250 4585 3300 4615
rect 3250 4565 3265 4585
rect 3285 4565 3300 4585
rect 3250 4535 3300 4565
rect 3250 4515 3265 4535
rect 3285 4515 3300 4535
rect 3250 4485 3300 4515
rect 3250 4465 3265 4485
rect 3285 4465 3300 4485
rect 3250 4435 3300 4465
rect 3250 4415 3265 4435
rect 3285 4415 3300 4435
rect 3250 4385 3300 4415
rect 3250 4365 3265 4385
rect 3285 4365 3300 4385
rect 3250 4350 3300 4365
rect 3400 4835 3450 4850
rect 3400 4815 3415 4835
rect 3435 4815 3450 4835
rect 3400 4785 3450 4815
rect 3400 4765 3415 4785
rect 3435 4765 3450 4785
rect 3400 4735 3450 4765
rect 3400 4715 3415 4735
rect 3435 4715 3450 4735
rect 3400 4685 3450 4715
rect 3400 4665 3415 4685
rect 3435 4665 3450 4685
rect 3400 4635 3450 4665
rect 3400 4615 3415 4635
rect 3435 4615 3450 4635
rect 3400 4585 3450 4615
rect 3400 4565 3415 4585
rect 3435 4565 3450 4585
rect 3400 4535 3450 4565
rect 3400 4515 3415 4535
rect 3435 4515 3450 4535
rect 3400 4485 3450 4515
rect 3400 4465 3415 4485
rect 3435 4465 3450 4485
rect 3400 4435 3450 4465
rect 3400 4415 3415 4435
rect 3435 4415 3450 4435
rect 3400 4385 3450 4415
rect 3400 4365 3415 4385
rect 3435 4365 3450 4385
rect 3400 4350 3450 4365
rect 3550 4835 3600 4850
rect 3550 4815 3565 4835
rect 3585 4815 3600 4835
rect 3550 4785 3600 4815
rect 3550 4765 3565 4785
rect 3585 4765 3600 4785
rect 3550 4735 3600 4765
rect 3550 4715 3565 4735
rect 3585 4715 3600 4735
rect 3550 4685 3600 4715
rect 3550 4665 3565 4685
rect 3585 4665 3600 4685
rect 3550 4635 3600 4665
rect 3550 4615 3565 4635
rect 3585 4615 3600 4635
rect 3550 4585 3600 4615
rect 3550 4565 3565 4585
rect 3585 4565 3600 4585
rect 3550 4535 3600 4565
rect 3550 4515 3565 4535
rect 3585 4515 3600 4535
rect 3550 4485 3600 4515
rect 3550 4465 3565 4485
rect 3585 4465 3600 4485
rect 3550 4435 3600 4465
rect 3550 4415 3565 4435
rect 3585 4415 3600 4435
rect 3550 4385 3600 4415
rect 3550 4365 3565 4385
rect 3585 4365 3600 4385
rect 3550 4350 3600 4365
rect 3700 4350 3750 4850
rect 3850 4350 3900 4850
rect 4000 4350 4050 4850
rect 4150 4835 4200 4850
rect 4150 4815 4165 4835
rect 4185 4815 4200 4835
rect 4150 4785 4200 4815
rect 4150 4765 4165 4785
rect 4185 4765 4200 4785
rect 4150 4735 4200 4765
rect 4150 4715 4165 4735
rect 4185 4715 4200 4735
rect 4150 4685 4200 4715
rect 4150 4665 4165 4685
rect 4185 4665 4200 4685
rect 4150 4635 4200 4665
rect 4150 4615 4165 4635
rect 4185 4615 4200 4635
rect 4150 4585 4200 4615
rect 4150 4565 4165 4585
rect 4185 4565 4200 4585
rect 4150 4535 4200 4565
rect 4150 4515 4165 4535
rect 4185 4515 4200 4535
rect 4150 4485 4200 4515
rect 4150 4465 4165 4485
rect 4185 4465 4200 4485
rect 4150 4435 4200 4465
rect 4150 4415 4165 4435
rect 4185 4415 4200 4435
rect 4150 4385 4200 4415
rect 4150 4365 4165 4385
rect 4185 4365 4200 4385
rect 4150 4350 4200 4365
rect 4300 4350 4350 4850
rect 4450 4350 4500 4850
rect 4600 4350 4650 4850
rect 4750 4835 4800 4850
rect 4750 4815 4765 4835
rect 4785 4815 4800 4835
rect 4750 4785 4800 4815
rect 4750 4765 4765 4785
rect 4785 4765 4800 4785
rect 4750 4735 4800 4765
rect 4750 4715 4765 4735
rect 4785 4715 4800 4735
rect 4750 4685 4800 4715
rect 4750 4665 4765 4685
rect 4785 4665 4800 4685
rect 4750 4635 4800 4665
rect 4750 4615 4765 4635
rect 4785 4615 4800 4635
rect 4750 4585 4800 4615
rect 4750 4565 4765 4585
rect 4785 4565 4800 4585
rect 4750 4535 4800 4565
rect 4750 4515 4765 4535
rect 4785 4515 4800 4535
rect 4750 4485 4800 4515
rect 4750 4465 4765 4485
rect 4785 4465 4800 4485
rect 4750 4435 4800 4465
rect 4750 4415 4765 4435
rect 4785 4415 4800 4435
rect 4750 4385 4800 4415
rect 4750 4365 4765 4385
rect 4785 4365 4800 4385
rect 4750 4350 4800 4365
rect 4900 4835 4950 4850
rect 4900 4815 4915 4835
rect 4935 4815 4950 4835
rect 4900 4785 4950 4815
rect 4900 4765 4915 4785
rect 4935 4765 4950 4785
rect 4900 4735 4950 4765
rect 4900 4715 4915 4735
rect 4935 4715 4950 4735
rect 4900 4685 4950 4715
rect 4900 4665 4915 4685
rect 4935 4665 4950 4685
rect 4900 4635 4950 4665
rect 4900 4615 4915 4635
rect 4935 4615 4950 4635
rect 4900 4585 4950 4615
rect 4900 4565 4915 4585
rect 4935 4565 4950 4585
rect 4900 4535 4950 4565
rect 4900 4515 4915 4535
rect 4935 4515 4950 4535
rect 4900 4485 4950 4515
rect 4900 4465 4915 4485
rect 4935 4465 4950 4485
rect 4900 4435 4950 4465
rect 4900 4415 4915 4435
rect 4935 4415 4950 4435
rect 4900 4385 4950 4415
rect 4900 4365 4915 4385
rect 4935 4365 4950 4385
rect 4900 4350 4950 4365
rect 5050 4835 5100 4850
rect 5050 4815 5065 4835
rect 5085 4815 5100 4835
rect 5050 4785 5100 4815
rect 5050 4765 5065 4785
rect 5085 4765 5100 4785
rect 5050 4735 5100 4765
rect 5050 4715 5065 4735
rect 5085 4715 5100 4735
rect 5050 4685 5100 4715
rect 5050 4665 5065 4685
rect 5085 4665 5100 4685
rect 5050 4635 5100 4665
rect 5050 4615 5065 4635
rect 5085 4615 5100 4635
rect 5050 4585 5100 4615
rect 5050 4565 5065 4585
rect 5085 4565 5100 4585
rect 5050 4535 5100 4565
rect 5050 4515 5065 4535
rect 5085 4515 5100 4535
rect 5050 4485 5100 4515
rect 5050 4465 5065 4485
rect 5085 4465 5100 4485
rect 5050 4435 5100 4465
rect 5050 4415 5065 4435
rect 5085 4415 5100 4435
rect 5050 4385 5100 4415
rect 5050 4365 5065 4385
rect 5085 4365 5100 4385
rect 5050 4350 5100 4365
rect 5200 4835 5250 4850
rect 5200 4815 5215 4835
rect 5235 4815 5250 4835
rect 5200 4785 5250 4815
rect 5200 4765 5215 4785
rect 5235 4765 5250 4785
rect 5200 4735 5250 4765
rect 5200 4715 5215 4735
rect 5235 4715 5250 4735
rect 5200 4685 5250 4715
rect 5200 4665 5215 4685
rect 5235 4665 5250 4685
rect 5200 4635 5250 4665
rect 5200 4615 5215 4635
rect 5235 4615 5250 4635
rect 5200 4585 5250 4615
rect 5200 4565 5215 4585
rect 5235 4565 5250 4585
rect 5200 4535 5250 4565
rect 5200 4515 5215 4535
rect 5235 4515 5250 4535
rect 5200 4485 5250 4515
rect 5200 4465 5215 4485
rect 5235 4465 5250 4485
rect 5200 4435 5250 4465
rect 5200 4415 5215 4435
rect 5235 4415 5250 4435
rect 5200 4385 5250 4415
rect 5200 4365 5215 4385
rect 5235 4365 5250 4385
rect 5200 4350 5250 4365
rect 5350 4835 5400 4850
rect 5350 4815 5365 4835
rect 5385 4815 5400 4835
rect 5350 4785 5400 4815
rect 5350 4765 5365 4785
rect 5385 4765 5400 4785
rect 5350 4735 5400 4765
rect 5350 4715 5365 4735
rect 5385 4715 5400 4735
rect 5350 4685 5400 4715
rect 5350 4665 5365 4685
rect 5385 4665 5400 4685
rect 5350 4635 5400 4665
rect 5350 4615 5365 4635
rect 5385 4615 5400 4635
rect 5350 4585 5400 4615
rect 5350 4565 5365 4585
rect 5385 4565 5400 4585
rect 5350 4535 5400 4565
rect 5350 4515 5365 4535
rect 5385 4515 5400 4535
rect 5350 4485 5400 4515
rect 5350 4465 5365 4485
rect 5385 4465 5400 4485
rect 5350 4435 5400 4465
rect 5350 4415 5365 4435
rect 5385 4415 5400 4435
rect 5350 4385 5400 4415
rect 5350 4365 5365 4385
rect 5385 4365 5400 4385
rect 5350 4350 5400 4365
rect 5500 4835 5550 4850
rect 5500 4815 5515 4835
rect 5535 4815 5550 4835
rect 5500 4785 5550 4815
rect 5500 4765 5515 4785
rect 5535 4765 5550 4785
rect 5500 4735 5550 4765
rect 5500 4715 5515 4735
rect 5535 4715 5550 4735
rect 5500 4685 5550 4715
rect 5500 4665 5515 4685
rect 5535 4665 5550 4685
rect 5500 4635 5550 4665
rect 5500 4615 5515 4635
rect 5535 4615 5550 4635
rect 5500 4585 5550 4615
rect 5500 4565 5515 4585
rect 5535 4565 5550 4585
rect 5500 4535 5550 4565
rect 5500 4515 5515 4535
rect 5535 4515 5550 4535
rect 5500 4485 5550 4515
rect 5500 4465 5515 4485
rect 5535 4465 5550 4485
rect 5500 4435 5550 4465
rect 5500 4415 5515 4435
rect 5535 4415 5550 4435
rect 5500 4385 5550 4415
rect 5500 4365 5515 4385
rect 5535 4365 5550 4385
rect 5500 4350 5550 4365
rect 5650 4835 5700 4850
rect 5650 4815 5665 4835
rect 5685 4815 5700 4835
rect 5650 4785 5700 4815
rect 5650 4765 5665 4785
rect 5685 4765 5700 4785
rect 5650 4735 5700 4765
rect 5650 4715 5665 4735
rect 5685 4715 5700 4735
rect 5650 4685 5700 4715
rect 5650 4665 5665 4685
rect 5685 4665 5700 4685
rect 5650 4635 5700 4665
rect 5650 4615 5665 4635
rect 5685 4615 5700 4635
rect 5650 4585 5700 4615
rect 5650 4565 5665 4585
rect 5685 4565 5700 4585
rect 5650 4535 5700 4565
rect 5650 4515 5665 4535
rect 5685 4515 5700 4535
rect 5650 4485 5700 4515
rect 5650 4465 5665 4485
rect 5685 4465 5700 4485
rect 5650 4435 5700 4465
rect 5650 4415 5665 4435
rect 5685 4415 5700 4435
rect 5650 4385 5700 4415
rect 5650 4365 5665 4385
rect 5685 4365 5700 4385
rect 5650 4350 5700 4365
rect 5800 4835 5850 4850
rect 5800 4815 5815 4835
rect 5835 4815 5850 4835
rect 5800 4785 5850 4815
rect 5800 4765 5815 4785
rect 5835 4765 5850 4785
rect 5800 4735 5850 4765
rect 5800 4715 5815 4735
rect 5835 4715 5850 4735
rect 5800 4685 5850 4715
rect 5800 4665 5815 4685
rect 5835 4665 5850 4685
rect 5800 4635 5850 4665
rect 5800 4615 5815 4635
rect 5835 4615 5850 4635
rect 5800 4585 5850 4615
rect 5800 4565 5815 4585
rect 5835 4565 5850 4585
rect 5800 4535 5850 4565
rect 5800 4515 5815 4535
rect 5835 4515 5850 4535
rect 5800 4485 5850 4515
rect 5800 4465 5815 4485
rect 5835 4465 5850 4485
rect 5800 4435 5850 4465
rect 5800 4415 5815 4435
rect 5835 4415 5850 4435
rect 5800 4385 5850 4415
rect 5800 4365 5815 4385
rect 5835 4365 5850 4385
rect 5800 4350 5850 4365
rect 5950 4835 6000 4850
rect 5950 4815 5965 4835
rect 5985 4815 6000 4835
rect 5950 4785 6000 4815
rect 5950 4765 5965 4785
rect 5985 4765 6000 4785
rect 5950 4735 6000 4765
rect 5950 4715 5965 4735
rect 5985 4715 6000 4735
rect 5950 4685 6000 4715
rect 5950 4665 5965 4685
rect 5985 4665 6000 4685
rect 5950 4635 6000 4665
rect 5950 4615 5965 4635
rect 5985 4615 6000 4635
rect 5950 4585 6000 4615
rect 5950 4565 5965 4585
rect 5985 4565 6000 4585
rect 5950 4535 6000 4565
rect 5950 4515 5965 4535
rect 5985 4515 6000 4535
rect 5950 4485 6000 4515
rect 5950 4465 5965 4485
rect 5985 4465 6000 4485
rect 5950 4435 6000 4465
rect 5950 4415 5965 4435
rect 5985 4415 6000 4435
rect 5950 4385 6000 4415
rect 5950 4365 5965 4385
rect 5985 4365 6000 4385
rect 5950 4350 6000 4365
rect 6100 4835 6150 4850
rect 6100 4815 6115 4835
rect 6135 4815 6150 4835
rect 6100 4785 6150 4815
rect 6100 4765 6115 4785
rect 6135 4765 6150 4785
rect 6100 4735 6150 4765
rect 6100 4715 6115 4735
rect 6135 4715 6150 4735
rect 6100 4685 6150 4715
rect 6100 4665 6115 4685
rect 6135 4665 6150 4685
rect 6100 4635 6150 4665
rect 6100 4615 6115 4635
rect 6135 4615 6150 4635
rect 6100 4585 6150 4615
rect 6100 4565 6115 4585
rect 6135 4565 6150 4585
rect 6100 4535 6150 4565
rect 6100 4515 6115 4535
rect 6135 4515 6150 4535
rect 6100 4485 6150 4515
rect 6100 4465 6115 4485
rect 6135 4465 6150 4485
rect 6100 4435 6150 4465
rect 6100 4415 6115 4435
rect 6135 4415 6150 4435
rect 6100 4385 6150 4415
rect 6100 4365 6115 4385
rect 6135 4365 6150 4385
rect 6100 4350 6150 4365
rect 6250 4835 6300 4850
rect 6250 4815 6265 4835
rect 6285 4815 6300 4835
rect 6250 4785 6300 4815
rect 6250 4765 6265 4785
rect 6285 4765 6300 4785
rect 6250 4735 6300 4765
rect 6250 4715 6265 4735
rect 6285 4715 6300 4735
rect 6250 4685 6300 4715
rect 6250 4665 6265 4685
rect 6285 4665 6300 4685
rect 6250 4635 6300 4665
rect 6250 4615 6265 4635
rect 6285 4615 6300 4635
rect 6250 4585 6300 4615
rect 6250 4565 6265 4585
rect 6285 4565 6300 4585
rect 6250 4535 6300 4565
rect 6250 4515 6265 4535
rect 6285 4515 6300 4535
rect 6250 4485 6300 4515
rect 6250 4465 6265 4485
rect 6285 4465 6300 4485
rect 6250 4435 6300 4465
rect 6250 4415 6265 4435
rect 6285 4415 6300 4435
rect 6250 4385 6300 4415
rect 6250 4365 6265 4385
rect 6285 4365 6300 4385
rect 6250 4350 6300 4365
rect 6400 4835 6450 4850
rect 6400 4815 6415 4835
rect 6435 4815 6450 4835
rect 6400 4785 6450 4815
rect 6400 4765 6415 4785
rect 6435 4765 6450 4785
rect 6400 4735 6450 4765
rect 6400 4715 6415 4735
rect 6435 4715 6450 4735
rect 6400 4685 6450 4715
rect 6400 4665 6415 4685
rect 6435 4665 6450 4685
rect 6400 4635 6450 4665
rect 6400 4615 6415 4635
rect 6435 4615 6450 4635
rect 6400 4585 6450 4615
rect 6400 4565 6415 4585
rect 6435 4565 6450 4585
rect 6400 4535 6450 4565
rect 6400 4515 6415 4535
rect 6435 4515 6450 4535
rect 6400 4485 6450 4515
rect 6400 4465 6415 4485
rect 6435 4465 6450 4485
rect 6400 4435 6450 4465
rect 6400 4415 6415 4435
rect 6435 4415 6450 4435
rect 6400 4385 6450 4415
rect 6400 4365 6415 4385
rect 6435 4365 6450 4385
rect 6400 4350 6450 4365
rect 6550 4835 6600 4850
rect 6550 4815 6565 4835
rect 6585 4815 6600 4835
rect 6550 4785 6600 4815
rect 6550 4765 6565 4785
rect 6585 4765 6600 4785
rect 6550 4735 6600 4765
rect 6550 4715 6565 4735
rect 6585 4715 6600 4735
rect 6550 4685 6600 4715
rect 6550 4665 6565 4685
rect 6585 4665 6600 4685
rect 6550 4635 6600 4665
rect 6550 4615 6565 4635
rect 6585 4615 6600 4635
rect 6550 4585 6600 4615
rect 6550 4565 6565 4585
rect 6585 4565 6600 4585
rect 6550 4535 6600 4565
rect 6550 4515 6565 4535
rect 6585 4515 6600 4535
rect 6550 4485 6600 4515
rect 6550 4465 6565 4485
rect 6585 4465 6600 4485
rect 6550 4435 6600 4465
rect 6550 4415 6565 4435
rect 6585 4415 6600 4435
rect 6550 4385 6600 4415
rect 6550 4365 6565 4385
rect 6585 4365 6600 4385
rect 6550 4350 6600 4365
rect 6700 4835 6750 4850
rect 6700 4815 6715 4835
rect 6735 4815 6750 4835
rect 6700 4785 6750 4815
rect 6700 4765 6715 4785
rect 6735 4765 6750 4785
rect 6700 4735 6750 4765
rect 6700 4715 6715 4735
rect 6735 4715 6750 4735
rect 6700 4685 6750 4715
rect 6700 4665 6715 4685
rect 6735 4665 6750 4685
rect 6700 4635 6750 4665
rect 6700 4615 6715 4635
rect 6735 4615 6750 4635
rect 6700 4585 6750 4615
rect 6700 4565 6715 4585
rect 6735 4565 6750 4585
rect 6700 4535 6750 4565
rect 6700 4515 6715 4535
rect 6735 4515 6750 4535
rect 6700 4485 6750 4515
rect 6700 4465 6715 4485
rect 6735 4465 6750 4485
rect 6700 4435 6750 4465
rect 6700 4415 6715 4435
rect 6735 4415 6750 4435
rect 6700 4385 6750 4415
rect 6700 4365 6715 4385
rect 6735 4365 6750 4385
rect 6700 4350 6750 4365
rect 6850 4835 6900 4850
rect 6850 4815 6865 4835
rect 6885 4815 6900 4835
rect 6850 4785 6900 4815
rect 6850 4765 6865 4785
rect 6885 4765 6900 4785
rect 6850 4735 6900 4765
rect 6850 4715 6865 4735
rect 6885 4715 6900 4735
rect 6850 4685 6900 4715
rect 6850 4665 6865 4685
rect 6885 4665 6900 4685
rect 6850 4635 6900 4665
rect 6850 4615 6865 4635
rect 6885 4615 6900 4635
rect 6850 4585 6900 4615
rect 6850 4565 6865 4585
rect 6885 4565 6900 4585
rect 6850 4535 6900 4565
rect 6850 4515 6865 4535
rect 6885 4515 6900 4535
rect 6850 4485 6900 4515
rect 6850 4465 6865 4485
rect 6885 4465 6900 4485
rect 6850 4435 6900 4465
rect 6850 4415 6865 4435
rect 6885 4415 6900 4435
rect 6850 4385 6900 4415
rect 6850 4365 6865 4385
rect 6885 4365 6900 4385
rect 6850 4350 6900 4365
rect 7000 4835 7050 4850
rect 7000 4815 7015 4835
rect 7035 4815 7050 4835
rect 7000 4785 7050 4815
rect 7000 4765 7015 4785
rect 7035 4765 7050 4785
rect 7000 4735 7050 4765
rect 7000 4715 7015 4735
rect 7035 4715 7050 4735
rect 7000 4685 7050 4715
rect 7000 4665 7015 4685
rect 7035 4665 7050 4685
rect 7000 4635 7050 4665
rect 7000 4615 7015 4635
rect 7035 4615 7050 4635
rect 7000 4585 7050 4615
rect 7000 4565 7015 4585
rect 7035 4565 7050 4585
rect 7000 4535 7050 4565
rect 7000 4515 7015 4535
rect 7035 4515 7050 4535
rect 7000 4485 7050 4515
rect 7000 4465 7015 4485
rect 7035 4465 7050 4485
rect 7000 4435 7050 4465
rect 7000 4415 7015 4435
rect 7035 4415 7050 4435
rect 7000 4385 7050 4415
rect 7000 4365 7015 4385
rect 7035 4365 7050 4385
rect 7000 4350 7050 4365
rect 7150 4835 7200 4850
rect 7150 4815 7165 4835
rect 7185 4815 7200 4835
rect 7150 4785 7200 4815
rect 7150 4765 7165 4785
rect 7185 4765 7200 4785
rect 7150 4735 7200 4765
rect 7150 4715 7165 4735
rect 7185 4715 7200 4735
rect 7150 4685 7200 4715
rect 7150 4665 7165 4685
rect 7185 4665 7200 4685
rect 7150 4635 7200 4665
rect 7150 4615 7165 4635
rect 7185 4615 7200 4635
rect 7150 4585 7200 4615
rect 7150 4565 7165 4585
rect 7185 4565 7200 4585
rect 7150 4535 7200 4565
rect 7150 4515 7165 4535
rect 7185 4515 7200 4535
rect 7150 4485 7200 4515
rect 7150 4465 7165 4485
rect 7185 4465 7200 4485
rect 7150 4435 7200 4465
rect 7150 4415 7165 4435
rect 7185 4415 7200 4435
rect 7150 4385 7200 4415
rect 7150 4365 7165 4385
rect 7185 4365 7200 4385
rect 7150 4350 7200 4365
rect 7300 4835 7350 4850
rect 7300 4815 7315 4835
rect 7335 4815 7350 4835
rect 7300 4785 7350 4815
rect 7300 4765 7315 4785
rect 7335 4765 7350 4785
rect 7300 4735 7350 4765
rect 7300 4715 7315 4735
rect 7335 4715 7350 4735
rect 7300 4685 7350 4715
rect 7300 4665 7315 4685
rect 7335 4665 7350 4685
rect 7300 4635 7350 4665
rect 7300 4615 7315 4635
rect 7335 4615 7350 4635
rect 7300 4585 7350 4615
rect 7300 4565 7315 4585
rect 7335 4565 7350 4585
rect 7300 4535 7350 4565
rect 7300 4515 7315 4535
rect 7335 4515 7350 4535
rect 7300 4485 7350 4515
rect 7300 4465 7315 4485
rect 7335 4465 7350 4485
rect 7300 4435 7350 4465
rect 7300 4415 7315 4435
rect 7335 4415 7350 4435
rect 7300 4385 7350 4415
rect 7300 4365 7315 4385
rect 7335 4365 7350 4385
rect 7300 4350 7350 4365
rect 7450 4835 7500 4850
rect 7450 4815 7465 4835
rect 7485 4815 7500 4835
rect 7450 4785 7500 4815
rect 7450 4765 7465 4785
rect 7485 4765 7500 4785
rect 7450 4735 7500 4765
rect 7450 4715 7465 4735
rect 7485 4715 7500 4735
rect 7450 4685 7500 4715
rect 7450 4665 7465 4685
rect 7485 4665 7500 4685
rect 7450 4635 7500 4665
rect 7450 4615 7465 4635
rect 7485 4615 7500 4635
rect 7450 4585 7500 4615
rect 7450 4565 7465 4585
rect 7485 4565 7500 4585
rect 7450 4535 7500 4565
rect 7450 4515 7465 4535
rect 7485 4515 7500 4535
rect 7450 4485 7500 4515
rect 7450 4465 7465 4485
rect 7485 4465 7500 4485
rect 7450 4435 7500 4465
rect 7450 4415 7465 4435
rect 7485 4415 7500 4435
rect 7450 4385 7500 4415
rect 7450 4365 7465 4385
rect 7485 4365 7500 4385
rect 7450 4350 7500 4365
rect 7600 4835 7650 4850
rect 7600 4815 7615 4835
rect 7635 4815 7650 4835
rect 7600 4785 7650 4815
rect 7600 4765 7615 4785
rect 7635 4765 7650 4785
rect 7600 4735 7650 4765
rect 7600 4715 7615 4735
rect 7635 4715 7650 4735
rect 7600 4685 7650 4715
rect 7600 4665 7615 4685
rect 7635 4665 7650 4685
rect 7600 4635 7650 4665
rect 7600 4615 7615 4635
rect 7635 4615 7650 4635
rect 7600 4585 7650 4615
rect 7600 4565 7615 4585
rect 7635 4565 7650 4585
rect 7600 4535 7650 4565
rect 7600 4515 7615 4535
rect 7635 4515 7650 4535
rect 7600 4485 7650 4515
rect 7600 4465 7615 4485
rect 7635 4465 7650 4485
rect 7600 4435 7650 4465
rect 7600 4415 7615 4435
rect 7635 4415 7650 4435
rect 7600 4385 7650 4415
rect 7600 4365 7615 4385
rect 7635 4365 7650 4385
rect 7600 4350 7650 4365
rect 7750 4835 7800 4850
rect 7750 4815 7765 4835
rect 7785 4815 7800 4835
rect 7750 4785 7800 4815
rect 7750 4765 7765 4785
rect 7785 4765 7800 4785
rect 7750 4735 7800 4765
rect 7750 4715 7765 4735
rect 7785 4715 7800 4735
rect 7750 4685 7800 4715
rect 7750 4665 7765 4685
rect 7785 4665 7800 4685
rect 7750 4635 7800 4665
rect 7750 4615 7765 4635
rect 7785 4615 7800 4635
rect 7750 4585 7800 4615
rect 7750 4565 7765 4585
rect 7785 4565 7800 4585
rect 7750 4535 7800 4565
rect 7750 4515 7765 4535
rect 7785 4515 7800 4535
rect 7750 4485 7800 4515
rect 7750 4465 7765 4485
rect 7785 4465 7800 4485
rect 7750 4435 7800 4465
rect 7750 4415 7765 4435
rect 7785 4415 7800 4435
rect 7750 4385 7800 4415
rect 7750 4365 7765 4385
rect 7785 4365 7800 4385
rect 7750 4350 7800 4365
rect 7900 4350 7950 4850
rect 8050 4350 8100 4850
rect 8200 4350 8250 4850
rect 8350 4835 8400 4850
rect 8350 4815 8365 4835
rect 8385 4815 8400 4835
rect 8350 4785 8400 4815
rect 8350 4765 8365 4785
rect 8385 4765 8400 4785
rect 8350 4735 8400 4765
rect 8350 4715 8365 4735
rect 8385 4715 8400 4735
rect 8350 4685 8400 4715
rect 8350 4665 8365 4685
rect 8385 4665 8400 4685
rect 8350 4635 8400 4665
rect 8350 4615 8365 4635
rect 8385 4615 8400 4635
rect 8350 4585 8400 4615
rect 8350 4565 8365 4585
rect 8385 4565 8400 4585
rect 8350 4535 8400 4565
rect 8350 4515 8365 4535
rect 8385 4515 8400 4535
rect 8350 4485 8400 4515
rect 8350 4465 8365 4485
rect 8385 4465 8400 4485
rect 8350 4435 8400 4465
rect 8350 4415 8365 4435
rect 8385 4415 8400 4435
rect 8350 4385 8400 4415
rect 8350 4365 8365 4385
rect 8385 4365 8400 4385
rect 8350 4350 8400 4365
rect 8500 4835 8550 4850
rect 8500 4815 8515 4835
rect 8535 4815 8550 4835
rect 8500 4785 8550 4815
rect 8500 4765 8515 4785
rect 8535 4765 8550 4785
rect 8500 4735 8550 4765
rect 8500 4715 8515 4735
rect 8535 4715 8550 4735
rect 8500 4685 8550 4715
rect 8500 4665 8515 4685
rect 8535 4665 8550 4685
rect 8500 4635 8550 4665
rect 8500 4615 8515 4635
rect 8535 4615 8550 4635
rect 8500 4585 8550 4615
rect 8500 4565 8515 4585
rect 8535 4565 8550 4585
rect 8500 4535 8550 4565
rect 8500 4515 8515 4535
rect 8535 4515 8550 4535
rect 8500 4485 8550 4515
rect 8500 4465 8515 4485
rect 8535 4465 8550 4485
rect 8500 4435 8550 4465
rect 8500 4415 8515 4435
rect 8535 4415 8550 4435
rect 8500 4385 8550 4415
rect 8500 4365 8515 4385
rect 8535 4365 8550 4385
rect 8500 4350 8550 4365
rect 8650 4835 8700 4850
rect 8650 4815 8665 4835
rect 8685 4815 8700 4835
rect 8650 4785 8700 4815
rect 8650 4765 8665 4785
rect 8685 4765 8700 4785
rect 8650 4735 8700 4765
rect 8650 4715 8665 4735
rect 8685 4715 8700 4735
rect 8650 4685 8700 4715
rect 8650 4665 8665 4685
rect 8685 4665 8700 4685
rect 8650 4635 8700 4665
rect 8650 4615 8665 4635
rect 8685 4615 8700 4635
rect 8650 4585 8700 4615
rect 8650 4565 8665 4585
rect 8685 4565 8700 4585
rect 8650 4535 8700 4565
rect 8650 4515 8665 4535
rect 8685 4515 8700 4535
rect 8650 4485 8700 4515
rect 8650 4465 8665 4485
rect 8685 4465 8700 4485
rect 8650 4435 8700 4465
rect 8650 4415 8665 4435
rect 8685 4415 8700 4435
rect 8650 4385 8700 4415
rect 8650 4365 8665 4385
rect 8685 4365 8700 4385
rect 8650 4350 8700 4365
rect 8800 4835 8850 4850
rect 8800 4815 8815 4835
rect 8835 4815 8850 4835
rect 8800 4785 8850 4815
rect 8800 4765 8815 4785
rect 8835 4765 8850 4785
rect 8800 4735 8850 4765
rect 8800 4715 8815 4735
rect 8835 4715 8850 4735
rect 8800 4685 8850 4715
rect 8800 4665 8815 4685
rect 8835 4665 8850 4685
rect 8800 4635 8850 4665
rect 8800 4615 8815 4635
rect 8835 4615 8850 4635
rect 8800 4585 8850 4615
rect 8800 4565 8815 4585
rect 8835 4565 8850 4585
rect 8800 4535 8850 4565
rect 8800 4515 8815 4535
rect 8835 4515 8850 4535
rect 8800 4485 8850 4515
rect 8800 4465 8815 4485
rect 8835 4465 8850 4485
rect 8800 4435 8850 4465
rect 8800 4415 8815 4435
rect 8835 4415 8850 4435
rect 8800 4385 8850 4415
rect 8800 4365 8815 4385
rect 8835 4365 8850 4385
rect 8800 4350 8850 4365
rect 8950 4835 9000 4850
rect 8950 4815 8965 4835
rect 8985 4815 9000 4835
rect 8950 4785 9000 4815
rect 8950 4765 8965 4785
rect 8985 4765 9000 4785
rect 8950 4735 9000 4765
rect 8950 4715 8965 4735
rect 8985 4715 9000 4735
rect 8950 4685 9000 4715
rect 8950 4665 8965 4685
rect 8985 4665 9000 4685
rect 8950 4635 9000 4665
rect 8950 4615 8965 4635
rect 8985 4615 9000 4635
rect 8950 4585 9000 4615
rect 8950 4565 8965 4585
rect 8985 4565 9000 4585
rect 8950 4535 9000 4565
rect 8950 4515 8965 4535
rect 8985 4515 9000 4535
rect 8950 4485 9000 4515
rect 8950 4465 8965 4485
rect 8985 4465 9000 4485
rect 8950 4435 9000 4465
rect 8950 4415 8965 4435
rect 8985 4415 9000 4435
rect 8950 4385 9000 4415
rect 8950 4365 8965 4385
rect 8985 4365 9000 4385
rect 8950 4350 9000 4365
rect 9100 4835 9150 4850
rect 9100 4815 9115 4835
rect 9135 4815 9150 4835
rect 9100 4785 9150 4815
rect 9100 4765 9115 4785
rect 9135 4765 9150 4785
rect 9100 4735 9150 4765
rect 9100 4715 9115 4735
rect 9135 4715 9150 4735
rect 9100 4685 9150 4715
rect 9100 4665 9115 4685
rect 9135 4665 9150 4685
rect 9100 4635 9150 4665
rect 9100 4615 9115 4635
rect 9135 4615 9150 4635
rect 9100 4585 9150 4615
rect 9100 4565 9115 4585
rect 9135 4565 9150 4585
rect 9100 4535 9150 4565
rect 9100 4515 9115 4535
rect 9135 4515 9150 4535
rect 9100 4485 9150 4515
rect 9100 4465 9115 4485
rect 9135 4465 9150 4485
rect 9100 4435 9150 4465
rect 9100 4415 9115 4435
rect 9135 4415 9150 4435
rect 9100 4385 9150 4415
rect 9100 4365 9115 4385
rect 9135 4365 9150 4385
rect 9100 4350 9150 4365
rect 9250 4835 9300 4850
rect 9250 4815 9265 4835
rect 9285 4815 9300 4835
rect 9250 4785 9300 4815
rect 9250 4765 9265 4785
rect 9285 4765 9300 4785
rect 9250 4735 9300 4765
rect 9250 4715 9265 4735
rect 9285 4715 9300 4735
rect 9250 4685 9300 4715
rect 9250 4665 9265 4685
rect 9285 4665 9300 4685
rect 9250 4635 9300 4665
rect 9250 4615 9265 4635
rect 9285 4615 9300 4635
rect 9250 4585 9300 4615
rect 9250 4565 9265 4585
rect 9285 4565 9300 4585
rect 9250 4535 9300 4565
rect 9250 4515 9265 4535
rect 9285 4515 9300 4535
rect 9250 4485 9300 4515
rect 9250 4465 9265 4485
rect 9285 4465 9300 4485
rect 9250 4435 9300 4465
rect 9250 4415 9265 4435
rect 9285 4415 9300 4435
rect 9250 4385 9300 4415
rect 9250 4365 9265 4385
rect 9285 4365 9300 4385
rect 9250 4350 9300 4365
rect 9400 4835 9450 4850
rect 9400 4815 9415 4835
rect 9435 4815 9450 4835
rect 9400 4785 9450 4815
rect 9400 4765 9415 4785
rect 9435 4765 9450 4785
rect 9400 4735 9450 4765
rect 9400 4715 9415 4735
rect 9435 4715 9450 4735
rect 9400 4685 9450 4715
rect 9400 4665 9415 4685
rect 9435 4665 9450 4685
rect 9400 4635 9450 4665
rect 9400 4615 9415 4635
rect 9435 4615 9450 4635
rect 9400 4585 9450 4615
rect 9400 4565 9415 4585
rect 9435 4565 9450 4585
rect 9400 4535 9450 4565
rect 9400 4515 9415 4535
rect 9435 4515 9450 4535
rect 9400 4485 9450 4515
rect 9400 4465 9415 4485
rect 9435 4465 9450 4485
rect 9400 4435 9450 4465
rect 9400 4415 9415 4435
rect 9435 4415 9450 4435
rect 9400 4385 9450 4415
rect 9400 4365 9415 4385
rect 9435 4365 9450 4385
rect 9400 4350 9450 4365
rect 9550 4835 9600 4850
rect 9550 4815 9565 4835
rect 9585 4815 9600 4835
rect 9550 4785 9600 4815
rect 9550 4765 9565 4785
rect 9585 4765 9600 4785
rect 9550 4735 9600 4765
rect 9550 4715 9565 4735
rect 9585 4715 9600 4735
rect 9550 4685 9600 4715
rect 9550 4665 9565 4685
rect 9585 4665 9600 4685
rect 9550 4635 9600 4665
rect 9550 4615 9565 4635
rect 9585 4615 9600 4635
rect 9550 4585 9600 4615
rect 9550 4565 9565 4585
rect 9585 4565 9600 4585
rect 9550 4535 9600 4565
rect 9550 4515 9565 4535
rect 9585 4515 9600 4535
rect 9550 4485 9600 4515
rect 9550 4465 9565 4485
rect 9585 4465 9600 4485
rect 9550 4435 9600 4465
rect 9550 4415 9565 4435
rect 9585 4415 9600 4435
rect 9550 4385 9600 4415
rect 9550 4365 9565 4385
rect 9585 4365 9600 4385
rect 9550 4350 9600 4365
rect 9700 4835 9750 4850
rect 9700 4815 9715 4835
rect 9735 4815 9750 4835
rect 9700 4785 9750 4815
rect 9700 4765 9715 4785
rect 9735 4765 9750 4785
rect 9700 4735 9750 4765
rect 9700 4715 9715 4735
rect 9735 4715 9750 4735
rect 9700 4685 9750 4715
rect 9700 4665 9715 4685
rect 9735 4665 9750 4685
rect 9700 4635 9750 4665
rect 9700 4615 9715 4635
rect 9735 4615 9750 4635
rect 9700 4585 9750 4615
rect 9700 4565 9715 4585
rect 9735 4565 9750 4585
rect 9700 4535 9750 4565
rect 9700 4515 9715 4535
rect 9735 4515 9750 4535
rect 9700 4485 9750 4515
rect 9700 4465 9715 4485
rect 9735 4465 9750 4485
rect 9700 4435 9750 4465
rect 9700 4415 9715 4435
rect 9735 4415 9750 4435
rect 9700 4385 9750 4415
rect 9700 4365 9715 4385
rect 9735 4365 9750 4385
rect 9700 4350 9750 4365
rect 9850 4835 9900 4850
rect 9850 4815 9865 4835
rect 9885 4815 9900 4835
rect 9850 4785 9900 4815
rect 9850 4765 9865 4785
rect 9885 4765 9900 4785
rect 9850 4735 9900 4765
rect 9850 4715 9865 4735
rect 9885 4715 9900 4735
rect 9850 4685 9900 4715
rect 9850 4665 9865 4685
rect 9885 4665 9900 4685
rect 9850 4635 9900 4665
rect 9850 4615 9865 4635
rect 9885 4615 9900 4635
rect 9850 4585 9900 4615
rect 9850 4565 9865 4585
rect 9885 4565 9900 4585
rect 9850 4535 9900 4565
rect 9850 4515 9865 4535
rect 9885 4515 9900 4535
rect 9850 4485 9900 4515
rect 9850 4465 9865 4485
rect 9885 4465 9900 4485
rect 9850 4435 9900 4465
rect 9850 4415 9865 4435
rect 9885 4415 9900 4435
rect 9850 4385 9900 4415
rect 9850 4365 9865 4385
rect 9885 4365 9900 4385
rect 9850 4350 9900 4365
rect 10000 4835 10050 4850
rect 10000 4815 10015 4835
rect 10035 4815 10050 4835
rect 10000 4785 10050 4815
rect 10000 4765 10015 4785
rect 10035 4765 10050 4785
rect 10000 4735 10050 4765
rect 10000 4715 10015 4735
rect 10035 4715 10050 4735
rect 10000 4685 10050 4715
rect 10000 4665 10015 4685
rect 10035 4665 10050 4685
rect 10000 4635 10050 4665
rect 10000 4615 10015 4635
rect 10035 4615 10050 4635
rect 10000 4585 10050 4615
rect 10000 4565 10015 4585
rect 10035 4565 10050 4585
rect 10000 4535 10050 4565
rect 10000 4515 10015 4535
rect 10035 4515 10050 4535
rect 10000 4485 10050 4515
rect 10000 4465 10015 4485
rect 10035 4465 10050 4485
rect 10000 4435 10050 4465
rect 10000 4415 10015 4435
rect 10035 4415 10050 4435
rect 10000 4385 10050 4415
rect 10000 4365 10015 4385
rect 10035 4365 10050 4385
rect 10000 4350 10050 4365
rect 10150 4835 10200 4850
rect 10150 4815 10165 4835
rect 10185 4815 10200 4835
rect 10150 4785 10200 4815
rect 10150 4765 10165 4785
rect 10185 4765 10200 4785
rect 10150 4735 10200 4765
rect 10150 4715 10165 4735
rect 10185 4715 10200 4735
rect 10150 4685 10200 4715
rect 10150 4665 10165 4685
rect 10185 4665 10200 4685
rect 10150 4635 10200 4665
rect 10150 4615 10165 4635
rect 10185 4615 10200 4635
rect 10150 4585 10200 4615
rect 10150 4565 10165 4585
rect 10185 4565 10200 4585
rect 10150 4535 10200 4565
rect 10150 4515 10165 4535
rect 10185 4515 10200 4535
rect 10150 4485 10200 4515
rect 10150 4465 10165 4485
rect 10185 4465 10200 4485
rect 10150 4435 10200 4465
rect 10150 4415 10165 4435
rect 10185 4415 10200 4435
rect 10150 4385 10200 4415
rect 10150 4365 10165 4385
rect 10185 4365 10200 4385
rect 10150 4350 10200 4365
rect 10300 4835 10350 4850
rect 10300 4815 10315 4835
rect 10335 4815 10350 4835
rect 10300 4785 10350 4815
rect 10300 4765 10315 4785
rect 10335 4765 10350 4785
rect 10300 4735 10350 4765
rect 10300 4715 10315 4735
rect 10335 4715 10350 4735
rect 10300 4685 10350 4715
rect 10300 4665 10315 4685
rect 10335 4665 10350 4685
rect 10300 4635 10350 4665
rect 10300 4615 10315 4635
rect 10335 4615 10350 4635
rect 10300 4585 10350 4615
rect 10300 4565 10315 4585
rect 10335 4565 10350 4585
rect 10300 4535 10350 4565
rect 10300 4515 10315 4535
rect 10335 4515 10350 4535
rect 10300 4485 10350 4515
rect 10300 4465 10315 4485
rect 10335 4465 10350 4485
rect 10300 4435 10350 4465
rect 10300 4415 10315 4435
rect 10335 4415 10350 4435
rect 10300 4385 10350 4415
rect 10300 4365 10315 4385
rect 10335 4365 10350 4385
rect 10300 4350 10350 4365
rect 10450 4835 10500 4850
rect 10450 4815 10465 4835
rect 10485 4815 10500 4835
rect 10450 4785 10500 4815
rect 10450 4765 10465 4785
rect 10485 4765 10500 4785
rect 10450 4735 10500 4765
rect 10450 4715 10465 4735
rect 10485 4715 10500 4735
rect 10450 4685 10500 4715
rect 10450 4665 10465 4685
rect 10485 4665 10500 4685
rect 10450 4635 10500 4665
rect 10450 4615 10465 4635
rect 10485 4615 10500 4635
rect 10450 4585 10500 4615
rect 10450 4565 10465 4585
rect 10485 4565 10500 4585
rect 10450 4535 10500 4565
rect 10450 4515 10465 4535
rect 10485 4515 10500 4535
rect 10450 4485 10500 4515
rect 10450 4465 10465 4485
rect 10485 4465 10500 4485
rect 10450 4435 10500 4465
rect 10450 4415 10465 4435
rect 10485 4415 10500 4435
rect 10450 4385 10500 4415
rect 10450 4365 10465 4385
rect 10485 4365 10500 4385
rect 10450 4350 10500 4365
rect 10600 4835 10650 4850
rect 10600 4815 10615 4835
rect 10635 4815 10650 4835
rect 10600 4785 10650 4815
rect 10600 4765 10615 4785
rect 10635 4765 10650 4785
rect 10600 4735 10650 4765
rect 10600 4715 10615 4735
rect 10635 4715 10650 4735
rect 10600 4685 10650 4715
rect 10600 4665 10615 4685
rect 10635 4665 10650 4685
rect 10600 4635 10650 4665
rect 10600 4615 10615 4635
rect 10635 4615 10650 4635
rect 10600 4585 10650 4615
rect 10600 4565 10615 4585
rect 10635 4565 10650 4585
rect 10600 4535 10650 4565
rect 10600 4515 10615 4535
rect 10635 4515 10650 4535
rect 10600 4485 10650 4515
rect 10600 4465 10615 4485
rect 10635 4465 10650 4485
rect 10600 4435 10650 4465
rect 10600 4415 10615 4435
rect 10635 4415 10650 4435
rect 10600 4385 10650 4415
rect 10600 4365 10615 4385
rect 10635 4365 10650 4385
rect 10600 4350 10650 4365
rect 10750 4835 10800 4850
rect 10750 4815 10765 4835
rect 10785 4815 10800 4835
rect 10750 4785 10800 4815
rect 10750 4765 10765 4785
rect 10785 4765 10800 4785
rect 10750 4735 10800 4765
rect 10750 4715 10765 4735
rect 10785 4715 10800 4735
rect 10750 4685 10800 4715
rect 10750 4665 10765 4685
rect 10785 4665 10800 4685
rect 10750 4635 10800 4665
rect 10750 4615 10765 4635
rect 10785 4615 10800 4635
rect 10750 4585 10800 4615
rect 10750 4565 10765 4585
rect 10785 4565 10800 4585
rect 10750 4535 10800 4565
rect 10750 4515 10765 4535
rect 10785 4515 10800 4535
rect 10750 4485 10800 4515
rect 10750 4465 10765 4485
rect 10785 4465 10800 4485
rect 10750 4435 10800 4465
rect 10750 4415 10765 4435
rect 10785 4415 10800 4435
rect 10750 4385 10800 4415
rect 10750 4365 10765 4385
rect 10785 4365 10800 4385
rect 10750 4350 10800 4365
rect 10900 4350 10950 4850
rect 11050 4350 11100 4850
rect 11200 4350 11250 4850
rect 11350 4835 11400 4850
rect 11350 4815 11365 4835
rect 11385 4815 11400 4835
rect 11350 4785 11400 4815
rect 11350 4765 11365 4785
rect 11385 4765 11400 4785
rect 11350 4735 11400 4765
rect 11350 4715 11365 4735
rect 11385 4715 11400 4735
rect 11350 4685 11400 4715
rect 11350 4665 11365 4685
rect 11385 4665 11400 4685
rect 11350 4635 11400 4665
rect 11350 4615 11365 4635
rect 11385 4615 11400 4635
rect 11350 4585 11400 4615
rect 11350 4565 11365 4585
rect 11385 4565 11400 4585
rect 11350 4535 11400 4565
rect 11350 4515 11365 4535
rect 11385 4515 11400 4535
rect 11350 4485 11400 4515
rect 11350 4465 11365 4485
rect 11385 4465 11400 4485
rect 11350 4435 11400 4465
rect 11350 4415 11365 4435
rect 11385 4415 11400 4435
rect 11350 4385 11400 4415
rect 11350 4365 11365 4385
rect 11385 4365 11400 4385
rect 11350 4350 11400 4365
rect 11500 4350 11550 4850
rect 11650 4350 11700 4850
rect 11800 4350 11850 4850
rect 11950 4835 12000 4850
rect 11950 4815 11965 4835
rect 11985 4815 12000 4835
rect 11950 4785 12000 4815
rect 11950 4765 11965 4785
rect 11985 4765 12000 4785
rect 11950 4735 12000 4765
rect 11950 4715 11965 4735
rect 11985 4715 12000 4735
rect 11950 4685 12000 4715
rect 11950 4665 11965 4685
rect 11985 4665 12000 4685
rect 11950 4635 12000 4665
rect 11950 4615 11965 4635
rect 11985 4615 12000 4635
rect 11950 4585 12000 4615
rect 11950 4565 11965 4585
rect 11985 4565 12000 4585
rect 11950 4535 12000 4565
rect 11950 4515 11965 4535
rect 11985 4515 12000 4535
rect 11950 4485 12000 4515
rect 11950 4465 11965 4485
rect 11985 4465 12000 4485
rect 11950 4435 12000 4465
rect 11950 4415 11965 4435
rect 11985 4415 12000 4435
rect 11950 4385 12000 4415
rect 11950 4365 11965 4385
rect 11985 4365 12000 4385
rect 11950 4350 12000 4365
rect 12100 4350 12150 4850
rect 12250 4350 12300 4850
rect 12400 4350 12450 4850
rect 12550 4835 12600 4850
rect 12550 4815 12565 4835
rect 12585 4815 12600 4835
rect 12550 4785 12600 4815
rect 12550 4765 12565 4785
rect 12585 4765 12600 4785
rect 12550 4735 12600 4765
rect 12550 4715 12565 4735
rect 12585 4715 12600 4735
rect 12550 4685 12600 4715
rect 12550 4665 12565 4685
rect 12585 4665 12600 4685
rect 12550 4635 12600 4665
rect 12550 4615 12565 4635
rect 12585 4615 12600 4635
rect 12550 4585 12600 4615
rect 12550 4565 12565 4585
rect 12585 4565 12600 4585
rect 12550 4535 12600 4565
rect 12550 4515 12565 4535
rect 12585 4515 12600 4535
rect 12550 4485 12600 4515
rect 12550 4465 12565 4485
rect 12585 4465 12600 4485
rect 12550 4435 12600 4465
rect 12550 4415 12565 4435
rect 12585 4415 12600 4435
rect 12550 4385 12600 4415
rect 12550 4365 12565 4385
rect 12585 4365 12600 4385
rect 12550 4350 12600 4365
rect 12700 4350 12750 4850
rect 12850 4350 12900 4850
rect 13000 4350 13050 4850
rect 13150 4835 13200 4850
rect 13150 4815 13165 4835
rect 13185 4815 13200 4835
rect 13150 4785 13200 4815
rect 13150 4765 13165 4785
rect 13185 4765 13200 4785
rect 13150 4735 13200 4765
rect 13150 4715 13165 4735
rect 13185 4715 13200 4735
rect 13150 4685 13200 4715
rect 13150 4665 13165 4685
rect 13185 4665 13200 4685
rect 13150 4635 13200 4665
rect 13150 4615 13165 4635
rect 13185 4615 13200 4635
rect 13150 4585 13200 4615
rect 13150 4565 13165 4585
rect 13185 4565 13200 4585
rect 13150 4535 13200 4565
rect 13150 4515 13165 4535
rect 13185 4515 13200 4535
rect 13150 4485 13200 4515
rect 13150 4465 13165 4485
rect 13185 4465 13200 4485
rect 13150 4435 13200 4465
rect 13150 4415 13165 4435
rect 13185 4415 13200 4435
rect 13150 4385 13200 4415
rect 13150 4365 13165 4385
rect 13185 4365 13200 4385
rect 13150 4350 13200 4365
rect 13300 4350 13350 4850
rect 13450 4350 13500 4850
rect 13600 4350 13650 4850
rect 13750 4835 13800 4850
rect 13750 4815 13765 4835
rect 13785 4815 13800 4835
rect 13750 4785 13800 4815
rect 13750 4765 13765 4785
rect 13785 4765 13800 4785
rect 13750 4735 13800 4765
rect 13750 4715 13765 4735
rect 13785 4715 13800 4735
rect 13750 4685 13800 4715
rect 13750 4665 13765 4685
rect 13785 4665 13800 4685
rect 13750 4635 13800 4665
rect 13750 4615 13765 4635
rect 13785 4615 13800 4635
rect 13750 4585 13800 4615
rect 13750 4565 13765 4585
rect 13785 4565 13800 4585
rect 13750 4535 13800 4565
rect 13750 4515 13765 4535
rect 13785 4515 13800 4535
rect 13750 4485 13800 4515
rect 13750 4465 13765 4485
rect 13785 4465 13800 4485
rect 13750 4435 13800 4465
rect 13750 4415 13765 4435
rect 13785 4415 13800 4435
rect 13750 4385 13800 4415
rect 13750 4365 13765 4385
rect 13785 4365 13800 4385
rect 13750 4350 13800 4365
rect 13900 4350 13950 4850
rect 14050 4350 14100 4850
rect 14200 4350 14250 4850
rect 14350 4835 14400 4850
rect 14350 4815 14365 4835
rect 14385 4815 14400 4835
rect 14350 4785 14400 4815
rect 14350 4765 14365 4785
rect 14385 4765 14400 4785
rect 14350 4735 14400 4765
rect 14350 4715 14365 4735
rect 14385 4715 14400 4735
rect 14350 4685 14400 4715
rect 14350 4665 14365 4685
rect 14385 4665 14400 4685
rect 14350 4635 14400 4665
rect 14350 4615 14365 4635
rect 14385 4615 14400 4635
rect 14350 4585 14400 4615
rect 14350 4565 14365 4585
rect 14385 4565 14400 4585
rect 14350 4535 14400 4565
rect 14350 4515 14365 4535
rect 14385 4515 14400 4535
rect 14350 4485 14400 4515
rect 14350 4465 14365 4485
rect 14385 4465 14400 4485
rect 14350 4435 14400 4465
rect 14350 4415 14365 4435
rect 14385 4415 14400 4435
rect 14350 4385 14400 4415
rect 14350 4365 14365 4385
rect 14385 4365 14400 4385
rect 14350 4350 14400 4365
rect 14500 4350 14550 4850
rect 14650 4350 14700 4850
rect 14800 4350 14850 4850
rect 14950 4835 15000 4850
rect 14950 4815 14965 4835
rect 14985 4815 15000 4835
rect 14950 4785 15000 4815
rect 14950 4765 14965 4785
rect 14985 4765 15000 4785
rect 14950 4735 15000 4765
rect 14950 4715 14965 4735
rect 14985 4715 15000 4735
rect 14950 4685 15000 4715
rect 14950 4665 14965 4685
rect 14985 4665 15000 4685
rect 14950 4635 15000 4665
rect 14950 4615 14965 4635
rect 14985 4615 15000 4635
rect 14950 4585 15000 4615
rect 14950 4565 14965 4585
rect 14985 4565 15000 4585
rect 14950 4535 15000 4565
rect 14950 4515 14965 4535
rect 14985 4515 15000 4535
rect 14950 4485 15000 4515
rect 14950 4465 14965 4485
rect 14985 4465 15000 4485
rect 14950 4435 15000 4465
rect 14950 4415 14965 4435
rect 14985 4415 15000 4435
rect 14950 4385 15000 4415
rect 14950 4365 14965 4385
rect 14985 4365 15000 4385
rect 14950 4350 15000 4365
rect 15100 4350 15150 4850
rect 15250 4350 15300 4850
rect 15400 4350 15450 4850
rect 15550 4835 15600 4850
rect 15550 4815 15565 4835
rect 15585 4815 15600 4835
rect 15550 4785 15600 4815
rect 15550 4765 15565 4785
rect 15585 4765 15600 4785
rect 15550 4735 15600 4765
rect 15550 4715 15565 4735
rect 15585 4715 15600 4735
rect 15550 4685 15600 4715
rect 15550 4665 15565 4685
rect 15585 4665 15600 4685
rect 15550 4635 15600 4665
rect 15550 4615 15565 4635
rect 15585 4615 15600 4635
rect 15550 4585 15600 4615
rect 15550 4565 15565 4585
rect 15585 4565 15600 4585
rect 15550 4535 15600 4565
rect 15550 4515 15565 4535
rect 15585 4515 15600 4535
rect 15550 4485 15600 4515
rect 15550 4465 15565 4485
rect 15585 4465 15600 4485
rect 15550 4435 15600 4465
rect 15550 4415 15565 4435
rect 15585 4415 15600 4435
rect 15550 4385 15600 4415
rect 15550 4365 15565 4385
rect 15585 4365 15600 4385
rect 15550 4350 15600 4365
rect 15700 4350 15750 4850
rect 15850 4350 15900 4850
rect 16000 4350 16050 4850
rect 16150 4835 16200 4850
rect 16150 4815 16165 4835
rect 16185 4815 16200 4835
rect 16150 4785 16200 4815
rect 16150 4765 16165 4785
rect 16185 4765 16200 4785
rect 16150 4735 16200 4765
rect 16150 4715 16165 4735
rect 16185 4715 16200 4735
rect 16150 4685 16200 4715
rect 16150 4665 16165 4685
rect 16185 4665 16200 4685
rect 16150 4635 16200 4665
rect 16150 4615 16165 4635
rect 16185 4615 16200 4635
rect 16150 4585 16200 4615
rect 16150 4565 16165 4585
rect 16185 4565 16200 4585
rect 16150 4535 16200 4565
rect 16150 4515 16165 4535
rect 16185 4515 16200 4535
rect 16150 4485 16200 4515
rect 16150 4465 16165 4485
rect 16185 4465 16200 4485
rect 16150 4435 16200 4465
rect 16150 4415 16165 4435
rect 16185 4415 16200 4435
rect 16150 4385 16200 4415
rect 16150 4365 16165 4385
rect 16185 4365 16200 4385
rect 16150 4350 16200 4365
rect 16300 4835 16350 4850
rect 16300 4815 16315 4835
rect 16335 4815 16350 4835
rect 16300 4785 16350 4815
rect 16300 4765 16315 4785
rect 16335 4765 16350 4785
rect 16300 4735 16350 4765
rect 16300 4715 16315 4735
rect 16335 4715 16350 4735
rect 16300 4685 16350 4715
rect 16300 4665 16315 4685
rect 16335 4665 16350 4685
rect 16300 4635 16350 4665
rect 16300 4615 16315 4635
rect 16335 4615 16350 4635
rect 16300 4585 16350 4615
rect 16300 4565 16315 4585
rect 16335 4565 16350 4585
rect 16300 4535 16350 4565
rect 16300 4515 16315 4535
rect 16335 4515 16350 4535
rect 16300 4485 16350 4515
rect 16300 4465 16315 4485
rect 16335 4465 16350 4485
rect 16300 4435 16350 4465
rect 16300 4415 16315 4435
rect 16335 4415 16350 4435
rect 16300 4385 16350 4415
rect 16300 4365 16315 4385
rect 16335 4365 16350 4385
rect 16300 4350 16350 4365
rect 16450 4835 16500 4850
rect 16450 4815 16465 4835
rect 16485 4815 16500 4835
rect 16450 4785 16500 4815
rect 16450 4765 16465 4785
rect 16485 4765 16500 4785
rect 16450 4735 16500 4765
rect 16450 4715 16465 4735
rect 16485 4715 16500 4735
rect 16450 4685 16500 4715
rect 16450 4665 16465 4685
rect 16485 4665 16500 4685
rect 16450 4635 16500 4665
rect 16450 4615 16465 4635
rect 16485 4615 16500 4635
rect 16450 4585 16500 4615
rect 16450 4565 16465 4585
rect 16485 4565 16500 4585
rect 16450 4535 16500 4565
rect 16450 4515 16465 4535
rect 16485 4515 16500 4535
rect 16450 4485 16500 4515
rect 16450 4465 16465 4485
rect 16485 4465 16500 4485
rect 16450 4435 16500 4465
rect 16450 4415 16465 4435
rect 16485 4415 16500 4435
rect 16450 4385 16500 4415
rect 16450 4365 16465 4385
rect 16485 4365 16500 4385
rect 16450 4350 16500 4365
rect 16600 4835 16650 4850
rect 16600 4815 16615 4835
rect 16635 4815 16650 4835
rect 16600 4785 16650 4815
rect 16600 4765 16615 4785
rect 16635 4765 16650 4785
rect 16600 4735 16650 4765
rect 16600 4715 16615 4735
rect 16635 4715 16650 4735
rect 16600 4685 16650 4715
rect 16600 4665 16615 4685
rect 16635 4665 16650 4685
rect 16600 4635 16650 4665
rect 16600 4615 16615 4635
rect 16635 4615 16650 4635
rect 16600 4585 16650 4615
rect 16600 4565 16615 4585
rect 16635 4565 16650 4585
rect 16600 4535 16650 4565
rect 16600 4515 16615 4535
rect 16635 4515 16650 4535
rect 16600 4485 16650 4515
rect 16600 4465 16615 4485
rect 16635 4465 16650 4485
rect 16600 4435 16650 4465
rect 16600 4415 16615 4435
rect 16635 4415 16650 4435
rect 16600 4385 16650 4415
rect 16600 4365 16615 4385
rect 16635 4365 16650 4385
rect 16600 4350 16650 4365
rect 16750 4835 16800 4850
rect 16750 4815 16765 4835
rect 16785 4815 16800 4835
rect 16750 4785 16800 4815
rect 16750 4765 16765 4785
rect 16785 4765 16800 4785
rect 16750 4735 16800 4765
rect 16750 4715 16765 4735
rect 16785 4715 16800 4735
rect 16750 4685 16800 4715
rect 16750 4665 16765 4685
rect 16785 4665 16800 4685
rect 16750 4635 16800 4665
rect 16750 4615 16765 4635
rect 16785 4615 16800 4635
rect 16750 4585 16800 4615
rect 16750 4565 16765 4585
rect 16785 4565 16800 4585
rect 16750 4535 16800 4565
rect 16750 4515 16765 4535
rect 16785 4515 16800 4535
rect 16750 4485 16800 4515
rect 16750 4465 16765 4485
rect 16785 4465 16800 4485
rect 16750 4435 16800 4465
rect 16750 4415 16765 4435
rect 16785 4415 16800 4435
rect 16750 4385 16800 4415
rect 16750 4365 16765 4385
rect 16785 4365 16800 4385
rect 16750 4350 16800 4365
rect 16900 4835 16950 4850
rect 16900 4815 16915 4835
rect 16935 4815 16950 4835
rect 16900 4785 16950 4815
rect 16900 4765 16915 4785
rect 16935 4765 16950 4785
rect 16900 4735 16950 4765
rect 16900 4715 16915 4735
rect 16935 4715 16950 4735
rect 16900 4685 16950 4715
rect 16900 4665 16915 4685
rect 16935 4665 16950 4685
rect 16900 4635 16950 4665
rect 16900 4615 16915 4635
rect 16935 4615 16950 4635
rect 16900 4585 16950 4615
rect 16900 4565 16915 4585
rect 16935 4565 16950 4585
rect 16900 4535 16950 4565
rect 16900 4515 16915 4535
rect 16935 4515 16950 4535
rect 16900 4485 16950 4515
rect 16900 4465 16915 4485
rect 16935 4465 16950 4485
rect 16900 4435 16950 4465
rect 16900 4415 16915 4435
rect 16935 4415 16950 4435
rect 16900 4385 16950 4415
rect 16900 4365 16915 4385
rect 16935 4365 16950 4385
rect 16900 4350 16950 4365
rect 17050 4835 17100 4850
rect 17050 4815 17065 4835
rect 17085 4815 17100 4835
rect 17050 4785 17100 4815
rect 17050 4765 17065 4785
rect 17085 4765 17100 4785
rect 17050 4735 17100 4765
rect 17050 4715 17065 4735
rect 17085 4715 17100 4735
rect 17050 4685 17100 4715
rect 17050 4665 17065 4685
rect 17085 4665 17100 4685
rect 17050 4635 17100 4665
rect 17050 4615 17065 4635
rect 17085 4615 17100 4635
rect 17050 4585 17100 4615
rect 17050 4565 17065 4585
rect 17085 4565 17100 4585
rect 17050 4535 17100 4565
rect 17050 4515 17065 4535
rect 17085 4515 17100 4535
rect 17050 4485 17100 4515
rect 17050 4465 17065 4485
rect 17085 4465 17100 4485
rect 17050 4435 17100 4465
rect 17050 4415 17065 4435
rect 17085 4415 17100 4435
rect 17050 4385 17100 4415
rect 17050 4365 17065 4385
rect 17085 4365 17100 4385
rect 17050 4350 17100 4365
rect 17200 4835 17250 4850
rect 17200 4815 17215 4835
rect 17235 4815 17250 4835
rect 17200 4785 17250 4815
rect 17200 4765 17215 4785
rect 17235 4765 17250 4785
rect 17200 4735 17250 4765
rect 17200 4715 17215 4735
rect 17235 4715 17250 4735
rect 17200 4685 17250 4715
rect 17200 4665 17215 4685
rect 17235 4665 17250 4685
rect 17200 4635 17250 4665
rect 17200 4615 17215 4635
rect 17235 4615 17250 4635
rect 17200 4585 17250 4615
rect 17200 4565 17215 4585
rect 17235 4565 17250 4585
rect 17200 4535 17250 4565
rect 17200 4515 17215 4535
rect 17235 4515 17250 4535
rect 17200 4485 17250 4515
rect 17200 4465 17215 4485
rect 17235 4465 17250 4485
rect 17200 4435 17250 4465
rect 17200 4415 17215 4435
rect 17235 4415 17250 4435
rect 17200 4385 17250 4415
rect 17200 4365 17215 4385
rect 17235 4365 17250 4385
rect 17200 4350 17250 4365
rect 17350 4835 17400 4850
rect 17350 4815 17365 4835
rect 17385 4815 17400 4835
rect 17350 4785 17400 4815
rect 17350 4765 17365 4785
rect 17385 4765 17400 4785
rect 17350 4735 17400 4765
rect 17350 4715 17365 4735
rect 17385 4715 17400 4735
rect 17350 4685 17400 4715
rect 17350 4665 17365 4685
rect 17385 4665 17400 4685
rect 17350 4635 17400 4665
rect 17350 4615 17365 4635
rect 17385 4615 17400 4635
rect 17350 4585 17400 4615
rect 17350 4565 17365 4585
rect 17385 4565 17400 4585
rect 17350 4535 17400 4565
rect 17350 4515 17365 4535
rect 17385 4515 17400 4535
rect 17350 4485 17400 4515
rect 17350 4465 17365 4485
rect 17385 4465 17400 4485
rect 17350 4435 17400 4465
rect 17350 4415 17365 4435
rect 17385 4415 17400 4435
rect 17350 4385 17400 4415
rect 17350 4365 17365 4385
rect 17385 4365 17400 4385
rect 17350 4350 17400 4365
rect 17500 4350 17550 4850
rect 17650 4350 17700 4850
rect 17800 4350 17850 4850
rect 17950 4835 18000 4850
rect 17950 4815 17965 4835
rect 17985 4815 18000 4835
rect 17950 4785 18000 4815
rect 17950 4765 17965 4785
rect 17985 4765 18000 4785
rect 17950 4735 18000 4765
rect 17950 4715 17965 4735
rect 17985 4715 18000 4735
rect 17950 4685 18000 4715
rect 17950 4665 17965 4685
rect 17985 4665 18000 4685
rect 17950 4635 18000 4665
rect 17950 4615 17965 4635
rect 17985 4615 18000 4635
rect 17950 4585 18000 4615
rect 17950 4565 17965 4585
rect 17985 4565 18000 4585
rect 17950 4535 18000 4565
rect 17950 4515 17965 4535
rect 17985 4515 18000 4535
rect 17950 4485 18000 4515
rect 17950 4465 17965 4485
rect 17985 4465 18000 4485
rect 17950 4435 18000 4465
rect 17950 4415 17965 4435
rect 17985 4415 18000 4435
rect 17950 4385 18000 4415
rect 17950 4365 17965 4385
rect 17985 4365 18000 4385
rect 17950 4350 18000 4365
rect 18100 4350 18150 4850
rect 18250 4350 18300 4850
rect 18400 4350 18450 4850
rect 18550 4835 18600 4850
rect 18550 4815 18565 4835
rect 18585 4815 18600 4835
rect 18550 4785 18600 4815
rect 18550 4765 18565 4785
rect 18585 4765 18600 4785
rect 18550 4735 18600 4765
rect 18550 4715 18565 4735
rect 18585 4715 18600 4735
rect 18550 4685 18600 4715
rect 18550 4665 18565 4685
rect 18585 4665 18600 4685
rect 18550 4635 18600 4665
rect 18550 4615 18565 4635
rect 18585 4615 18600 4635
rect 18550 4585 18600 4615
rect 18550 4565 18565 4585
rect 18585 4565 18600 4585
rect 18550 4535 18600 4565
rect 18550 4515 18565 4535
rect 18585 4515 18600 4535
rect 18550 4485 18600 4515
rect 18550 4465 18565 4485
rect 18585 4465 18600 4485
rect 18550 4435 18600 4465
rect 18550 4415 18565 4435
rect 18585 4415 18600 4435
rect 18550 4385 18600 4415
rect 18550 4365 18565 4385
rect 18585 4365 18600 4385
rect 18550 4350 18600 4365
rect 18700 4835 18750 4850
rect 18700 4815 18715 4835
rect 18735 4815 18750 4835
rect 18700 4785 18750 4815
rect 18700 4765 18715 4785
rect 18735 4765 18750 4785
rect 18700 4735 18750 4765
rect 18700 4715 18715 4735
rect 18735 4715 18750 4735
rect 18700 4685 18750 4715
rect 18700 4665 18715 4685
rect 18735 4665 18750 4685
rect 18700 4635 18750 4665
rect 18700 4615 18715 4635
rect 18735 4615 18750 4635
rect 18700 4585 18750 4615
rect 18700 4565 18715 4585
rect 18735 4565 18750 4585
rect 18700 4535 18750 4565
rect 18700 4515 18715 4535
rect 18735 4515 18750 4535
rect 18700 4485 18750 4515
rect 18700 4465 18715 4485
rect 18735 4465 18750 4485
rect 18700 4435 18750 4465
rect 18700 4415 18715 4435
rect 18735 4415 18750 4435
rect 18700 4385 18750 4415
rect 18700 4365 18715 4385
rect 18735 4365 18750 4385
rect 18700 4350 18750 4365
rect 18850 4835 18900 4850
rect 18850 4815 18865 4835
rect 18885 4815 18900 4835
rect 18850 4785 18900 4815
rect 18850 4765 18865 4785
rect 18885 4765 18900 4785
rect 18850 4735 18900 4765
rect 18850 4715 18865 4735
rect 18885 4715 18900 4735
rect 18850 4685 18900 4715
rect 18850 4665 18865 4685
rect 18885 4665 18900 4685
rect 18850 4635 18900 4665
rect 18850 4615 18865 4635
rect 18885 4615 18900 4635
rect 18850 4585 18900 4615
rect 18850 4565 18865 4585
rect 18885 4565 18900 4585
rect 18850 4535 18900 4565
rect 18850 4515 18865 4535
rect 18885 4515 18900 4535
rect 18850 4485 18900 4515
rect 18850 4465 18865 4485
rect 18885 4465 18900 4485
rect 18850 4435 18900 4465
rect 18850 4415 18865 4435
rect 18885 4415 18900 4435
rect 18850 4385 18900 4415
rect 18850 4365 18865 4385
rect 18885 4365 18900 4385
rect 18850 4350 18900 4365
rect 19000 4835 19050 4850
rect 19000 4815 19015 4835
rect 19035 4815 19050 4835
rect 19000 4785 19050 4815
rect 19000 4765 19015 4785
rect 19035 4765 19050 4785
rect 19000 4735 19050 4765
rect 19000 4715 19015 4735
rect 19035 4715 19050 4735
rect 19000 4685 19050 4715
rect 19000 4665 19015 4685
rect 19035 4665 19050 4685
rect 19000 4635 19050 4665
rect 19000 4615 19015 4635
rect 19035 4615 19050 4635
rect 19000 4585 19050 4615
rect 19000 4565 19015 4585
rect 19035 4565 19050 4585
rect 19000 4535 19050 4565
rect 19000 4515 19015 4535
rect 19035 4515 19050 4535
rect 19000 4485 19050 4515
rect 19000 4465 19015 4485
rect 19035 4465 19050 4485
rect 19000 4435 19050 4465
rect 19000 4415 19015 4435
rect 19035 4415 19050 4435
rect 19000 4385 19050 4415
rect 19000 4365 19015 4385
rect 19035 4365 19050 4385
rect 19000 4350 19050 4365
rect 19150 4835 19200 4850
rect 19150 4815 19165 4835
rect 19185 4815 19200 4835
rect 19150 4785 19200 4815
rect 19150 4765 19165 4785
rect 19185 4765 19200 4785
rect 19150 4735 19200 4765
rect 19150 4715 19165 4735
rect 19185 4715 19200 4735
rect 19150 4685 19200 4715
rect 19150 4665 19165 4685
rect 19185 4665 19200 4685
rect 19150 4635 19200 4665
rect 19150 4615 19165 4635
rect 19185 4615 19200 4635
rect 19150 4585 19200 4615
rect 19150 4565 19165 4585
rect 19185 4565 19200 4585
rect 19150 4535 19200 4565
rect 19150 4515 19165 4535
rect 19185 4515 19200 4535
rect 19150 4485 19200 4515
rect 19150 4465 19165 4485
rect 19185 4465 19200 4485
rect 19150 4435 19200 4465
rect 19150 4415 19165 4435
rect 19185 4415 19200 4435
rect 19150 4385 19200 4415
rect 19150 4365 19165 4385
rect 19185 4365 19200 4385
rect 19150 4350 19200 4365
rect 19300 4835 19350 4850
rect 19300 4815 19315 4835
rect 19335 4815 19350 4835
rect 19300 4785 19350 4815
rect 19300 4765 19315 4785
rect 19335 4765 19350 4785
rect 19300 4735 19350 4765
rect 19300 4715 19315 4735
rect 19335 4715 19350 4735
rect 19300 4685 19350 4715
rect 19300 4665 19315 4685
rect 19335 4665 19350 4685
rect 19300 4635 19350 4665
rect 19300 4615 19315 4635
rect 19335 4615 19350 4635
rect 19300 4585 19350 4615
rect 19300 4565 19315 4585
rect 19335 4565 19350 4585
rect 19300 4535 19350 4565
rect 19300 4515 19315 4535
rect 19335 4515 19350 4535
rect 19300 4485 19350 4515
rect 19300 4465 19315 4485
rect 19335 4465 19350 4485
rect 19300 4435 19350 4465
rect 19300 4415 19315 4435
rect 19335 4415 19350 4435
rect 19300 4385 19350 4415
rect 19300 4365 19315 4385
rect 19335 4365 19350 4385
rect 19300 4350 19350 4365
rect 19450 4835 19500 4850
rect 19450 4815 19465 4835
rect 19485 4815 19500 4835
rect 19450 4785 19500 4815
rect 19450 4765 19465 4785
rect 19485 4765 19500 4785
rect 19450 4735 19500 4765
rect 19450 4715 19465 4735
rect 19485 4715 19500 4735
rect 19450 4685 19500 4715
rect 19450 4665 19465 4685
rect 19485 4665 19500 4685
rect 19450 4635 19500 4665
rect 19450 4615 19465 4635
rect 19485 4615 19500 4635
rect 19450 4585 19500 4615
rect 19450 4565 19465 4585
rect 19485 4565 19500 4585
rect 19450 4535 19500 4565
rect 19450 4515 19465 4535
rect 19485 4515 19500 4535
rect 19450 4485 19500 4515
rect 19450 4465 19465 4485
rect 19485 4465 19500 4485
rect 19450 4435 19500 4465
rect 19450 4415 19465 4435
rect 19485 4415 19500 4435
rect 19450 4385 19500 4415
rect 19450 4365 19465 4385
rect 19485 4365 19500 4385
rect 19450 4350 19500 4365
rect 19600 4835 19650 4850
rect 19600 4815 19615 4835
rect 19635 4815 19650 4835
rect 19600 4785 19650 4815
rect 19600 4765 19615 4785
rect 19635 4765 19650 4785
rect 19600 4735 19650 4765
rect 19600 4715 19615 4735
rect 19635 4715 19650 4735
rect 19600 4685 19650 4715
rect 19600 4665 19615 4685
rect 19635 4665 19650 4685
rect 19600 4635 19650 4665
rect 19600 4615 19615 4635
rect 19635 4615 19650 4635
rect 19600 4585 19650 4615
rect 19600 4565 19615 4585
rect 19635 4565 19650 4585
rect 19600 4535 19650 4565
rect 19600 4515 19615 4535
rect 19635 4515 19650 4535
rect 19600 4485 19650 4515
rect 19600 4465 19615 4485
rect 19635 4465 19650 4485
rect 19600 4435 19650 4465
rect 19600 4415 19615 4435
rect 19635 4415 19650 4435
rect 19600 4385 19650 4415
rect 19600 4365 19615 4385
rect 19635 4365 19650 4385
rect 19600 4350 19650 4365
rect 19750 4835 19800 4850
rect 19750 4815 19765 4835
rect 19785 4815 19800 4835
rect 19750 4785 19800 4815
rect 19750 4765 19765 4785
rect 19785 4765 19800 4785
rect 19750 4735 19800 4765
rect 19750 4715 19765 4735
rect 19785 4715 19800 4735
rect 19750 4685 19800 4715
rect 19750 4665 19765 4685
rect 19785 4665 19800 4685
rect 19750 4635 19800 4665
rect 19750 4615 19765 4635
rect 19785 4615 19800 4635
rect 19750 4585 19800 4615
rect 19750 4565 19765 4585
rect 19785 4565 19800 4585
rect 19750 4535 19800 4565
rect 19750 4515 19765 4535
rect 19785 4515 19800 4535
rect 19750 4485 19800 4515
rect 19750 4465 19765 4485
rect 19785 4465 19800 4485
rect 19750 4435 19800 4465
rect 19750 4415 19765 4435
rect 19785 4415 19800 4435
rect 19750 4385 19800 4415
rect 19750 4365 19765 4385
rect 19785 4365 19800 4385
rect 19750 4350 19800 4365
rect 19900 4350 19950 4850
rect 20050 4350 20100 4850
rect 20200 4350 20250 4850
rect 20350 4835 20400 4850
rect 20350 4815 20365 4835
rect 20385 4815 20400 4835
rect 20350 4785 20400 4815
rect 20350 4765 20365 4785
rect 20385 4765 20400 4785
rect 20350 4735 20400 4765
rect 20350 4715 20365 4735
rect 20385 4715 20400 4735
rect 20350 4685 20400 4715
rect 20350 4665 20365 4685
rect 20385 4665 20400 4685
rect 20350 4635 20400 4665
rect 20350 4615 20365 4635
rect 20385 4615 20400 4635
rect 20350 4585 20400 4615
rect 20350 4565 20365 4585
rect 20385 4565 20400 4585
rect 20350 4535 20400 4565
rect 20350 4515 20365 4535
rect 20385 4515 20400 4535
rect 20350 4485 20400 4515
rect 20350 4465 20365 4485
rect 20385 4465 20400 4485
rect 20350 4435 20400 4465
rect 20350 4415 20365 4435
rect 20385 4415 20400 4435
rect 20350 4385 20400 4415
rect 20350 4365 20365 4385
rect 20385 4365 20400 4385
rect 20350 4350 20400 4365
rect 20500 4350 20550 4850
rect 20650 4350 20700 4850
rect 20800 4350 20850 4850
rect 20950 4835 21000 4850
rect 20950 4815 20965 4835
rect 20985 4815 21000 4835
rect 20950 4785 21000 4815
rect 20950 4765 20965 4785
rect 20985 4765 21000 4785
rect 20950 4735 21000 4765
rect 20950 4715 20965 4735
rect 20985 4715 21000 4735
rect 20950 4685 21000 4715
rect 20950 4665 20965 4685
rect 20985 4665 21000 4685
rect 20950 4635 21000 4665
rect 20950 4615 20965 4635
rect 20985 4615 21000 4635
rect 20950 4585 21000 4615
rect 20950 4565 20965 4585
rect 20985 4565 21000 4585
rect 20950 4535 21000 4565
rect 20950 4515 20965 4535
rect 20985 4515 21000 4535
rect 20950 4485 21000 4515
rect 20950 4465 20965 4485
rect 20985 4465 21000 4485
rect 20950 4435 21000 4465
rect 20950 4415 20965 4435
rect 20985 4415 21000 4435
rect 20950 4385 21000 4415
rect 20950 4365 20965 4385
rect 20985 4365 21000 4385
rect 20950 4350 21000 4365
rect 21100 4350 21150 4850
rect 21250 4350 21300 4850
rect 21400 4835 21450 4850
rect 21400 4815 21415 4835
rect 21435 4815 21450 4835
rect 21400 4785 21450 4815
rect 21400 4765 21415 4785
rect 21435 4765 21450 4785
rect 21400 4735 21450 4765
rect 21400 4715 21415 4735
rect 21435 4715 21450 4735
rect 21400 4685 21450 4715
rect 21400 4665 21415 4685
rect 21435 4665 21450 4685
rect 21400 4635 21450 4665
rect 21400 4615 21415 4635
rect 21435 4615 21450 4635
rect 21400 4585 21450 4615
rect 21400 4565 21415 4585
rect 21435 4565 21450 4585
rect 21400 4535 21450 4565
rect 21400 4515 21415 4535
rect 21435 4515 21450 4535
rect 21400 4485 21450 4515
rect 21400 4465 21415 4485
rect 21435 4465 21450 4485
rect 21400 4435 21450 4465
rect 21400 4415 21415 4435
rect 21435 4415 21450 4435
rect 21400 4385 21450 4415
rect 21400 4365 21415 4385
rect 21435 4365 21450 4385
rect 21400 4350 21450 4365
rect 21550 4350 21600 4850
rect 21700 4350 21750 4850
rect 21850 4835 21900 4850
rect 21850 4815 21865 4835
rect 21885 4815 21900 4835
rect 21850 4785 21900 4815
rect 21850 4765 21865 4785
rect 21885 4765 21900 4785
rect 21850 4735 21900 4765
rect 21850 4715 21865 4735
rect 21885 4715 21900 4735
rect 21850 4685 21900 4715
rect 21850 4665 21865 4685
rect 21885 4665 21900 4685
rect 21850 4635 21900 4665
rect 21850 4615 21865 4635
rect 21885 4615 21900 4635
rect 21850 4585 21900 4615
rect 21850 4565 21865 4585
rect 21885 4565 21900 4585
rect 21850 4535 21900 4565
rect 21850 4515 21865 4535
rect 21885 4515 21900 4535
rect 21850 4485 21900 4515
rect 21850 4465 21865 4485
rect 21885 4465 21900 4485
rect 21850 4435 21900 4465
rect 21850 4415 21865 4435
rect 21885 4415 21900 4435
rect 21850 4385 21900 4415
rect 21850 4365 21865 4385
rect 21885 4365 21900 4385
rect 21850 4350 21900 4365
rect 22000 4350 22050 4850
rect 22150 4350 22200 4850
rect 22300 4350 22350 4850
rect 22450 4835 22500 4850
rect 22450 4815 22465 4835
rect 22485 4815 22500 4835
rect 22450 4785 22500 4815
rect 22450 4765 22465 4785
rect 22485 4765 22500 4785
rect 22450 4735 22500 4765
rect 22450 4715 22465 4735
rect 22485 4715 22500 4735
rect 22450 4685 22500 4715
rect 22450 4665 22465 4685
rect 22485 4665 22500 4685
rect 22450 4635 22500 4665
rect 22450 4615 22465 4635
rect 22485 4615 22500 4635
rect 22450 4585 22500 4615
rect 22450 4565 22465 4585
rect 22485 4565 22500 4585
rect 22450 4535 22500 4565
rect 22450 4515 22465 4535
rect 22485 4515 22500 4535
rect 22450 4485 22500 4515
rect 22450 4465 22465 4485
rect 22485 4465 22500 4485
rect 22450 4435 22500 4465
rect 22450 4415 22465 4435
rect 22485 4415 22500 4435
rect 22450 4385 22500 4415
rect 22450 4365 22465 4385
rect 22485 4365 22500 4385
rect 22450 4350 22500 4365
rect 22600 4350 22650 4850
rect 22750 4350 22800 4850
rect 22900 4350 22950 4850
rect 23050 4835 23100 4850
rect 23050 4815 23065 4835
rect 23085 4815 23100 4835
rect 23050 4785 23100 4815
rect 23050 4765 23065 4785
rect 23085 4765 23100 4785
rect 23050 4735 23100 4765
rect 23050 4715 23065 4735
rect 23085 4715 23100 4735
rect 23050 4685 23100 4715
rect 23050 4665 23065 4685
rect 23085 4665 23100 4685
rect 23050 4635 23100 4665
rect 23050 4615 23065 4635
rect 23085 4615 23100 4635
rect 23050 4585 23100 4615
rect 23050 4565 23065 4585
rect 23085 4565 23100 4585
rect 23050 4535 23100 4565
rect 23050 4515 23065 4535
rect 23085 4515 23100 4535
rect 23050 4485 23100 4515
rect 23050 4465 23065 4485
rect 23085 4465 23100 4485
rect 23050 4435 23100 4465
rect 23050 4415 23065 4435
rect 23085 4415 23100 4435
rect 23050 4385 23100 4415
rect 23050 4365 23065 4385
rect 23085 4365 23100 4385
rect 23050 4350 23100 4365
rect 23200 4350 23250 4850
rect 23350 4350 23400 4850
rect 23500 4835 23550 4850
rect 23500 4815 23515 4835
rect 23535 4815 23550 4835
rect 23500 4785 23550 4815
rect 23500 4765 23515 4785
rect 23535 4765 23550 4785
rect 23500 4735 23550 4765
rect 23500 4715 23515 4735
rect 23535 4715 23550 4735
rect 23500 4685 23550 4715
rect 23500 4665 23515 4685
rect 23535 4665 23550 4685
rect 23500 4635 23550 4665
rect 23500 4615 23515 4635
rect 23535 4615 23550 4635
rect 23500 4585 23550 4615
rect 23500 4565 23515 4585
rect 23535 4565 23550 4585
rect 23500 4535 23550 4565
rect 23500 4515 23515 4535
rect 23535 4515 23550 4535
rect 23500 4485 23550 4515
rect 23500 4465 23515 4485
rect 23535 4465 23550 4485
rect 23500 4435 23550 4465
rect 23500 4415 23515 4435
rect 23535 4415 23550 4435
rect 23500 4385 23550 4415
rect 23500 4365 23515 4385
rect 23535 4365 23550 4385
rect 23500 4350 23550 4365
rect 23650 4350 23700 4850
rect 23800 4350 23850 4850
rect 23950 4835 24000 4850
rect 23950 4815 23965 4835
rect 23985 4815 24000 4835
rect 23950 4785 24000 4815
rect 23950 4765 23965 4785
rect 23985 4765 24000 4785
rect 23950 4735 24000 4765
rect 23950 4715 23965 4735
rect 23985 4715 24000 4735
rect 23950 4685 24000 4715
rect 23950 4665 23965 4685
rect 23985 4665 24000 4685
rect 23950 4635 24000 4665
rect 23950 4615 23965 4635
rect 23985 4615 24000 4635
rect 23950 4585 24000 4615
rect 23950 4565 23965 4585
rect 23985 4565 24000 4585
rect 23950 4535 24000 4565
rect 23950 4515 23965 4535
rect 23985 4515 24000 4535
rect 23950 4485 24000 4515
rect 23950 4465 23965 4485
rect 23985 4465 24000 4485
rect 23950 4435 24000 4465
rect 23950 4415 23965 4435
rect 23985 4415 24000 4435
rect 23950 4385 24000 4415
rect 23950 4365 23965 4385
rect 23985 4365 24000 4385
rect 23950 4350 24000 4365
rect 24100 4350 24150 4850
rect 24250 4350 24300 4850
rect 24400 4350 24450 4850
rect 24550 4835 24600 4850
rect 24550 4815 24565 4835
rect 24585 4815 24600 4835
rect 24550 4785 24600 4815
rect 24550 4765 24565 4785
rect 24585 4765 24600 4785
rect 24550 4735 24600 4765
rect 24550 4715 24565 4735
rect 24585 4715 24600 4735
rect 24550 4685 24600 4715
rect 24550 4665 24565 4685
rect 24585 4665 24600 4685
rect 24550 4635 24600 4665
rect 24550 4615 24565 4635
rect 24585 4615 24600 4635
rect 24550 4585 24600 4615
rect 24550 4565 24565 4585
rect 24585 4565 24600 4585
rect 24550 4535 24600 4565
rect 24550 4515 24565 4535
rect 24585 4515 24600 4535
rect 24550 4485 24600 4515
rect 24550 4465 24565 4485
rect 24585 4465 24600 4485
rect 24550 4435 24600 4465
rect 24550 4415 24565 4435
rect 24585 4415 24600 4435
rect 24550 4385 24600 4415
rect 24550 4365 24565 4385
rect 24585 4365 24600 4385
rect 24550 4350 24600 4365
rect 24700 4350 24750 4850
rect 24850 4350 24900 4850
rect 25000 4350 25050 4850
rect 25150 4835 25200 4850
rect 25150 4815 25165 4835
rect 25185 4815 25200 4835
rect 25150 4785 25200 4815
rect 25150 4765 25165 4785
rect 25185 4765 25200 4785
rect 25150 4735 25200 4765
rect 25150 4715 25165 4735
rect 25185 4715 25200 4735
rect 25150 4685 25200 4715
rect 25150 4665 25165 4685
rect 25185 4665 25200 4685
rect 25150 4635 25200 4665
rect 25150 4615 25165 4635
rect 25185 4615 25200 4635
rect 25150 4585 25200 4615
rect 25150 4565 25165 4585
rect 25185 4565 25200 4585
rect 25150 4535 25200 4565
rect 25150 4515 25165 4535
rect 25185 4515 25200 4535
rect 25150 4485 25200 4515
rect 25150 4465 25165 4485
rect 25185 4465 25200 4485
rect 25150 4435 25200 4465
rect 25150 4415 25165 4435
rect 25185 4415 25200 4435
rect 25150 4385 25200 4415
rect 25150 4365 25165 4385
rect 25185 4365 25200 4385
rect 25150 4350 25200 4365
rect 25300 4350 25350 4850
rect 25450 4350 25500 4850
rect 25600 4835 25650 4850
rect 25600 4815 25615 4835
rect 25635 4815 25650 4835
rect 25600 4785 25650 4815
rect 25600 4765 25615 4785
rect 25635 4765 25650 4785
rect 25600 4735 25650 4765
rect 25600 4715 25615 4735
rect 25635 4715 25650 4735
rect 25600 4685 25650 4715
rect 25600 4665 25615 4685
rect 25635 4665 25650 4685
rect 25600 4635 25650 4665
rect 25600 4615 25615 4635
rect 25635 4615 25650 4635
rect 25600 4585 25650 4615
rect 25600 4565 25615 4585
rect 25635 4565 25650 4585
rect 25600 4535 25650 4565
rect 25600 4515 25615 4535
rect 25635 4515 25650 4535
rect 25600 4485 25650 4515
rect 25600 4465 25615 4485
rect 25635 4465 25650 4485
rect 25600 4435 25650 4465
rect 25600 4415 25615 4435
rect 25635 4415 25650 4435
rect 25600 4385 25650 4415
rect 25600 4365 25615 4385
rect 25635 4365 25650 4385
rect 25600 4350 25650 4365
rect 25750 4350 25800 4850
rect 25900 4350 25950 4850
rect 26050 4835 26100 4850
rect 26050 4815 26065 4835
rect 26085 4815 26100 4835
rect 26050 4785 26100 4815
rect 26050 4765 26065 4785
rect 26085 4765 26100 4785
rect 26050 4735 26100 4765
rect 26050 4715 26065 4735
rect 26085 4715 26100 4735
rect 26050 4685 26100 4715
rect 26050 4665 26065 4685
rect 26085 4665 26100 4685
rect 26050 4635 26100 4665
rect 26050 4615 26065 4635
rect 26085 4615 26100 4635
rect 26050 4585 26100 4615
rect 26050 4565 26065 4585
rect 26085 4565 26100 4585
rect 26050 4535 26100 4565
rect 26050 4515 26065 4535
rect 26085 4515 26100 4535
rect 26050 4485 26100 4515
rect 26050 4465 26065 4485
rect 26085 4465 26100 4485
rect 26050 4435 26100 4465
rect 26050 4415 26065 4435
rect 26085 4415 26100 4435
rect 26050 4385 26100 4415
rect 26050 4365 26065 4385
rect 26085 4365 26100 4385
rect 26050 4350 26100 4365
rect 26200 4350 26250 4850
rect 26350 4350 26400 4850
rect 26500 4350 26550 4850
rect 26650 4835 26700 4850
rect 26650 4815 26665 4835
rect 26685 4815 26700 4835
rect 26650 4785 26700 4815
rect 26650 4765 26665 4785
rect 26685 4765 26700 4785
rect 26650 4735 26700 4765
rect 26650 4715 26665 4735
rect 26685 4715 26700 4735
rect 26650 4685 26700 4715
rect 26650 4665 26665 4685
rect 26685 4665 26700 4685
rect 26650 4635 26700 4665
rect 26650 4615 26665 4635
rect 26685 4615 26700 4635
rect 26650 4585 26700 4615
rect 26650 4565 26665 4585
rect 26685 4565 26700 4585
rect 26650 4535 26700 4565
rect 26650 4515 26665 4535
rect 26685 4515 26700 4535
rect 26650 4485 26700 4515
rect 26650 4465 26665 4485
rect 26685 4465 26700 4485
rect 26650 4435 26700 4465
rect 26650 4415 26665 4435
rect 26685 4415 26700 4435
rect 26650 4385 26700 4415
rect 26650 4365 26665 4385
rect 26685 4365 26700 4385
rect 26650 4350 26700 4365
rect 26800 4350 26850 4850
rect 26950 4350 27000 4850
rect 27100 4350 27150 4850
rect 27250 4835 27300 4850
rect 27250 4815 27265 4835
rect 27285 4815 27300 4835
rect 27250 4785 27300 4815
rect 27250 4765 27265 4785
rect 27285 4765 27300 4785
rect 27250 4735 27300 4765
rect 27250 4715 27265 4735
rect 27285 4715 27300 4735
rect 27250 4685 27300 4715
rect 27250 4665 27265 4685
rect 27285 4665 27300 4685
rect 27250 4635 27300 4665
rect 27250 4615 27265 4635
rect 27285 4615 27300 4635
rect 27250 4585 27300 4615
rect 27250 4565 27265 4585
rect 27285 4565 27300 4585
rect 27250 4535 27300 4565
rect 27250 4515 27265 4535
rect 27285 4515 27300 4535
rect 27250 4485 27300 4515
rect 27250 4465 27265 4485
rect 27285 4465 27300 4485
rect 27250 4435 27300 4465
rect 27250 4415 27265 4435
rect 27285 4415 27300 4435
rect 27250 4385 27300 4415
rect 27250 4365 27265 4385
rect 27285 4365 27300 4385
rect 27250 4350 27300 4365
rect 27400 4350 27450 4850
rect 27550 4350 27600 4850
rect 27700 4835 27750 4850
rect 27700 4815 27715 4835
rect 27735 4815 27750 4835
rect 27700 4785 27750 4815
rect 27700 4765 27715 4785
rect 27735 4765 27750 4785
rect 27700 4735 27750 4765
rect 27700 4715 27715 4735
rect 27735 4715 27750 4735
rect 27700 4685 27750 4715
rect 27700 4665 27715 4685
rect 27735 4665 27750 4685
rect 27700 4635 27750 4665
rect 27700 4615 27715 4635
rect 27735 4615 27750 4635
rect 27700 4585 27750 4615
rect 27700 4565 27715 4585
rect 27735 4565 27750 4585
rect 27700 4535 27750 4565
rect 27700 4515 27715 4535
rect 27735 4515 27750 4535
rect 27700 4485 27750 4515
rect 27700 4465 27715 4485
rect 27735 4465 27750 4485
rect 27700 4435 27750 4465
rect 27700 4415 27715 4435
rect 27735 4415 27750 4435
rect 27700 4385 27750 4415
rect 27700 4365 27715 4385
rect 27735 4365 27750 4385
rect 27700 4350 27750 4365
rect 27850 4350 27900 4850
rect 28000 4350 28050 4850
rect 28150 4835 28200 4850
rect 28150 4815 28165 4835
rect 28185 4815 28200 4835
rect 28150 4785 28200 4815
rect 28150 4765 28165 4785
rect 28185 4765 28200 4785
rect 28150 4735 28200 4765
rect 28150 4715 28165 4735
rect 28185 4715 28200 4735
rect 28150 4685 28200 4715
rect 28150 4665 28165 4685
rect 28185 4665 28200 4685
rect 28150 4635 28200 4665
rect 28150 4615 28165 4635
rect 28185 4615 28200 4635
rect 28150 4585 28200 4615
rect 28150 4565 28165 4585
rect 28185 4565 28200 4585
rect 28150 4535 28200 4565
rect 28150 4515 28165 4535
rect 28185 4515 28200 4535
rect 28150 4485 28200 4515
rect 28150 4465 28165 4485
rect 28185 4465 28200 4485
rect 28150 4435 28200 4465
rect 28150 4415 28165 4435
rect 28185 4415 28200 4435
rect 28150 4385 28200 4415
rect 28150 4365 28165 4385
rect 28185 4365 28200 4385
rect 28150 4350 28200 4365
rect 28300 4350 28350 4850
rect 28450 4350 28500 4850
rect 28600 4350 28650 4850
rect 28750 4835 28800 4850
rect 28750 4815 28765 4835
rect 28785 4815 28800 4835
rect 28750 4785 28800 4815
rect 28750 4765 28765 4785
rect 28785 4765 28800 4785
rect 28750 4735 28800 4765
rect 28750 4715 28765 4735
rect 28785 4715 28800 4735
rect 28750 4685 28800 4715
rect 28750 4665 28765 4685
rect 28785 4665 28800 4685
rect 28750 4635 28800 4665
rect 28750 4615 28765 4635
rect 28785 4615 28800 4635
rect 28750 4585 28800 4615
rect 28750 4565 28765 4585
rect 28785 4565 28800 4585
rect 28750 4535 28800 4565
rect 28750 4515 28765 4535
rect 28785 4515 28800 4535
rect 28750 4485 28800 4515
rect 28750 4465 28765 4485
rect 28785 4465 28800 4485
rect 28750 4435 28800 4465
rect 28750 4415 28765 4435
rect 28785 4415 28800 4435
rect 28750 4385 28800 4415
rect 28750 4365 28765 4385
rect 28785 4365 28800 4385
rect 28750 4350 28800 4365
rect 28900 4350 28950 4850
rect 29050 4350 29100 4850
rect 29200 4350 29250 4850
rect 29350 4835 29400 4850
rect 29350 4815 29365 4835
rect 29385 4815 29400 4835
rect 29350 4785 29400 4815
rect 29350 4765 29365 4785
rect 29385 4765 29400 4785
rect 29350 4735 29400 4765
rect 29350 4715 29365 4735
rect 29385 4715 29400 4735
rect 29350 4685 29400 4715
rect 29350 4665 29365 4685
rect 29385 4665 29400 4685
rect 29350 4635 29400 4665
rect 29350 4615 29365 4635
rect 29385 4615 29400 4635
rect 29350 4585 29400 4615
rect 29350 4565 29365 4585
rect 29385 4565 29400 4585
rect 29350 4535 29400 4565
rect 29350 4515 29365 4535
rect 29385 4515 29400 4535
rect 29350 4485 29400 4515
rect 29350 4465 29365 4485
rect 29385 4465 29400 4485
rect 29350 4435 29400 4465
rect 29350 4415 29365 4435
rect 29385 4415 29400 4435
rect 29350 4385 29400 4415
rect 29350 4365 29365 4385
rect 29385 4365 29400 4385
rect 29350 4350 29400 4365
rect 29500 4835 29550 4850
rect 29500 4815 29515 4835
rect 29535 4815 29550 4835
rect 29500 4785 29550 4815
rect 29500 4765 29515 4785
rect 29535 4765 29550 4785
rect 29500 4735 29550 4765
rect 29500 4715 29515 4735
rect 29535 4715 29550 4735
rect 29500 4685 29550 4715
rect 29500 4665 29515 4685
rect 29535 4665 29550 4685
rect 29500 4635 29550 4665
rect 29500 4615 29515 4635
rect 29535 4615 29550 4635
rect 29500 4585 29550 4615
rect 29500 4565 29515 4585
rect 29535 4565 29550 4585
rect 29500 4535 29550 4565
rect 29500 4515 29515 4535
rect 29535 4515 29550 4535
rect 29500 4485 29550 4515
rect 29500 4465 29515 4485
rect 29535 4465 29550 4485
rect 29500 4435 29550 4465
rect 29500 4415 29515 4435
rect 29535 4415 29550 4435
rect 29500 4385 29550 4415
rect 29500 4365 29515 4385
rect 29535 4365 29550 4385
rect 29500 4350 29550 4365
rect 29650 4835 29700 4850
rect 29650 4815 29665 4835
rect 29685 4815 29700 4835
rect 29650 4785 29700 4815
rect 29650 4765 29665 4785
rect 29685 4765 29700 4785
rect 29650 4735 29700 4765
rect 29650 4715 29665 4735
rect 29685 4715 29700 4735
rect 29650 4685 29700 4715
rect 29650 4665 29665 4685
rect 29685 4665 29700 4685
rect 29650 4635 29700 4665
rect 29650 4615 29665 4635
rect 29685 4615 29700 4635
rect 29650 4585 29700 4615
rect 29650 4565 29665 4585
rect 29685 4565 29700 4585
rect 29650 4535 29700 4565
rect 29650 4515 29665 4535
rect 29685 4515 29700 4535
rect 29650 4485 29700 4515
rect 29650 4465 29665 4485
rect 29685 4465 29700 4485
rect 29650 4435 29700 4465
rect 29650 4415 29665 4435
rect 29685 4415 29700 4435
rect 29650 4385 29700 4415
rect 29650 4365 29665 4385
rect 29685 4365 29700 4385
rect 29650 4350 29700 4365
rect 29800 4835 29850 4850
rect 29800 4815 29815 4835
rect 29835 4815 29850 4835
rect 29800 4785 29850 4815
rect 29800 4765 29815 4785
rect 29835 4765 29850 4785
rect 29800 4735 29850 4765
rect 29800 4715 29815 4735
rect 29835 4715 29850 4735
rect 29800 4685 29850 4715
rect 29800 4665 29815 4685
rect 29835 4665 29850 4685
rect 29800 4635 29850 4665
rect 29800 4615 29815 4635
rect 29835 4615 29850 4635
rect 29800 4585 29850 4615
rect 29800 4565 29815 4585
rect 29835 4565 29850 4585
rect 29800 4535 29850 4565
rect 29800 4515 29815 4535
rect 29835 4515 29850 4535
rect 29800 4485 29850 4515
rect 29800 4465 29815 4485
rect 29835 4465 29850 4485
rect 29800 4435 29850 4465
rect 29800 4415 29815 4435
rect 29835 4415 29850 4435
rect 29800 4385 29850 4415
rect 29800 4365 29815 4385
rect 29835 4365 29850 4385
rect 29800 4350 29850 4365
rect 29950 4835 30000 4850
rect 29950 4815 29965 4835
rect 29985 4815 30000 4835
rect 29950 4785 30000 4815
rect 29950 4765 29965 4785
rect 29985 4765 30000 4785
rect 29950 4735 30000 4765
rect 29950 4715 29965 4735
rect 29985 4715 30000 4735
rect 29950 4685 30000 4715
rect 29950 4665 29965 4685
rect 29985 4665 30000 4685
rect 29950 4635 30000 4665
rect 29950 4615 29965 4635
rect 29985 4615 30000 4635
rect 29950 4585 30000 4615
rect 29950 4565 29965 4585
rect 29985 4565 30000 4585
rect 29950 4535 30000 4565
rect 29950 4515 29965 4535
rect 29985 4515 30000 4535
rect 29950 4485 30000 4515
rect 29950 4465 29965 4485
rect 29985 4465 30000 4485
rect 29950 4435 30000 4465
rect 29950 4415 29965 4435
rect 29985 4415 30000 4435
rect 29950 4385 30000 4415
rect 29950 4365 29965 4385
rect 29985 4365 30000 4385
rect 29950 4350 30000 4365
rect 30100 4835 30150 4850
rect 30100 4815 30115 4835
rect 30135 4815 30150 4835
rect 30100 4785 30150 4815
rect 30100 4765 30115 4785
rect 30135 4765 30150 4785
rect 30100 4735 30150 4765
rect 30100 4715 30115 4735
rect 30135 4715 30150 4735
rect 30100 4685 30150 4715
rect 30100 4665 30115 4685
rect 30135 4665 30150 4685
rect 30100 4635 30150 4665
rect 30100 4615 30115 4635
rect 30135 4615 30150 4635
rect 30100 4585 30150 4615
rect 30100 4565 30115 4585
rect 30135 4565 30150 4585
rect 30100 4535 30150 4565
rect 30100 4515 30115 4535
rect 30135 4515 30150 4535
rect 30100 4485 30150 4515
rect 30100 4465 30115 4485
rect 30135 4465 30150 4485
rect 30100 4435 30150 4465
rect 30100 4415 30115 4435
rect 30135 4415 30150 4435
rect 30100 4385 30150 4415
rect 30100 4365 30115 4385
rect 30135 4365 30150 4385
rect 30100 4350 30150 4365
rect 30250 4835 30300 4850
rect 30250 4815 30265 4835
rect 30285 4815 30300 4835
rect 30250 4785 30300 4815
rect 30250 4765 30265 4785
rect 30285 4765 30300 4785
rect 30250 4735 30300 4765
rect 30250 4715 30265 4735
rect 30285 4715 30300 4735
rect 30250 4685 30300 4715
rect 30250 4665 30265 4685
rect 30285 4665 30300 4685
rect 30250 4635 30300 4665
rect 30250 4615 30265 4635
rect 30285 4615 30300 4635
rect 30250 4585 30300 4615
rect 30250 4565 30265 4585
rect 30285 4565 30300 4585
rect 30250 4535 30300 4565
rect 30250 4515 30265 4535
rect 30285 4515 30300 4535
rect 30250 4485 30300 4515
rect 30250 4465 30265 4485
rect 30285 4465 30300 4485
rect 30250 4435 30300 4465
rect 30250 4415 30265 4435
rect 30285 4415 30300 4435
rect 30250 4385 30300 4415
rect 30250 4365 30265 4385
rect 30285 4365 30300 4385
rect 30250 4350 30300 4365
rect 30400 4835 30450 4850
rect 30400 4815 30415 4835
rect 30435 4815 30450 4835
rect 30400 4785 30450 4815
rect 30400 4765 30415 4785
rect 30435 4765 30450 4785
rect 30400 4735 30450 4765
rect 30400 4715 30415 4735
rect 30435 4715 30450 4735
rect 30400 4685 30450 4715
rect 30400 4665 30415 4685
rect 30435 4665 30450 4685
rect 30400 4635 30450 4665
rect 30400 4615 30415 4635
rect 30435 4615 30450 4635
rect 30400 4585 30450 4615
rect 30400 4565 30415 4585
rect 30435 4565 30450 4585
rect 30400 4535 30450 4565
rect 30400 4515 30415 4535
rect 30435 4515 30450 4535
rect 30400 4485 30450 4515
rect 30400 4465 30415 4485
rect 30435 4465 30450 4485
rect 30400 4435 30450 4465
rect 30400 4415 30415 4435
rect 30435 4415 30450 4435
rect 30400 4385 30450 4415
rect 30400 4365 30415 4385
rect 30435 4365 30450 4385
rect 30400 4350 30450 4365
rect 30550 4835 30600 4850
rect 30550 4815 30565 4835
rect 30585 4815 30600 4835
rect 30550 4785 30600 4815
rect 30550 4765 30565 4785
rect 30585 4765 30600 4785
rect 30550 4735 30600 4765
rect 30550 4715 30565 4735
rect 30585 4715 30600 4735
rect 30550 4685 30600 4715
rect 30550 4665 30565 4685
rect 30585 4665 30600 4685
rect 30550 4635 30600 4665
rect 30550 4615 30565 4635
rect 30585 4615 30600 4635
rect 30550 4585 30600 4615
rect 30550 4565 30565 4585
rect 30585 4565 30600 4585
rect 30550 4535 30600 4565
rect 30550 4515 30565 4535
rect 30585 4515 30600 4535
rect 30550 4485 30600 4515
rect 30550 4465 30565 4485
rect 30585 4465 30600 4485
rect 30550 4435 30600 4465
rect 30550 4415 30565 4435
rect 30585 4415 30600 4435
rect 30550 4385 30600 4415
rect 30550 4365 30565 4385
rect 30585 4365 30600 4385
rect 30550 4350 30600 4365
rect 30700 4835 30750 4850
rect 30700 4815 30715 4835
rect 30735 4815 30750 4835
rect 30700 4785 30750 4815
rect 30700 4765 30715 4785
rect 30735 4765 30750 4785
rect 30700 4735 30750 4765
rect 30700 4715 30715 4735
rect 30735 4715 30750 4735
rect 30700 4685 30750 4715
rect 30700 4665 30715 4685
rect 30735 4665 30750 4685
rect 30700 4635 30750 4665
rect 30700 4615 30715 4635
rect 30735 4615 30750 4635
rect 30700 4585 30750 4615
rect 30700 4565 30715 4585
rect 30735 4565 30750 4585
rect 30700 4535 30750 4565
rect 30700 4515 30715 4535
rect 30735 4515 30750 4535
rect 30700 4485 30750 4515
rect 30700 4465 30715 4485
rect 30735 4465 30750 4485
rect 30700 4435 30750 4465
rect 30700 4415 30715 4435
rect 30735 4415 30750 4435
rect 30700 4385 30750 4415
rect 30700 4365 30715 4385
rect 30735 4365 30750 4385
rect 30700 4350 30750 4365
rect 30850 4835 30900 4850
rect 30850 4815 30865 4835
rect 30885 4815 30900 4835
rect 30850 4785 30900 4815
rect 30850 4765 30865 4785
rect 30885 4765 30900 4785
rect 30850 4735 30900 4765
rect 30850 4715 30865 4735
rect 30885 4715 30900 4735
rect 30850 4685 30900 4715
rect 30850 4665 30865 4685
rect 30885 4665 30900 4685
rect 30850 4635 30900 4665
rect 30850 4615 30865 4635
rect 30885 4615 30900 4635
rect 30850 4585 30900 4615
rect 30850 4565 30865 4585
rect 30885 4565 30900 4585
rect 30850 4535 30900 4565
rect 30850 4515 30865 4535
rect 30885 4515 30900 4535
rect 30850 4485 30900 4515
rect 30850 4465 30865 4485
rect 30885 4465 30900 4485
rect 30850 4435 30900 4465
rect 30850 4415 30865 4435
rect 30885 4415 30900 4435
rect 30850 4385 30900 4415
rect 30850 4365 30865 4385
rect 30885 4365 30900 4385
rect 30850 4350 30900 4365
rect 31000 4835 31050 4850
rect 31000 4815 31015 4835
rect 31035 4815 31050 4835
rect 31000 4785 31050 4815
rect 31000 4765 31015 4785
rect 31035 4765 31050 4785
rect 31000 4735 31050 4765
rect 31000 4715 31015 4735
rect 31035 4715 31050 4735
rect 31000 4685 31050 4715
rect 31000 4665 31015 4685
rect 31035 4665 31050 4685
rect 31000 4635 31050 4665
rect 31000 4615 31015 4635
rect 31035 4615 31050 4635
rect 31000 4585 31050 4615
rect 31000 4565 31015 4585
rect 31035 4565 31050 4585
rect 31000 4535 31050 4565
rect 31000 4515 31015 4535
rect 31035 4515 31050 4535
rect 31000 4485 31050 4515
rect 31000 4465 31015 4485
rect 31035 4465 31050 4485
rect 31000 4435 31050 4465
rect 31000 4415 31015 4435
rect 31035 4415 31050 4435
rect 31000 4385 31050 4415
rect 31000 4365 31015 4385
rect 31035 4365 31050 4385
rect 31000 4350 31050 4365
rect 31150 4835 31200 4850
rect 31150 4815 31165 4835
rect 31185 4815 31200 4835
rect 31150 4785 31200 4815
rect 31150 4765 31165 4785
rect 31185 4765 31200 4785
rect 31150 4735 31200 4765
rect 31150 4715 31165 4735
rect 31185 4715 31200 4735
rect 31150 4685 31200 4715
rect 31150 4665 31165 4685
rect 31185 4665 31200 4685
rect 31150 4635 31200 4665
rect 31150 4615 31165 4635
rect 31185 4615 31200 4635
rect 31150 4585 31200 4615
rect 31150 4565 31165 4585
rect 31185 4565 31200 4585
rect 31150 4535 31200 4565
rect 31150 4515 31165 4535
rect 31185 4515 31200 4535
rect 31150 4485 31200 4515
rect 31150 4465 31165 4485
rect 31185 4465 31200 4485
rect 31150 4435 31200 4465
rect 31150 4415 31165 4435
rect 31185 4415 31200 4435
rect 31150 4385 31200 4415
rect 31150 4365 31165 4385
rect 31185 4365 31200 4385
rect 31150 4350 31200 4365
rect 31300 4835 31350 4850
rect 31300 4815 31315 4835
rect 31335 4815 31350 4835
rect 31300 4785 31350 4815
rect 31300 4765 31315 4785
rect 31335 4765 31350 4785
rect 31300 4735 31350 4765
rect 31300 4715 31315 4735
rect 31335 4715 31350 4735
rect 31300 4685 31350 4715
rect 31300 4665 31315 4685
rect 31335 4665 31350 4685
rect 31300 4635 31350 4665
rect 31300 4615 31315 4635
rect 31335 4615 31350 4635
rect 31300 4585 31350 4615
rect 31300 4565 31315 4585
rect 31335 4565 31350 4585
rect 31300 4535 31350 4565
rect 31300 4515 31315 4535
rect 31335 4515 31350 4535
rect 31300 4485 31350 4515
rect 31300 4465 31315 4485
rect 31335 4465 31350 4485
rect 31300 4435 31350 4465
rect 31300 4415 31315 4435
rect 31335 4415 31350 4435
rect 31300 4385 31350 4415
rect 31300 4365 31315 4385
rect 31335 4365 31350 4385
rect 31300 4350 31350 4365
rect 31450 4835 31500 4850
rect 31450 4815 31465 4835
rect 31485 4815 31500 4835
rect 31450 4785 31500 4815
rect 31450 4765 31465 4785
rect 31485 4765 31500 4785
rect 31450 4735 31500 4765
rect 31450 4715 31465 4735
rect 31485 4715 31500 4735
rect 31450 4685 31500 4715
rect 31450 4665 31465 4685
rect 31485 4665 31500 4685
rect 31450 4635 31500 4665
rect 31450 4615 31465 4635
rect 31485 4615 31500 4635
rect 31450 4585 31500 4615
rect 31450 4565 31465 4585
rect 31485 4565 31500 4585
rect 31450 4535 31500 4565
rect 31450 4515 31465 4535
rect 31485 4515 31500 4535
rect 31450 4485 31500 4515
rect 31450 4465 31465 4485
rect 31485 4465 31500 4485
rect 31450 4435 31500 4465
rect 31450 4415 31465 4435
rect 31485 4415 31500 4435
rect 31450 4385 31500 4415
rect 31450 4365 31465 4385
rect 31485 4365 31500 4385
rect 31450 4350 31500 4365
rect 31600 4350 31650 4850
rect 31750 4350 31800 4850
rect 31900 4350 31950 4850
rect 32050 4835 32100 4850
rect 32050 4815 32065 4835
rect 32085 4815 32100 4835
rect 32050 4785 32100 4815
rect 32050 4765 32065 4785
rect 32085 4765 32100 4785
rect 32050 4735 32100 4765
rect 32050 4715 32065 4735
rect 32085 4715 32100 4735
rect 32050 4685 32100 4715
rect 32050 4665 32065 4685
rect 32085 4665 32100 4685
rect 32050 4635 32100 4665
rect 32050 4615 32065 4635
rect 32085 4615 32100 4635
rect 32050 4585 32100 4615
rect 32050 4565 32065 4585
rect 32085 4565 32100 4585
rect 32050 4535 32100 4565
rect 32050 4515 32065 4535
rect 32085 4515 32100 4535
rect 32050 4485 32100 4515
rect 32050 4465 32065 4485
rect 32085 4465 32100 4485
rect 32050 4435 32100 4465
rect 32050 4415 32065 4435
rect 32085 4415 32100 4435
rect 32050 4385 32100 4415
rect 32050 4365 32065 4385
rect 32085 4365 32100 4385
rect 32050 4350 32100 4365
rect -650 4185 -600 4200
rect -650 4165 -635 4185
rect -615 4165 -600 4185
rect -650 4135 -600 4165
rect -650 4115 -635 4135
rect -615 4115 -600 4135
rect -650 4085 -600 4115
rect -650 4065 -635 4085
rect -615 4065 -600 4085
rect -650 4035 -600 4065
rect -650 4015 -635 4035
rect -615 4015 -600 4035
rect -650 3985 -600 4015
rect -650 3965 -635 3985
rect -615 3965 -600 3985
rect -650 3935 -600 3965
rect -650 3915 -635 3935
rect -615 3915 -600 3935
rect -650 3885 -600 3915
rect -650 3865 -635 3885
rect -615 3865 -600 3885
rect -650 3835 -600 3865
rect -650 3815 -635 3835
rect -615 3815 -600 3835
rect -650 3785 -600 3815
rect -650 3765 -635 3785
rect -615 3765 -600 3785
rect -650 3735 -600 3765
rect -650 3715 -635 3735
rect -615 3715 -600 3735
rect -650 3700 -600 3715
rect -500 4185 -450 4200
rect -500 4165 -485 4185
rect -465 4165 -450 4185
rect -500 4135 -450 4165
rect -500 4115 -485 4135
rect -465 4115 -450 4135
rect -500 4085 -450 4115
rect -500 4065 -485 4085
rect -465 4065 -450 4085
rect -500 4035 -450 4065
rect -500 4015 -485 4035
rect -465 4015 -450 4035
rect -500 3985 -450 4015
rect -500 3965 -485 3985
rect -465 3965 -450 3985
rect -500 3935 -450 3965
rect -500 3915 -485 3935
rect -465 3915 -450 3935
rect -500 3885 -450 3915
rect -500 3865 -485 3885
rect -465 3865 -450 3885
rect -500 3835 -450 3865
rect -500 3815 -485 3835
rect -465 3815 -450 3835
rect -500 3785 -450 3815
rect -500 3765 -485 3785
rect -465 3765 -450 3785
rect -500 3735 -450 3765
rect -500 3715 -485 3735
rect -465 3715 -450 3735
rect -500 3700 -450 3715
rect -350 4185 -300 4200
rect -350 4165 -335 4185
rect -315 4165 -300 4185
rect -350 4135 -300 4165
rect -350 4115 -335 4135
rect -315 4115 -300 4135
rect -350 4085 -300 4115
rect -350 4065 -335 4085
rect -315 4065 -300 4085
rect -350 4035 -300 4065
rect -350 4015 -335 4035
rect -315 4015 -300 4035
rect -350 3985 -300 4015
rect -350 3965 -335 3985
rect -315 3965 -300 3985
rect -350 3935 -300 3965
rect -350 3915 -335 3935
rect -315 3915 -300 3935
rect -350 3885 -300 3915
rect -350 3865 -335 3885
rect -315 3865 -300 3885
rect -350 3835 -300 3865
rect -350 3815 -335 3835
rect -315 3815 -300 3835
rect -350 3785 -300 3815
rect -350 3765 -335 3785
rect -315 3765 -300 3785
rect -350 3735 -300 3765
rect -350 3715 -335 3735
rect -315 3715 -300 3735
rect -350 3700 -300 3715
rect -200 4185 -150 4200
rect -200 4165 -185 4185
rect -165 4165 -150 4185
rect -200 4135 -150 4165
rect -200 4115 -185 4135
rect -165 4115 -150 4135
rect -200 4085 -150 4115
rect -200 4065 -185 4085
rect -165 4065 -150 4085
rect -200 4035 -150 4065
rect -200 4015 -185 4035
rect -165 4015 -150 4035
rect -200 3985 -150 4015
rect -200 3965 -185 3985
rect -165 3965 -150 3985
rect -200 3935 -150 3965
rect -200 3915 -185 3935
rect -165 3915 -150 3935
rect -200 3885 -150 3915
rect -200 3865 -185 3885
rect -165 3865 -150 3885
rect -200 3835 -150 3865
rect -200 3815 -185 3835
rect -165 3815 -150 3835
rect -200 3785 -150 3815
rect -200 3765 -185 3785
rect -165 3765 -150 3785
rect -200 3735 -150 3765
rect -200 3715 -185 3735
rect -165 3715 -150 3735
rect -200 3700 -150 3715
rect -50 4185 0 4200
rect -50 4165 -35 4185
rect -15 4165 0 4185
rect -50 4135 0 4165
rect -50 4115 -35 4135
rect -15 4115 0 4135
rect -50 4085 0 4115
rect -50 4065 -35 4085
rect -15 4065 0 4085
rect -50 4035 0 4065
rect -50 4015 -35 4035
rect -15 4015 0 4035
rect -50 3985 0 4015
rect -50 3965 -35 3985
rect -15 3965 0 3985
rect -50 3935 0 3965
rect -50 3915 -35 3935
rect -15 3915 0 3935
rect -50 3885 0 3915
rect -50 3865 -35 3885
rect -15 3865 0 3885
rect -50 3835 0 3865
rect -50 3815 -35 3835
rect -15 3815 0 3835
rect -50 3785 0 3815
rect -50 3765 -35 3785
rect -15 3765 0 3785
rect -50 3735 0 3765
rect -50 3715 -35 3735
rect -15 3715 0 3735
rect -50 3700 0 3715
rect 100 3700 150 4200
rect 250 3700 300 4200
rect 400 3700 450 4200
rect 550 4185 600 4200
rect 550 4165 565 4185
rect 585 4165 600 4185
rect 550 4135 600 4165
rect 550 4115 565 4135
rect 585 4115 600 4135
rect 550 4085 600 4115
rect 550 4065 565 4085
rect 585 4065 600 4085
rect 550 4035 600 4065
rect 550 4015 565 4035
rect 585 4015 600 4035
rect 550 3985 600 4015
rect 550 3965 565 3985
rect 585 3965 600 3985
rect 550 3935 600 3965
rect 550 3915 565 3935
rect 585 3915 600 3935
rect 550 3885 600 3915
rect 550 3865 565 3885
rect 585 3865 600 3885
rect 550 3835 600 3865
rect 550 3815 565 3835
rect 585 3815 600 3835
rect 550 3785 600 3815
rect 550 3765 565 3785
rect 585 3765 600 3785
rect 550 3735 600 3765
rect 550 3715 565 3735
rect 585 3715 600 3735
rect 550 3700 600 3715
rect 700 4185 750 4200
rect 700 4165 715 4185
rect 735 4165 750 4185
rect 700 4135 750 4165
rect 700 4115 715 4135
rect 735 4115 750 4135
rect 700 4085 750 4115
rect 700 4065 715 4085
rect 735 4065 750 4085
rect 700 4035 750 4065
rect 700 4015 715 4035
rect 735 4015 750 4035
rect 700 3985 750 4015
rect 700 3965 715 3985
rect 735 3965 750 3985
rect 700 3935 750 3965
rect 700 3915 715 3935
rect 735 3915 750 3935
rect 700 3885 750 3915
rect 700 3865 715 3885
rect 735 3865 750 3885
rect 700 3835 750 3865
rect 700 3815 715 3835
rect 735 3815 750 3835
rect 700 3785 750 3815
rect 700 3765 715 3785
rect 735 3765 750 3785
rect 700 3735 750 3765
rect 700 3715 715 3735
rect 735 3715 750 3735
rect 700 3700 750 3715
rect 850 4185 900 4200
rect 850 4165 865 4185
rect 885 4165 900 4185
rect 850 4135 900 4165
rect 850 4115 865 4135
rect 885 4115 900 4135
rect 850 4085 900 4115
rect 850 4065 865 4085
rect 885 4065 900 4085
rect 850 4035 900 4065
rect 850 4015 865 4035
rect 885 4015 900 4035
rect 850 3985 900 4015
rect 850 3965 865 3985
rect 885 3965 900 3985
rect 850 3935 900 3965
rect 850 3915 865 3935
rect 885 3915 900 3935
rect 850 3885 900 3915
rect 850 3865 865 3885
rect 885 3865 900 3885
rect 850 3835 900 3865
rect 850 3815 865 3835
rect 885 3815 900 3835
rect 850 3785 900 3815
rect 850 3765 865 3785
rect 885 3765 900 3785
rect 850 3735 900 3765
rect 850 3715 865 3735
rect 885 3715 900 3735
rect 850 3700 900 3715
rect 1000 4185 1050 4200
rect 1000 4165 1015 4185
rect 1035 4165 1050 4185
rect 1000 4135 1050 4165
rect 1000 4115 1015 4135
rect 1035 4115 1050 4135
rect 1000 4085 1050 4115
rect 1000 4065 1015 4085
rect 1035 4065 1050 4085
rect 1000 4035 1050 4065
rect 1000 4015 1015 4035
rect 1035 4015 1050 4035
rect 1000 3985 1050 4015
rect 1000 3965 1015 3985
rect 1035 3965 1050 3985
rect 1000 3935 1050 3965
rect 1000 3915 1015 3935
rect 1035 3915 1050 3935
rect 1000 3885 1050 3915
rect 1000 3865 1015 3885
rect 1035 3865 1050 3885
rect 1000 3835 1050 3865
rect 1000 3815 1015 3835
rect 1035 3815 1050 3835
rect 1000 3785 1050 3815
rect 1000 3765 1015 3785
rect 1035 3765 1050 3785
rect 1000 3735 1050 3765
rect 1000 3715 1015 3735
rect 1035 3715 1050 3735
rect 1000 3700 1050 3715
rect 1150 4185 1200 4200
rect 1150 4165 1165 4185
rect 1185 4165 1200 4185
rect 1150 4135 1200 4165
rect 1150 4115 1165 4135
rect 1185 4115 1200 4135
rect 1150 4085 1200 4115
rect 1150 4065 1165 4085
rect 1185 4065 1200 4085
rect 1150 4035 1200 4065
rect 1150 4015 1165 4035
rect 1185 4015 1200 4035
rect 1150 3985 1200 4015
rect 1150 3965 1165 3985
rect 1185 3965 1200 3985
rect 1150 3935 1200 3965
rect 1150 3915 1165 3935
rect 1185 3915 1200 3935
rect 1150 3885 1200 3915
rect 1150 3865 1165 3885
rect 1185 3865 1200 3885
rect 1150 3835 1200 3865
rect 1150 3815 1165 3835
rect 1185 3815 1200 3835
rect 1150 3785 1200 3815
rect 1150 3765 1165 3785
rect 1185 3765 1200 3785
rect 1150 3735 1200 3765
rect 1150 3715 1165 3735
rect 1185 3715 1200 3735
rect 1150 3700 1200 3715
rect 1300 4185 1350 4200
rect 1300 4165 1315 4185
rect 1335 4165 1350 4185
rect 1300 4135 1350 4165
rect 1300 4115 1315 4135
rect 1335 4115 1350 4135
rect 1300 4085 1350 4115
rect 1300 4065 1315 4085
rect 1335 4065 1350 4085
rect 1300 4035 1350 4065
rect 1300 4015 1315 4035
rect 1335 4015 1350 4035
rect 1300 3985 1350 4015
rect 1300 3965 1315 3985
rect 1335 3965 1350 3985
rect 1300 3935 1350 3965
rect 1300 3915 1315 3935
rect 1335 3915 1350 3935
rect 1300 3885 1350 3915
rect 1300 3865 1315 3885
rect 1335 3865 1350 3885
rect 1300 3835 1350 3865
rect 1300 3815 1315 3835
rect 1335 3815 1350 3835
rect 1300 3785 1350 3815
rect 1300 3765 1315 3785
rect 1335 3765 1350 3785
rect 1300 3735 1350 3765
rect 1300 3715 1315 3735
rect 1335 3715 1350 3735
rect 1300 3700 1350 3715
rect 1450 4185 1500 4200
rect 1450 4165 1465 4185
rect 1485 4165 1500 4185
rect 1450 4135 1500 4165
rect 1450 4115 1465 4135
rect 1485 4115 1500 4135
rect 1450 4085 1500 4115
rect 1450 4065 1465 4085
rect 1485 4065 1500 4085
rect 1450 4035 1500 4065
rect 1450 4015 1465 4035
rect 1485 4015 1500 4035
rect 1450 3985 1500 4015
rect 1450 3965 1465 3985
rect 1485 3965 1500 3985
rect 1450 3935 1500 3965
rect 1450 3915 1465 3935
rect 1485 3915 1500 3935
rect 1450 3885 1500 3915
rect 1450 3865 1465 3885
rect 1485 3865 1500 3885
rect 1450 3835 1500 3865
rect 1450 3815 1465 3835
rect 1485 3815 1500 3835
rect 1450 3785 1500 3815
rect 1450 3765 1465 3785
rect 1485 3765 1500 3785
rect 1450 3735 1500 3765
rect 1450 3715 1465 3735
rect 1485 3715 1500 3735
rect 1450 3700 1500 3715
rect 1600 4185 1650 4200
rect 1600 4165 1615 4185
rect 1635 4165 1650 4185
rect 1600 4135 1650 4165
rect 1600 4115 1615 4135
rect 1635 4115 1650 4135
rect 1600 4085 1650 4115
rect 1600 4065 1615 4085
rect 1635 4065 1650 4085
rect 1600 4035 1650 4065
rect 1600 4015 1615 4035
rect 1635 4015 1650 4035
rect 1600 3985 1650 4015
rect 1600 3965 1615 3985
rect 1635 3965 1650 3985
rect 1600 3935 1650 3965
rect 1600 3915 1615 3935
rect 1635 3915 1650 3935
rect 1600 3885 1650 3915
rect 1600 3865 1615 3885
rect 1635 3865 1650 3885
rect 1600 3835 1650 3865
rect 1600 3815 1615 3835
rect 1635 3815 1650 3835
rect 1600 3785 1650 3815
rect 1600 3765 1615 3785
rect 1635 3765 1650 3785
rect 1600 3735 1650 3765
rect 1600 3715 1615 3735
rect 1635 3715 1650 3735
rect 1600 3700 1650 3715
rect 1750 4185 1800 4200
rect 1750 4165 1765 4185
rect 1785 4165 1800 4185
rect 1750 4135 1800 4165
rect 1750 4115 1765 4135
rect 1785 4115 1800 4135
rect 1750 4085 1800 4115
rect 1750 4065 1765 4085
rect 1785 4065 1800 4085
rect 1750 4035 1800 4065
rect 1750 4015 1765 4035
rect 1785 4015 1800 4035
rect 1750 3985 1800 4015
rect 1750 3965 1765 3985
rect 1785 3965 1800 3985
rect 1750 3935 1800 3965
rect 1750 3915 1765 3935
rect 1785 3915 1800 3935
rect 1750 3885 1800 3915
rect 1750 3865 1765 3885
rect 1785 3865 1800 3885
rect 1750 3835 1800 3865
rect 1750 3815 1765 3835
rect 1785 3815 1800 3835
rect 1750 3785 1800 3815
rect 1750 3765 1765 3785
rect 1785 3765 1800 3785
rect 1750 3735 1800 3765
rect 1750 3715 1765 3735
rect 1785 3715 1800 3735
rect 1750 3700 1800 3715
rect 1900 4185 1950 4200
rect 1900 4165 1915 4185
rect 1935 4165 1950 4185
rect 1900 4135 1950 4165
rect 1900 4115 1915 4135
rect 1935 4115 1950 4135
rect 1900 4085 1950 4115
rect 1900 4065 1915 4085
rect 1935 4065 1950 4085
rect 1900 4035 1950 4065
rect 1900 4015 1915 4035
rect 1935 4015 1950 4035
rect 1900 3985 1950 4015
rect 1900 3965 1915 3985
rect 1935 3965 1950 3985
rect 1900 3935 1950 3965
rect 1900 3915 1915 3935
rect 1935 3915 1950 3935
rect 1900 3885 1950 3915
rect 1900 3865 1915 3885
rect 1935 3865 1950 3885
rect 1900 3835 1950 3865
rect 1900 3815 1915 3835
rect 1935 3815 1950 3835
rect 1900 3785 1950 3815
rect 1900 3765 1915 3785
rect 1935 3765 1950 3785
rect 1900 3735 1950 3765
rect 1900 3715 1915 3735
rect 1935 3715 1950 3735
rect 1900 3700 1950 3715
rect 2050 4185 2100 4200
rect 2050 4165 2065 4185
rect 2085 4165 2100 4185
rect 2050 4135 2100 4165
rect 2050 4115 2065 4135
rect 2085 4115 2100 4135
rect 2050 4085 2100 4115
rect 2050 4065 2065 4085
rect 2085 4065 2100 4085
rect 2050 4035 2100 4065
rect 2050 4015 2065 4035
rect 2085 4015 2100 4035
rect 2050 3985 2100 4015
rect 2050 3965 2065 3985
rect 2085 3965 2100 3985
rect 2050 3935 2100 3965
rect 2050 3915 2065 3935
rect 2085 3915 2100 3935
rect 2050 3885 2100 3915
rect 2050 3865 2065 3885
rect 2085 3865 2100 3885
rect 2050 3835 2100 3865
rect 2050 3815 2065 3835
rect 2085 3815 2100 3835
rect 2050 3785 2100 3815
rect 2050 3765 2065 3785
rect 2085 3765 2100 3785
rect 2050 3735 2100 3765
rect 2050 3715 2065 3735
rect 2085 3715 2100 3735
rect 2050 3700 2100 3715
rect 2200 4185 2250 4200
rect 2200 4165 2215 4185
rect 2235 4165 2250 4185
rect 2200 4135 2250 4165
rect 2200 4115 2215 4135
rect 2235 4115 2250 4135
rect 2200 4085 2250 4115
rect 2200 4065 2215 4085
rect 2235 4065 2250 4085
rect 2200 4035 2250 4065
rect 2200 4015 2215 4035
rect 2235 4015 2250 4035
rect 2200 3985 2250 4015
rect 2200 3965 2215 3985
rect 2235 3965 2250 3985
rect 2200 3935 2250 3965
rect 2200 3915 2215 3935
rect 2235 3915 2250 3935
rect 2200 3885 2250 3915
rect 2200 3865 2215 3885
rect 2235 3865 2250 3885
rect 2200 3835 2250 3865
rect 2200 3815 2215 3835
rect 2235 3815 2250 3835
rect 2200 3785 2250 3815
rect 2200 3765 2215 3785
rect 2235 3765 2250 3785
rect 2200 3735 2250 3765
rect 2200 3715 2215 3735
rect 2235 3715 2250 3735
rect 2200 3700 2250 3715
rect 2350 4185 2400 4200
rect 2350 4165 2365 4185
rect 2385 4165 2400 4185
rect 2350 4135 2400 4165
rect 2350 4115 2365 4135
rect 2385 4115 2400 4135
rect 2350 4085 2400 4115
rect 2350 4065 2365 4085
rect 2385 4065 2400 4085
rect 2350 4035 2400 4065
rect 2350 4015 2365 4035
rect 2385 4015 2400 4035
rect 2350 3985 2400 4015
rect 2350 3965 2365 3985
rect 2385 3965 2400 3985
rect 2350 3935 2400 3965
rect 2350 3915 2365 3935
rect 2385 3915 2400 3935
rect 2350 3885 2400 3915
rect 2350 3865 2365 3885
rect 2385 3865 2400 3885
rect 2350 3835 2400 3865
rect 2350 3815 2365 3835
rect 2385 3815 2400 3835
rect 2350 3785 2400 3815
rect 2350 3765 2365 3785
rect 2385 3765 2400 3785
rect 2350 3735 2400 3765
rect 2350 3715 2365 3735
rect 2385 3715 2400 3735
rect 2350 3700 2400 3715
rect 2500 4185 2550 4200
rect 2500 4165 2515 4185
rect 2535 4165 2550 4185
rect 2500 4135 2550 4165
rect 2500 4115 2515 4135
rect 2535 4115 2550 4135
rect 2500 4085 2550 4115
rect 2500 4065 2515 4085
rect 2535 4065 2550 4085
rect 2500 4035 2550 4065
rect 2500 4015 2515 4035
rect 2535 4015 2550 4035
rect 2500 3985 2550 4015
rect 2500 3965 2515 3985
rect 2535 3965 2550 3985
rect 2500 3935 2550 3965
rect 2500 3915 2515 3935
rect 2535 3915 2550 3935
rect 2500 3885 2550 3915
rect 2500 3865 2515 3885
rect 2535 3865 2550 3885
rect 2500 3835 2550 3865
rect 2500 3815 2515 3835
rect 2535 3815 2550 3835
rect 2500 3785 2550 3815
rect 2500 3765 2515 3785
rect 2535 3765 2550 3785
rect 2500 3735 2550 3765
rect 2500 3715 2515 3735
rect 2535 3715 2550 3735
rect 2500 3700 2550 3715
rect 2650 4185 2700 4200
rect 2650 4165 2665 4185
rect 2685 4165 2700 4185
rect 2650 4135 2700 4165
rect 2650 4115 2665 4135
rect 2685 4115 2700 4135
rect 2650 4085 2700 4115
rect 2650 4065 2665 4085
rect 2685 4065 2700 4085
rect 2650 4035 2700 4065
rect 2650 4015 2665 4035
rect 2685 4015 2700 4035
rect 2650 3985 2700 4015
rect 2650 3965 2665 3985
rect 2685 3965 2700 3985
rect 2650 3935 2700 3965
rect 2650 3915 2665 3935
rect 2685 3915 2700 3935
rect 2650 3885 2700 3915
rect 2650 3865 2665 3885
rect 2685 3865 2700 3885
rect 2650 3835 2700 3865
rect 2650 3815 2665 3835
rect 2685 3815 2700 3835
rect 2650 3785 2700 3815
rect 2650 3765 2665 3785
rect 2685 3765 2700 3785
rect 2650 3735 2700 3765
rect 2650 3715 2665 3735
rect 2685 3715 2700 3735
rect 2650 3700 2700 3715
rect 2800 4185 2850 4200
rect 2800 4165 2815 4185
rect 2835 4165 2850 4185
rect 2800 4135 2850 4165
rect 2800 4115 2815 4135
rect 2835 4115 2850 4135
rect 2800 4085 2850 4115
rect 2800 4065 2815 4085
rect 2835 4065 2850 4085
rect 2800 4035 2850 4065
rect 2800 4015 2815 4035
rect 2835 4015 2850 4035
rect 2800 3985 2850 4015
rect 2800 3965 2815 3985
rect 2835 3965 2850 3985
rect 2800 3935 2850 3965
rect 2800 3915 2815 3935
rect 2835 3915 2850 3935
rect 2800 3885 2850 3915
rect 2800 3865 2815 3885
rect 2835 3865 2850 3885
rect 2800 3835 2850 3865
rect 2800 3815 2815 3835
rect 2835 3815 2850 3835
rect 2800 3785 2850 3815
rect 2800 3765 2815 3785
rect 2835 3765 2850 3785
rect 2800 3735 2850 3765
rect 2800 3715 2815 3735
rect 2835 3715 2850 3735
rect 2800 3700 2850 3715
rect 2950 4185 3000 4200
rect 2950 4165 2965 4185
rect 2985 4165 3000 4185
rect 2950 4135 3000 4165
rect 2950 4115 2965 4135
rect 2985 4115 3000 4135
rect 2950 4085 3000 4115
rect 2950 4065 2965 4085
rect 2985 4065 3000 4085
rect 2950 4035 3000 4065
rect 2950 4015 2965 4035
rect 2985 4015 3000 4035
rect 2950 3985 3000 4015
rect 2950 3965 2965 3985
rect 2985 3965 3000 3985
rect 2950 3935 3000 3965
rect 2950 3915 2965 3935
rect 2985 3915 3000 3935
rect 2950 3885 3000 3915
rect 2950 3865 2965 3885
rect 2985 3865 3000 3885
rect 2950 3835 3000 3865
rect 2950 3815 2965 3835
rect 2985 3815 3000 3835
rect 2950 3785 3000 3815
rect 2950 3765 2965 3785
rect 2985 3765 3000 3785
rect 2950 3735 3000 3765
rect 2950 3715 2965 3735
rect 2985 3715 3000 3735
rect 2950 3700 3000 3715
rect 3100 4185 3150 4200
rect 3100 4165 3115 4185
rect 3135 4165 3150 4185
rect 3100 4135 3150 4165
rect 3100 4115 3115 4135
rect 3135 4115 3150 4135
rect 3100 4085 3150 4115
rect 3100 4065 3115 4085
rect 3135 4065 3150 4085
rect 3100 4035 3150 4065
rect 3100 4015 3115 4035
rect 3135 4015 3150 4035
rect 3100 3985 3150 4015
rect 3100 3965 3115 3985
rect 3135 3965 3150 3985
rect 3100 3935 3150 3965
rect 3100 3915 3115 3935
rect 3135 3915 3150 3935
rect 3100 3885 3150 3915
rect 3100 3865 3115 3885
rect 3135 3865 3150 3885
rect 3100 3835 3150 3865
rect 3100 3815 3115 3835
rect 3135 3815 3150 3835
rect 3100 3785 3150 3815
rect 3100 3765 3115 3785
rect 3135 3765 3150 3785
rect 3100 3735 3150 3765
rect 3100 3715 3115 3735
rect 3135 3715 3150 3735
rect 3100 3700 3150 3715
rect 3250 4185 3300 4200
rect 3250 4165 3265 4185
rect 3285 4165 3300 4185
rect 3250 4135 3300 4165
rect 3250 4115 3265 4135
rect 3285 4115 3300 4135
rect 3250 4085 3300 4115
rect 3250 4065 3265 4085
rect 3285 4065 3300 4085
rect 3250 4035 3300 4065
rect 3250 4015 3265 4035
rect 3285 4015 3300 4035
rect 3250 3985 3300 4015
rect 3250 3965 3265 3985
rect 3285 3965 3300 3985
rect 3250 3935 3300 3965
rect 3250 3915 3265 3935
rect 3285 3915 3300 3935
rect 3250 3885 3300 3915
rect 3250 3865 3265 3885
rect 3285 3865 3300 3885
rect 3250 3835 3300 3865
rect 3250 3815 3265 3835
rect 3285 3815 3300 3835
rect 3250 3785 3300 3815
rect 3250 3765 3265 3785
rect 3285 3765 3300 3785
rect 3250 3735 3300 3765
rect 3250 3715 3265 3735
rect 3285 3715 3300 3735
rect 3250 3700 3300 3715
rect 3400 4185 3450 4200
rect 3400 4165 3415 4185
rect 3435 4165 3450 4185
rect 3400 4135 3450 4165
rect 3400 4115 3415 4135
rect 3435 4115 3450 4135
rect 3400 4085 3450 4115
rect 3400 4065 3415 4085
rect 3435 4065 3450 4085
rect 3400 4035 3450 4065
rect 3400 4015 3415 4035
rect 3435 4015 3450 4035
rect 3400 3985 3450 4015
rect 3400 3965 3415 3985
rect 3435 3965 3450 3985
rect 3400 3935 3450 3965
rect 3400 3915 3415 3935
rect 3435 3915 3450 3935
rect 3400 3885 3450 3915
rect 3400 3865 3415 3885
rect 3435 3865 3450 3885
rect 3400 3835 3450 3865
rect 3400 3815 3415 3835
rect 3435 3815 3450 3835
rect 3400 3785 3450 3815
rect 3400 3765 3415 3785
rect 3435 3765 3450 3785
rect 3400 3735 3450 3765
rect 3400 3715 3415 3735
rect 3435 3715 3450 3735
rect 3400 3700 3450 3715
rect 3550 4185 3600 4200
rect 3550 4165 3565 4185
rect 3585 4165 3600 4185
rect 3550 4135 3600 4165
rect 3550 4115 3565 4135
rect 3585 4115 3600 4135
rect 3550 4085 3600 4115
rect 3550 4065 3565 4085
rect 3585 4065 3600 4085
rect 3550 4035 3600 4065
rect 3550 4015 3565 4035
rect 3585 4015 3600 4035
rect 3550 3985 3600 4015
rect 3550 3965 3565 3985
rect 3585 3965 3600 3985
rect 3550 3935 3600 3965
rect 3550 3915 3565 3935
rect 3585 3915 3600 3935
rect 3550 3885 3600 3915
rect 3550 3865 3565 3885
rect 3585 3865 3600 3885
rect 3550 3835 3600 3865
rect 3550 3815 3565 3835
rect 3585 3815 3600 3835
rect 3550 3785 3600 3815
rect 3550 3765 3565 3785
rect 3585 3765 3600 3785
rect 3550 3735 3600 3765
rect 3550 3715 3565 3735
rect 3585 3715 3600 3735
rect 3550 3700 3600 3715
rect 3700 3700 3750 4200
rect 3850 3700 3900 4200
rect 4000 3700 4050 4200
rect 4150 4185 4200 4200
rect 4150 4165 4165 4185
rect 4185 4165 4200 4185
rect 4150 4135 4200 4165
rect 4150 4115 4165 4135
rect 4185 4115 4200 4135
rect 4150 4085 4200 4115
rect 4150 4065 4165 4085
rect 4185 4065 4200 4085
rect 4150 4035 4200 4065
rect 4150 4015 4165 4035
rect 4185 4015 4200 4035
rect 4150 3985 4200 4015
rect 4150 3965 4165 3985
rect 4185 3965 4200 3985
rect 4150 3935 4200 3965
rect 4150 3915 4165 3935
rect 4185 3915 4200 3935
rect 4150 3885 4200 3915
rect 4150 3865 4165 3885
rect 4185 3865 4200 3885
rect 4150 3835 4200 3865
rect 4150 3815 4165 3835
rect 4185 3815 4200 3835
rect 4150 3785 4200 3815
rect 4150 3765 4165 3785
rect 4185 3765 4200 3785
rect 4150 3735 4200 3765
rect 4150 3715 4165 3735
rect 4185 3715 4200 3735
rect 4150 3700 4200 3715
rect 4300 3700 4350 4200
rect 4450 3700 4500 4200
rect 4600 3700 4650 4200
rect 4750 4185 4800 4200
rect 4750 4165 4765 4185
rect 4785 4165 4800 4185
rect 4750 4135 4800 4165
rect 4750 4115 4765 4135
rect 4785 4115 4800 4135
rect 4750 4085 4800 4115
rect 4750 4065 4765 4085
rect 4785 4065 4800 4085
rect 4750 4035 4800 4065
rect 4750 4015 4765 4035
rect 4785 4015 4800 4035
rect 4750 3985 4800 4015
rect 4750 3965 4765 3985
rect 4785 3965 4800 3985
rect 4750 3935 4800 3965
rect 4750 3915 4765 3935
rect 4785 3915 4800 3935
rect 4750 3885 4800 3915
rect 4750 3865 4765 3885
rect 4785 3865 4800 3885
rect 4750 3835 4800 3865
rect 4750 3815 4765 3835
rect 4785 3815 4800 3835
rect 4750 3785 4800 3815
rect 4750 3765 4765 3785
rect 4785 3765 4800 3785
rect 4750 3735 4800 3765
rect 4750 3715 4765 3735
rect 4785 3715 4800 3735
rect 4750 3700 4800 3715
rect 4900 4185 4950 4200
rect 4900 4165 4915 4185
rect 4935 4165 4950 4185
rect 4900 4135 4950 4165
rect 4900 4115 4915 4135
rect 4935 4115 4950 4135
rect 4900 4085 4950 4115
rect 4900 4065 4915 4085
rect 4935 4065 4950 4085
rect 4900 4035 4950 4065
rect 4900 4015 4915 4035
rect 4935 4015 4950 4035
rect 4900 3985 4950 4015
rect 4900 3965 4915 3985
rect 4935 3965 4950 3985
rect 4900 3935 4950 3965
rect 4900 3915 4915 3935
rect 4935 3915 4950 3935
rect 4900 3885 4950 3915
rect 4900 3865 4915 3885
rect 4935 3865 4950 3885
rect 4900 3835 4950 3865
rect 4900 3815 4915 3835
rect 4935 3815 4950 3835
rect 4900 3785 4950 3815
rect 4900 3765 4915 3785
rect 4935 3765 4950 3785
rect 4900 3735 4950 3765
rect 4900 3715 4915 3735
rect 4935 3715 4950 3735
rect 4900 3700 4950 3715
rect 5050 4185 5100 4200
rect 5050 4165 5065 4185
rect 5085 4165 5100 4185
rect 5050 4135 5100 4165
rect 5050 4115 5065 4135
rect 5085 4115 5100 4135
rect 5050 4085 5100 4115
rect 5050 4065 5065 4085
rect 5085 4065 5100 4085
rect 5050 4035 5100 4065
rect 5050 4015 5065 4035
rect 5085 4015 5100 4035
rect 5050 3985 5100 4015
rect 5050 3965 5065 3985
rect 5085 3965 5100 3985
rect 5050 3935 5100 3965
rect 5050 3915 5065 3935
rect 5085 3915 5100 3935
rect 5050 3885 5100 3915
rect 5050 3865 5065 3885
rect 5085 3865 5100 3885
rect 5050 3835 5100 3865
rect 5050 3815 5065 3835
rect 5085 3815 5100 3835
rect 5050 3785 5100 3815
rect 5050 3765 5065 3785
rect 5085 3765 5100 3785
rect 5050 3735 5100 3765
rect 5050 3715 5065 3735
rect 5085 3715 5100 3735
rect 5050 3700 5100 3715
rect 5200 4185 5250 4200
rect 5200 4165 5215 4185
rect 5235 4165 5250 4185
rect 5200 4135 5250 4165
rect 5200 4115 5215 4135
rect 5235 4115 5250 4135
rect 5200 4085 5250 4115
rect 5200 4065 5215 4085
rect 5235 4065 5250 4085
rect 5200 4035 5250 4065
rect 5200 4015 5215 4035
rect 5235 4015 5250 4035
rect 5200 3985 5250 4015
rect 5200 3965 5215 3985
rect 5235 3965 5250 3985
rect 5200 3935 5250 3965
rect 5200 3915 5215 3935
rect 5235 3915 5250 3935
rect 5200 3885 5250 3915
rect 5200 3865 5215 3885
rect 5235 3865 5250 3885
rect 5200 3835 5250 3865
rect 5200 3815 5215 3835
rect 5235 3815 5250 3835
rect 5200 3785 5250 3815
rect 5200 3765 5215 3785
rect 5235 3765 5250 3785
rect 5200 3735 5250 3765
rect 5200 3715 5215 3735
rect 5235 3715 5250 3735
rect 5200 3700 5250 3715
rect 5350 4185 5400 4200
rect 5350 4165 5365 4185
rect 5385 4165 5400 4185
rect 5350 4135 5400 4165
rect 5350 4115 5365 4135
rect 5385 4115 5400 4135
rect 5350 4085 5400 4115
rect 5350 4065 5365 4085
rect 5385 4065 5400 4085
rect 5350 4035 5400 4065
rect 5350 4015 5365 4035
rect 5385 4015 5400 4035
rect 5350 3985 5400 4015
rect 5350 3965 5365 3985
rect 5385 3965 5400 3985
rect 5350 3935 5400 3965
rect 5350 3915 5365 3935
rect 5385 3915 5400 3935
rect 5350 3885 5400 3915
rect 5350 3865 5365 3885
rect 5385 3865 5400 3885
rect 5350 3835 5400 3865
rect 5350 3815 5365 3835
rect 5385 3815 5400 3835
rect 5350 3785 5400 3815
rect 5350 3765 5365 3785
rect 5385 3765 5400 3785
rect 5350 3735 5400 3765
rect 5350 3715 5365 3735
rect 5385 3715 5400 3735
rect 5350 3700 5400 3715
rect 5500 4185 5550 4200
rect 5500 4165 5515 4185
rect 5535 4165 5550 4185
rect 5500 4135 5550 4165
rect 5500 4115 5515 4135
rect 5535 4115 5550 4135
rect 5500 4085 5550 4115
rect 5500 4065 5515 4085
rect 5535 4065 5550 4085
rect 5500 4035 5550 4065
rect 5500 4015 5515 4035
rect 5535 4015 5550 4035
rect 5500 3985 5550 4015
rect 5500 3965 5515 3985
rect 5535 3965 5550 3985
rect 5500 3935 5550 3965
rect 5500 3915 5515 3935
rect 5535 3915 5550 3935
rect 5500 3885 5550 3915
rect 5500 3865 5515 3885
rect 5535 3865 5550 3885
rect 5500 3835 5550 3865
rect 5500 3815 5515 3835
rect 5535 3815 5550 3835
rect 5500 3785 5550 3815
rect 5500 3765 5515 3785
rect 5535 3765 5550 3785
rect 5500 3735 5550 3765
rect 5500 3715 5515 3735
rect 5535 3715 5550 3735
rect 5500 3700 5550 3715
rect 5650 4185 5700 4200
rect 5650 4165 5665 4185
rect 5685 4165 5700 4185
rect 5650 4135 5700 4165
rect 5650 4115 5665 4135
rect 5685 4115 5700 4135
rect 5650 4085 5700 4115
rect 5650 4065 5665 4085
rect 5685 4065 5700 4085
rect 5650 4035 5700 4065
rect 5650 4015 5665 4035
rect 5685 4015 5700 4035
rect 5650 3985 5700 4015
rect 5650 3965 5665 3985
rect 5685 3965 5700 3985
rect 5650 3935 5700 3965
rect 5650 3915 5665 3935
rect 5685 3915 5700 3935
rect 5650 3885 5700 3915
rect 5650 3865 5665 3885
rect 5685 3865 5700 3885
rect 5650 3835 5700 3865
rect 5650 3815 5665 3835
rect 5685 3815 5700 3835
rect 5650 3785 5700 3815
rect 5650 3765 5665 3785
rect 5685 3765 5700 3785
rect 5650 3735 5700 3765
rect 5650 3715 5665 3735
rect 5685 3715 5700 3735
rect 5650 3700 5700 3715
rect 5800 4185 5850 4200
rect 5800 4165 5815 4185
rect 5835 4165 5850 4185
rect 5800 4135 5850 4165
rect 5800 4115 5815 4135
rect 5835 4115 5850 4135
rect 5800 4085 5850 4115
rect 5800 4065 5815 4085
rect 5835 4065 5850 4085
rect 5800 4035 5850 4065
rect 5800 4015 5815 4035
rect 5835 4015 5850 4035
rect 5800 3985 5850 4015
rect 5800 3965 5815 3985
rect 5835 3965 5850 3985
rect 5800 3935 5850 3965
rect 5800 3915 5815 3935
rect 5835 3915 5850 3935
rect 5800 3885 5850 3915
rect 5800 3865 5815 3885
rect 5835 3865 5850 3885
rect 5800 3835 5850 3865
rect 5800 3815 5815 3835
rect 5835 3815 5850 3835
rect 5800 3785 5850 3815
rect 5800 3765 5815 3785
rect 5835 3765 5850 3785
rect 5800 3735 5850 3765
rect 5800 3715 5815 3735
rect 5835 3715 5850 3735
rect 5800 3700 5850 3715
rect 5950 4185 6000 4200
rect 5950 4165 5965 4185
rect 5985 4165 6000 4185
rect 5950 4135 6000 4165
rect 5950 4115 5965 4135
rect 5985 4115 6000 4135
rect 5950 4085 6000 4115
rect 5950 4065 5965 4085
rect 5985 4065 6000 4085
rect 5950 4035 6000 4065
rect 5950 4015 5965 4035
rect 5985 4015 6000 4035
rect 5950 3985 6000 4015
rect 5950 3965 5965 3985
rect 5985 3965 6000 3985
rect 5950 3935 6000 3965
rect 5950 3915 5965 3935
rect 5985 3915 6000 3935
rect 5950 3885 6000 3915
rect 5950 3865 5965 3885
rect 5985 3865 6000 3885
rect 5950 3835 6000 3865
rect 5950 3815 5965 3835
rect 5985 3815 6000 3835
rect 5950 3785 6000 3815
rect 5950 3765 5965 3785
rect 5985 3765 6000 3785
rect 5950 3735 6000 3765
rect 5950 3715 5965 3735
rect 5985 3715 6000 3735
rect 5950 3700 6000 3715
rect 6100 4185 6150 4200
rect 6100 4165 6115 4185
rect 6135 4165 6150 4185
rect 6100 4135 6150 4165
rect 6100 4115 6115 4135
rect 6135 4115 6150 4135
rect 6100 4085 6150 4115
rect 6100 4065 6115 4085
rect 6135 4065 6150 4085
rect 6100 4035 6150 4065
rect 6100 4015 6115 4035
rect 6135 4015 6150 4035
rect 6100 3985 6150 4015
rect 6100 3965 6115 3985
rect 6135 3965 6150 3985
rect 6100 3935 6150 3965
rect 6100 3915 6115 3935
rect 6135 3915 6150 3935
rect 6100 3885 6150 3915
rect 6100 3865 6115 3885
rect 6135 3865 6150 3885
rect 6100 3835 6150 3865
rect 6100 3815 6115 3835
rect 6135 3815 6150 3835
rect 6100 3785 6150 3815
rect 6100 3765 6115 3785
rect 6135 3765 6150 3785
rect 6100 3735 6150 3765
rect 6100 3715 6115 3735
rect 6135 3715 6150 3735
rect 6100 3700 6150 3715
rect 6250 4185 6300 4200
rect 6250 4165 6265 4185
rect 6285 4165 6300 4185
rect 6250 4135 6300 4165
rect 6250 4115 6265 4135
rect 6285 4115 6300 4135
rect 6250 4085 6300 4115
rect 6250 4065 6265 4085
rect 6285 4065 6300 4085
rect 6250 4035 6300 4065
rect 6250 4015 6265 4035
rect 6285 4015 6300 4035
rect 6250 3985 6300 4015
rect 6250 3965 6265 3985
rect 6285 3965 6300 3985
rect 6250 3935 6300 3965
rect 6250 3915 6265 3935
rect 6285 3915 6300 3935
rect 6250 3885 6300 3915
rect 6250 3865 6265 3885
rect 6285 3865 6300 3885
rect 6250 3835 6300 3865
rect 6250 3815 6265 3835
rect 6285 3815 6300 3835
rect 6250 3785 6300 3815
rect 6250 3765 6265 3785
rect 6285 3765 6300 3785
rect 6250 3735 6300 3765
rect 6250 3715 6265 3735
rect 6285 3715 6300 3735
rect 6250 3700 6300 3715
rect 6400 4185 6450 4200
rect 6400 4165 6415 4185
rect 6435 4165 6450 4185
rect 6400 4135 6450 4165
rect 6400 4115 6415 4135
rect 6435 4115 6450 4135
rect 6400 4085 6450 4115
rect 6400 4065 6415 4085
rect 6435 4065 6450 4085
rect 6400 4035 6450 4065
rect 6400 4015 6415 4035
rect 6435 4015 6450 4035
rect 6400 3985 6450 4015
rect 6400 3965 6415 3985
rect 6435 3965 6450 3985
rect 6400 3935 6450 3965
rect 6400 3915 6415 3935
rect 6435 3915 6450 3935
rect 6400 3885 6450 3915
rect 6400 3865 6415 3885
rect 6435 3865 6450 3885
rect 6400 3835 6450 3865
rect 6400 3815 6415 3835
rect 6435 3815 6450 3835
rect 6400 3785 6450 3815
rect 6400 3765 6415 3785
rect 6435 3765 6450 3785
rect 6400 3735 6450 3765
rect 6400 3715 6415 3735
rect 6435 3715 6450 3735
rect 6400 3700 6450 3715
rect 6550 4185 6600 4200
rect 6550 4165 6565 4185
rect 6585 4165 6600 4185
rect 6550 4135 6600 4165
rect 6550 4115 6565 4135
rect 6585 4115 6600 4135
rect 6550 4085 6600 4115
rect 6550 4065 6565 4085
rect 6585 4065 6600 4085
rect 6550 4035 6600 4065
rect 6550 4015 6565 4035
rect 6585 4015 6600 4035
rect 6550 3985 6600 4015
rect 6550 3965 6565 3985
rect 6585 3965 6600 3985
rect 6550 3935 6600 3965
rect 6550 3915 6565 3935
rect 6585 3915 6600 3935
rect 6550 3885 6600 3915
rect 6550 3865 6565 3885
rect 6585 3865 6600 3885
rect 6550 3835 6600 3865
rect 6550 3815 6565 3835
rect 6585 3815 6600 3835
rect 6550 3785 6600 3815
rect 6550 3765 6565 3785
rect 6585 3765 6600 3785
rect 6550 3735 6600 3765
rect 6550 3715 6565 3735
rect 6585 3715 6600 3735
rect 6550 3700 6600 3715
rect 6700 4185 6750 4200
rect 6700 4165 6715 4185
rect 6735 4165 6750 4185
rect 6700 4135 6750 4165
rect 6700 4115 6715 4135
rect 6735 4115 6750 4135
rect 6700 4085 6750 4115
rect 6700 4065 6715 4085
rect 6735 4065 6750 4085
rect 6700 4035 6750 4065
rect 6700 4015 6715 4035
rect 6735 4015 6750 4035
rect 6700 3985 6750 4015
rect 6700 3965 6715 3985
rect 6735 3965 6750 3985
rect 6700 3935 6750 3965
rect 6700 3915 6715 3935
rect 6735 3915 6750 3935
rect 6700 3885 6750 3915
rect 6700 3865 6715 3885
rect 6735 3865 6750 3885
rect 6700 3835 6750 3865
rect 6700 3815 6715 3835
rect 6735 3815 6750 3835
rect 6700 3785 6750 3815
rect 6700 3765 6715 3785
rect 6735 3765 6750 3785
rect 6700 3735 6750 3765
rect 6700 3715 6715 3735
rect 6735 3715 6750 3735
rect 6700 3700 6750 3715
rect 6850 4185 6900 4200
rect 6850 4165 6865 4185
rect 6885 4165 6900 4185
rect 6850 4135 6900 4165
rect 6850 4115 6865 4135
rect 6885 4115 6900 4135
rect 6850 4085 6900 4115
rect 6850 4065 6865 4085
rect 6885 4065 6900 4085
rect 6850 4035 6900 4065
rect 6850 4015 6865 4035
rect 6885 4015 6900 4035
rect 6850 3985 6900 4015
rect 6850 3965 6865 3985
rect 6885 3965 6900 3985
rect 6850 3935 6900 3965
rect 6850 3915 6865 3935
rect 6885 3915 6900 3935
rect 6850 3885 6900 3915
rect 6850 3865 6865 3885
rect 6885 3865 6900 3885
rect 6850 3835 6900 3865
rect 6850 3815 6865 3835
rect 6885 3815 6900 3835
rect 6850 3785 6900 3815
rect 6850 3765 6865 3785
rect 6885 3765 6900 3785
rect 6850 3735 6900 3765
rect 6850 3715 6865 3735
rect 6885 3715 6900 3735
rect 6850 3700 6900 3715
rect 7000 4185 7050 4200
rect 7000 4165 7015 4185
rect 7035 4165 7050 4185
rect 7000 4135 7050 4165
rect 7000 4115 7015 4135
rect 7035 4115 7050 4135
rect 7000 4085 7050 4115
rect 7000 4065 7015 4085
rect 7035 4065 7050 4085
rect 7000 4035 7050 4065
rect 7000 4015 7015 4035
rect 7035 4015 7050 4035
rect 7000 3985 7050 4015
rect 7000 3965 7015 3985
rect 7035 3965 7050 3985
rect 7000 3935 7050 3965
rect 7000 3915 7015 3935
rect 7035 3915 7050 3935
rect 7000 3885 7050 3915
rect 7000 3865 7015 3885
rect 7035 3865 7050 3885
rect 7000 3835 7050 3865
rect 7000 3815 7015 3835
rect 7035 3815 7050 3835
rect 7000 3785 7050 3815
rect 7000 3765 7015 3785
rect 7035 3765 7050 3785
rect 7000 3735 7050 3765
rect 7000 3715 7015 3735
rect 7035 3715 7050 3735
rect 7000 3700 7050 3715
rect 7150 4185 7200 4200
rect 7150 4165 7165 4185
rect 7185 4165 7200 4185
rect 7150 4135 7200 4165
rect 7150 4115 7165 4135
rect 7185 4115 7200 4135
rect 7150 4085 7200 4115
rect 7150 4065 7165 4085
rect 7185 4065 7200 4085
rect 7150 4035 7200 4065
rect 7150 4015 7165 4035
rect 7185 4015 7200 4035
rect 7150 3985 7200 4015
rect 7150 3965 7165 3985
rect 7185 3965 7200 3985
rect 7150 3935 7200 3965
rect 7150 3915 7165 3935
rect 7185 3915 7200 3935
rect 7150 3885 7200 3915
rect 7150 3865 7165 3885
rect 7185 3865 7200 3885
rect 7150 3835 7200 3865
rect 7150 3815 7165 3835
rect 7185 3815 7200 3835
rect 7150 3785 7200 3815
rect 7150 3765 7165 3785
rect 7185 3765 7200 3785
rect 7150 3735 7200 3765
rect 7150 3715 7165 3735
rect 7185 3715 7200 3735
rect 7150 3700 7200 3715
rect 7300 4185 7350 4200
rect 7300 4165 7315 4185
rect 7335 4165 7350 4185
rect 7300 4135 7350 4165
rect 7300 4115 7315 4135
rect 7335 4115 7350 4135
rect 7300 4085 7350 4115
rect 7300 4065 7315 4085
rect 7335 4065 7350 4085
rect 7300 4035 7350 4065
rect 7300 4015 7315 4035
rect 7335 4015 7350 4035
rect 7300 3985 7350 4015
rect 7300 3965 7315 3985
rect 7335 3965 7350 3985
rect 7300 3935 7350 3965
rect 7300 3915 7315 3935
rect 7335 3915 7350 3935
rect 7300 3885 7350 3915
rect 7300 3865 7315 3885
rect 7335 3865 7350 3885
rect 7300 3835 7350 3865
rect 7300 3815 7315 3835
rect 7335 3815 7350 3835
rect 7300 3785 7350 3815
rect 7300 3765 7315 3785
rect 7335 3765 7350 3785
rect 7300 3735 7350 3765
rect 7300 3715 7315 3735
rect 7335 3715 7350 3735
rect 7300 3700 7350 3715
rect 7450 4185 7500 4200
rect 7450 4165 7465 4185
rect 7485 4165 7500 4185
rect 7450 4135 7500 4165
rect 7450 4115 7465 4135
rect 7485 4115 7500 4135
rect 7450 4085 7500 4115
rect 7450 4065 7465 4085
rect 7485 4065 7500 4085
rect 7450 4035 7500 4065
rect 7450 4015 7465 4035
rect 7485 4015 7500 4035
rect 7450 3985 7500 4015
rect 7450 3965 7465 3985
rect 7485 3965 7500 3985
rect 7450 3935 7500 3965
rect 7450 3915 7465 3935
rect 7485 3915 7500 3935
rect 7450 3885 7500 3915
rect 7450 3865 7465 3885
rect 7485 3865 7500 3885
rect 7450 3835 7500 3865
rect 7450 3815 7465 3835
rect 7485 3815 7500 3835
rect 7450 3785 7500 3815
rect 7450 3765 7465 3785
rect 7485 3765 7500 3785
rect 7450 3735 7500 3765
rect 7450 3715 7465 3735
rect 7485 3715 7500 3735
rect 7450 3700 7500 3715
rect 7600 4185 7650 4200
rect 7600 4165 7615 4185
rect 7635 4165 7650 4185
rect 7600 4135 7650 4165
rect 7600 4115 7615 4135
rect 7635 4115 7650 4135
rect 7600 4085 7650 4115
rect 7600 4065 7615 4085
rect 7635 4065 7650 4085
rect 7600 4035 7650 4065
rect 7600 4015 7615 4035
rect 7635 4015 7650 4035
rect 7600 3985 7650 4015
rect 7600 3965 7615 3985
rect 7635 3965 7650 3985
rect 7600 3935 7650 3965
rect 7600 3915 7615 3935
rect 7635 3915 7650 3935
rect 7600 3885 7650 3915
rect 7600 3865 7615 3885
rect 7635 3865 7650 3885
rect 7600 3835 7650 3865
rect 7600 3815 7615 3835
rect 7635 3815 7650 3835
rect 7600 3785 7650 3815
rect 7600 3765 7615 3785
rect 7635 3765 7650 3785
rect 7600 3735 7650 3765
rect 7600 3715 7615 3735
rect 7635 3715 7650 3735
rect 7600 3700 7650 3715
rect 7750 4185 7800 4200
rect 7750 4165 7765 4185
rect 7785 4165 7800 4185
rect 7750 4135 7800 4165
rect 7750 4115 7765 4135
rect 7785 4115 7800 4135
rect 7750 4085 7800 4115
rect 7750 4065 7765 4085
rect 7785 4065 7800 4085
rect 7750 4035 7800 4065
rect 7750 4015 7765 4035
rect 7785 4015 7800 4035
rect 7750 3985 7800 4015
rect 7750 3965 7765 3985
rect 7785 3965 7800 3985
rect 7750 3935 7800 3965
rect 7750 3915 7765 3935
rect 7785 3915 7800 3935
rect 7750 3885 7800 3915
rect 7750 3865 7765 3885
rect 7785 3865 7800 3885
rect 7750 3835 7800 3865
rect 7750 3815 7765 3835
rect 7785 3815 7800 3835
rect 7750 3785 7800 3815
rect 7750 3765 7765 3785
rect 7785 3765 7800 3785
rect 7750 3735 7800 3765
rect 7750 3715 7765 3735
rect 7785 3715 7800 3735
rect 7750 3700 7800 3715
rect 7900 3700 7950 4200
rect 8050 3700 8100 4200
rect 8200 3700 8250 4200
rect 8350 4185 8400 4200
rect 8350 4165 8365 4185
rect 8385 4165 8400 4185
rect 8350 4135 8400 4165
rect 8350 4115 8365 4135
rect 8385 4115 8400 4135
rect 8350 4085 8400 4115
rect 8350 4065 8365 4085
rect 8385 4065 8400 4085
rect 8350 4035 8400 4065
rect 8350 4015 8365 4035
rect 8385 4015 8400 4035
rect 8350 3985 8400 4015
rect 8350 3965 8365 3985
rect 8385 3965 8400 3985
rect 8350 3935 8400 3965
rect 8350 3915 8365 3935
rect 8385 3915 8400 3935
rect 8350 3885 8400 3915
rect 8350 3865 8365 3885
rect 8385 3865 8400 3885
rect 8350 3835 8400 3865
rect 8350 3815 8365 3835
rect 8385 3815 8400 3835
rect 8350 3785 8400 3815
rect 8350 3765 8365 3785
rect 8385 3765 8400 3785
rect 8350 3735 8400 3765
rect 8350 3715 8365 3735
rect 8385 3715 8400 3735
rect 8350 3700 8400 3715
rect 8500 4185 8550 4200
rect 8500 4165 8515 4185
rect 8535 4165 8550 4185
rect 8500 4135 8550 4165
rect 8500 4115 8515 4135
rect 8535 4115 8550 4135
rect 8500 4085 8550 4115
rect 8500 4065 8515 4085
rect 8535 4065 8550 4085
rect 8500 4035 8550 4065
rect 8500 4015 8515 4035
rect 8535 4015 8550 4035
rect 8500 3985 8550 4015
rect 8500 3965 8515 3985
rect 8535 3965 8550 3985
rect 8500 3935 8550 3965
rect 8500 3915 8515 3935
rect 8535 3915 8550 3935
rect 8500 3885 8550 3915
rect 8500 3865 8515 3885
rect 8535 3865 8550 3885
rect 8500 3835 8550 3865
rect 8500 3815 8515 3835
rect 8535 3815 8550 3835
rect 8500 3785 8550 3815
rect 8500 3765 8515 3785
rect 8535 3765 8550 3785
rect 8500 3735 8550 3765
rect 8500 3715 8515 3735
rect 8535 3715 8550 3735
rect 8500 3700 8550 3715
rect 8650 4185 8700 4200
rect 8650 4165 8665 4185
rect 8685 4165 8700 4185
rect 8650 4135 8700 4165
rect 8650 4115 8665 4135
rect 8685 4115 8700 4135
rect 8650 4085 8700 4115
rect 8650 4065 8665 4085
rect 8685 4065 8700 4085
rect 8650 4035 8700 4065
rect 8650 4015 8665 4035
rect 8685 4015 8700 4035
rect 8650 3985 8700 4015
rect 8650 3965 8665 3985
rect 8685 3965 8700 3985
rect 8650 3935 8700 3965
rect 8650 3915 8665 3935
rect 8685 3915 8700 3935
rect 8650 3885 8700 3915
rect 8650 3865 8665 3885
rect 8685 3865 8700 3885
rect 8650 3835 8700 3865
rect 8650 3815 8665 3835
rect 8685 3815 8700 3835
rect 8650 3785 8700 3815
rect 8650 3765 8665 3785
rect 8685 3765 8700 3785
rect 8650 3735 8700 3765
rect 8650 3715 8665 3735
rect 8685 3715 8700 3735
rect 8650 3700 8700 3715
rect 8800 4185 8850 4200
rect 8800 4165 8815 4185
rect 8835 4165 8850 4185
rect 8800 4135 8850 4165
rect 8800 4115 8815 4135
rect 8835 4115 8850 4135
rect 8800 4085 8850 4115
rect 8800 4065 8815 4085
rect 8835 4065 8850 4085
rect 8800 4035 8850 4065
rect 8800 4015 8815 4035
rect 8835 4015 8850 4035
rect 8800 3985 8850 4015
rect 8800 3965 8815 3985
rect 8835 3965 8850 3985
rect 8800 3935 8850 3965
rect 8800 3915 8815 3935
rect 8835 3915 8850 3935
rect 8800 3885 8850 3915
rect 8800 3865 8815 3885
rect 8835 3865 8850 3885
rect 8800 3835 8850 3865
rect 8800 3815 8815 3835
rect 8835 3815 8850 3835
rect 8800 3785 8850 3815
rect 8800 3765 8815 3785
rect 8835 3765 8850 3785
rect 8800 3735 8850 3765
rect 8800 3715 8815 3735
rect 8835 3715 8850 3735
rect 8800 3700 8850 3715
rect 8950 4185 9000 4200
rect 8950 4165 8965 4185
rect 8985 4165 9000 4185
rect 8950 4135 9000 4165
rect 8950 4115 8965 4135
rect 8985 4115 9000 4135
rect 8950 4085 9000 4115
rect 8950 4065 8965 4085
rect 8985 4065 9000 4085
rect 8950 4035 9000 4065
rect 8950 4015 8965 4035
rect 8985 4015 9000 4035
rect 8950 3985 9000 4015
rect 8950 3965 8965 3985
rect 8985 3965 9000 3985
rect 8950 3935 9000 3965
rect 8950 3915 8965 3935
rect 8985 3915 9000 3935
rect 8950 3885 9000 3915
rect 8950 3865 8965 3885
rect 8985 3865 9000 3885
rect 8950 3835 9000 3865
rect 8950 3815 8965 3835
rect 8985 3815 9000 3835
rect 8950 3785 9000 3815
rect 8950 3765 8965 3785
rect 8985 3765 9000 3785
rect 8950 3735 9000 3765
rect 8950 3715 8965 3735
rect 8985 3715 9000 3735
rect 8950 3700 9000 3715
rect 9100 4185 9150 4200
rect 9100 4165 9115 4185
rect 9135 4165 9150 4185
rect 9100 4135 9150 4165
rect 9100 4115 9115 4135
rect 9135 4115 9150 4135
rect 9100 4085 9150 4115
rect 9100 4065 9115 4085
rect 9135 4065 9150 4085
rect 9100 4035 9150 4065
rect 9100 4015 9115 4035
rect 9135 4015 9150 4035
rect 9100 3985 9150 4015
rect 9100 3965 9115 3985
rect 9135 3965 9150 3985
rect 9100 3935 9150 3965
rect 9100 3915 9115 3935
rect 9135 3915 9150 3935
rect 9100 3885 9150 3915
rect 9100 3865 9115 3885
rect 9135 3865 9150 3885
rect 9100 3835 9150 3865
rect 9100 3815 9115 3835
rect 9135 3815 9150 3835
rect 9100 3785 9150 3815
rect 9100 3765 9115 3785
rect 9135 3765 9150 3785
rect 9100 3735 9150 3765
rect 9100 3715 9115 3735
rect 9135 3715 9150 3735
rect 9100 3700 9150 3715
rect 9250 4185 9300 4200
rect 9250 4165 9265 4185
rect 9285 4165 9300 4185
rect 9250 4135 9300 4165
rect 9250 4115 9265 4135
rect 9285 4115 9300 4135
rect 9250 4085 9300 4115
rect 9250 4065 9265 4085
rect 9285 4065 9300 4085
rect 9250 4035 9300 4065
rect 9250 4015 9265 4035
rect 9285 4015 9300 4035
rect 9250 3985 9300 4015
rect 9250 3965 9265 3985
rect 9285 3965 9300 3985
rect 9250 3935 9300 3965
rect 9250 3915 9265 3935
rect 9285 3915 9300 3935
rect 9250 3885 9300 3915
rect 9250 3865 9265 3885
rect 9285 3865 9300 3885
rect 9250 3835 9300 3865
rect 9250 3815 9265 3835
rect 9285 3815 9300 3835
rect 9250 3785 9300 3815
rect 9250 3765 9265 3785
rect 9285 3765 9300 3785
rect 9250 3735 9300 3765
rect 9250 3715 9265 3735
rect 9285 3715 9300 3735
rect 9250 3700 9300 3715
rect 9400 4185 9450 4200
rect 9400 4165 9415 4185
rect 9435 4165 9450 4185
rect 9400 4135 9450 4165
rect 9400 4115 9415 4135
rect 9435 4115 9450 4135
rect 9400 4085 9450 4115
rect 9400 4065 9415 4085
rect 9435 4065 9450 4085
rect 9400 4035 9450 4065
rect 9400 4015 9415 4035
rect 9435 4015 9450 4035
rect 9400 3985 9450 4015
rect 9400 3965 9415 3985
rect 9435 3965 9450 3985
rect 9400 3935 9450 3965
rect 9400 3915 9415 3935
rect 9435 3915 9450 3935
rect 9400 3885 9450 3915
rect 9400 3865 9415 3885
rect 9435 3865 9450 3885
rect 9400 3835 9450 3865
rect 9400 3815 9415 3835
rect 9435 3815 9450 3835
rect 9400 3785 9450 3815
rect 9400 3765 9415 3785
rect 9435 3765 9450 3785
rect 9400 3735 9450 3765
rect 9400 3715 9415 3735
rect 9435 3715 9450 3735
rect 9400 3700 9450 3715
rect 9550 4185 9600 4200
rect 9550 4165 9565 4185
rect 9585 4165 9600 4185
rect 9550 4135 9600 4165
rect 9550 4115 9565 4135
rect 9585 4115 9600 4135
rect 9550 4085 9600 4115
rect 9550 4065 9565 4085
rect 9585 4065 9600 4085
rect 9550 4035 9600 4065
rect 9550 4015 9565 4035
rect 9585 4015 9600 4035
rect 9550 3985 9600 4015
rect 9550 3965 9565 3985
rect 9585 3965 9600 3985
rect 9550 3935 9600 3965
rect 9550 3915 9565 3935
rect 9585 3915 9600 3935
rect 9550 3885 9600 3915
rect 9550 3865 9565 3885
rect 9585 3865 9600 3885
rect 9550 3835 9600 3865
rect 9550 3815 9565 3835
rect 9585 3815 9600 3835
rect 9550 3785 9600 3815
rect 9550 3765 9565 3785
rect 9585 3765 9600 3785
rect 9550 3735 9600 3765
rect 9550 3715 9565 3735
rect 9585 3715 9600 3735
rect 9550 3700 9600 3715
rect 9700 4185 9750 4200
rect 9700 4165 9715 4185
rect 9735 4165 9750 4185
rect 9700 4135 9750 4165
rect 9700 4115 9715 4135
rect 9735 4115 9750 4135
rect 9700 4085 9750 4115
rect 9700 4065 9715 4085
rect 9735 4065 9750 4085
rect 9700 4035 9750 4065
rect 9700 4015 9715 4035
rect 9735 4015 9750 4035
rect 9700 3985 9750 4015
rect 9700 3965 9715 3985
rect 9735 3965 9750 3985
rect 9700 3935 9750 3965
rect 9700 3915 9715 3935
rect 9735 3915 9750 3935
rect 9700 3885 9750 3915
rect 9700 3865 9715 3885
rect 9735 3865 9750 3885
rect 9700 3835 9750 3865
rect 9700 3815 9715 3835
rect 9735 3815 9750 3835
rect 9700 3785 9750 3815
rect 9700 3765 9715 3785
rect 9735 3765 9750 3785
rect 9700 3735 9750 3765
rect 9700 3715 9715 3735
rect 9735 3715 9750 3735
rect 9700 3700 9750 3715
rect 9850 4185 9900 4200
rect 9850 4165 9865 4185
rect 9885 4165 9900 4185
rect 9850 4135 9900 4165
rect 9850 4115 9865 4135
rect 9885 4115 9900 4135
rect 9850 4085 9900 4115
rect 9850 4065 9865 4085
rect 9885 4065 9900 4085
rect 9850 4035 9900 4065
rect 9850 4015 9865 4035
rect 9885 4015 9900 4035
rect 9850 3985 9900 4015
rect 9850 3965 9865 3985
rect 9885 3965 9900 3985
rect 9850 3935 9900 3965
rect 9850 3915 9865 3935
rect 9885 3915 9900 3935
rect 9850 3885 9900 3915
rect 9850 3865 9865 3885
rect 9885 3865 9900 3885
rect 9850 3835 9900 3865
rect 9850 3815 9865 3835
rect 9885 3815 9900 3835
rect 9850 3785 9900 3815
rect 9850 3765 9865 3785
rect 9885 3765 9900 3785
rect 9850 3735 9900 3765
rect 9850 3715 9865 3735
rect 9885 3715 9900 3735
rect 9850 3700 9900 3715
rect 10000 4185 10050 4200
rect 10000 4165 10015 4185
rect 10035 4165 10050 4185
rect 10000 4135 10050 4165
rect 10000 4115 10015 4135
rect 10035 4115 10050 4135
rect 10000 4085 10050 4115
rect 10000 4065 10015 4085
rect 10035 4065 10050 4085
rect 10000 4035 10050 4065
rect 10000 4015 10015 4035
rect 10035 4015 10050 4035
rect 10000 3985 10050 4015
rect 10000 3965 10015 3985
rect 10035 3965 10050 3985
rect 10000 3935 10050 3965
rect 10000 3915 10015 3935
rect 10035 3915 10050 3935
rect 10000 3885 10050 3915
rect 10000 3865 10015 3885
rect 10035 3865 10050 3885
rect 10000 3835 10050 3865
rect 10000 3815 10015 3835
rect 10035 3815 10050 3835
rect 10000 3785 10050 3815
rect 10000 3765 10015 3785
rect 10035 3765 10050 3785
rect 10000 3735 10050 3765
rect 10000 3715 10015 3735
rect 10035 3715 10050 3735
rect 10000 3700 10050 3715
rect 10150 4185 10200 4200
rect 10150 4165 10165 4185
rect 10185 4165 10200 4185
rect 10150 4135 10200 4165
rect 10150 4115 10165 4135
rect 10185 4115 10200 4135
rect 10150 4085 10200 4115
rect 10150 4065 10165 4085
rect 10185 4065 10200 4085
rect 10150 4035 10200 4065
rect 10150 4015 10165 4035
rect 10185 4015 10200 4035
rect 10150 3985 10200 4015
rect 10150 3965 10165 3985
rect 10185 3965 10200 3985
rect 10150 3935 10200 3965
rect 10150 3915 10165 3935
rect 10185 3915 10200 3935
rect 10150 3885 10200 3915
rect 10150 3865 10165 3885
rect 10185 3865 10200 3885
rect 10150 3835 10200 3865
rect 10150 3815 10165 3835
rect 10185 3815 10200 3835
rect 10150 3785 10200 3815
rect 10150 3765 10165 3785
rect 10185 3765 10200 3785
rect 10150 3735 10200 3765
rect 10150 3715 10165 3735
rect 10185 3715 10200 3735
rect 10150 3700 10200 3715
rect 10300 4185 10350 4200
rect 10300 4165 10315 4185
rect 10335 4165 10350 4185
rect 10300 4135 10350 4165
rect 10300 4115 10315 4135
rect 10335 4115 10350 4135
rect 10300 4085 10350 4115
rect 10300 4065 10315 4085
rect 10335 4065 10350 4085
rect 10300 4035 10350 4065
rect 10300 4015 10315 4035
rect 10335 4015 10350 4035
rect 10300 3985 10350 4015
rect 10300 3965 10315 3985
rect 10335 3965 10350 3985
rect 10300 3935 10350 3965
rect 10300 3915 10315 3935
rect 10335 3915 10350 3935
rect 10300 3885 10350 3915
rect 10300 3865 10315 3885
rect 10335 3865 10350 3885
rect 10300 3835 10350 3865
rect 10300 3815 10315 3835
rect 10335 3815 10350 3835
rect 10300 3785 10350 3815
rect 10300 3765 10315 3785
rect 10335 3765 10350 3785
rect 10300 3735 10350 3765
rect 10300 3715 10315 3735
rect 10335 3715 10350 3735
rect 10300 3700 10350 3715
rect 10450 4185 10500 4200
rect 10450 4165 10465 4185
rect 10485 4165 10500 4185
rect 10450 4135 10500 4165
rect 10450 4115 10465 4135
rect 10485 4115 10500 4135
rect 10450 4085 10500 4115
rect 10450 4065 10465 4085
rect 10485 4065 10500 4085
rect 10450 4035 10500 4065
rect 10450 4015 10465 4035
rect 10485 4015 10500 4035
rect 10450 3985 10500 4015
rect 10450 3965 10465 3985
rect 10485 3965 10500 3985
rect 10450 3935 10500 3965
rect 10450 3915 10465 3935
rect 10485 3915 10500 3935
rect 10450 3885 10500 3915
rect 10450 3865 10465 3885
rect 10485 3865 10500 3885
rect 10450 3835 10500 3865
rect 10450 3815 10465 3835
rect 10485 3815 10500 3835
rect 10450 3785 10500 3815
rect 10450 3765 10465 3785
rect 10485 3765 10500 3785
rect 10450 3735 10500 3765
rect 10450 3715 10465 3735
rect 10485 3715 10500 3735
rect 10450 3700 10500 3715
rect 10600 4185 10650 4200
rect 10600 4165 10615 4185
rect 10635 4165 10650 4185
rect 10600 4135 10650 4165
rect 10600 4115 10615 4135
rect 10635 4115 10650 4135
rect 10600 4085 10650 4115
rect 10600 4065 10615 4085
rect 10635 4065 10650 4085
rect 10600 4035 10650 4065
rect 10600 4015 10615 4035
rect 10635 4015 10650 4035
rect 10600 3985 10650 4015
rect 10600 3965 10615 3985
rect 10635 3965 10650 3985
rect 10600 3935 10650 3965
rect 10600 3915 10615 3935
rect 10635 3915 10650 3935
rect 10600 3885 10650 3915
rect 10600 3865 10615 3885
rect 10635 3865 10650 3885
rect 10600 3835 10650 3865
rect 10600 3815 10615 3835
rect 10635 3815 10650 3835
rect 10600 3785 10650 3815
rect 10600 3765 10615 3785
rect 10635 3765 10650 3785
rect 10600 3735 10650 3765
rect 10600 3715 10615 3735
rect 10635 3715 10650 3735
rect 10600 3700 10650 3715
rect 10750 4185 10800 4200
rect 10750 4165 10765 4185
rect 10785 4165 10800 4185
rect 10750 4135 10800 4165
rect 10750 4115 10765 4135
rect 10785 4115 10800 4135
rect 10750 4085 10800 4115
rect 10750 4065 10765 4085
rect 10785 4065 10800 4085
rect 10750 4035 10800 4065
rect 10750 4015 10765 4035
rect 10785 4015 10800 4035
rect 10750 3985 10800 4015
rect 10750 3965 10765 3985
rect 10785 3965 10800 3985
rect 10750 3935 10800 3965
rect 10750 3915 10765 3935
rect 10785 3915 10800 3935
rect 10750 3885 10800 3915
rect 10750 3865 10765 3885
rect 10785 3865 10800 3885
rect 10750 3835 10800 3865
rect 10750 3815 10765 3835
rect 10785 3815 10800 3835
rect 10750 3785 10800 3815
rect 10750 3765 10765 3785
rect 10785 3765 10800 3785
rect 10750 3735 10800 3765
rect 10750 3715 10765 3735
rect 10785 3715 10800 3735
rect 10750 3700 10800 3715
rect 10900 3700 10950 4200
rect 11050 3700 11100 4200
rect 11200 3700 11250 4200
rect 11350 4185 11400 4200
rect 11350 4165 11365 4185
rect 11385 4165 11400 4185
rect 11350 4135 11400 4165
rect 11350 4115 11365 4135
rect 11385 4115 11400 4135
rect 11350 4085 11400 4115
rect 11350 4065 11365 4085
rect 11385 4065 11400 4085
rect 11350 4035 11400 4065
rect 11350 4015 11365 4035
rect 11385 4015 11400 4035
rect 11350 3985 11400 4015
rect 11350 3965 11365 3985
rect 11385 3965 11400 3985
rect 11350 3935 11400 3965
rect 11350 3915 11365 3935
rect 11385 3915 11400 3935
rect 11350 3885 11400 3915
rect 11350 3865 11365 3885
rect 11385 3865 11400 3885
rect 11350 3835 11400 3865
rect 11350 3815 11365 3835
rect 11385 3815 11400 3835
rect 11350 3785 11400 3815
rect 11350 3765 11365 3785
rect 11385 3765 11400 3785
rect 11350 3735 11400 3765
rect 11350 3715 11365 3735
rect 11385 3715 11400 3735
rect 11350 3700 11400 3715
rect 11500 3700 11550 4200
rect 11650 3700 11700 4200
rect 11800 3700 11850 4200
rect 11950 4185 12000 4200
rect 11950 4165 11965 4185
rect 11985 4165 12000 4185
rect 11950 4135 12000 4165
rect 11950 4115 11965 4135
rect 11985 4115 12000 4135
rect 11950 4085 12000 4115
rect 11950 4065 11965 4085
rect 11985 4065 12000 4085
rect 11950 4035 12000 4065
rect 11950 4015 11965 4035
rect 11985 4015 12000 4035
rect 11950 3985 12000 4015
rect 11950 3965 11965 3985
rect 11985 3965 12000 3985
rect 11950 3935 12000 3965
rect 11950 3915 11965 3935
rect 11985 3915 12000 3935
rect 11950 3885 12000 3915
rect 11950 3865 11965 3885
rect 11985 3865 12000 3885
rect 11950 3835 12000 3865
rect 11950 3815 11965 3835
rect 11985 3815 12000 3835
rect 11950 3785 12000 3815
rect 11950 3765 11965 3785
rect 11985 3765 12000 3785
rect 11950 3735 12000 3765
rect 11950 3715 11965 3735
rect 11985 3715 12000 3735
rect 11950 3700 12000 3715
rect 12100 3700 12150 4200
rect 12250 3700 12300 4200
rect 12400 3700 12450 4200
rect 12550 4185 12600 4200
rect 12550 4165 12565 4185
rect 12585 4165 12600 4185
rect 12550 4135 12600 4165
rect 12550 4115 12565 4135
rect 12585 4115 12600 4135
rect 12550 4085 12600 4115
rect 12550 4065 12565 4085
rect 12585 4065 12600 4085
rect 12550 4035 12600 4065
rect 12550 4015 12565 4035
rect 12585 4015 12600 4035
rect 12550 3985 12600 4015
rect 12550 3965 12565 3985
rect 12585 3965 12600 3985
rect 12550 3935 12600 3965
rect 12550 3915 12565 3935
rect 12585 3915 12600 3935
rect 12550 3885 12600 3915
rect 12550 3865 12565 3885
rect 12585 3865 12600 3885
rect 12550 3835 12600 3865
rect 12550 3815 12565 3835
rect 12585 3815 12600 3835
rect 12550 3785 12600 3815
rect 12550 3765 12565 3785
rect 12585 3765 12600 3785
rect 12550 3735 12600 3765
rect 12550 3715 12565 3735
rect 12585 3715 12600 3735
rect 12550 3700 12600 3715
rect 12700 3700 12750 4200
rect 12850 3700 12900 4200
rect 13000 3700 13050 4200
rect 13150 4185 13200 4200
rect 13150 4165 13165 4185
rect 13185 4165 13200 4185
rect 13150 4135 13200 4165
rect 13150 4115 13165 4135
rect 13185 4115 13200 4135
rect 13150 4085 13200 4115
rect 13150 4065 13165 4085
rect 13185 4065 13200 4085
rect 13150 4035 13200 4065
rect 13150 4015 13165 4035
rect 13185 4015 13200 4035
rect 13150 3985 13200 4015
rect 13150 3965 13165 3985
rect 13185 3965 13200 3985
rect 13150 3935 13200 3965
rect 13150 3915 13165 3935
rect 13185 3915 13200 3935
rect 13150 3885 13200 3915
rect 13150 3865 13165 3885
rect 13185 3865 13200 3885
rect 13150 3835 13200 3865
rect 13150 3815 13165 3835
rect 13185 3815 13200 3835
rect 13150 3785 13200 3815
rect 13150 3765 13165 3785
rect 13185 3765 13200 3785
rect 13150 3735 13200 3765
rect 13150 3715 13165 3735
rect 13185 3715 13200 3735
rect 13150 3700 13200 3715
rect 13300 3700 13350 4200
rect 13450 3700 13500 4200
rect 13600 3700 13650 4200
rect 13750 4185 13800 4200
rect 13750 4165 13765 4185
rect 13785 4165 13800 4185
rect 13750 4135 13800 4165
rect 13750 4115 13765 4135
rect 13785 4115 13800 4135
rect 13750 4085 13800 4115
rect 13750 4065 13765 4085
rect 13785 4065 13800 4085
rect 13750 4035 13800 4065
rect 13750 4015 13765 4035
rect 13785 4015 13800 4035
rect 13750 3985 13800 4015
rect 13750 3965 13765 3985
rect 13785 3965 13800 3985
rect 13750 3935 13800 3965
rect 13750 3915 13765 3935
rect 13785 3915 13800 3935
rect 13750 3885 13800 3915
rect 13750 3865 13765 3885
rect 13785 3865 13800 3885
rect 13750 3835 13800 3865
rect 13750 3815 13765 3835
rect 13785 3815 13800 3835
rect 13750 3785 13800 3815
rect 13750 3765 13765 3785
rect 13785 3765 13800 3785
rect 13750 3735 13800 3765
rect 13750 3715 13765 3735
rect 13785 3715 13800 3735
rect 13750 3700 13800 3715
rect 13900 3700 13950 4200
rect 14050 3700 14100 4200
rect 14200 3700 14250 4200
rect 14350 4185 14400 4200
rect 14350 4165 14365 4185
rect 14385 4165 14400 4185
rect 14350 4135 14400 4165
rect 14350 4115 14365 4135
rect 14385 4115 14400 4135
rect 14350 4085 14400 4115
rect 14350 4065 14365 4085
rect 14385 4065 14400 4085
rect 14350 4035 14400 4065
rect 14350 4015 14365 4035
rect 14385 4015 14400 4035
rect 14350 3985 14400 4015
rect 14350 3965 14365 3985
rect 14385 3965 14400 3985
rect 14350 3935 14400 3965
rect 14350 3915 14365 3935
rect 14385 3915 14400 3935
rect 14350 3885 14400 3915
rect 14350 3865 14365 3885
rect 14385 3865 14400 3885
rect 14350 3835 14400 3865
rect 14350 3815 14365 3835
rect 14385 3815 14400 3835
rect 14350 3785 14400 3815
rect 14350 3765 14365 3785
rect 14385 3765 14400 3785
rect 14350 3735 14400 3765
rect 14350 3715 14365 3735
rect 14385 3715 14400 3735
rect 14350 3700 14400 3715
rect 14500 3700 14550 4200
rect 14650 3700 14700 4200
rect 14800 3700 14850 4200
rect 14950 4185 15000 4200
rect 14950 4165 14965 4185
rect 14985 4165 15000 4185
rect 14950 4135 15000 4165
rect 14950 4115 14965 4135
rect 14985 4115 15000 4135
rect 14950 4085 15000 4115
rect 14950 4065 14965 4085
rect 14985 4065 15000 4085
rect 14950 4035 15000 4065
rect 14950 4015 14965 4035
rect 14985 4015 15000 4035
rect 14950 3985 15000 4015
rect 14950 3965 14965 3985
rect 14985 3965 15000 3985
rect 14950 3935 15000 3965
rect 14950 3915 14965 3935
rect 14985 3915 15000 3935
rect 14950 3885 15000 3915
rect 14950 3865 14965 3885
rect 14985 3865 15000 3885
rect 14950 3835 15000 3865
rect 14950 3815 14965 3835
rect 14985 3815 15000 3835
rect 14950 3785 15000 3815
rect 14950 3765 14965 3785
rect 14985 3765 15000 3785
rect 14950 3735 15000 3765
rect 14950 3715 14965 3735
rect 14985 3715 15000 3735
rect 14950 3700 15000 3715
rect 15100 3700 15150 4200
rect 15250 3700 15300 4200
rect 15400 3700 15450 4200
rect 15550 4185 15600 4200
rect 15550 4165 15565 4185
rect 15585 4165 15600 4185
rect 15550 4135 15600 4165
rect 15550 4115 15565 4135
rect 15585 4115 15600 4135
rect 15550 4085 15600 4115
rect 15550 4065 15565 4085
rect 15585 4065 15600 4085
rect 15550 4035 15600 4065
rect 15550 4015 15565 4035
rect 15585 4015 15600 4035
rect 15550 3985 15600 4015
rect 15550 3965 15565 3985
rect 15585 3965 15600 3985
rect 15550 3935 15600 3965
rect 15550 3915 15565 3935
rect 15585 3915 15600 3935
rect 15550 3885 15600 3915
rect 15550 3865 15565 3885
rect 15585 3865 15600 3885
rect 15550 3835 15600 3865
rect 15550 3815 15565 3835
rect 15585 3815 15600 3835
rect 15550 3785 15600 3815
rect 15550 3765 15565 3785
rect 15585 3765 15600 3785
rect 15550 3735 15600 3765
rect 15550 3715 15565 3735
rect 15585 3715 15600 3735
rect 15550 3700 15600 3715
rect 15700 3700 15750 4200
rect 15850 3700 15900 4200
rect 16000 3700 16050 4200
rect 16150 4185 16200 4200
rect 16150 4165 16165 4185
rect 16185 4165 16200 4185
rect 16150 4135 16200 4165
rect 16150 4115 16165 4135
rect 16185 4115 16200 4135
rect 16150 4085 16200 4115
rect 16150 4065 16165 4085
rect 16185 4065 16200 4085
rect 16150 4035 16200 4065
rect 16150 4015 16165 4035
rect 16185 4015 16200 4035
rect 16150 3985 16200 4015
rect 16150 3965 16165 3985
rect 16185 3965 16200 3985
rect 16150 3935 16200 3965
rect 16150 3915 16165 3935
rect 16185 3915 16200 3935
rect 16150 3885 16200 3915
rect 16150 3865 16165 3885
rect 16185 3865 16200 3885
rect 16150 3835 16200 3865
rect 16150 3815 16165 3835
rect 16185 3815 16200 3835
rect 16150 3785 16200 3815
rect 16150 3765 16165 3785
rect 16185 3765 16200 3785
rect 16150 3735 16200 3765
rect 16150 3715 16165 3735
rect 16185 3715 16200 3735
rect 16150 3700 16200 3715
rect 16300 4185 16350 4200
rect 16300 4165 16315 4185
rect 16335 4165 16350 4185
rect 16300 4135 16350 4165
rect 16300 4115 16315 4135
rect 16335 4115 16350 4135
rect 16300 4085 16350 4115
rect 16300 4065 16315 4085
rect 16335 4065 16350 4085
rect 16300 4035 16350 4065
rect 16300 4015 16315 4035
rect 16335 4015 16350 4035
rect 16300 3985 16350 4015
rect 16300 3965 16315 3985
rect 16335 3965 16350 3985
rect 16300 3935 16350 3965
rect 16300 3915 16315 3935
rect 16335 3915 16350 3935
rect 16300 3885 16350 3915
rect 16300 3865 16315 3885
rect 16335 3865 16350 3885
rect 16300 3835 16350 3865
rect 16300 3815 16315 3835
rect 16335 3815 16350 3835
rect 16300 3785 16350 3815
rect 16300 3765 16315 3785
rect 16335 3765 16350 3785
rect 16300 3735 16350 3765
rect 16300 3715 16315 3735
rect 16335 3715 16350 3735
rect 16300 3700 16350 3715
rect 16450 4185 16500 4200
rect 16450 4165 16465 4185
rect 16485 4165 16500 4185
rect 16450 4135 16500 4165
rect 16450 4115 16465 4135
rect 16485 4115 16500 4135
rect 16450 4085 16500 4115
rect 16450 4065 16465 4085
rect 16485 4065 16500 4085
rect 16450 4035 16500 4065
rect 16450 4015 16465 4035
rect 16485 4015 16500 4035
rect 16450 3985 16500 4015
rect 16450 3965 16465 3985
rect 16485 3965 16500 3985
rect 16450 3935 16500 3965
rect 16450 3915 16465 3935
rect 16485 3915 16500 3935
rect 16450 3885 16500 3915
rect 16450 3865 16465 3885
rect 16485 3865 16500 3885
rect 16450 3835 16500 3865
rect 16450 3815 16465 3835
rect 16485 3815 16500 3835
rect 16450 3785 16500 3815
rect 16450 3765 16465 3785
rect 16485 3765 16500 3785
rect 16450 3735 16500 3765
rect 16450 3715 16465 3735
rect 16485 3715 16500 3735
rect 16450 3700 16500 3715
rect 16600 4185 16650 4200
rect 16600 4165 16615 4185
rect 16635 4165 16650 4185
rect 16600 4135 16650 4165
rect 16600 4115 16615 4135
rect 16635 4115 16650 4135
rect 16600 4085 16650 4115
rect 16600 4065 16615 4085
rect 16635 4065 16650 4085
rect 16600 4035 16650 4065
rect 16600 4015 16615 4035
rect 16635 4015 16650 4035
rect 16600 3985 16650 4015
rect 16600 3965 16615 3985
rect 16635 3965 16650 3985
rect 16600 3935 16650 3965
rect 16600 3915 16615 3935
rect 16635 3915 16650 3935
rect 16600 3885 16650 3915
rect 16600 3865 16615 3885
rect 16635 3865 16650 3885
rect 16600 3835 16650 3865
rect 16600 3815 16615 3835
rect 16635 3815 16650 3835
rect 16600 3785 16650 3815
rect 16600 3765 16615 3785
rect 16635 3765 16650 3785
rect 16600 3735 16650 3765
rect 16600 3715 16615 3735
rect 16635 3715 16650 3735
rect 16600 3700 16650 3715
rect 16750 4185 16800 4200
rect 16750 4165 16765 4185
rect 16785 4165 16800 4185
rect 16750 4135 16800 4165
rect 16750 4115 16765 4135
rect 16785 4115 16800 4135
rect 16750 4085 16800 4115
rect 16750 4065 16765 4085
rect 16785 4065 16800 4085
rect 16750 4035 16800 4065
rect 16750 4015 16765 4035
rect 16785 4015 16800 4035
rect 16750 3985 16800 4015
rect 16750 3965 16765 3985
rect 16785 3965 16800 3985
rect 16750 3935 16800 3965
rect 16750 3915 16765 3935
rect 16785 3915 16800 3935
rect 16750 3885 16800 3915
rect 16750 3865 16765 3885
rect 16785 3865 16800 3885
rect 16750 3835 16800 3865
rect 16750 3815 16765 3835
rect 16785 3815 16800 3835
rect 16750 3785 16800 3815
rect 16750 3765 16765 3785
rect 16785 3765 16800 3785
rect 16750 3735 16800 3765
rect 16750 3715 16765 3735
rect 16785 3715 16800 3735
rect 16750 3700 16800 3715
rect 16900 4185 16950 4200
rect 16900 4165 16915 4185
rect 16935 4165 16950 4185
rect 16900 4135 16950 4165
rect 16900 4115 16915 4135
rect 16935 4115 16950 4135
rect 16900 4085 16950 4115
rect 16900 4065 16915 4085
rect 16935 4065 16950 4085
rect 16900 4035 16950 4065
rect 16900 4015 16915 4035
rect 16935 4015 16950 4035
rect 16900 3985 16950 4015
rect 16900 3965 16915 3985
rect 16935 3965 16950 3985
rect 16900 3935 16950 3965
rect 16900 3915 16915 3935
rect 16935 3915 16950 3935
rect 16900 3885 16950 3915
rect 16900 3865 16915 3885
rect 16935 3865 16950 3885
rect 16900 3835 16950 3865
rect 16900 3815 16915 3835
rect 16935 3815 16950 3835
rect 16900 3785 16950 3815
rect 16900 3765 16915 3785
rect 16935 3765 16950 3785
rect 16900 3735 16950 3765
rect 16900 3715 16915 3735
rect 16935 3715 16950 3735
rect 16900 3700 16950 3715
rect 17050 4185 17100 4200
rect 17050 4165 17065 4185
rect 17085 4165 17100 4185
rect 17050 4135 17100 4165
rect 17050 4115 17065 4135
rect 17085 4115 17100 4135
rect 17050 4085 17100 4115
rect 17050 4065 17065 4085
rect 17085 4065 17100 4085
rect 17050 4035 17100 4065
rect 17050 4015 17065 4035
rect 17085 4015 17100 4035
rect 17050 3985 17100 4015
rect 17050 3965 17065 3985
rect 17085 3965 17100 3985
rect 17050 3935 17100 3965
rect 17050 3915 17065 3935
rect 17085 3915 17100 3935
rect 17050 3885 17100 3915
rect 17050 3865 17065 3885
rect 17085 3865 17100 3885
rect 17050 3835 17100 3865
rect 17050 3815 17065 3835
rect 17085 3815 17100 3835
rect 17050 3785 17100 3815
rect 17050 3765 17065 3785
rect 17085 3765 17100 3785
rect 17050 3735 17100 3765
rect 17050 3715 17065 3735
rect 17085 3715 17100 3735
rect 17050 3700 17100 3715
rect 17200 4185 17250 4200
rect 17200 4165 17215 4185
rect 17235 4165 17250 4185
rect 17200 4135 17250 4165
rect 17200 4115 17215 4135
rect 17235 4115 17250 4135
rect 17200 4085 17250 4115
rect 17200 4065 17215 4085
rect 17235 4065 17250 4085
rect 17200 4035 17250 4065
rect 17200 4015 17215 4035
rect 17235 4015 17250 4035
rect 17200 3985 17250 4015
rect 17200 3965 17215 3985
rect 17235 3965 17250 3985
rect 17200 3935 17250 3965
rect 17200 3915 17215 3935
rect 17235 3915 17250 3935
rect 17200 3885 17250 3915
rect 17200 3865 17215 3885
rect 17235 3865 17250 3885
rect 17200 3835 17250 3865
rect 17200 3815 17215 3835
rect 17235 3815 17250 3835
rect 17200 3785 17250 3815
rect 17200 3765 17215 3785
rect 17235 3765 17250 3785
rect 17200 3735 17250 3765
rect 17200 3715 17215 3735
rect 17235 3715 17250 3735
rect 17200 3700 17250 3715
rect 17350 4185 17400 4200
rect 17350 4165 17365 4185
rect 17385 4165 17400 4185
rect 17350 4135 17400 4165
rect 17350 4115 17365 4135
rect 17385 4115 17400 4135
rect 17350 4085 17400 4115
rect 17350 4065 17365 4085
rect 17385 4065 17400 4085
rect 17350 4035 17400 4065
rect 17350 4015 17365 4035
rect 17385 4015 17400 4035
rect 17350 3985 17400 4015
rect 17350 3965 17365 3985
rect 17385 3965 17400 3985
rect 17350 3935 17400 3965
rect 17350 3915 17365 3935
rect 17385 3915 17400 3935
rect 17350 3885 17400 3915
rect 17350 3865 17365 3885
rect 17385 3865 17400 3885
rect 17350 3835 17400 3865
rect 17350 3815 17365 3835
rect 17385 3815 17400 3835
rect 17350 3785 17400 3815
rect 17350 3765 17365 3785
rect 17385 3765 17400 3785
rect 17350 3735 17400 3765
rect 17350 3715 17365 3735
rect 17385 3715 17400 3735
rect 17350 3700 17400 3715
rect 17500 3700 17550 4200
rect 17650 3700 17700 4200
rect 17800 3700 17850 4200
rect 17950 4185 18000 4200
rect 17950 4165 17965 4185
rect 17985 4165 18000 4185
rect 17950 4135 18000 4165
rect 17950 4115 17965 4135
rect 17985 4115 18000 4135
rect 17950 4085 18000 4115
rect 17950 4065 17965 4085
rect 17985 4065 18000 4085
rect 17950 4035 18000 4065
rect 17950 4015 17965 4035
rect 17985 4015 18000 4035
rect 17950 3985 18000 4015
rect 17950 3965 17965 3985
rect 17985 3965 18000 3985
rect 17950 3935 18000 3965
rect 17950 3915 17965 3935
rect 17985 3915 18000 3935
rect 17950 3885 18000 3915
rect 17950 3865 17965 3885
rect 17985 3865 18000 3885
rect 17950 3835 18000 3865
rect 17950 3815 17965 3835
rect 17985 3815 18000 3835
rect 17950 3785 18000 3815
rect 17950 3765 17965 3785
rect 17985 3765 18000 3785
rect 17950 3735 18000 3765
rect 17950 3715 17965 3735
rect 17985 3715 18000 3735
rect 17950 3700 18000 3715
rect 18100 3700 18150 4200
rect 18250 3700 18300 4200
rect 18400 3700 18450 4200
rect 18550 4185 18600 4200
rect 18550 4165 18565 4185
rect 18585 4165 18600 4185
rect 18550 4135 18600 4165
rect 18550 4115 18565 4135
rect 18585 4115 18600 4135
rect 18550 4085 18600 4115
rect 18550 4065 18565 4085
rect 18585 4065 18600 4085
rect 18550 4035 18600 4065
rect 18550 4015 18565 4035
rect 18585 4015 18600 4035
rect 18550 3985 18600 4015
rect 18550 3965 18565 3985
rect 18585 3965 18600 3985
rect 18550 3935 18600 3965
rect 18550 3915 18565 3935
rect 18585 3915 18600 3935
rect 18550 3885 18600 3915
rect 18550 3865 18565 3885
rect 18585 3865 18600 3885
rect 18550 3835 18600 3865
rect 18550 3815 18565 3835
rect 18585 3815 18600 3835
rect 18550 3785 18600 3815
rect 18550 3765 18565 3785
rect 18585 3765 18600 3785
rect 18550 3735 18600 3765
rect 18550 3715 18565 3735
rect 18585 3715 18600 3735
rect 18550 3700 18600 3715
rect 18700 4185 18750 4200
rect 18700 4165 18715 4185
rect 18735 4165 18750 4185
rect 18700 4135 18750 4165
rect 18700 4115 18715 4135
rect 18735 4115 18750 4135
rect 18700 4085 18750 4115
rect 18700 4065 18715 4085
rect 18735 4065 18750 4085
rect 18700 4035 18750 4065
rect 18700 4015 18715 4035
rect 18735 4015 18750 4035
rect 18700 3985 18750 4015
rect 18700 3965 18715 3985
rect 18735 3965 18750 3985
rect 18700 3935 18750 3965
rect 18700 3915 18715 3935
rect 18735 3915 18750 3935
rect 18700 3885 18750 3915
rect 18700 3865 18715 3885
rect 18735 3865 18750 3885
rect 18700 3835 18750 3865
rect 18700 3815 18715 3835
rect 18735 3815 18750 3835
rect 18700 3785 18750 3815
rect 18700 3765 18715 3785
rect 18735 3765 18750 3785
rect 18700 3735 18750 3765
rect 18700 3715 18715 3735
rect 18735 3715 18750 3735
rect 18700 3700 18750 3715
rect 18850 4185 18900 4200
rect 18850 4165 18865 4185
rect 18885 4165 18900 4185
rect 18850 4135 18900 4165
rect 18850 4115 18865 4135
rect 18885 4115 18900 4135
rect 18850 4085 18900 4115
rect 18850 4065 18865 4085
rect 18885 4065 18900 4085
rect 18850 4035 18900 4065
rect 18850 4015 18865 4035
rect 18885 4015 18900 4035
rect 18850 3985 18900 4015
rect 18850 3965 18865 3985
rect 18885 3965 18900 3985
rect 18850 3935 18900 3965
rect 18850 3915 18865 3935
rect 18885 3915 18900 3935
rect 18850 3885 18900 3915
rect 18850 3865 18865 3885
rect 18885 3865 18900 3885
rect 18850 3835 18900 3865
rect 18850 3815 18865 3835
rect 18885 3815 18900 3835
rect 18850 3785 18900 3815
rect 18850 3765 18865 3785
rect 18885 3765 18900 3785
rect 18850 3735 18900 3765
rect 18850 3715 18865 3735
rect 18885 3715 18900 3735
rect 18850 3700 18900 3715
rect 19000 4185 19050 4200
rect 19000 4165 19015 4185
rect 19035 4165 19050 4185
rect 19000 4135 19050 4165
rect 19000 4115 19015 4135
rect 19035 4115 19050 4135
rect 19000 4085 19050 4115
rect 19000 4065 19015 4085
rect 19035 4065 19050 4085
rect 19000 4035 19050 4065
rect 19000 4015 19015 4035
rect 19035 4015 19050 4035
rect 19000 3985 19050 4015
rect 19000 3965 19015 3985
rect 19035 3965 19050 3985
rect 19000 3935 19050 3965
rect 19000 3915 19015 3935
rect 19035 3915 19050 3935
rect 19000 3885 19050 3915
rect 19000 3865 19015 3885
rect 19035 3865 19050 3885
rect 19000 3835 19050 3865
rect 19000 3815 19015 3835
rect 19035 3815 19050 3835
rect 19000 3785 19050 3815
rect 19000 3765 19015 3785
rect 19035 3765 19050 3785
rect 19000 3735 19050 3765
rect 19000 3715 19015 3735
rect 19035 3715 19050 3735
rect 19000 3700 19050 3715
rect 19150 4185 19200 4200
rect 19150 4165 19165 4185
rect 19185 4165 19200 4185
rect 19150 4135 19200 4165
rect 19150 4115 19165 4135
rect 19185 4115 19200 4135
rect 19150 4085 19200 4115
rect 19150 4065 19165 4085
rect 19185 4065 19200 4085
rect 19150 4035 19200 4065
rect 19150 4015 19165 4035
rect 19185 4015 19200 4035
rect 19150 3985 19200 4015
rect 19150 3965 19165 3985
rect 19185 3965 19200 3985
rect 19150 3935 19200 3965
rect 19150 3915 19165 3935
rect 19185 3915 19200 3935
rect 19150 3885 19200 3915
rect 19150 3865 19165 3885
rect 19185 3865 19200 3885
rect 19150 3835 19200 3865
rect 19150 3815 19165 3835
rect 19185 3815 19200 3835
rect 19150 3785 19200 3815
rect 19150 3765 19165 3785
rect 19185 3765 19200 3785
rect 19150 3735 19200 3765
rect 19150 3715 19165 3735
rect 19185 3715 19200 3735
rect 19150 3700 19200 3715
rect 19300 4185 19350 4200
rect 19300 4165 19315 4185
rect 19335 4165 19350 4185
rect 19300 4135 19350 4165
rect 19300 4115 19315 4135
rect 19335 4115 19350 4135
rect 19300 4085 19350 4115
rect 19300 4065 19315 4085
rect 19335 4065 19350 4085
rect 19300 4035 19350 4065
rect 19300 4015 19315 4035
rect 19335 4015 19350 4035
rect 19300 3985 19350 4015
rect 19300 3965 19315 3985
rect 19335 3965 19350 3985
rect 19300 3935 19350 3965
rect 19300 3915 19315 3935
rect 19335 3915 19350 3935
rect 19300 3885 19350 3915
rect 19300 3865 19315 3885
rect 19335 3865 19350 3885
rect 19300 3835 19350 3865
rect 19300 3815 19315 3835
rect 19335 3815 19350 3835
rect 19300 3785 19350 3815
rect 19300 3765 19315 3785
rect 19335 3765 19350 3785
rect 19300 3735 19350 3765
rect 19300 3715 19315 3735
rect 19335 3715 19350 3735
rect 19300 3700 19350 3715
rect 19450 4185 19500 4200
rect 19450 4165 19465 4185
rect 19485 4165 19500 4185
rect 19450 4135 19500 4165
rect 19450 4115 19465 4135
rect 19485 4115 19500 4135
rect 19450 4085 19500 4115
rect 19450 4065 19465 4085
rect 19485 4065 19500 4085
rect 19450 4035 19500 4065
rect 19450 4015 19465 4035
rect 19485 4015 19500 4035
rect 19450 3985 19500 4015
rect 19450 3965 19465 3985
rect 19485 3965 19500 3985
rect 19450 3935 19500 3965
rect 19450 3915 19465 3935
rect 19485 3915 19500 3935
rect 19450 3885 19500 3915
rect 19450 3865 19465 3885
rect 19485 3865 19500 3885
rect 19450 3835 19500 3865
rect 19450 3815 19465 3835
rect 19485 3815 19500 3835
rect 19450 3785 19500 3815
rect 19450 3765 19465 3785
rect 19485 3765 19500 3785
rect 19450 3735 19500 3765
rect 19450 3715 19465 3735
rect 19485 3715 19500 3735
rect 19450 3700 19500 3715
rect 19600 4185 19650 4200
rect 19600 4165 19615 4185
rect 19635 4165 19650 4185
rect 19600 4135 19650 4165
rect 19600 4115 19615 4135
rect 19635 4115 19650 4135
rect 19600 4085 19650 4115
rect 19600 4065 19615 4085
rect 19635 4065 19650 4085
rect 19600 4035 19650 4065
rect 19600 4015 19615 4035
rect 19635 4015 19650 4035
rect 19600 3985 19650 4015
rect 19600 3965 19615 3985
rect 19635 3965 19650 3985
rect 19600 3935 19650 3965
rect 19600 3915 19615 3935
rect 19635 3915 19650 3935
rect 19600 3885 19650 3915
rect 19600 3865 19615 3885
rect 19635 3865 19650 3885
rect 19600 3835 19650 3865
rect 19600 3815 19615 3835
rect 19635 3815 19650 3835
rect 19600 3785 19650 3815
rect 19600 3765 19615 3785
rect 19635 3765 19650 3785
rect 19600 3735 19650 3765
rect 19600 3715 19615 3735
rect 19635 3715 19650 3735
rect 19600 3700 19650 3715
rect 19750 4185 19800 4200
rect 19750 4165 19765 4185
rect 19785 4165 19800 4185
rect 19750 4135 19800 4165
rect 19750 4115 19765 4135
rect 19785 4115 19800 4135
rect 19750 4085 19800 4115
rect 19750 4065 19765 4085
rect 19785 4065 19800 4085
rect 19750 4035 19800 4065
rect 19750 4015 19765 4035
rect 19785 4015 19800 4035
rect 19750 3985 19800 4015
rect 19750 3965 19765 3985
rect 19785 3965 19800 3985
rect 19750 3935 19800 3965
rect 19750 3915 19765 3935
rect 19785 3915 19800 3935
rect 19750 3885 19800 3915
rect 19750 3865 19765 3885
rect 19785 3865 19800 3885
rect 19750 3835 19800 3865
rect 19750 3815 19765 3835
rect 19785 3815 19800 3835
rect 19750 3785 19800 3815
rect 19750 3765 19765 3785
rect 19785 3765 19800 3785
rect 19750 3735 19800 3765
rect 19750 3715 19765 3735
rect 19785 3715 19800 3735
rect 19750 3700 19800 3715
rect 19900 3700 19950 4200
rect 20050 3700 20100 4200
rect 20200 3700 20250 4200
rect 20350 4185 20400 4200
rect 20350 4165 20365 4185
rect 20385 4165 20400 4185
rect 20350 4135 20400 4165
rect 20350 4115 20365 4135
rect 20385 4115 20400 4135
rect 20350 4085 20400 4115
rect 20350 4065 20365 4085
rect 20385 4065 20400 4085
rect 20350 4035 20400 4065
rect 20350 4015 20365 4035
rect 20385 4015 20400 4035
rect 20350 3985 20400 4015
rect 20350 3965 20365 3985
rect 20385 3965 20400 3985
rect 20350 3935 20400 3965
rect 20350 3915 20365 3935
rect 20385 3915 20400 3935
rect 20350 3885 20400 3915
rect 20350 3865 20365 3885
rect 20385 3865 20400 3885
rect 20350 3835 20400 3865
rect 20350 3815 20365 3835
rect 20385 3815 20400 3835
rect 20350 3785 20400 3815
rect 20350 3765 20365 3785
rect 20385 3765 20400 3785
rect 20350 3735 20400 3765
rect 20350 3715 20365 3735
rect 20385 3715 20400 3735
rect 20350 3700 20400 3715
rect 20500 3700 20550 4200
rect 20650 3700 20700 4200
rect 20800 3700 20850 4200
rect 20950 4185 21000 4200
rect 20950 4165 20965 4185
rect 20985 4165 21000 4185
rect 20950 4135 21000 4165
rect 20950 4115 20965 4135
rect 20985 4115 21000 4135
rect 20950 4085 21000 4115
rect 20950 4065 20965 4085
rect 20985 4065 21000 4085
rect 20950 4035 21000 4065
rect 20950 4015 20965 4035
rect 20985 4015 21000 4035
rect 20950 3985 21000 4015
rect 20950 3965 20965 3985
rect 20985 3965 21000 3985
rect 20950 3935 21000 3965
rect 20950 3915 20965 3935
rect 20985 3915 21000 3935
rect 20950 3885 21000 3915
rect 20950 3865 20965 3885
rect 20985 3865 21000 3885
rect 20950 3835 21000 3865
rect 20950 3815 20965 3835
rect 20985 3815 21000 3835
rect 20950 3785 21000 3815
rect 20950 3765 20965 3785
rect 20985 3765 21000 3785
rect 20950 3735 21000 3765
rect 20950 3715 20965 3735
rect 20985 3715 21000 3735
rect 20950 3700 21000 3715
rect 21100 3700 21150 4200
rect 21250 3700 21300 4200
rect 21400 4185 21450 4200
rect 21400 4165 21415 4185
rect 21435 4165 21450 4185
rect 21400 4135 21450 4165
rect 21400 4115 21415 4135
rect 21435 4115 21450 4135
rect 21400 4085 21450 4115
rect 21400 4065 21415 4085
rect 21435 4065 21450 4085
rect 21400 4035 21450 4065
rect 21400 4015 21415 4035
rect 21435 4015 21450 4035
rect 21400 3985 21450 4015
rect 21400 3965 21415 3985
rect 21435 3965 21450 3985
rect 21400 3935 21450 3965
rect 21400 3915 21415 3935
rect 21435 3915 21450 3935
rect 21400 3885 21450 3915
rect 21400 3865 21415 3885
rect 21435 3865 21450 3885
rect 21400 3835 21450 3865
rect 21400 3815 21415 3835
rect 21435 3815 21450 3835
rect 21400 3785 21450 3815
rect 21400 3765 21415 3785
rect 21435 3765 21450 3785
rect 21400 3735 21450 3765
rect 21400 3715 21415 3735
rect 21435 3715 21450 3735
rect 21400 3700 21450 3715
rect 21550 3700 21600 4200
rect 21700 3700 21750 4200
rect 21850 4185 21900 4200
rect 21850 4165 21865 4185
rect 21885 4165 21900 4185
rect 21850 4135 21900 4165
rect 21850 4115 21865 4135
rect 21885 4115 21900 4135
rect 21850 4085 21900 4115
rect 21850 4065 21865 4085
rect 21885 4065 21900 4085
rect 21850 4035 21900 4065
rect 21850 4015 21865 4035
rect 21885 4015 21900 4035
rect 21850 3985 21900 4015
rect 21850 3965 21865 3985
rect 21885 3965 21900 3985
rect 21850 3935 21900 3965
rect 21850 3915 21865 3935
rect 21885 3915 21900 3935
rect 21850 3885 21900 3915
rect 21850 3865 21865 3885
rect 21885 3865 21900 3885
rect 21850 3835 21900 3865
rect 21850 3815 21865 3835
rect 21885 3815 21900 3835
rect 21850 3785 21900 3815
rect 21850 3765 21865 3785
rect 21885 3765 21900 3785
rect 21850 3735 21900 3765
rect 21850 3715 21865 3735
rect 21885 3715 21900 3735
rect 21850 3700 21900 3715
rect 22000 3700 22050 4200
rect 22150 3700 22200 4200
rect 22300 3700 22350 4200
rect 22450 4185 22500 4200
rect 22450 4165 22465 4185
rect 22485 4165 22500 4185
rect 22450 4135 22500 4165
rect 22450 4115 22465 4135
rect 22485 4115 22500 4135
rect 22450 4085 22500 4115
rect 22450 4065 22465 4085
rect 22485 4065 22500 4085
rect 22450 4035 22500 4065
rect 22450 4015 22465 4035
rect 22485 4015 22500 4035
rect 22450 3985 22500 4015
rect 22450 3965 22465 3985
rect 22485 3965 22500 3985
rect 22450 3935 22500 3965
rect 22450 3915 22465 3935
rect 22485 3915 22500 3935
rect 22450 3885 22500 3915
rect 22450 3865 22465 3885
rect 22485 3865 22500 3885
rect 22450 3835 22500 3865
rect 22450 3815 22465 3835
rect 22485 3815 22500 3835
rect 22450 3785 22500 3815
rect 22450 3765 22465 3785
rect 22485 3765 22500 3785
rect 22450 3735 22500 3765
rect 22450 3715 22465 3735
rect 22485 3715 22500 3735
rect 22450 3700 22500 3715
rect 22600 3700 22650 4200
rect 22750 3700 22800 4200
rect 22900 3700 22950 4200
rect 23050 4185 23100 4200
rect 23050 4165 23065 4185
rect 23085 4165 23100 4185
rect 23050 4135 23100 4165
rect 23050 4115 23065 4135
rect 23085 4115 23100 4135
rect 23050 4085 23100 4115
rect 23050 4065 23065 4085
rect 23085 4065 23100 4085
rect 23050 4035 23100 4065
rect 23050 4015 23065 4035
rect 23085 4015 23100 4035
rect 23050 3985 23100 4015
rect 23050 3965 23065 3985
rect 23085 3965 23100 3985
rect 23050 3935 23100 3965
rect 23050 3915 23065 3935
rect 23085 3915 23100 3935
rect 23050 3885 23100 3915
rect 23050 3865 23065 3885
rect 23085 3865 23100 3885
rect 23050 3835 23100 3865
rect 23050 3815 23065 3835
rect 23085 3815 23100 3835
rect 23050 3785 23100 3815
rect 23050 3765 23065 3785
rect 23085 3765 23100 3785
rect 23050 3735 23100 3765
rect 23050 3715 23065 3735
rect 23085 3715 23100 3735
rect 23050 3700 23100 3715
rect 23200 3700 23250 4200
rect 23350 3700 23400 4200
rect 23500 4185 23550 4200
rect 23500 4165 23515 4185
rect 23535 4165 23550 4185
rect 23500 4135 23550 4165
rect 23500 4115 23515 4135
rect 23535 4115 23550 4135
rect 23500 4085 23550 4115
rect 23500 4065 23515 4085
rect 23535 4065 23550 4085
rect 23500 4035 23550 4065
rect 23500 4015 23515 4035
rect 23535 4015 23550 4035
rect 23500 3985 23550 4015
rect 23500 3965 23515 3985
rect 23535 3965 23550 3985
rect 23500 3935 23550 3965
rect 23500 3915 23515 3935
rect 23535 3915 23550 3935
rect 23500 3885 23550 3915
rect 23500 3865 23515 3885
rect 23535 3865 23550 3885
rect 23500 3835 23550 3865
rect 23500 3815 23515 3835
rect 23535 3815 23550 3835
rect 23500 3785 23550 3815
rect 23500 3765 23515 3785
rect 23535 3765 23550 3785
rect 23500 3735 23550 3765
rect 23500 3715 23515 3735
rect 23535 3715 23550 3735
rect 23500 3700 23550 3715
rect 23650 3700 23700 4200
rect 23800 3700 23850 4200
rect 23950 4185 24000 4200
rect 23950 4165 23965 4185
rect 23985 4165 24000 4185
rect 23950 4135 24000 4165
rect 23950 4115 23965 4135
rect 23985 4115 24000 4135
rect 23950 4085 24000 4115
rect 23950 4065 23965 4085
rect 23985 4065 24000 4085
rect 23950 4035 24000 4065
rect 23950 4015 23965 4035
rect 23985 4015 24000 4035
rect 23950 3985 24000 4015
rect 23950 3965 23965 3985
rect 23985 3965 24000 3985
rect 23950 3935 24000 3965
rect 23950 3915 23965 3935
rect 23985 3915 24000 3935
rect 23950 3885 24000 3915
rect 23950 3865 23965 3885
rect 23985 3865 24000 3885
rect 23950 3835 24000 3865
rect 23950 3815 23965 3835
rect 23985 3815 24000 3835
rect 23950 3785 24000 3815
rect 23950 3765 23965 3785
rect 23985 3765 24000 3785
rect 23950 3735 24000 3765
rect 23950 3715 23965 3735
rect 23985 3715 24000 3735
rect 23950 3700 24000 3715
rect 24100 3700 24150 4200
rect 24250 3700 24300 4200
rect 24400 3700 24450 4200
rect 24550 4185 24600 4200
rect 24550 4165 24565 4185
rect 24585 4165 24600 4185
rect 24550 4135 24600 4165
rect 24550 4115 24565 4135
rect 24585 4115 24600 4135
rect 24550 4085 24600 4115
rect 24550 4065 24565 4085
rect 24585 4065 24600 4085
rect 24550 4035 24600 4065
rect 24550 4015 24565 4035
rect 24585 4015 24600 4035
rect 24550 3985 24600 4015
rect 24550 3965 24565 3985
rect 24585 3965 24600 3985
rect 24550 3935 24600 3965
rect 24550 3915 24565 3935
rect 24585 3915 24600 3935
rect 24550 3885 24600 3915
rect 24550 3865 24565 3885
rect 24585 3865 24600 3885
rect 24550 3835 24600 3865
rect 24550 3815 24565 3835
rect 24585 3815 24600 3835
rect 24550 3785 24600 3815
rect 24550 3765 24565 3785
rect 24585 3765 24600 3785
rect 24550 3735 24600 3765
rect 24550 3715 24565 3735
rect 24585 3715 24600 3735
rect 24550 3700 24600 3715
rect 24700 3700 24750 4200
rect 24850 3700 24900 4200
rect 25000 3700 25050 4200
rect 25150 4185 25200 4200
rect 25150 4165 25165 4185
rect 25185 4165 25200 4185
rect 25150 4135 25200 4165
rect 25150 4115 25165 4135
rect 25185 4115 25200 4135
rect 25150 4085 25200 4115
rect 25150 4065 25165 4085
rect 25185 4065 25200 4085
rect 25150 4035 25200 4065
rect 25150 4015 25165 4035
rect 25185 4015 25200 4035
rect 25150 3985 25200 4015
rect 25150 3965 25165 3985
rect 25185 3965 25200 3985
rect 25150 3935 25200 3965
rect 25150 3915 25165 3935
rect 25185 3915 25200 3935
rect 25150 3885 25200 3915
rect 25150 3865 25165 3885
rect 25185 3865 25200 3885
rect 25150 3835 25200 3865
rect 25150 3815 25165 3835
rect 25185 3815 25200 3835
rect 25150 3785 25200 3815
rect 25150 3765 25165 3785
rect 25185 3765 25200 3785
rect 25150 3735 25200 3765
rect 25150 3715 25165 3735
rect 25185 3715 25200 3735
rect 25150 3700 25200 3715
rect 25300 3700 25350 4200
rect 25450 3700 25500 4200
rect 25600 4185 25650 4200
rect 25600 4165 25615 4185
rect 25635 4165 25650 4185
rect 25600 4135 25650 4165
rect 25600 4115 25615 4135
rect 25635 4115 25650 4135
rect 25600 4085 25650 4115
rect 25600 4065 25615 4085
rect 25635 4065 25650 4085
rect 25600 4035 25650 4065
rect 25600 4015 25615 4035
rect 25635 4015 25650 4035
rect 25600 3985 25650 4015
rect 25600 3965 25615 3985
rect 25635 3965 25650 3985
rect 25600 3935 25650 3965
rect 25600 3915 25615 3935
rect 25635 3915 25650 3935
rect 25600 3885 25650 3915
rect 25600 3865 25615 3885
rect 25635 3865 25650 3885
rect 25600 3835 25650 3865
rect 25600 3815 25615 3835
rect 25635 3815 25650 3835
rect 25600 3785 25650 3815
rect 25600 3765 25615 3785
rect 25635 3765 25650 3785
rect 25600 3735 25650 3765
rect 25600 3715 25615 3735
rect 25635 3715 25650 3735
rect 25600 3700 25650 3715
rect 25750 3700 25800 4200
rect 25900 3700 25950 4200
rect 26050 4185 26100 4200
rect 26050 4165 26065 4185
rect 26085 4165 26100 4185
rect 26050 4135 26100 4165
rect 26050 4115 26065 4135
rect 26085 4115 26100 4135
rect 26050 4085 26100 4115
rect 26050 4065 26065 4085
rect 26085 4065 26100 4085
rect 26050 4035 26100 4065
rect 26050 4015 26065 4035
rect 26085 4015 26100 4035
rect 26050 3985 26100 4015
rect 26050 3965 26065 3985
rect 26085 3965 26100 3985
rect 26050 3935 26100 3965
rect 26050 3915 26065 3935
rect 26085 3915 26100 3935
rect 26050 3885 26100 3915
rect 26050 3865 26065 3885
rect 26085 3865 26100 3885
rect 26050 3835 26100 3865
rect 26050 3815 26065 3835
rect 26085 3815 26100 3835
rect 26050 3785 26100 3815
rect 26050 3765 26065 3785
rect 26085 3765 26100 3785
rect 26050 3735 26100 3765
rect 26050 3715 26065 3735
rect 26085 3715 26100 3735
rect 26050 3700 26100 3715
rect 26200 3700 26250 4200
rect 26350 3700 26400 4200
rect 26500 3700 26550 4200
rect 26650 4185 26700 4200
rect 26650 4165 26665 4185
rect 26685 4165 26700 4185
rect 26650 4135 26700 4165
rect 26650 4115 26665 4135
rect 26685 4115 26700 4135
rect 26650 4085 26700 4115
rect 26650 4065 26665 4085
rect 26685 4065 26700 4085
rect 26650 4035 26700 4065
rect 26650 4015 26665 4035
rect 26685 4015 26700 4035
rect 26650 3985 26700 4015
rect 26650 3965 26665 3985
rect 26685 3965 26700 3985
rect 26650 3935 26700 3965
rect 26650 3915 26665 3935
rect 26685 3915 26700 3935
rect 26650 3885 26700 3915
rect 26650 3865 26665 3885
rect 26685 3865 26700 3885
rect 26650 3835 26700 3865
rect 26650 3815 26665 3835
rect 26685 3815 26700 3835
rect 26650 3785 26700 3815
rect 26650 3765 26665 3785
rect 26685 3765 26700 3785
rect 26650 3735 26700 3765
rect 26650 3715 26665 3735
rect 26685 3715 26700 3735
rect 26650 3700 26700 3715
rect 26800 3700 26850 4200
rect 26950 3700 27000 4200
rect 27100 3700 27150 4200
rect 27250 4185 27300 4200
rect 27250 4165 27265 4185
rect 27285 4165 27300 4185
rect 27250 4135 27300 4165
rect 27250 4115 27265 4135
rect 27285 4115 27300 4135
rect 27250 4085 27300 4115
rect 27250 4065 27265 4085
rect 27285 4065 27300 4085
rect 27250 4035 27300 4065
rect 27250 4015 27265 4035
rect 27285 4015 27300 4035
rect 27250 3985 27300 4015
rect 27250 3965 27265 3985
rect 27285 3965 27300 3985
rect 27250 3935 27300 3965
rect 27250 3915 27265 3935
rect 27285 3915 27300 3935
rect 27250 3885 27300 3915
rect 27250 3865 27265 3885
rect 27285 3865 27300 3885
rect 27250 3835 27300 3865
rect 27250 3815 27265 3835
rect 27285 3815 27300 3835
rect 27250 3785 27300 3815
rect 27250 3765 27265 3785
rect 27285 3765 27300 3785
rect 27250 3735 27300 3765
rect 27250 3715 27265 3735
rect 27285 3715 27300 3735
rect 27250 3700 27300 3715
rect 27400 3700 27450 4200
rect 27550 3700 27600 4200
rect 27700 4185 27750 4200
rect 27700 4165 27715 4185
rect 27735 4165 27750 4185
rect 27700 4135 27750 4165
rect 27700 4115 27715 4135
rect 27735 4115 27750 4135
rect 27700 4085 27750 4115
rect 27700 4065 27715 4085
rect 27735 4065 27750 4085
rect 27700 4035 27750 4065
rect 27700 4015 27715 4035
rect 27735 4015 27750 4035
rect 27700 3985 27750 4015
rect 27700 3965 27715 3985
rect 27735 3965 27750 3985
rect 27700 3935 27750 3965
rect 27700 3915 27715 3935
rect 27735 3915 27750 3935
rect 27700 3885 27750 3915
rect 27700 3865 27715 3885
rect 27735 3865 27750 3885
rect 27700 3835 27750 3865
rect 27700 3815 27715 3835
rect 27735 3815 27750 3835
rect 27700 3785 27750 3815
rect 27700 3765 27715 3785
rect 27735 3765 27750 3785
rect 27700 3735 27750 3765
rect 27700 3715 27715 3735
rect 27735 3715 27750 3735
rect 27700 3700 27750 3715
rect 27850 3700 27900 4200
rect 28000 3700 28050 4200
rect 28150 4185 28200 4200
rect 28150 4165 28165 4185
rect 28185 4165 28200 4185
rect 28150 4135 28200 4165
rect 28150 4115 28165 4135
rect 28185 4115 28200 4135
rect 28150 4085 28200 4115
rect 28150 4065 28165 4085
rect 28185 4065 28200 4085
rect 28150 4035 28200 4065
rect 28150 4015 28165 4035
rect 28185 4015 28200 4035
rect 28150 3985 28200 4015
rect 28150 3965 28165 3985
rect 28185 3965 28200 3985
rect 28150 3935 28200 3965
rect 28150 3915 28165 3935
rect 28185 3915 28200 3935
rect 28150 3885 28200 3915
rect 28150 3865 28165 3885
rect 28185 3865 28200 3885
rect 28150 3835 28200 3865
rect 28150 3815 28165 3835
rect 28185 3815 28200 3835
rect 28150 3785 28200 3815
rect 28150 3765 28165 3785
rect 28185 3765 28200 3785
rect 28150 3735 28200 3765
rect 28150 3715 28165 3735
rect 28185 3715 28200 3735
rect 28150 3700 28200 3715
rect 28300 3700 28350 4200
rect 28450 3700 28500 4200
rect 28600 3700 28650 4200
rect 28750 4185 28800 4200
rect 28750 4165 28765 4185
rect 28785 4165 28800 4185
rect 28750 4135 28800 4165
rect 28750 4115 28765 4135
rect 28785 4115 28800 4135
rect 28750 4085 28800 4115
rect 28750 4065 28765 4085
rect 28785 4065 28800 4085
rect 28750 4035 28800 4065
rect 28750 4015 28765 4035
rect 28785 4015 28800 4035
rect 28750 3985 28800 4015
rect 28750 3965 28765 3985
rect 28785 3965 28800 3985
rect 28750 3935 28800 3965
rect 28750 3915 28765 3935
rect 28785 3915 28800 3935
rect 28750 3885 28800 3915
rect 28750 3865 28765 3885
rect 28785 3865 28800 3885
rect 28750 3835 28800 3865
rect 28750 3815 28765 3835
rect 28785 3815 28800 3835
rect 28750 3785 28800 3815
rect 28750 3765 28765 3785
rect 28785 3765 28800 3785
rect 28750 3735 28800 3765
rect 28750 3715 28765 3735
rect 28785 3715 28800 3735
rect 28750 3700 28800 3715
rect 28900 3700 28950 4200
rect 29050 3700 29100 4200
rect 29200 3700 29250 4200
rect 29350 4185 29400 4200
rect 29350 4165 29365 4185
rect 29385 4165 29400 4185
rect 29350 4135 29400 4165
rect 29350 4115 29365 4135
rect 29385 4115 29400 4135
rect 29350 4085 29400 4115
rect 29350 4065 29365 4085
rect 29385 4065 29400 4085
rect 29350 4035 29400 4065
rect 29350 4015 29365 4035
rect 29385 4015 29400 4035
rect 29350 3985 29400 4015
rect 29350 3965 29365 3985
rect 29385 3965 29400 3985
rect 29350 3935 29400 3965
rect 29350 3915 29365 3935
rect 29385 3915 29400 3935
rect 29350 3885 29400 3915
rect 29350 3865 29365 3885
rect 29385 3865 29400 3885
rect 29350 3835 29400 3865
rect 29350 3815 29365 3835
rect 29385 3815 29400 3835
rect 29350 3785 29400 3815
rect 29350 3765 29365 3785
rect 29385 3765 29400 3785
rect 29350 3735 29400 3765
rect 29350 3715 29365 3735
rect 29385 3715 29400 3735
rect 29350 3700 29400 3715
rect 29500 4185 29550 4200
rect 29500 4165 29515 4185
rect 29535 4165 29550 4185
rect 29500 4135 29550 4165
rect 29500 4115 29515 4135
rect 29535 4115 29550 4135
rect 29500 4085 29550 4115
rect 29500 4065 29515 4085
rect 29535 4065 29550 4085
rect 29500 4035 29550 4065
rect 29500 4015 29515 4035
rect 29535 4015 29550 4035
rect 29500 3985 29550 4015
rect 29500 3965 29515 3985
rect 29535 3965 29550 3985
rect 29500 3935 29550 3965
rect 29500 3915 29515 3935
rect 29535 3915 29550 3935
rect 29500 3885 29550 3915
rect 29500 3865 29515 3885
rect 29535 3865 29550 3885
rect 29500 3835 29550 3865
rect 29500 3815 29515 3835
rect 29535 3815 29550 3835
rect 29500 3785 29550 3815
rect 29500 3765 29515 3785
rect 29535 3765 29550 3785
rect 29500 3735 29550 3765
rect 29500 3715 29515 3735
rect 29535 3715 29550 3735
rect 29500 3700 29550 3715
rect 29650 4185 29700 4200
rect 29650 4165 29665 4185
rect 29685 4165 29700 4185
rect 29650 4135 29700 4165
rect 29650 4115 29665 4135
rect 29685 4115 29700 4135
rect 29650 4085 29700 4115
rect 29650 4065 29665 4085
rect 29685 4065 29700 4085
rect 29650 4035 29700 4065
rect 29650 4015 29665 4035
rect 29685 4015 29700 4035
rect 29650 3985 29700 4015
rect 29650 3965 29665 3985
rect 29685 3965 29700 3985
rect 29650 3935 29700 3965
rect 29650 3915 29665 3935
rect 29685 3915 29700 3935
rect 29650 3885 29700 3915
rect 29650 3865 29665 3885
rect 29685 3865 29700 3885
rect 29650 3835 29700 3865
rect 29650 3815 29665 3835
rect 29685 3815 29700 3835
rect 29650 3785 29700 3815
rect 29650 3765 29665 3785
rect 29685 3765 29700 3785
rect 29650 3735 29700 3765
rect 29650 3715 29665 3735
rect 29685 3715 29700 3735
rect 29650 3700 29700 3715
rect 29800 4185 29850 4200
rect 29800 4165 29815 4185
rect 29835 4165 29850 4185
rect 29800 4135 29850 4165
rect 29800 4115 29815 4135
rect 29835 4115 29850 4135
rect 29800 4085 29850 4115
rect 29800 4065 29815 4085
rect 29835 4065 29850 4085
rect 29800 4035 29850 4065
rect 29800 4015 29815 4035
rect 29835 4015 29850 4035
rect 29800 3985 29850 4015
rect 29800 3965 29815 3985
rect 29835 3965 29850 3985
rect 29800 3935 29850 3965
rect 29800 3915 29815 3935
rect 29835 3915 29850 3935
rect 29800 3885 29850 3915
rect 29800 3865 29815 3885
rect 29835 3865 29850 3885
rect 29800 3835 29850 3865
rect 29800 3815 29815 3835
rect 29835 3815 29850 3835
rect 29800 3785 29850 3815
rect 29800 3765 29815 3785
rect 29835 3765 29850 3785
rect 29800 3735 29850 3765
rect 29800 3715 29815 3735
rect 29835 3715 29850 3735
rect 29800 3700 29850 3715
rect 29950 4185 30000 4200
rect 29950 4165 29965 4185
rect 29985 4165 30000 4185
rect 29950 4135 30000 4165
rect 29950 4115 29965 4135
rect 29985 4115 30000 4135
rect 29950 4085 30000 4115
rect 29950 4065 29965 4085
rect 29985 4065 30000 4085
rect 29950 4035 30000 4065
rect 29950 4015 29965 4035
rect 29985 4015 30000 4035
rect 29950 3985 30000 4015
rect 29950 3965 29965 3985
rect 29985 3965 30000 3985
rect 29950 3935 30000 3965
rect 29950 3915 29965 3935
rect 29985 3915 30000 3935
rect 29950 3885 30000 3915
rect 29950 3865 29965 3885
rect 29985 3865 30000 3885
rect 29950 3835 30000 3865
rect 29950 3815 29965 3835
rect 29985 3815 30000 3835
rect 29950 3785 30000 3815
rect 29950 3765 29965 3785
rect 29985 3765 30000 3785
rect 29950 3735 30000 3765
rect 29950 3715 29965 3735
rect 29985 3715 30000 3735
rect 29950 3700 30000 3715
rect 30100 4185 30150 4200
rect 30100 4165 30115 4185
rect 30135 4165 30150 4185
rect 30100 4135 30150 4165
rect 30100 4115 30115 4135
rect 30135 4115 30150 4135
rect 30100 4085 30150 4115
rect 30100 4065 30115 4085
rect 30135 4065 30150 4085
rect 30100 4035 30150 4065
rect 30100 4015 30115 4035
rect 30135 4015 30150 4035
rect 30100 3985 30150 4015
rect 30100 3965 30115 3985
rect 30135 3965 30150 3985
rect 30100 3935 30150 3965
rect 30100 3915 30115 3935
rect 30135 3915 30150 3935
rect 30100 3885 30150 3915
rect 30100 3865 30115 3885
rect 30135 3865 30150 3885
rect 30100 3835 30150 3865
rect 30100 3815 30115 3835
rect 30135 3815 30150 3835
rect 30100 3785 30150 3815
rect 30100 3765 30115 3785
rect 30135 3765 30150 3785
rect 30100 3735 30150 3765
rect 30100 3715 30115 3735
rect 30135 3715 30150 3735
rect 30100 3700 30150 3715
rect 30250 4185 30300 4200
rect 30250 4165 30265 4185
rect 30285 4165 30300 4185
rect 30250 4135 30300 4165
rect 30250 4115 30265 4135
rect 30285 4115 30300 4135
rect 30250 4085 30300 4115
rect 30250 4065 30265 4085
rect 30285 4065 30300 4085
rect 30250 4035 30300 4065
rect 30250 4015 30265 4035
rect 30285 4015 30300 4035
rect 30250 3985 30300 4015
rect 30250 3965 30265 3985
rect 30285 3965 30300 3985
rect 30250 3935 30300 3965
rect 30250 3915 30265 3935
rect 30285 3915 30300 3935
rect 30250 3885 30300 3915
rect 30250 3865 30265 3885
rect 30285 3865 30300 3885
rect 30250 3835 30300 3865
rect 30250 3815 30265 3835
rect 30285 3815 30300 3835
rect 30250 3785 30300 3815
rect 30250 3765 30265 3785
rect 30285 3765 30300 3785
rect 30250 3735 30300 3765
rect 30250 3715 30265 3735
rect 30285 3715 30300 3735
rect 30250 3700 30300 3715
rect 30400 4185 30450 4200
rect 30400 4165 30415 4185
rect 30435 4165 30450 4185
rect 30400 4135 30450 4165
rect 30400 4115 30415 4135
rect 30435 4115 30450 4135
rect 30400 4085 30450 4115
rect 30400 4065 30415 4085
rect 30435 4065 30450 4085
rect 30400 4035 30450 4065
rect 30400 4015 30415 4035
rect 30435 4015 30450 4035
rect 30400 3985 30450 4015
rect 30400 3965 30415 3985
rect 30435 3965 30450 3985
rect 30400 3935 30450 3965
rect 30400 3915 30415 3935
rect 30435 3915 30450 3935
rect 30400 3885 30450 3915
rect 30400 3865 30415 3885
rect 30435 3865 30450 3885
rect 30400 3835 30450 3865
rect 30400 3815 30415 3835
rect 30435 3815 30450 3835
rect 30400 3785 30450 3815
rect 30400 3765 30415 3785
rect 30435 3765 30450 3785
rect 30400 3735 30450 3765
rect 30400 3715 30415 3735
rect 30435 3715 30450 3735
rect 30400 3700 30450 3715
rect 30550 4185 30600 4200
rect 30550 4165 30565 4185
rect 30585 4165 30600 4185
rect 30550 4135 30600 4165
rect 30550 4115 30565 4135
rect 30585 4115 30600 4135
rect 30550 4085 30600 4115
rect 30550 4065 30565 4085
rect 30585 4065 30600 4085
rect 30550 4035 30600 4065
rect 30550 4015 30565 4035
rect 30585 4015 30600 4035
rect 30550 3985 30600 4015
rect 30550 3965 30565 3985
rect 30585 3965 30600 3985
rect 30550 3935 30600 3965
rect 30550 3915 30565 3935
rect 30585 3915 30600 3935
rect 30550 3885 30600 3915
rect 30550 3865 30565 3885
rect 30585 3865 30600 3885
rect 30550 3835 30600 3865
rect 30550 3815 30565 3835
rect 30585 3815 30600 3835
rect 30550 3785 30600 3815
rect 30550 3765 30565 3785
rect 30585 3765 30600 3785
rect 30550 3735 30600 3765
rect 30550 3715 30565 3735
rect 30585 3715 30600 3735
rect 30550 3700 30600 3715
rect 30700 4185 30750 4200
rect 30700 4165 30715 4185
rect 30735 4165 30750 4185
rect 30700 4135 30750 4165
rect 30700 4115 30715 4135
rect 30735 4115 30750 4135
rect 30700 4085 30750 4115
rect 30700 4065 30715 4085
rect 30735 4065 30750 4085
rect 30700 4035 30750 4065
rect 30700 4015 30715 4035
rect 30735 4015 30750 4035
rect 30700 3985 30750 4015
rect 30700 3965 30715 3985
rect 30735 3965 30750 3985
rect 30700 3935 30750 3965
rect 30700 3915 30715 3935
rect 30735 3915 30750 3935
rect 30700 3885 30750 3915
rect 30700 3865 30715 3885
rect 30735 3865 30750 3885
rect 30700 3835 30750 3865
rect 30700 3815 30715 3835
rect 30735 3815 30750 3835
rect 30700 3785 30750 3815
rect 30700 3765 30715 3785
rect 30735 3765 30750 3785
rect 30700 3735 30750 3765
rect 30700 3715 30715 3735
rect 30735 3715 30750 3735
rect 30700 3700 30750 3715
rect 30850 4185 30900 4200
rect 30850 4165 30865 4185
rect 30885 4165 30900 4185
rect 30850 4135 30900 4165
rect 30850 4115 30865 4135
rect 30885 4115 30900 4135
rect 30850 4085 30900 4115
rect 30850 4065 30865 4085
rect 30885 4065 30900 4085
rect 30850 4035 30900 4065
rect 30850 4015 30865 4035
rect 30885 4015 30900 4035
rect 30850 3985 30900 4015
rect 30850 3965 30865 3985
rect 30885 3965 30900 3985
rect 30850 3935 30900 3965
rect 30850 3915 30865 3935
rect 30885 3915 30900 3935
rect 30850 3885 30900 3915
rect 30850 3865 30865 3885
rect 30885 3865 30900 3885
rect 30850 3835 30900 3865
rect 30850 3815 30865 3835
rect 30885 3815 30900 3835
rect 30850 3785 30900 3815
rect 30850 3765 30865 3785
rect 30885 3765 30900 3785
rect 30850 3735 30900 3765
rect 30850 3715 30865 3735
rect 30885 3715 30900 3735
rect 30850 3700 30900 3715
rect 31000 4185 31050 4200
rect 31000 4165 31015 4185
rect 31035 4165 31050 4185
rect 31000 4135 31050 4165
rect 31000 4115 31015 4135
rect 31035 4115 31050 4135
rect 31000 4085 31050 4115
rect 31000 4065 31015 4085
rect 31035 4065 31050 4085
rect 31000 4035 31050 4065
rect 31000 4015 31015 4035
rect 31035 4015 31050 4035
rect 31000 3985 31050 4015
rect 31000 3965 31015 3985
rect 31035 3965 31050 3985
rect 31000 3935 31050 3965
rect 31000 3915 31015 3935
rect 31035 3915 31050 3935
rect 31000 3885 31050 3915
rect 31000 3865 31015 3885
rect 31035 3865 31050 3885
rect 31000 3835 31050 3865
rect 31000 3815 31015 3835
rect 31035 3815 31050 3835
rect 31000 3785 31050 3815
rect 31000 3765 31015 3785
rect 31035 3765 31050 3785
rect 31000 3735 31050 3765
rect 31000 3715 31015 3735
rect 31035 3715 31050 3735
rect 31000 3700 31050 3715
rect 31150 4185 31200 4200
rect 31150 4165 31165 4185
rect 31185 4165 31200 4185
rect 31150 4135 31200 4165
rect 31150 4115 31165 4135
rect 31185 4115 31200 4135
rect 31150 4085 31200 4115
rect 31150 4065 31165 4085
rect 31185 4065 31200 4085
rect 31150 4035 31200 4065
rect 31150 4015 31165 4035
rect 31185 4015 31200 4035
rect 31150 3985 31200 4015
rect 31150 3965 31165 3985
rect 31185 3965 31200 3985
rect 31150 3935 31200 3965
rect 31150 3915 31165 3935
rect 31185 3915 31200 3935
rect 31150 3885 31200 3915
rect 31150 3865 31165 3885
rect 31185 3865 31200 3885
rect 31150 3835 31200 3865
rect 31150 3815 31165 3835
rect 31185 3815 31200 3835
rect 31150 3785 31200 3815
rect 31150 3765 31165 3785
rect 31185 3765 31200 3785
rect 31150 3735 31200 3765
rect 31150 3715 31165 3735
rect 31185 3715 31200 3735
rect 31150 3700 31200 3715
rect 31300 4185 31350 4200
rect 31300 4165 31315 4185
rect 31335 4165 31350 4185
rect 31300 4135 31350 4165
rect 31300 4115 31315 4135
rect 31335 4115 31350 4135
rect 31300 4085 31350 4115
rect 31300 4065 31315 4085
rect 31335 4065 31350 4085
rect 31300 4035 31350 4065
rect 31300 4015 31315 4035
rect 31335 4015 31350 4035
rect 31300 3985 31350 4015
rect 31300 3965 31315 3985
rect 31335 3965 31350 3985
rect 31300 3935 31350 3965
rect 31300 3915 31315 3935
rect 31335 3915 31350 3935
rect 31300 3885 31350 3915
rect 31300 3865 31315 3885
rect 31335 3865 31350 3885
rect 31300 3835 31350 3865
rect 31300 3815 31315 3835
rect 31335 3815 31350 3835
rect 31300 3785 31350 3815
rect 31300 3765 31315 3785
rect 31335 3765 31350 3785
rect 31300 3735 31350 3765
rect 31300 3715 31315 3735
rect 31335 3715 31350 3735
rect 31300 3700 31350 3715
rect 31450 4185 31500 4200
rect 31450 4165 31465 4185
rect 31485 4165 31500 4185
rect 31450 4135 31500 4165
rect 31450 4115 31465 4135
rect 31485 4115 31500 4135
rect 31450 4085 31500 4115
rect 31450 4065 31465 4085
rect 31485 4065 31500 4085
rect 31450 4035 31500 4065
rect 31450 4015 31465 4035
rect 31485 4015 31500 4035
rect 31450 3985 31500 4015
rect 31450 3965 31465 3985
rect 31485 3965 31500 3985
rect 31450 3935 31500 3965
rect 31450 3915 31465 3935
rect 31485 3915 31500 3935
rect 31450 3885 31500 3915
rect 31450 3865 31465 3885
rect 31485 3865 31500 3885
rect 31450 3835 31500 3865
rect 31450 3815 31465 3835
rect 31485 3815 31500 3835
rect 31450 3785 31500 3815
rect 31450 3765 31465 3785
rect 31485 3765 31500 3785
rect 31450 3735 31500 3765
rect 31450 3715 31465 3735
rect 31485 3715 31500 3735
rect 31450 3700 31500 3715
rect 31600 3700 31650 4200
rect 31750 3700 31800 4200
rect 31900 3700 31950 4200
rect 32050 4185 32100 4200
rect 32050 4165 32065 4185
rect 32085 4165 32100 4185
rect 32050 4135 32100 4165
rect 32050 4115 32065 4135
rect 32085 4115 32100 4135
rect 32050 4085 32100 4115
rect 32050 4065 32065 4085
rect 32085 4065 32100 4085
rect 32050 4035 32100 4065
rect 32050 4015 32065 4035
rect 32085 4015 32100 4035
rect 32050 3985 32100 4015
rect 32050 3965 32065 3985
rect 32085 3965 32100 3985
rect 32050 3935 32100 3965
rect 32050 3915 32065 3935
rect 32085 3915 32100 3935
rect 32050 3885 32100 3915
rect 32050 3865 32065 3885
rect 32085 3865 32100 3885
rect 32050 3835 32100 3865
rect 32050 3815 32065 3835
rect 32085 3815 32100 3835
rect 32050 3785 32100 3815
rect 32050 3765 32065 3785
rect 32085 3765 32100 3785
rect 32050 3735 32100 3765
rect 32050 3715 32065 3735
rect 32085 3715 32100 3735
rect 32050 3700 32100 3715
rect -650 3535 -600 3550
rect -650 3515 -635 3535
rect -615 3515 -600 3535
rect -650 3485 -600 3515
rect -650 3465 -635 3485
rect -615 3465 -600 3485
rect -650 3435 -600 3465
rect -650 3415 -635 3435
rect -615 3415 -600 3435
rect -650 3385 -600 3415
rect -650 3365 -635 3385
rect -615 3365 -600 3385
rect -650 3335 -600 3365
rect -650 3315 -635 3335
rect -615 3315 -600 3335
rect -650 3285 -600 3315
rect -650 3265 -635 3285
rect -615 3265 -600 3285
rect -650 3235 -600 3265
rect -650 3215 -635 3235
rect -615 3215 -600 3235
rect -650 3185 -600 3215
rect -650 3165 -635 3185
rect -615 3165 -600 3185
rect -650 3135 -600 3165
rect -650 3115 -635 3135
rect -615 3115 -600 3135
rect -650 3085 -600 3115
rect -650 3065 -635 3085
rect -615 3065 -600 3085
rect -650 3050 -600 3065
rect -500 3535 -450 3550
rect -500 3515 -485 3535
rect -465 3515 -450 3535
rect -500 3485 -450 3515
rect -500 3465 -485 3485
rect -465 3465 -450 3485
rect -500 3435 -450 3465
rect -500 3415 -485 3435
rect -465 3415 -450 3435
rect -500 3385 -450 3415
rect -500 3365 -485 3385
rect -465 3365 -450 3385
rect -500 3335 -450 3365
rect -500 3315 -485 3335
rect -465 3315 -450 3335
rect -500 3285 -450 3315
rect -500 3265 -485 3285
rect -465 3265 -450 3285
rect -500 3235 -450 3265
rect -500 3215 -485 3235
rect -465 3215 -450 3235
rect -500 3185 -450 3215
rect -500 3165 -485 3185
rect -465 3165 -450 3185
rect -500 3135 -450 3165
rect -500 3115 -485 3135
rect -465 3115 -450 3135
rect -500 3085 -450 3115
rect -500 3065 -485 3085
rect -465 3065 -450 3085
rect -500 3050 -450 3065
rect -350 3535 -300 3550
rect -350 3515 -335 3535
rect -315 3515 -300 3535
rect -350 3485 -300 3515
rect -350 3465 -335 3485
rect -315 3465 -300 3485
rect -350 3435 -300 3465
rect -350 3415 -335 3435
rect -315 3415 -300 3435
rect -350 3385 -300 3415
rect -350 3365 -335 3385
rect -315 3365 -300 3385
rect -350 3335 -300 3365
rect -350 3315 -335 3335
rect -315 3315 -300 3335
rect -350 3285 -300 3315
rect -350 3265 -335 3285
rect -315 3265 -300 3285
rect -350 3235 -300 3265
rect -350 3215 -335 3235
rect -315 3215 -300 3235
rect -350 3185 -300 3215
rect -350 3165 -335 3185
rect -315 3165 -300 3185
rect -350 3135 -300 3165
rect -350 3115 -335 3135
rect -315 3115 -300 3135
rect -350 3085 -300 3115
rect -350 3065 -335 3085
rect -315 3065 -300 3085
rect -350 3050 -300 3065
rect -200 3535 -150 3550
rect -200 3515 -185 3535
rect -165 3515 -150 3535
rect -200 3485 -150 3515
rect -200 3465 -185 3485
rect -165 3465 -150 3485
rect -200 3435 -150 3465
rect -200 3415 -185 3435
rect -165 3415 -150 3435
rect -200 3385 -150 3415
rect -200 3365 -185 3385
rect -165 3365 -150 3385
rect -200 3335 -150 3365
rect -200 3315 -185 3335
rect -165 3315 -150 3335
rect -200 3285 -150 3315
rect -200 3265 -185 3285
rect -165 3265 -150 3285
rect -200 3235 -150 3265
rect -200 3215 -185 3235
rect -165 3215 -150 3235
rect -200 3185 -150 3215
rect -200 3165 -185 3185
rect -165 3165 -150 3185
rect -200 3135 -150 3165
rect -200 3115 -185 3135
rect -165 3115 -150 3135
rect -200 3085 -150 3115
rect -200 3065 -185 3085
rect -165 3065 -150 3085
rect -200 3050 -150 3065
rect -50 3535 0 3550
rect -50 3515 -35 3535
rect -15 3515 0 3535
rect -50 3485 0 3515
rect -50 3465 -35 3485
rect -15 3465 0 3485
rect -50 3435 0 3465
rect -50 3415 -35 3435
rect -15 3415 0 3435
rect -50 3385 0 3415
rect -50 3365 -35 3385
rect -15 3365 0 3385
rect -50 3335 0 3365
rect -50 3315 -35 3335
rect -15 3315 0 3335
rect -50 3285 0 3315
rect -50 3265 -35 3285
rect -15 3265 0 3285
rect -50 3235 0 3265
rect -50 3215 -35 3235
rect -15 3215 0 3235
rect -50 3185 0 3215
rect -50 3165 -35 3185
rect -15 3165 0 3185
rect -50 3135 0 3165
rect -50 3115 -35 3135
rect -15 3115 0 3135
rect -50 3085 0 3115
rect -50 3065 -35 3085
rect -15 3065 0 3085
rect -50 3050 0 3065
rect 100 3050 150 3550
rect 250 3050 300 3550
rect 400 3050 450 3550
rect 550 3535 600 3550
rect 550 3515 565 3535
rect 585 3515 600 3535
rect 550 3485 600 3515
rect 550 3465 565 3485
rect 585 3465 600 3485
rect 550 3435 600 3465
rect 550 3415 565 3435
rect 585 3415 600 3435
rect 550 3385 600 3415
rect 550 3365 565 3385
rect 585 3365 600 3385
rect 550 3335 600 3365
rect 550 3315 565 3335
rect 585 3315 600 3335
rect 550 3285 600 3315
rect 550 3265 565 3285
rect 585 3265 600 3285
rect 550 3235 600 3265
rect 550 3215 565 3235
rect 585 3215 600 3235
rect 550 3185 600 3215
rect 550 3165 565 3185
rect 585 3165 600 3185
rect 550 3135 600 3165
rect 550 3115 565 3135
rect 585 3115 600 3135
rect 550 3085 600 3115
rect 550 3065 565 3085
rect 585 3065 600 3085
rect 550 3050 600 3065
rect 700 3535 750 3550
rect 700 3515 715 3535
rect 735 3515 750 3535
rect 700 3485 750 3515
rect 700 3465 715 3485
rect 735 3465 750 3485
rect 700 3435 750 3465
rect 700 3415 715 3435
rect 735 3415 750 3435
rect 700 3385 750 3415
rect 700 3365 715 3385
rect 735 3365 750 3385
rect 700 3335 750 3365
rect 700 3315 715 3335
rect 735 3315 750 3335
rect 700 3285 750 3315
rect 700 3265 715 3285
rect 735 3265 750 3285
rect 700 3235 750 3265
rect 700 3215 715 3235
rect 735 3215 750 3235
rect 700 3185 750 3215
rect 700 3165 715 3185
rect 735 3165 750 3185
rect 700 3135 750 3165
rect 700 3115 715 3135
rect 735 3115 750 3135
rect 700 3085 750 3115
rect 700 3065 715 3085
rect 735 3065 750 3085
rect 700 3050 750 3065
rect 850 3535 900 3550
rect 850 3515 865 3535
rect 885 3515 900 3535
rect 850 3485 900 3515
rect 850 3465 865 3485
rect 885 3465 900 3485
rect 850 3435 900 3465
rect 850 3415 865 3435
rect 885 3415 900 3435
rect 850 3385 900 3415
rect 850 3365 865 3385
rect 885 3365 900 3385
rect 850 3335 900 3365
rect 850 3315 865 3335
rect 885 3315 900 3335
rect 850 3285 900 3315
rect 850 3265 865 3285
rect 885 3265 900 3285
rect 850 3235 900 3265
rect 850 3215 865 3235
rect 885 3215 900 3235
rect 850 3185 900 3215
rect 850 3165 865 3185
rect 885 3165 900 3185
rect 850 3135 900 3165
rect 850 3115 865 3135
rect 885 3115 900 3135
rect 850 3085 900 3115
rect 850 3065 865 3085
rect 885 3065 900 3085
rect 850 3050 900 3065
rect 1000 3535 1050 3550
rect 1000 3515 1015 3535
rect 1035 3515 1050 3535
rect 1000 3485 1050 3515
rect 1000 3465 1015 3485
rect 1035 3465 1050 3485
rect 1000 3435 1050 3465
rect 1000 3415 1015 3435
rect 1035 3415 1050 3435
rect 1000 3385 1050 3415
rect 1000 3365 1015 3385
rect 1035 3365 1050 3385
rect 1000 3335 1050 3365
rect 1000 3315 1015 3335
rect 1035 3315 1050 3335
rect 1000 3285 1050 3315
rect 1000 3265 1015 3285
rect 1035 3265 1050 3285
rect 1000 3235 1050 3265
rect 1000 3215 1015 3235
rect 1035 3215 1050 3235
rect 1000 3185 1050 3215
rect 1000 3165 1015 3185
rect 1035 3165 1050 3185
rect 1000 3135 1050 3165
rect 1000 3115 1015 3135
rect 1035 3115 1050 3135
rect 1000 3085 1050 3115
rect 1000 3065 1015 3085
rect 1035 3065 1050 3085
rect 1000 3050 1050 3065
rect 1150 3535 1200 3550
rect 1150 3515 1165 3535
rect 1185 3515 1200 3535
rect 1150 3485 1200 3515
rect 1150 3465 1165 3485
rect 1185 3465 1200 3485
rect 1150 3435 1200 3465
rect 1150 3415 1165 3435
rect 1185 3415 1200 3435
rect 1150 3385 1200 3415
rect 1150 3365 1165 3385
rect 1185 3365 1200 3385
rect 1150 3335 1200 3365
rect 1150 3315 1165 3335
rect 1185 3315 1200 3335
rect 1150 3285 1200 3315
rect 1150 3265 1165 3285
rect 1185 3265 1200 3285
rect 1150 3235 1200 3265
rect 1150 3215 1165 3235
rect 1185 3215 1200 3235
rect 1150 3185 1200 3215
rect 1150 3165 1165 3185
rect 1185 3165 1200 3185
rect 1150 3135 1200 3165
rect 1150 3115 1165 3135
rect 1185 3115 1200 3135
rect 1150 3085 1200 3115
rect 1150 3065 1165 3085
rect 1185 3065 1200 3085
rect 1150 3050 1200 3065
rect 1300 3535 1350 3550
rect 1300 3515 1315 3535
rect 1335 3515 1350 3535
rect 1300 3485 1350 3515
rect 1300 3465 1315 3485
rect 1335 3465 1350 3485
rect 1300 3435 1350 3465
rect 1300 3415 1315 3435
rect 1335 3415 1350 3435
rect 1300 3385 1350 3415
rect 1300 3365 1315 3385
rect 1335 3365 1350 3385
rect 1300 3335 1350 3365
rect 1300 3315 1315 3335
rect 1335 3315 1350 3335
rect 1300 3285 1350 3315
rect 1300 3265 1315 3285
rect 1335 3265 1350 3285
rect 1300 3235 1350 3265
rect 1300 3215 1315 3235
rect 1335 3215 1350 3235
rect 1300 3185 1350 3215
rect 1300 3165 1315 3185
rect 1335 3165 1350 3185
rect 1300 3135 1350 3165
rect 1300 3115 1315 3135
rect 1335 3115 1350 3135
rect 1300 3085 1350 3115
rect 1300 3065 1315 3085
rect 1335 3065 1350 3085
rect 1300 3050 1350 3065
rect 1450 3535 1500 3550
rect 1450 3515 1465 3535
rect 1485 3515 1500 3535
rect 1450 3485 1500 3515
rect 1450 3465 1465 3485
rect 1485 3465 1500 3485
rect 1450 3435 1500 3465
rect 1450 3415 1465 3435
rect 1485 3415 1500 3435
rect 1450 3385 1500 3415
rect 1450 3365 1465 3385
rect 1485 3365 1500 3385
rect 1450 3335 1500 3365
rect 1450 3315 1465 3335
rect 1485 3315 1500 3335
rect 1450 3285 1500 3315
rect 1450 3265 1465 3285
rect 1485 3265 1500 3285
rect 1450 3235 1500 3265
rect 1450 3215 1465 3235
rect 1485 3215 1500 3235
rect 1450 3185 1500 3215
rect 1450 3165 1465 3185
rect 1485 3165 1500 3185
rect 1450 3135 1500 3165
rect 1450 3115 1465 3135
rect 1485 3115 1500 3135
rect 1450 3085 1500 3115
rect 1450 3065 1465 3085
rect 1485 3065 1500 3085
rect 1450 3050 1500 3065
rect 1600 3535 1650 3550
rect 1600 3515 1615 3535
rect 1635 3515 1650 3535
rect 1600 3485 1650 3515
rect 1600 3465 1615 3485
rect 1635 3465 1650 3485
rect 1600 3435 1650 3465
rect 1600 3415 1615 3435
rect 1635 3415 1650 3435
rect 1600 3385 1650 3415
rect 1600 3365 1615 3385
rect 1635 3365 1650 3385
rect 1600 3335 1650 3365
rect 1600 3315 1615 3335
rect 1635 3315 1650 3335
rect 1600 3285 1650 3315
rect 1600 3265 1615 3285
rect 1635 3265 1650 3285
rect 1600 3235 1650 3265
rect 1600 3215 1615 3235
rect 1635 3215 1650 3235
rect 1600 3185 1650 3215
rect 1600 3165 1615 3185
rect 1635 3165 1650 3185
rect 1600 3135 1650 3165
rect 1600 3115 1615 3135
rect 1635 3115 1650 3135
rect 1600 3085 1650 3115
rect 1600 3065 1615 3085
rect 1635 3065 1650 3085
rect 1600 3050 1650 3065
rect 1750 3535 1800 3550
rect 1750 3515 1765 3535
rect 1785 3515 1800 3535
rect 1750 3485 1800 3515
rect 1750 3465 1765 3485
rect 1785 3465 1800 3485
rect 1750 3435 1800 3465
rect 1750 3415 1765 3435
rect 1785 3415 1800 3435
rect 1750 3385 1800 3415
rect 1750 3365 1765 3385
rect 1785 3365 1800 3385
rect 1750 3335 1800 3365
rect 1750 3315 1765 3335
rect 1785 3315 1800 3335
rect 1750 3285 1800 3315
rect 1750 3265 1765 3285
rect 1785 3265 1800 3285
rect 1750 3235 1800 3265
rect 1750 3215 1765 3235
rect 1785 3215 1800 3235
rect 1750 3185 1800 3215
rect 1750 3165 1765 3185
rect 1785 3165 1800 3185
rect 1750 3135 1800 3165
rect 1750 3115 1765 3135
rect 1785 3115 1800 3135
rect 1750 3085 1800 3115
rect 1750 3065 1765 3085
rect 1785 3065 1800 3085
rect 1750 3050 1800 3065
rect 1900 3535 1950 3550
rect 1900 3515 1915 3535
rect 1935 3515 1950 3535
rect 1900 3485 1950 3515
rect 1900 3465 1915 3485
rect 1935 3465 1950 3485
rect 1900 3435 1950 3465
rect 1900 3415 1915 3435
rect 1935 3415 1950 3435
rect 1900 3385 1950 3415
rect 1900 3365 1915 3385
rect 1935 3365 1950 3385
rect 1900 3335 1950 3365
rect 1900 3315 1915 3335
rect 1935 3315 1950 3335
rect 1900 3285 1950 3315
rect 1900 3265 1915 3285
rect 1935 3265 1950 3285
rect 1900 3235 1950 3265
rect 1900 3215 1915 3235
rect 1935 3215 1950 3235
rect 1900 3185 1950 3215
rect 1900 3165 1915 3185
rect 1935 3165 1950 3185
rect 1900 3135 1950 3165
rect 1900 3115 1915 3135
rect 1935 3115 1950 3135
rect 1900 3085 1950 3115
rect 1900 3065 1915 3085
rect 1935 3065 1950 3085
rect 1900 3050 1950 3065
rect 2050 3535 2100 3550
rect 2050 3515 2065 3535
rect 2085 3515 2100 3535
rect 2050 3485 2100 3515
rect 2050 3465 2065 3485
rect 2085 3465 2100 3485
rect 2050 3435 2100 3465
rect 2050 3415 2065 3435
rect 2085 3415 2100 3435
rect 2050 3385 2100 3415
rect 2050 3365 2065 3385
rect 2085 3365 2100 3385
rect 2050 3335 2100 3365
rect 2050 3315 2065 3335
rect 2085 3315 2100 3335
rect 2050 3285 2100 3315
rect 2050 3265 2065 3285
rect 2085 3265 2100 3285
rect 2050 3235 2100 3265
rect 2050 3215 2065 3235
rect 2085 3215 2100 3235
rect 2050 3185 2100 3215
rect 2050 3165 2065 3185
rect 2085 3165 2100 3185
rect 2050 3135 2100 3165
rect 2050 3115 2065 3135
rect 2085 3115 2100 3135
rect 2050 3085 2100 3115
rect 2050 3065 2065 3085
rect 2085 3065 2100 3085
rect 2050 3050 2100 3065
rect 2200 3535 2250 3550
rect 2200 3515 2215 3535
rect 2235 3515 2250 3535
rect 2200 3485 2250 3515
rect 2200 3465 2215 3485
rect 2235 3465 2250 3485
rect 2200 3435 2250 3465
rect 2200 3415 2215 3435
rect 2235 3415 2250 3435
rect 2200 3385 2250 3415
rect 2200 3365 2215 3385
rect 2235 3365 2250 3385
rect 2200 3335 2250 3365
rect 2200 3315 2215 3335
rect 2235 3315 2250 3335
rect 2200 3285 2250 3315
rect 2200 3265 2215 3285
rect 2235 3265 2250 3285
rect 2200 3235 2250 3265
rect 2200 3215 2215 3235
rect 2235 3215 2250 3235
rect 2200 3185 2250 3215
rect 2200 3165 2215 3185
rect 2235 3165 2250 3185
rect 2200 3135 2250 3165
rect 2200 3115 2215 3135
rect 2235 3115 2250 3135
rect 2200 3085 2250 3115
rect 2200 3065 2215 3085
rect 2235 3065 2250 3085
rect 2200 3050 2250 3065
rect 2350 3535 2400 3550
rect 2350 3515 2365 3535
rect 2385 3515 2400 3535
rect 2350 3485 2400 3515
rect 2350 3465 2365 3485
rect 2385 3465 2400 3485
rect 2350 3435 2400 3465
rect 2350 3415 2365 3435
rect 2385 3415 2400 3435
rect 2350 3385 2400 3415
rect 2350 3365 2365 3385
rect 2385 3365 2400 3385
rect 2350 3335 2400 3365
rect 2350 3315 2365 3335
rect 2385 3315 2400 3335
rect 2350 3285 2400 3315
rect 2350 3265 2365 3285
rect 2385 3265 2400 3285
rect 2350 3235 2400 3265
rect 2350 3215 2365 3235
rect 2385 3215 2400 3235
rect 2350 3185 2400 3215
rect 2350 3165 2365 3185
rect 2385 3165 2400 3185
rect 2350 3135 2400 3165
rect 2350 3115 2365 3135
rect 2385 3115 2400 3135
rect 2350 3085 2400 3115
rect 2350 3065 2365 3085
rect 2385 3065 2400 3085
rect 2350 3050 2400 3065
rect 2500 3535 2550 3550
rect 2500 3515 2515 3535
rect 2535 3515 2550 3535
rect 2500 3485 2550 3515
rect 2500 3465 2515 3485
rect 2535 3465 2550 3485
rect 2500 3435 2550 3465
rect 2500 3415 2515 3435
rect 2535 3415 2550 3435
rect 2500 3385 2550 3415
rect 2500 3365 2515 3385
rect 2535 3365 2550 3385
rect 2500 3335 2550 3365
rect 2500 3315 2515 3335
rect 2535 3315 2550 3335
rect 2500 3285 2550 3315
rect 2500 3265 2515 3285
rect 2535 3265 2550 3285
rect 2500 3235 2550 3265
rect 2500 3215 2515 3235
rect 2535 3215 2550 3235
rect 2500 3185 2550 3215
rect 2500 3165 2515 3185
rect 2535 3165 2550 3185
rect 2500 3135 2550 3165
rect 2500 3115 2515 3135
rect 2535 3115 2550 3135
rect 2500 3085 2550 3115
rect 2500 3065 2515 3085
rect 2535 3065 2550 3085
rect 2500 3050 2550 3065
rect 2650 3535 2700 3550
rect 2650 3515 2665 3535
rect 2685 3515 2700 3535
rect 2650 3485 2700 3515
rect 2650 3465 2665 3485
rect 2685 3465 2700 3485
rect 2650 3435 2700 3465
rect 2650 3415 2665 3435
rect 2685 3415 2700 3435
rect 2650 3385 2700 3415
rect 2650 3365 2665 3385
rect 2685 3365 2700 3385
rect 2650 3335 2700 3365
rect 2650 3315 2665 3335
rect 2685 3315 2700 3335
rect 2650 3285 2700 3315
rect 2650 3265 2665 3285
rect 2685 3265 2700 3285
rect 2650 3235 2700 3265
rect 2650 3215 2665 3235
rect 2685 3215 2700 3235
rect 2650 3185 2700 3215
rect 2650 3165 2665 3185
rect 2685 3165 2700 3185
rect 2650 3135 2700 3165
rect 2650 3115 2665 3135
rect 2685 3115 2700 3135
rect 2650 3085 2700 3115
rect 2650 3065 2665 3085
rect 2685 3065 2700 3085
rect 2650 3050 2700 3065
rect 2800 3535 2850 3550
rect 2800 3515 2815 3535
rect 2835 3515 2850 3535
rect 2800 3485 2850 3515
rect 2800 3465 2815 3485
rect 2835 3465 2850 3485
rect 2800 3435 2850 3465
rect 2800 3415 2815 3435
rect 2835 3415 2850 3435
rect 2800 3385 2850 3415
rect 2800 3365 2815 3385
rect 2835 3365 2850 3385
rect 2800 3335 2850 3365
rect 2800 3315 2815 3335
rect 2835 3315 2850 3335
rect 2800 3285 2850 3315
rect 2800 3265 2815 3285
rect 2835 3265 2850 3285
rect 2800 3235 2850 3265
rect 2800 3215 2815 3235
rect 2835 3215 2850 3235
rect 2800 3185 2850 3215
rect 2800 3165 2815 3185
rect 2835 3165 2850 3185
rect 2800 3135 2850 3165
rect 2800 3115 2815 3135
rect 2835 3115 2850 3135
rect 2800 3085 2850 3115
rect 2800 3065 2815 3085
rect 2835 3065 2850 3085
rect 2800 3050 2850 3065
rect 2950 3535 3000 3550
rect 2950 3515 2965 3535
rect 2985 3515 3000 3535
rect 2950 3485 3000 3515
rect 2950 3465 2965 3485
rect 2985 3465 3000 3485
rect 2950 3435 3000 3465
rect 2950 3415 2965 3435
rect 2985 3415 3000 3435
rect 2950 3385 3000 3415
rect 2950 3365 2965 3385
rect 2985 3365 3000 3385
rect 2950 3335 3000 3365
rect 2950 3315 2965 3335
rect 2985 3315 3000 3335
rect 2950 3285 3000 3315
rect 2950 3265 2965 3285
rect 2985 3265 3000 3285
rect 2950 3235 3000 3265
rect 2950 3215 2965 3235
rect 2985 3215 3000 3235
rect 2950 3185 3000 3215
rect 2950 3165 2965 3185
rect 2985 3165 3000 3185
rect 2950 3135 3000 3165
rect 2950 3115 2965 3135
rect 2985 3115 3000 3135
rect 2950 3085 3000 3115
rect 2950 3065 2965 3085
rect 2985 3065 3000 3085
rect 2950 3050 3000 3065
rect 3100 3535 3150 3550
rect 3100 3515 3115 3535
rect 3135 3515 3150 3535
rect 3100 3485 3150 3515
rect 3100 3465 3115 3485
rect 3135 3465 3150 3485
rect 3100 3435 3150 3465
rect 3100 3415 3115 3435
rect 3135 3415 3150 3435
rect 3100 3385 3150 3415
rect 3100 3365 3115 3385
rect 3135 3365 3150 3385
rect 3100 3335 3150 3365
rect 3100 3315 3115 3335
rect 3135 3315 3150 3335
rect 3100 3285 3150 3315
rect 3100 3265 3115 3285
rect 3135 3265 3150 3285
rect 3100 3235 3150 3265
rect 3100 3215 3115 3235
rect 3135 3215 3150 3235
rect 3100 3185 3150 3215
rect 3100 3165 3115 3185
rect 3135 3165 3150 3185
rect 3100 3135 3150 3165
rect 3100 3115 3115 3135
rect 3135 3115 3150 3135
rect 3100 3085 3150 3115
rect 3100 3065 3115 3085
rect 3135 3065 3150 3085
rect 3100 3050 3150 3065
rect 3250 3535 3300 3550
rect 3250 3515 3265 3535
rect 3285 3515 3300 3535
rect 3250 3485 3300 3515
rect 3250 3465 3265 3485
rect 3285 3465 3300 3485
rect 3250 3435 3300 3465
rect 3250 3415 3265 3435
rect 3285 3415 3300 3435
rect 3250 3385 3300 3415
rect 3250 3365 3265 3385
rect 3285 3365 3300 3385
rect 3250 3335 3300 3365
rect 3250 3315 3265 3335
rect 3285 3315 3300 3335
rect 3250 3285 3300 3315
rect 3250 3265 3265 3285
rect 3285 3265 3300 3285
rect 3250 3235 3300 3265
rect 3250 3215 3265 3235
rect 3285 3215 3300 3235
rect 3250 3185 3300 3215
rect 3250 3165 3265 3185
rect 3285 3165 3300 3185
rect 3250 3135 3300 3165
rect 3250 3115 3265 3135
rect 3285 3115 3300 3135
rect 3250 3085 3300 3115
rect 3250 3065 3265 3085
rect 3285 3065 3300 3085
rect 3250 3050 3300 3065
rect 3400 3535 3450 3550
rect 3400 3515 3415 3535
rect 3435 3515 3450 3535
rect 3400 3485 3450 3515
rect 3400 3465 3415 3485
rect 3435 3465 3450 3485
rect 3400 3435 3450 3465
rect 3400 3415 3415 3435
rect 3435 3415 3450 3435
rect 3400 3385 3450 3415
rect 3400 3365 3415 3385
rect 3435 3365 3450 3385
rect 3400 3335 3450 3365
rect 3400 3315 3415 3335
rect 3435 3315 3450 3335
rect 3400 3285 3450 3315
rect 3400 3265 3415 3285
rect 3435 3265 3450 3285
rect 3400 3235 3450 3265
rect 3400 3215 3415 3235
rect 3435 3215 3450 3235
rect 3400 3185 3450 3215
rect 3400 3165 3415 3185
rect 3435 3165 3450 3185
rect 3400 3135 3450 3165
rect 3400 3115 3415 3135
rect 3435 3115 3450 3135
rect 3400 3085 3450 3115
rect 3400 3065 3415 3085
rect 3435 3065 3450 3085
rect 3400 3050 3450 3065
rect 3550 3535 3600 3550
rect 3550 3515 3565 3535
rect 3585 3515 3600 3535
rect 3550 3485 3600 3515
rect 3550 3465 3565 3485
rect 3585 3465 3600 3485
rect 3550 3435 3600 3465
rect 3550 3415 3565 3435
rect 3585 3415 3600 3435
rect 3550 3385 3600 3415
rect 3550 3365 3565 3385
rect 3585 3365 3600 3385
rect 3550 3335 3600 3365
rect 3550 3315 3565 3335
rect 3585 3315 3600 3335
rect 3550 3285 3600 3315
rect 3550 3265 3565 3285
rect 3585 3265 3600 3285
rect 3550 3235 3600 3265
rect 3550 3215 3565 3235
rect 3585 3215 3600 3235
rect 3550 3185 3600 3215
rect 3550 3165 3565 3185
rect 3585 3165 3600 3185
rect 3550 3135 3600 3165
rect 3550 3115 3565 3135
rect 3585 3115 3600 3135
rect 3550 3085 3600 3115
rect 3550 3065 3565 3085
rect 3585 3065 3600 3085
rect 3550 3050 3600 3065
rect 3700 3050 3750 3550
rect 3850 3050 3900 3550
rect 4000 3050 4050 3550
rect 4150 3535 4200 3550
rect 4150 3515 4165 3535
rect 4185 3515 4200 3535
rect 4150 3485 4200 3515
rect 4150 3465 4165 3485
rect 4185 3465 4200 3485
rect 4150 3435 4200 3465
rect 4150 3415 4165 3435
rect 4185 3415 4200 3435
rect 4150 3385 4200 3415
rect 4150 3365 4165 3385
rect 4185 3365 4200 3385
rect 4150 3335 4200 3365
rect 4150 3315 4165 3335
rect 4185 3315 4200 3335
rect 4150 3285 4200 3315
rect 4150 3265 4165 3285
rect 4185 3265 4200 3285
rect 4150 3235 4200 3265
rect 4150 3215 4165 3235
rect 4185 3215 4200 3235
rect 4150 3185 4200 3215
rect 4150 3165 4165 3185
rect 4185 3165 4200 3185
rect 4150 3135 4200 3165
rect 4150 3115 4165 3135
rect 4185 3115 4200 3135
rect 4150 3085 4200 3115
rect 4150 3065 4165 3085
rect 4185 3065 4200 3085
rect 4150 3050 4200 3065
rect 4300 3050 4350 3550
rect 4450 3050 4500 3550
rect 4600 3050 4650 3550
rect 4750 3535 4800 3550
rect 4750 3515 4765 3535
rect 4785 3515 4800 3535
rect 4750 3485 4800 3515
rect 4750 3465 4765 3485
rect 4785 3465 4800 3485
rect 4750 3435 4800 3465
rect 4750 3415 4765 3435
rect 4785 3415 4800 3435
rect 4750 3385 4800 3415
rect 4750 3365 4765 3385
rect 4785 3365 4800 3385
rect 4750 3335 4800 3365
rect 4750 3315 4765 3335
rect 4785 3315 4800 3335
rect 4750 3285 4800 3315
rect 4750 3265 4765 3285
rect 4785 3265 4800 3285
rect 4750 3235 4800 3265
rect 4750 3215 4765 3235
rect 4785 3215 4800 3235
rect 4750 3185 4800 3215
rect 4750 3165 4765 3185
rect 4785 3165 4800 3185
rect 4750 3135 4800 3165
rect 4750 3115 4765 3135
rect 4785 3115 4800 3135
rect 4750 3085 4800 3115
rect 4750 3065 4765 3085
rect 4785 3065 4800 3085
rect 4750 3050 4800 3065
rect 4900 3535 4950 3550
rect 4900 3515 4915 3535
rect 4935 3515 4950 3535
rect 4900 3485 4950 3515
rect 4900 3465 4915 3485
rect 4935 3465 4950 3485
rect 4900 3435 4950 3465
rect 4900 3415 4915 3435
rect 4935 3415 4950 3435
rect 4900 3385 4950 3415
rect 4900 3365 4915 3385
rect 4935 3365 4950 3385
rect 4900 3335 4950 3365
rect 4900 3315 4915 3335
rect 4935 3315 4950 3335
rect 4900 3285 4950 3315
rect 4900 3265 4915 3285
rect 4935 3265 4950 3285
rect 4900 3235 4950 3265
rect 4900 3215 4915 3235
rect 4935 3215 4950 3235
rect 4900 3185 4950 3215
rect 4900 3165 4915 3185
rect 4935 3165 4950 3185
rect 4900 3135 4950 3165
rect 4900 3115 4915 3135
rect 4935 3115 4950 3135
rect 4900 3085 4950 3115
rect 4900 3065 4915 3085
rect 4935 3065 4950 3085
rect 4900 3050 4950 3065
rect 5050 3535 5100 3550
rect 5050 3515 5065 3535
rect 5085 3515 5100 3535
rect 5050 3485 5100 3515
rect 5050 3465 5065 3485
rect 5085 3465 5100 3485
rect 5050 3435 5100 3465
rect 5050 3415 5065 3435
rect 5085 3415 5100 3435
rect 5050 3385 5100 3415
rect 5050 3365 5065 3385
rect 5085 3365 5100 3385
rect 5050 3335 5100 3365
rect 5050 3315 5065 3335
rect 5085 3315 5100 3335
rect 5050 3285 5100 3315
rect 5050 3265 5065 3285
rect 5085 3265 5100 3285
rect 5050 3235 5100 3265
rect 5050 3215 5065 3235
rect 5085 3215 5100 3235
rect 5050 3185 5100 3215
rect 5050 3165 5065 3185
rect 5085 3165 5100 3185
rect 5050 3135 5100 3165
rect 5050 3115 5065 3135
rect 5085 3115 5100 3135
rect 5050 3085 5100 3115
rect 5050 3065 5065 3085
rect 5085 3065 5100 3085
rect 5050 3050 5100 3065
rect 5200 3535 5250 3550
rect 5200 3515 5215 3535
rect 5235 3515 5250 3535
rect 5200 3485 5250 3515
rect 5200 3465 5215 3485
rect 5235 3465 5250 3485
rect 5200 3435 5250 3465
rect 5200 3415 5215 3435
rect 5235 3415 5250 3435
rect 5200 3385 5250 3415
rect 5200 3365 5215 3385
rect 5235 3365 5250 3385
rect 5200 3335 5250 3365
rect 5200 3315 5215 3335
rect 5235 3315 5250 3335
rect 5200 3285 5250 3315
rect 5200 3265 5215 3285
rect 5235 3265 5250 3285
rect 5200 3235 5250 3265
rect 5200 3215 5215 3235
rect 5235 3215 5250 3235
rect 5200 3185 5250 3215
rect 5200 3165 5215 3185
rect 5235 3165 5250 3185
rect 5200 3135 5250 3165
rect 5200 3115 5215 3135
rect 5235 3115 5250 3135
rect 5200 3085 5250 3115
rect 5200 3065 5215 3085
rect 5235 3065 5250 3085
rect 5200 3050 5250 3065
rect 5350 3535 5400 3550
rect 5350 3515 5365 3535
rect 5385 3515 5400 3535
rect 5350 3485 5400 3515
rect 5350 3465 5365 3485
rect 5385 3465 5400 3485
rect 5350 3435 5400 3465
rect 5350 3415 5365 3435
rect 5385 3415 5400 3435
rect 5350 3385 5400 3415
rect 5350 3365 5365 3385
rect 5385 3365 5400 3385
rect 5350 3335 5400 3365
rect 5350 3315 5365 3335
rect 5385 3315 5400 3335
rect 5350 3285 5400 3315
rect 5350 3265 5365 3285
rect 5385 3265 5400 3285
rect 5350 3235 5400 3265
rect 5350 3215 5365 3235
rect 5385 3215 5400 3235
rect 5350 3185 5400 3215
rect 5350 3165 5365 3185
rect 5385 3165 5400 3185
rect 5350 3135 5400 3165
rect 5350 3115 5365 3135
rect 5385 3115 5400 3135
rect 5350 3085 5400 3115
rect 5350 3065 5365 3085
rect 5385 3065 5400 3085
rect 5350 3050 5400 3065
rect 5500 3535 5550 3550
rect 5500 3515 5515 3535
rect 5535 3515 5550 3535
rect 5500 3485 5550 3515
rect 5500 3465 5515 3485
rect 5535 3465 5550 3485
rect 5500 3435 5550 3465
rect 5500 3415 5515 3435
rect 5535 3415 5550 3435
rect 5500 3385 5550 3415
rect 5500 3365 5515 3385
rect 5535 3365 5550 3385
rect 5500 3335 5550 3365
rect 5500 3315 5515 3335
rect 5535 3315 5550 3335
rect 5500 3285 5550 3315
rect 5500 3265 5515 3285
rect 5535 3265 5550 3285
rect 5500 3235 5550 3265
rect 5500 3215 5515 3235
rect 5535 3215 5550 3235
rect 5500 3185 5550 3215
rect 5500 3165 5515 3185
rect 5535 3165 5550 3185
rect 5500 3135 5550 3165
rect 5500 3115 5515 3135
rect 5535 3115 5550 3135
rect 5500 3085 5550 3115
rect 5500 3065 5515 3085
rect 5535 3065 5550 3085
rect 5500 3050 5550 3065
rect 5650 3535 5700 3550
rect 5650 3515 5665 3535
rect 5685 3515 5700 3535
rect 5650 3485 5700 3515
rect 5650 3465 5665 3485
rect 5685 3465 5700 3485
rect 5650 3435 5700 3465
rect 5650 3415 5665 3435
rect 5685 3415 5700 3435
rect 5650 3385 5700 3415
rect 5650 3365 5665 3385
rect 5685 3365 5700 3385
rect 5650 3335 5700 3365
rect 5650 3315 5665 3335
rect 5685 3315 5700 3335
rect 5650 3285 5700 3315
rect 5650 3265 5665 3285
rect 5685 3265 5700 3285
rect 5650 3235 5700 3265
rect 5650 3215 5665 3235
rect 5685 3215 5700 3235
rect 5650 3185 5700 3215
rect 5650 3165 5665 3185
rect 5685 3165 5700 3185
rect 5650 3135 5700 3165
rect 5650 3115 5665 3135
rect 5685 3115 5700 3135
rect 5650 3085 5700 3115
rect 5650 3065 5665 3085
rect 5685 3065 5700 3085
rect 5650 3050 5700 3065
rect 5800 3535 5850 3550
rect 5800 3515 5815 3535
rect 5835 3515 5850 3535
rect 5800 3485 5850 3515
rect 5800 3465 5815 3485
rect 5835 3465 5850 3485
rect 5800 3435 5850 3465
rect 5800 3415 5815 3435
rect 5835 3415 5850 3435
rect 5800 3385 5850 3415
rect 5800 3365 5815 3385
rect 5835 3365 5850 3385
rect 5800 3335 5850 3365
rect 5800 3315 5815 3335
rect 5835 3315 5850 3335
rect 5800 3285 5850 3315
rect 5800 3265 5815 3285
rect 5835 3265 5850 3285
rect 5800 3235 5850 3265
rect 5800 3215 5815 3235
rect 5835 3215 5850 3235
rect 5800 3185 5850 3215
rect 5800 3165 5815 3185
rect 5835 3165 5850 3185
rect 5800 3135 5850 3165
rect 5800 3115 5815 3135
rect 5835 3115 5850 3135
rect 5800 3085 5850 3115
rect 5800 3065 5815 3085
rect 5835 3065 5850 3085
rect 5800 3050 5850 3065
rect 5950 3535 6000 3550
rect 5950 3515 5965 3535
rect 5985 3515 6000 3535
rect 5950 3485 6000 3515
rect 5950 3465 5965 3485
rect 5985 3465 6000 3485
rect 5950 3435 6000 3465
rect 5950 3415 5965 3435
rect 5985 3415 6000 3435
rect 5950 3385 6000 3415
rect 5950 3365 5965 3385
rect 5985 3365 6000 3385
rect 5950 3335 6000 3365
rect 5950 3315 5965 3335
rect 5985 3315 6000 3335
rect 5950 3285 6000 3315
rect 5950 3265 5965 3285
rect 5985 3265 6000 3285
rect 5950 3235 6000 3265
rect 5950 3215 5965 3235
rect 5985 3215 6000 3235
rect 5950 3185 6000 3215
rect 5950 3165 5965 3185
rect 5985 3165 6000 3185
rect 5950 3135 6000 3165
rect 5950 3115 5965 3135
rect 5985 3115 6000 3135
rect 5950 3085 6000 3115
rect 5950 3065 5965 3085
rect 5985 3065 6000 3085
rect 5950 3050 6000 3065
rect 6100 3535 6150 3550
rect 6100 3515 6115 3535
rect 6135 3515 6150 3535
rect 6100 3485 6150 3515
rect 6100 3465 6115 3485
rect 6135 3465 6150 3485
rect 6100 3435 6150 3465
rect 6100 3415 6115 3435
rect 6135 3415 6150 3435
rect 6100 3385 6150 3415
rect 6100 3365 6115 3385
rect 6135 3365 6150 3385
rect 6100 3335 6150 3365
rect 6100 3315 6115 3335
rect 6135 3315 6150 3335
rect 6100 3285 6150 3315
rect 6100 3265 6115 3285
rect 6135 3265 6150 3285
rect 6100 3235 6150 3265
rect 6100 3215 6115 3235
rect 6135 3215 6150 3235
rect 6100 3185 6150 3215
rect 6100 3165 6115 3185
rect 6135 3165 6150 3185
rect 6100 3135 6150 3165
rect 6100 3115 6115 3135
rect 6135 3115 6150 3135
rect 6100 3085 6150 3115
rect 6100 3065 6115 3085
rect 6135 3065 6150 3085
rect 6100 3050 6150 3065
rect 6250 3535 6300 3550
rect 6250 3515 6265 3535
rect 6285 3515 6300 3535
rect 6250 3485 6300 3515
rect 6250 3465 6265 3485
rect 6285 3465 6300 3485
rect 6250 3435 6300 3465
rect 6250 3415 6265 3435
rect 6285 3415 6300 3435
rect 6250 3385 6300 3415
rect 6250 3365 6265 3385
rect 6285 3365 6300 3385
rect 6250 3335 6300 3365
rect 6250 3315 6265 3335
rect 6285 3315 6300 3335
rect 6250 3285 6300 3315
rect 6250 3265 6265 3285
rect 6285 3265 6300 3285
rect 6250 3235 6300 3265
rect 6250 3215 6265 3235
rect 6285 3215 6300 3235
rect 6250 3185 6300 3215
rect 6250 3165 6265 3185
rect 6285 3165 6300 3185
rect 6250 3135 6300 3165
rect 6250 3115 6265 3135
rect 6285 3115 6300 3135
rect 6250 3085 6300 3115
rect 6250 3065 6265 3085
rect 6285 3065 6300 3085
rect 6250 3050 6300 3065
rect 6400 3535 6450 3550
rect 6400 3515 6415 3535
rect 6435 3515 6450 3535
rect 6400 3485 6450 3515
rect 6400 3465 6415 3485
rect 6435 3465 6450 3485
rect 6400 3435 6450 3465
rect 6400 3415 6415 3435
rect 6435 3415 6450 3435
rect 6400 3385 6450 3415
rect 6400 3365 6415 3385
rect 6435 3365 6450 3385
rect 6400 3335 6450 3365
rect 6400 3315 6415 3335
rect 6435 3315 6450 3335
rect 6400 3285 6450 3315
rect 6400 3265 6415 3285
rect 6435 3265 6450 3285
rect 6400 3235 6450 3265
rect 6400 3215 6415 3235
rect 6435 3215 6450 3235
rect 6400 3185 6450 3215
rect 6400 3165 6415 3185
rect 6435 3165 6450 3185
rect 6400 3135 6450 3165
rect 6400 3115 6415 3135
rect 6435 3115 6450 3135
rect 6400 3085 6450 3115
rect 6400 3065 6415 3085
rect 6435 3065 6450 3085
rect 6400 3050 6450 3065
rect 6550 3535 6600 3550
rect 6550 3515 6565 3535
rect 6585 3515 6600 3535
rect 6550 3485 6600 3515
rect 6550 3465 6565 3485
rect 6585 3465 6600 3485
rect 6550 3435 6600 3465
rect 6550 3415 6565 3435
rect 6585 3415 6600 3435
rect 6550 3385 6600 3415
rect 6550 3365 6565 3385
rect 6585 3365 6600 3385
rect 6550 3335 6600 3365
rect 6550 3315 6565 3335
rect 6585 3315 6600 3335
rect 6550 3285 6600 3315
rect 6550 3265 6565 3285
rect 6585 3265 6600 3285
rect 6550 3235 6600 3265
rect 6550 3215 6565 3235
rect 6585 3215 6600 3235
rect 6550 3185 6600 3215
rect 6550 3165 6565 3185
rect 6585 3165 6600 3185
rect 6550 3135 6600 3165
rect 6550 3115 6565 3135
rect 6585 3115 6600 3135
rect 6550 3085 6600 3115
rect 6550 3065 6565 3085
rect 6585 3065 6600 3085
rect 6550 3050 6600 3065
rect 6700 3535 6750 3550
rect 6700 3515 6715 3535
rect 6735 3515 6750 3535
rect 6700 3485 6750 3515
rect 6700 3465 6715 3485
rect 6735 3465 6750 3485
rect 6700 3435 6750 3465
rect 6700 3415 6715 3435
rect 6735 3415 6750 3435
rect 6700 3385 6750 3415
rect 6700 3365 6715 3385
rect 6735 3365 6750 3385
rect 6700 3335 6750 3365
rect 6700 3315 6715 3335
rect 6735 3315 6750 3335
rect 6700 3285 6750 3315
rect 6700 3265 6715 3285
rect 6735 3265 6750 3285
rect 6700 3235 6750 3265
rect 6700 3215 6715 3235
rect 6735 3215 6750 3235
rect 6700 3185 6750 3215
rect 6700 3165 6715 3185
rect 6735 3165 6750 3185
rect 6700 3135 6750 3165
rect 6700 3115 6715 3135
rect 6735 3115 6750 3135
rect 6700 3085 6750 3115
rect 6700 3065 6715 3085
rect 6735 3065 6750 3085
rect 6700 3050 6750 3065
rect 6850 3535 6900 3550
rect 6850 3515 6865 3535
rect 6885 3515 6900 3535
rect 6850 3485 6900 3515
rect 6850 3465 6865 3485
rect 6885 3465 6900 3485
rect 6850 3435 6900 3465
rect 6850 3415 6865 3435
rect 6885 3415 6900 3435
rect 6850 3385 6900 3415
rect 6850 3365 6865 3385
rect 6885 3365 6900 3385
rect 6850 3335 6900 3365
rect 6850 3315 6865 3335
rect 6885 3315 6900 3335
rect 6850 3285 6900 3315
rect 6850 3265 6865 3285
rect 6885 3265 6900 3285
rect 6850 3235 6900 3265
rect 6850 3215 6865 3235
rect 6885 3215 6900 3235
rect 6850 3185 6900 3215
rect 6850 3165 6865 3185
rect 6885 3165 6900 3185
rect 6850 3135 6900 3165
rect 6850 3115 6865 3135
rect 6885 3115 6900 3135
rect 6850 3085 6900 3115
rect 6850 3065 6865 3085
rect 6885 3065 6900 3085
rect 6850 3050 6900 3065
rect 7000 3535 7050 3550
rect 7000 3515 7015 3535
rect 7035 3515 7050 3535
rect 7000 3485 7050 3515
rect 7000 3465 7015 3485
rect 7035 3465 7050 3485
rect 7000 3435 7050 3465
rect 7000 3415 7015 3435
rect 7035 3415 7050 3435
rect 7000 3385 7050 3415
rect 7000 3365 7015 3385
rect 7035 3365 7050 3385
rect 7000 3335 7050 3365
rect 7000 3315 7015 3335
rect 7035 3315 7050 3335
rect 7000 3285 7050 3315
rect 7000 3265 7015 3285
rect 7035 3265 7050 3285
rect 7000 3235 7050 3265
rect 7000 3215 7015 3235
rect 7035 3215 7050 3235
rect 7000 3185 7050 3215
rect 7000 3165 7015 3185
rect 7035 3165 7050 3185
rect 7000 3135 7050 3165
rect 7000 3115 7015 3135
rect 7035 3115 7050 3135
rect 7000 3085 7050 3115
rect 7000 3065 7015 3085
rect 7035 3065 7050 3085
rect 7000 3050 7050 3065
rect 7150 3535 7200 3550
rect 7150 3515 7165 3535
rect 7185 3515 7200 3535
rect 7150 3485 7200 3515
rect 7150 3465 7165 3485
rect 7185 3465 7200 3485
rect 7150 3435 7200 3465
rect 7150 3415 7165 3435
rect 7185 3415 7200 3435
rect 7150 3385 7200 3415
rect 7150 3365 7165 3385
rect 7185 3365 7200 3385
rect 7150 3335 7200 3365
rect 7150 3315 7165 3335
rect 7185 3315 7200 3335
rect 7150 3285 7200 3315
rect 7150 3265 7165 3285
rect 7185 3265 7200 3285
rect 7150 3235 7200 3265
rect 7150 3215 7165 3235
rect 7185 3215 7200 3235
rect 7150 3185 7200 3215
rect 7150 3165 7165 3185
rect 7185 3165 7200 3185
rect 7150 3135 7200 3165
rect 7150 3115 7165 3135
rect 7185 3115 7200 3135
rect 7150 3085 7200 3115
rect 7150 3065 7165 3085
rect 7185 3065 7200 3085
rect 7150 3050 7200 3065
rect 7300 3535 7350 3550
rect 7300 3515 7315 3535
rect 7335 3515 7350 3535
rect 7300 3485 7350 3515
rect 7300 3465 7315 3485
rect 7335 3465 7350 3485
rect 7300 3435 7350 3465
rect 7300 3415 7315 3435
rect 7335 3415 7350 3435
rect 7300 3385 7350 3415
rect 7300 3365 7315 3385
rect 7335 3365 7350 3385
rect 7300 3335 7350 3365
rect 7300 3315 7315 3335
rect 7335 3315 7350 3335
rect 7300 3285 7350 3315
rect 7300 3265 7315 3285
rect 7335 3265 7350 3285
rect 7300 3235 7350 3265
rect 7300 3215 7315 3235
rect 7335 3215 7350 3235
rect 7300 3185 7350 3215
rect 7300 3165 7315 3185
rect 7335 3165 7350 3185
rect 7300 3135 7350 3165
rect 7300 3115 7315 3135
rect 7335 3115 7350 3135
rect 7300 3085 7350 3115
rect 7300 3065 7315 3085
rect 7335 3065 7350 3085
rect 7300 3050 7350 3065
rect 7450 3535 7500 3550
rect 7450 3515 7465 3535
rect 7485 3515 7500 3535
rect 7450 3485 7500 3515
rect 7450 3465 7465 3485
rect 7485 3465 7500 3485
rect 7450 3435 7500 3465
rect 7450 3415 7465 3435
rect 7485 3415 7500 3435
rect 7450 3385 7500 3415
rect 7450 3365 7465 3385
rect 7485 3365 7500 3385
rect 7450 3335 7500 3365
rect 7450 3315 7465 3335
rect 7485 3315 7500 3335
rect 7450 3285 7500 3315
rect 7450 3265 7465 3285
rect 7485 3265 7500 3285
rect 7450 3235 7500 3265
rect 7450 3215 7465 3235
rect 7485 3215 7500 3235
rect 7450 3185 7500 3215
rect 7450 3165 7465 3185
rect 7485 3165 7500 3185
rect 7450 3135 7500 3165
rect 7450 3115 7465 3135
rect 7485 3115 7500 3135
rect 7450 3085 7500 3115
rect 7450 3065 7465 3085
rect 7485 3065 7500 3085
rect 7450 3050 7500 3065
rect 7600 3535 7650 3550
rect 7600 3515 7615 3535
rect 7635 3515 7650 3535
rect 7600 3485 7650 3515
rect 7600 3465 7615 3485
rect 7635 3465 7650 3485
rect 7600 3435 7650 3465
rect 7600 3415 7615 3435
rect 7635 3415 7650 3435
rect 7600 3385 7650 3415
rect 7600 3365 7615 3385
rect 7635 3365 7650 3385
rect 7600 3335 7650 3365
rect 7600 3315 7615 3335
rect 7635 3315 7650 3335
rect 7600 3285 7650 3315
rect 7600 3265 7615 3285
rect 7635 3265 7650 3285
rect 7600 3235 7650 3265
rect 7600 3215 7615 3235
rect 7635 3215 7650 3235
rect 7600 3185 7650 3215
rect 7600 3165 7615 3185
rect 7635 3165 7650 3185
rect 7600 3135 7650 3165
rect 7600 3115 7615 3135
rect 7635 3115 7650 3135
rect 7600 3085 7650 3115
rect 7600 3065 7615 3085
rect 7635 3065 7650 3085
rect 7600 3050 7650 3065
rect 7750 3535 7800 3550
rect 7750 3515 7765 3535
rect 7785 3515 7800 3535
rect 7750 3485 7800 3515
rect 7750 3465 7765 3485
rect 7785 3465 7800 3485
rect 7750 3435 7800 3465
rect 7750 3415 7765 3435
rect 7785 3415 7800 3435
rect 7750 3385 7800 3415
rect 7750 3365 7765 3385
rect 7785 3365 7800 3385
rect 7750 3335 7800 3365
rect 7750 3315 7765 3335
rect 7785 3315 7800 3335
rect 7750 3285 7800 3315
rect 7750 3265 7765 3285
rect 7785 3265 7800 3285
rect 7750 3235 7800 3265
rect 7750 3215 7765 3235
rect 7785 3215 7800 3235
rect 7750 3185 7800 3215
rect 7750 3165 7765 3185
rect 7785 3165 7800 3185
rect 7750 3135 7800 3165
rect 7750 3115 7765 3135
rect 7785 3115 7800 3135
rect 7750 3085 7800 3115
rect 7750 3065 7765 3085
rect 7785 3065 7800 3085
rect 7750 3050 7800 3065
rect 7900 3050 7950 3550
rect 8050 3050 8100 3550
rect 8200 3050 8250 3550
rect 8350 3535 8400 3550
rect 8350 3515 8365 3535
rect 8385 3515 8400 3535
rect 8350 3485 8400 3515
rect 8350 3465 8365 3485
rect 8385 3465 8400 3485
rect 8350 3435 8400 3465
rect 8350 3415 8365 3435
rect 8385 3415 8400 3435
rect 8350 3385 8400 3415
rect 8350 3365 8365 3385
rect 8385 3365 8400 3385
rect 8350 3335 8400 3365
rect 8350 3315 8365 3335
rect 8385 3315 8400 3335
rect 8350 3285 8400 3315
rect 8350 3265 8365 3285
rect 8385 3265 8400 3285
rect 8350 3235 8400 3265
rect 8350 3215 8365 3235
rect 8385 3215 8400 3235
rect 8350 3185 8400 3215
rect 8350 3165 8365 3185
rect 8385 3165 8400 3185
rect 8350 3135 8400 3165
rect 8350 3115 8365 3135
rect 8385 3115 8400 3135
rect 8350 3085 8400 3115
rect 8350 3065 8365 3085
rect 8385 3065 8400 3085
rect 8350 3050 8400 3065
rect 8500 3535 8550 3550
rect 8500 3515 8515 3535
rect 8535 3515 8550 3535
rect 8500 3485 8550 3515
rect 8500 3465 8515 3485
rect 8535 3465 8550 3485
rect 8500 3435 8550 3465
rect 8500 3415 8515 3435
rect 8535 3415 8550 3435
rect 8500 3385 8550 3415
rect 8500 3365 8515 3385
rect 8535 3365 8550 3385
rect 8500 3335 8550 3365
rect 8500 3315 8515 3335
rect 8535 3315 8550 3335
rect 8500 3285 8550 3315
rect 8500 3265 8515 3285
rect 8535 3265 8550 3285
rect 8500 3235 8550 3265
rect 8500 3215 8515 3235
rect 8535 3215 8550 3235
rect 8500 3185 8550 3215
rect 8500 3165 8515 3185
rect 8535 3165 8550 3185
rect 8500 3135 8550 3165
rect 8500 3115 8515 3135
rect 8535 3115 8550 3135
rect 8500 3085 8550 3115
rect 8500 3065 8515 3085
rect 8535 3065 8550 3085
rect 8500 3050 8550 3065
rect 8650 3535 8700 3550
rect 8650 3515 8665 3535
rect 8685 3515 8700 3535
rect 8650 3485 8700 3515
rect 8650 3465 8665 3485
rect 8685 3465 8700 3485
rect 8650 3435 8700 3465
rect 8650 3415 8665 3435
rect 8685 3415 8700 3435
rect 8650 3385 8700 3415
rect 8650 3365 8665 3385
rect 8685 3365 8700 3385
rect 8650 3335 8700 3365
rect 8650 3315 8665 3335
rect 8685 3315 8700 3335
rect 8650 3285 8700 3315
rect 8650 3265 8665 3285
rect 8685 3265 8700 3285
rect 8650 3235 8700 3265
rect 8650 3215 8665 3235
rect 8685 3215 8700 3235
rect 8650 3185 8700 3215
rect 8650 3165 8665 3185
rect 8685 3165 8700 3185
rect 8650 3135 8700 3165
rect 8650 3115 8665 3135
rect 8685 3115 8700 3135
rect 8650 3085 8700 3115
rect 8650 3065 8665 3085
rect 8685 3065 8700 3085
rect 8650 3050 8700 3065
rect 8800 3535 8850 3550
rect 8800 3515 8815 3535
rect 8835 3515 8850 3535
rect 8800 3485 8850 3515
rect 8800 3465 8815 3485
rect 8835 3465 8850 3485
rect 8800 3435 8850 3465
rect 8800 3415 8815 3435
rect 8835 3415 8850 3435
rect 8800 3385 8850 3415
rect 8800 3365 8815 3385
rect 8835 3365 8850 3385
rect 8800 3335 8850 3365
rect 8800 3315 8815 3335
rect 8835 3315 8850 3335
rect 8800 3285 8850 3315
rect 8800 3265 8815 3285
rect 8835 3265 8850 3285
rect 8800 3235 8850 3265
rect 8800 3215 8815 3235
rect 8835 3215 8850 3235
rect 8800 3185 8850 3215
rect 8800 3165 8815 3185
rect 8835 3165 8850 3185
rect 8800 3135 8850 3165
rect 8800 3115 8815 3135
rect 8835 3115 8850 3135
rect 8800 3085 8850 3115
rect 8800 3065 8815 3085
rect 8835 3065 8850 3085
rect 8800 3050 8850 3065
rect 8950 3535 9000 3550
rect 8950 3515 8965 3535
rect 8985 3515 9000 3535
rect 8950 3485 9000 3515
rect 8950 3465 8965 3485
rect 8985 3465 9000 3485
rect 8950 3435 9000 3465
rect 8950 3415 8965 3435
rect 8985 3415 9000 3435
rect 8950 3385 9000 3415
rect 8950 3365 8965 3385
rect 8985 3365 9000 3385
rect 8950 3335 9000 3365
rect 8950 3315 8965 3335
rect 8985 3315 9000 3335
rect 8950 3285 9000 3315
rect 8950 3265 8965 3285
rect 8985 3265 9000 3285
rect 8950 3235 9000 3265
rect 8950 3215 8965 3235
rect 8985 3215 9000 3235
rect 8950 3185 9000 3215
rect 8950 3165 8965 3185
rect 8985 3165 9000 3185
rect 8950 3135 9000 3165
rect 8950 3115 8965 3135
rect 8985 3115 9000 3135
rect 8950 3085 9000 3115
rect 8950 3065 8965 3085
rect 8985 3065 9000 3085
rect 8950 3050 9000 3065
rect 9100 3535 9150 3550
rect 9100 3515 9115 3535
rect 9135 3515 9150 3535
rect 9100 3485 9150 3515
rect 9100 3465 9115 3485
rect 9135 3465 9150 3485
rect 9100 3435 9150 3465
rect 9100 3415 9115 3435
rect 9135 3415 9150 3435
rect 9100 3385 9150 3415
rect 9100 3365 9115 3385
rect 9135 3365 9150 3385
rect 9100 3335 9150 3365
rect 9100 3315 9115 3335
rect 9135 3315 9150 3335
rect 9100 3285 9150 3315
rect 9100 3265 9115 3285
rect 9135 3265 9150 3285
rect 9100 3235 9150 3265
rect 9100 3215 9115 3235
rect 9135 3215 9150 3235
rect 9100 3185 9150 3215
rect 9100 3165 9115 3185
rect 9135 3165 9150 3185
rect 9100 3135 9150 3165
rect 9100 3115 9115 3135
rect 9135 3115 9150 3135
rect 9100 3085 9150 3115
rect 9100 3065 9115 3085
rect 9135 3065 9150 3085
rect 9100 3050 9150 3065
rect 9250 3535 9300 3550
rect 9250 3515 9265 3535
rect 9285 3515 9300 3535
rect 9250 3485 9300 3515
rect 9250 3465 9265 3485
rect 9285 3465 9300 3485
rect 9250 3435 9300 3465
rect 9250 3415 9265 3435
rect 9285 3415 9300 3435
rect 9250 3385 9300 3415
rect 9250 3365 9265 3385
rect 9285 3365 9300 3385
rect 9250 3335 9300 3365
rect 9250 3315 9265 3335
rect 9285 3315 9300 3335
rect 9250 3285 9300 3315
rect 9250 3265 9265 3285
rect 9285 3265 9300 3285
rect 9250 3235 9300 3265
rect 9250 3215 9265 3235
rect 9285 3215 9300 3235
rect 9250 3185 9300 3215
rect 9250 3165 9265 3185
rect 9285 3165 9300 3185
rect 9250 3135 9300 3165
rect 9250 3115 9265 3135
rect 9285 3115 9300 3135
rect 9250 3085 9300 3115
rect 9250 3065 9265 3085
rect 9285 3065 9300 3085
rect 9250 3050 9300 3065
rect 9400 3535 9450 3550
rect 9400 3515 9415 3535
rect 9435 3515 9450 3535
rect 9400 3485 9450 3515
rect 9400 3465 9415 3485
rect 9435 3465 9450 3485
rect 9400 3435 9450 3465
rect 9400 3415 9415 3435
rect 9435 3415 9450 3435
rect 9400 3385 9450 3415
rect 9400 3365 9415 3385
rect 9435 3365 9450 3385
rect 9400 3335 9450 3365
rect 9400 3315 9415 3335
rect 9435 3315 9450 3335
rect 9400 3285 9450 3315
rect 9400 3265 9415 3285
rect 9435 3265 9450 3285
rect 9400 3235 9450 3265
rect 9400 3215 9415 3235
rect 9435 3215 9450 3235
rect 9400 3185 9450 3215
rect 9400 3165 9415 3185
rect 9435 3165 9450 3185
rect 9400 3135 9450 3165
rect 9400 3115 9415 3135
rect 9435 3115 9450 3135
rect 9400 3085 9450 3115
rect 9400 3065 9415 3085
rect 9435 3065 9450 3085
rect 9400 3050 9450 3065
rect 9550 3535 9600 3550
rect 9550 3515 9565 3535
rect 9585 3515 9600 3535
rect 9550 3485 9600 3515
rect 9550 3465 9565 3485
rect 9585 3465 9600 3485
rect 9550 3435 9600 3465
rect 9550 3415 9565 3435
rect 9585 3415 9600 3435
rect 9550 3385 9600 3415
rect 9550 3365 9565 3385
rect 9585 3365 9600 3385
rect 9550 3335 9600 3365
rect 9550 3315 9565 3335
rect 9585 3315 9600 3335
rect 9550 3285 9600 3315
rect 9550 3265 9565 3285
rect 9585 3265 9600 3285
rect 9550 3235 9600 3265
rect 9550 3215 9565 3235
rect 9585 3215 9600 3235
rect 9550 3185 9600 3215
rect 9550 3165 9565 3185
rect 9585 3165 9600 3185
rect 9550 3135 9600 3165
rect 9550 3115 9565 3135
rect 9585 3115 9600 3135
rect 9550 3085 9600 3115
rect 9550 3065 9565 3085
rect 9585 3065 9600 3085
rect 9550 3050 9600 3065
rect 9700 3535 9750 3550
rect 9700 3515 9715 3535
rect 9735 3515 9750 3535
rect 9700 3485 9750 3515
rect 9700 3465 9715 3485
rect 9735 3465 9750 3485
rect 9700 3435 9750 3465
rect 9700 3415 9715 3435
rect 9735 3415 9750 3435
rect 9700 3385 9750 3415
rect 9700 3365 9715 3385
rect 9735 3365 9750 3385
rect 9700 3335 9750 3365
rect 9700 3315 9715 3335
rect 9735 3315 9750 3335
rect 9700 3285 9750 3315
rect 9700 3265 9715 3285
rect 9735 3265 9750 3285
rect 9700 3235 9750 3265
rect 9700 3215 9715 3235
rect 9735 3215 9750 3235
rect 9700 3185 9750 3215
rect 9700 3165 9715 3185
rect 9735 3165 9750 3185
rect 9700 3135 9750 3165
rect 9700 3115 9715 3135
rect 9735 3115 9750 3135
rect 9700 3085 9750 3115
rect 9700 3065 9715 3085
rect 9735 3065 9750 3085
rect 9700 3050 9750 3065
rect 9850 3535 9900 3550
rect 9850 3515 9865 3535
rect 9885 3515 9900 3535
rect 9850 3485 9900 3515
rect 9850 3465 9865 3485
rect 9885 3465 9900 3485
rect 9850 3435 9900 3465
rect 9850 3415 9865 3435
rect 9885 3415 9900 3435
rect 9850 3385 9900 3415
rect 9850 3365 9865 3385
rect 9885 3365 9900 3385
rect 9850 3335 9900 3365
rect 9850 3315 9865 3335
rect 9885 3315 9900 3335
rect 9850 3285 9900 3315
rect 9850 3265 9865 3285
rect 9885 3265 9900 3285
rect 9850 3235 9900 3265
rect 9850 3215 9865 3235
rect 9885 3215 9900 3235
rect 9850 3185 9900 3215
rect 9850 3165 9865 3185
rect 9885 3165 9900 3185
rect 9850 3135 9900 3165
rect 9850 3115 9865 3135
rect 9885 3115 9900 3135
rect 9850 3085 9900 3115
rect 9850 3065 9865 3085
rect 9885 3065 9900 3085
rect 9850 3050 9900 3065
rect 10000 3535 10050 3550
rect 10000 3515 10015 3535
rect 10035 3515 10050 3535
rect 10000 3485 10050 3515
rect 10000 3465 10015 3485
rect 10035 3465 10050 3485
rect 10000 3435 10050 3465
rect 10000 3415 10015 3435
rect 10035 3415 10050 3435
rect 10000 3385 10050 3415
rect 10000 3365 10015 3385
rect 10035 3365 10050 3385
rect 10000 3335 10050 3365
rect 10000 3315 10015 3335
rect 10035 3315 10050 3335
rect 10000 3285 10050 3315
rect 10000 3265 10015 3285
rect 10035 3265 10050 3285
rect 10000 3235 10050 3265
rect 10000 3215 10015 3235
rect 10035 3215 10050 3235
rect 10000 3185 10050 3215
rect 10000 3165 10015 3185
rect 10035 3165 10050 3185
rect 10000 3135 10050 3165
rect 10000 3115 10015 3135
rect 10035 3115 10050 3135
rect 10000 3085 10050 3115
rect 10000 3065 10015 3085
rect 10035 3065 10050 3085
rect 10000 3050 10050 3065
rect 10150 3535 10200 3550
rect 10150 3515 10165 3535
rect 10185 3515 10200 3535
rect 10150 3485 10200 3515
rect 10150 3465 10165 3485
rect 10185 3465 10200 3485
rect 10150 3435 10200 3465
rect 10150 3415 10165 3435
rect 10185 3415 10200 3435
rect 10150 3385 10200 3415
rect 10150 3365 10165 3385
rect 10185 3365 10200 3385
rect 10150 3335 10200 3365
rect 10150 3315 10165 3335
rect 10185 3315 10200 3335
rect 10150 3285 10200 3315
rect 10150 3265 10165 3285
rect 10185 3265 10200 3285
rect 10150 3235 10200 3265
rect 10150 3215 10165 3235
rect 10185 3215 10200 3235
rect 10150 3185 10200 3215
rect 10150 3165 10165 3185
rect 10185 3165 10200 3185
rect 10150 3135 10200 3165
rect 10150 3115 10165 3135
rect 10185 3115 10200 3135
rect 10150 3085 10200 3115
rect 10150 3065 10165 3085
rect 10185 3065 10200 3085
rect 10150 3050 10200 3065
rect 10300 3535 10350 3550
rect 10300 3515 10315 3535
rect 10335 3515 10350 3535
rect 10300 3485 10350 3515
rect 10300 3465 10315 3485
rect 10335 3465 10350 3485
rect 10300 3435 10350 3465
rect 10300 3415 10315 3435
rect 10335 3415 10350 3435
rect 10300 3385 10350 3415
rect 10300 3365 10315 3385
rect 10335 3365 10350 3385
rect 10300 3335 10350 3365
rect 10300 3315 10315 3335
rect 10335 3315 10350 3335
rect 10300 3285 10350 3315
rect 10300 3265 10315 3285
rect 10335 3265 10350 3285
rect 10300 3235 10350 3265
rect 10300 3215 10315 3235
rect 10335 3215 10350 3235
rect 10300 3185 10350 3215
rect 10300 3165 10315 3185
rect 10335 3165 10350 3185
rect 10300 3135 10350 3165
rect 10300 3115 10315 3135
rect 10335 3115 10350 3135
rect 10300 3085 10350 3115
rect 10300 3065 10315 3085
rect 10335 3065 10350 3085
rect 10300 3050 10350 3065
rect 10450 3535 10500 3550
rect 10450 3515 10465 3535
rect 10485 3515 10500 3535
rect 10450 3485 10500 3515
rect 10450 3465 10465 3485
rect 10485 3465 10500 3485
rect 10450 3435 10500 3465
rect 10450 3415 10465 3435
rect 10485 3415 10500 3435
rect 10450 3385 10500 3415
rect 10450 3365 10465 3385
rect 10485 3365 10500 3385
rect 10450 3335 10500 3365
rect 10450 3315 10465 3335
rect 10485 3315 10500 3335
rect 10450 3285 10500 3315
rect 10450 3265 10465 3285
rect 10485 3265 10500 3285
rect 10450 3235 10500 3265
rect 10450 3215 10465 3235
rect 10485 3215 10500 3235
rect 10450 3185 10500 3215
rect 10450 3165 10465 3185
rect 10485 3165 10500 3185
rect 10450 3135 10500 3165
rect 10450 3115 10465 3135
rect 10485 3115 10500 3135
rect 10450 3085 10500 3115
rect 10450 3065 10465 3085
rect 10485 3065 10500 3085
rect 10450 3050 10500 3065
rect 10600 3535 10650 3550
rect 10600 3515 10615 3535
rect 10635 3515 10650 3535
rect 10600 3485 10650 3515
rect 10600 3465 10615 3485
rect 10635 3465 10650 3485
rect 10600 3435 10650 3465
rect 10600 3415 10615 3435
rect 10635 3415 10650 3435
rect 10600 3385 10650 3415
rect 10600 3365 10615 3385
rect 10635 3365 10650 3385
rect 10600 3335 10650 3365
rect 10600 3315 10615 3335
rect 10635 3315 10650 3335
rect 10600 3285 10650 3315
rect 10600 3265 10615 3285
rect 10635 3265 10650 3285
rect 10600 3235 10650 3265
rect 10600 3215 10615 3235
rect 10635 3215 10650 3235
rect 10600 3185 10650 3215
rect 10600 3165 10615 3185
rect 10635 3165 10650 3185
rect 10600 3135 10650 3165
rect 10600 3115 10615 3135
rect 10635 3115 10650 3135
rect 10600 3085 10650 3115
rect 10600 3065 10615 3085
rect 10635 3065 10650 3085
rect 10600 3050 10650 3065
rect 10750 3535 10800 3550
rect 10750 3515 10765 3535
rect 10785 3515 10800 3535
rect 10750 3485 10800 3515
rect 10750 3465 10765 3485
rect 10785 3465 10800 3485
rect 10750 3435 10800 3465
rect 10750 3415 10765 3435
rect 10785 3415 10800 3435
rect 10750 3385 10800 3415
rect 10750 3365 10765 3385
rect 10785 3365 10800 3385
rect 10750 3335 10800 3365
rect 10750 3315 10765 3335
rect 10785 3315 10800 3335
rect 10750 3285 10800 3315
rect 10750 3265 10765 3285
rect 10785 3265 10800 3285
rect 10750 3235 10800 3265
rect 10750 3215 10765 3235
rect 10785 3215 10800 3235
rect 10750 3185 10800 3215
rect 10750 3165 10765 3185
rect 10785 3165 10800 3185
rect 10750 3135 10800 3165
rect 10750 3115 10765 3135
rect 10785 3115 10800 3135
rect 10750 3085 10800 3115
rect 10750 3065 10765 3085
rect 10785 3065 10800 3085
rect 10750 3050 10800 3065
rect 10900 3050 10950 3550
rect 11050 3050 11100 3550
rect 11200 3050 11250 3550
rect 11350 3535 11400 3550
rect 11350 3515 11365 3535
rect 11385 3515 11400 3535
rect 11350 3485 11400 3515
rect 11350 3465 11365 3485
rect 11385 3465 11400 3485
rect 11350 3435 11400 3465
rect 11350 3415 11365 3435
rect 11385 3415 11400 3435
rect 11350 3385 11400 3415
rect 11350 3365 11365 3385
rect 11385 3365 11400 3385
rect 11350 3335 11400 3365
rect 11350 3315 11365 3335
rect 11385 3315 11400 3335
rect 11350 3285 11400 3315
rect 11350 3265 11365 3285
rect 11385 3265 11400 3285
rect 11350 3235 11400 3265
rect 11350 3215 11365 3235
rect 11385 3215 11400 3235
rect 11350 3185 11400 3215
rect 11350 3165 11365 3185
rect 11385 3165 11400 3185
rect 11350 3135 11400 3165
rect 11350 3115 11365 3135
rect 11385 3115 11400 3135
rect 11350 3085 11400 3115
rect 11350 3065 11365 3085
rect 11385 3065 11400 3085
rect 11350 3050 11400 3065
rect 11500 3050 11550 3550
rect 11650 3050 11700 3550
rect 11800 3050 11850 3550
rect 11950 3535 12000 3550
rect 11950 3515 11965 3535
rect 11985 3515 12000 3535
rect 11950 3485 12000 3515
rect 11950 3465 11965 3485
rect 11985 3465 12000 3485
rect 11950 3435 12000 3465
rect 11950 3415 11965 3435
rect 11985 3415 12000 3435
rect 11950 3385 12000 3415
rect 11950 3365 11965 3385
rect 11985 3365 12000 3385
rect 11950 3335 12000 3365
rect 11950 3315 11965 3335
rect 11985 3315 12000 3335
rect 11950 3285 12000 3315
rect 11950 3265 11965 3285
rect 11985 3265 12000 3285
rect 11950 3235 12000 3265
rect 11950 3215 11965 3235
rect 11985 3215 12000 3235
rect 11950 3185 12000 3215
rect 11950 3165 11965 3185
rect 11985 3165 12000 3185
rect 11950 3135 12000 3165
rect 11950 3115 11965 3135
rect 11985 3115 12000 3135
rect 11950 3085 12000 3115
rect 11950 3065 11965 3085
rect 11985 3065 12000 3085
rect 11950 3050 12000 3065
rect 12100 3050 12150 3550
rect 12250 3050 12300 3550
rect 12400 3050 12450 3550
rect 12550 3535 12600 3550
rect 12550 3515 12565 3535
rect 12585 3515 12600 3535
rect 12550 3485 12600 3515
rect 12550 3465 12565 3485
rect 12585 3465 12600 3485
rect 12550 3435 12600 3465
rect 12550 3415 12565 3435
rect 12585 3415 12600 3435
rect 12550 3385 12600 3415
rect 12550 3365 12565 3385
rect 12585 3365 12600 3385
rect 12550 3335 12600 3365
rect 12550 3315 12565 3335
rect 12585 3315 12600 3335
rect 12550 3285 12600 3315
rect 12550 3265 12565 3285
rect 12585 3265 12600 3285
rect 12550 3235 12600 3265
rect 12550 3215 12565 3235
rect 12585 3215 12600 3235
rect 12550 3185 12600 3215
rect 12550 3165 12565 3185
rect 12585 3165 12600 3185
rect 12550 3135 12600 3165
rect 12550 3115 12565 3135
rect 12585 3115 12600 3135
rect 12550 3085 12600 3115
rect 12550 3065 12565 3085
rect 12585 3065 12600 3085
rect 12550 3050 12600 3065
rect 12700 3050 12750 3550
rect 12850 3050 12900 3550
rect 13000 3050 13050 3550
rect 13150 3535 13200 3550
rect 13150 3515 13165 3535
rect 13185 3515 13200 3535
rect 13150 3485 13200 3515
rect 13150 3465 13165 3485
rect 13185 3465 13200 3485
rect 13150 3435 13200 3465
rect 13150 3415 13165 3435
rect 13185 3415 13200 3435
rect 13150 3385 13200 3415
rect 13150 3365 13165 3385
rect 13185 3365 13200 3385
rect 13150 3335 13200 3365
rect 13150 3315 13165 3335
rect 13185 3315 13200 3335
rect 13150 3285 13200 3315
rect 13150 3265 13165 3285
rect 13185 3265 13200 3285
rect 13150 3235 13200 3265
rect 13150 3215 13165 3235
rect 13185 3215 13200 3235
rect 13150 3185 13200 3215
rect 13150 3165 13165 3185
rect 13185 3165 13200 3185
rect 13150 3135 13200 3165
rect 13150 3115 13165 3135
rect 13185 3115 13200 3135
rect 13150 3085 13200 3115
rect 13150 3065 13165 3085
rect 13185 3065 13200 3085
rect 13150 3050 13200 3065
rect 13300 3050 13350 3550
rect 13450 3050 13500 3550
rect 13600 3050 13650 3550
rect 13750 3535 13800 3550
rect 13750 3515 13765 3535
rect 13785 3515 13800 3535
rect 13750 3485 13800 3515
rect 13750 3465 13765 3485
rect 13785 3465 13800 3485
rect 13750 3435 13800 3465
rect 13750 3415 13765 3435
rect 13785 3415 13800 3435
rect 13750 3385 13800 3415
rect 13750 3365 13765 3385
rect 13785 3365 13800 3385
rect 13750 3335 13800 3365
rect 13750 3315 13765 3335
rect 13785 3315 13800 3335
rect 13750 3285 13800 3315
rect 13750 3265 13765 3285
rect 13785 3265 13800 3285
rect 13750 3235 13800 3265
rect 13750 3215 13765 3235
rect 13785 3215 13800 3235
rect 13750 3185 13800 3215
rect 13750 3165 13765 3185
rect 13785 3165 13800 3185
rect 13750 3135 13800 3165
rect 13750 3115 13765 3135
rect 13785 3115 13800 3135
rect 13750 3085 13800 3115
rect 13750 3065 13765 3085
rect 13785 3065 13800 3085
rect 13750 3050 13800 3065
rect 13900 3050 13950 3550
rect 14050 3050 14100 3550
rect 14200 3050 14250 3550
rect 14350 3535 14400 3550
rect 14350 3515 14365 3535
rect 14385 3515 14400 3535
rect 14350 3485 14400 3515
rect 14350 3465 14365 3485
rect 14385 3465 14400 3485
rect 14350 3435 14400 3465
rect 14350 3415 14365 3435
rect 14385 3415 14400 3435
rect 14350 3385 14400 3415
rect 14350 3365 14365 3385
rect 14385 3365 14400 3385
rect 14350 3335 14400 3365
rect 14350 3315 14365 3335
rect 14385 3315 14400 3335
rect 14350 3285 14400 3315
rect 14350 3265 14365 3285
rect 14385 3265 14400 3285
rect 14350 3235 14400 3265
rect 14350 3215 14365 3235
rect 14385 3215 14400 3235
rect 14350 3185 14400 3215
rect 14350 3165 14365 3185
rect 14385 3165 14400 3185
rect 14350 3135 14400 3165
rect 14350 3115 14365 3135
rect 14385 3115 14400 3135
rect 14350 3085 14400 3115
rect 14350 3065 14365 3085
rect 14385 3065 14400 3085
rect 14350 3050 14400 3065
rect 14500 3050 14550 3550
rect 14650 3050 14700 3550
rect 14800 3050 14850 3550
rect 14950 3535 15000 3550
rect 14950 3515 14965 3535
rect 14985 3515 15000 3535
rect 14950 3485 15000 3515
rect 14950 3465 14965 3485
rect 14985 3465 15000 3485
rect 14950 3435 15000 3465
rect 14950 3415 14965 3435
rect 14985 3415 15000 3435
rect 14950 3385 15000 3415
rect 14950 3365 14965 3385
rect 14985 3365 15000 3385
rect 14950 3335 15000 3365
rect 14950 3315 14965 3335
rect 14985 3315 15000 3335
rect 14950 3285 15000 3315
rect 14950 3265 14965 3285
rect 14985 3265 15000 3285
rect 14950 3235 15000 3265
rect 14950 3215 14965 3235
rect 14985 3215 15000 3235
rect 14950 3185 15000 3215
rect 14950 3165 14965 3185
rect 14985 3165 15000 3185
rect 14950 3135 15000 3165
rect 14950 3115 14965 3135
rect 14985 3115 15000 3135
rect 14950 3085 15000 3115
rect 14950 3065 14965 3085
rect 14985 3065 15000 3085
rect 14950 3050 15000 3065
rect 15100 3050 15150 3550
rect 15250 3050 15300 3550
rect 15400 3050 15450 3550
rect 15550 3535 15600 3550
rect 15550 3515 15565 3535
rect 15585 3515 15600 3535
rect 15550 3485 15600 3515
rect 15550 3465 15565 3485
rect 15585 3465 15600 3485
rect 15550 3435 15600 3465
rect 15550 3415 15565 3435
rect 15585 3415 15600 3435
rect 15550 3385 15600 3415
rect 15550 3365 15565 3385
rect 15585 3365 15600 3385
rect 15550 3335 15600 3365
rect 15550 3315 15565 3335
rect 15585 3315 15600 3335
rect 15550 3285 15600 3315
rect 15550 3265 15565 3285
rect 15585 3265 15600 3285
rect 15550 3235 15600 3265
rect 15550 3215 15565 3235
rect 15585 3215 15600 3235
rect 15550 3185 15600 3215
rect 15550 3165 15565 3185
rect 15585 3165 15600 3185
rect 15550 3135 15600 3165
rect 15550 3115 15565 3135
rect 15585 3115 15600 3135
rect 15550 3085 15600 3115
rect 15550 3065 15565 3085
rect 15585 3065 15600 3085
rect 15550 3050 15600 3065
rect 15700 3050 15750 3550
rect 15850 3050 15900 3550
rect 16000 3050 16050 3550
rect 16150 3535 16200 3550
rect 16150 3515 16165 3535
rect 16185 3515 16200 3535
rect 16150 3485 16200 3515
rect 16150 3465 16165 3485
rect 16185 3465 16200 3485
rect 16150 3435 16200 3465
rect 16150 3415 16165 3435
rect 16185 3415 16200 3435
rect 16150 3385 16200 3415
rect 16150 3365 16165 3385
rect 16185 3365 16200 3385
rect 16150 3335 16200 3365
rect 16150 3315 16165 3335
rect 16185 3315 16200 3335
rect 16150 3285 16200 3315
rect 16150 3265 16165 3285
rect 16185 3265 16200 3285
rect 16150 3235 16200 3265
rect 16150 3215 16165 3235
rect 16185 3215 16200 3235
rect 16150 3185 16200 3215
rect 16150 3165 16165 3185
rect 16185 3165 16200 3185
rect 16150 3135 16200 3165
rect 16150 3115 16165 3135
rect 16185 3115 16200 3135
rect 16150 3085 16200 3115
rect 16150 3065 16165 3085
rect 16185 3065 16200 3085
rect 16150 3050 16200 3065
rect 16300 3535 16350 3550
rect 16300 3515 16315 3535
rect 16335 3515 16350 3535
rect 16300 3485 16350 3515
rect 16300 3465 16315 3485
rect 16335 3465 16350 3485
rect 16300 3435 16350 3465
rect 16300 3415 16315 3435
rect 16335 3415 16350 3435
rect 16300 3385 16350 3415
rect 16300 3365 16315 3385
rect 16335 3365 16350 3385
rect 16300 3335 16350 3365
rect 16300 3315 16315 3335
rect 16335 3315 16350 3335
rect 16300 3285 16350 3315
rect 16300 3265 16315 3285
rect 16335 3265 16350 3285
rect 16300 3235 16350 3265
rect 16300 3215 16315 3235
rect 16335 3215 16350 3235
rect 16300 3185 16350 3215
rect 16300 3165 16315 3185
rect 16335 3165 16350 3185
rect 16300 3135 16350 3165
rect 16300 3115 16315 3135
rect 16335 3115 16350 3135
rect 16300 3085 16350 3115
rect 16300 3065 16315 3085
rect 16335 3065 16350 3085
rect 16300 3050 16350 3065
rect 16450 3535 16500 3550
rect 16450 3515 16465 3535
rect 16485 3515 16500 3535
rect 16450 3485 16500 3515
rect 16450 3465 16465 3485
rect 16485 3465 16500 3485
rect 16450 3435 16500 3465
rect 16450 3415 16465 3435
rect 16485 3415 16500 3435
rect 16450 3385 16500 3415
rect 16450 3365 16465 3385
rect 16485 3365 16500 3385
rect 16450 3335 16500 3365
rect 16450 3315 16465 3335
rect 16485 3315 16500 3335
rect 16450 3285 16500 3315
rect 16450 3265 16465 3285
rect 16485 3265 16500 3285
rect 16450 3235 16500 3265
rect 16450 3215 16465 3235
rect 16485 3215 16500 3235
rect 16450 3185 16500 3215
rect 16450 3165 16465 3185
rect 16485 3165 16500 3185
rect 16450 3135 16500 3165
rect 16450 3115 16465 3135
rect 16485 3115 16500 3135
rect 16450 3085 16500 3115
rect 16450 3065 16465 3085
rect 16485 3065 16500 3085
rect 16450 3050 16500 3065
rect 16600 3535 16650 3550
rect 16600 3515 16615 3535
rect 16635 3515 16650 3535
rect 16600 3485 16650 3515
rect 16600 3465 16615 3485
rect 16635 3465 16650 3485
rect 16600 3435 16650 3465
rect 16600 3415 16615 3435
rect 16635 3415 16650 3435
rect 16600 3385 16650 3415
rect 16600 3365 16615 3385
rect 16635 3365 16650 3385
rect 16600 3335 16650 3365
rect 16600 3315 16615 3335
rect 16635 3315 16650 3335
rect 16600 3285 16650 3315
rect 16600 3265 16615 3285
rect 16635 3265 16650 3285
rect 16600 3235 16650 3265
rect 16600 3215 16615 3235
rect 16635 3215 16650 3235
rect 16600 3185 16650 3215
rect 16600 3165 16615 3185
rect 16635 3165 16650 3185
rect 16600 3135 16650 3165
rect 16600 3115 16615 3135
rect 16635 3115 16650 3135
rect 16600 3085 16650 3115
rect 16600 3065 16615 3085
rect 16635 3065 16650 3085
rect 16600 3050 16650 3065
rect 16750 3535 16800 3550
rect 16750 3515 16765 3535
rect 16785 3515 16800 3535
rect 16750 3485 16800 3515
rect 16750 3465 16765 3485
rect 16785 3465 16800 3485
rect 16750 3435 16800 3465
rect 16750 3415 16765 3435
rect 16785 3415 16800 3435
rect 16750 3385 16800 3415
rect 16750 3365 16765 3385
rect 16785 3365 16800 3385
rect 16750 3335 16800 3365
rect 16750 3315 16765 3335
rect 16785 3315 16800 3335
rect 16750 3285 16800 3315
rect 16750 3265 16765 3285
rect 16785 3265 16800 3285
rect 16750 3235 16800 3265
rect 16750 3215 16765 3235
rect 16785 3215 16800 3235
rect 16750 3185 16800 3215
rect 16750 3165 16765 3185
rect 16785 3165 16800 3185
rect 16750 3135 16800 3165
rect 16750 3115 16765 3135
rect 16785 3115 16800 3135
rect 16750 3085 16800 3115
rect 16750 3065 16765 3085
rect 16785 3065 16800 3085
rect 16750 3050 16800 3065
rect 16900 3535 16950 3550
rect 16900 3515 16915 3535
rect 16935 3515 16950 3535
rect 16900 3485 16950 3515
rect 16900 3465 16915 3485
rect 16935 3465 16950 3485
rect 16900 3435 16950 3465
rect 16900 3415 16915 3435
rect 16935 3415 16950 3435
rect 16900 3385 16950 3415
rect 16900 3365 16915 3385
rect 16935 3365 16950 3385
rect 16900 3335 16950 3365
rect 16900 3315 16915 3335
rect 16935 3315 16950 3335
rect 16900 3285 16950 3315
rect 16900 3265 16915 3285
rect 16935 3265 16950 3285
rect 16900 3235 16950 3265
rect 16900 3215 16915 3235
rect 16935 3215 16950 3235
rect 16900 3185 16950 3215
rect 16900 3165 16915 3185
rect 16935 3165 16950 3185
rect 16900 3135 16950 3165
rect 16900 3115 16915 3135
rect 16935 3115 16950 3135
rect 16900 3085 16950 3115
rect 16900 3065 16915 3085
rect 16935 3065 16950 3085
rect 16900 3050 16950 3065
rect 17050 3535 17100 3550
rect 17050 3515 17065 3535
rect 17085 3515 17100 3535
rect 17050 3485 17100 3515
rect 17050 3465 17065 3485
rect 17085 3465 17100 3485
rect 17050 3435 17100 3465
rect 17050 3415 17065 3435
rect 17085 3415 17100 3435
rect 17050 3385 17100 3415
rect 17050 3365 17065 3385
rect 17085 3365 17100 3385
rect 17050 3335 17100 3365
rect 17050 3315 17065 3335
rect 17085 3315 17100 3335
rect 17050 3285 17100 3315
rect 17050 3265 17065 3285
rect 17085 3265 17100 3285
rect 17050 3235 17100 3265
rect 17050 3215 17065 3235
rect 17085 3215 17100 3235
rect 17050 3185 17100 3215
rect 17050 3165 17065 3185
rect 17085 3165 17100 3185
rect 17050 3135 17100 3165
rect 17050 3115 17065 3135
rect 17085 3115 17100 3135
rect 17050 3085 17100 3115
rect 17050 3065 17065 3085
rect 17085 3065 17100 3085
rect 17050 3050 17100 3065
rect 17200 3535 17250 3550
rect 17200 3515 17215 3535
rect 17235 3515 17250 3535
rect 17200 3485 17250 3515
rect 17200 3465 17215 3485
rect 17235 3465 17250 3485
rect 17200 3435 17250 3465
rect 17200 3415 17215 3435
rect 17235 3415 17250 3435
rect 17200 3385 17250 3415
rect 17200 3365 17215 3385
rect 17235 3365 17250 3385
rect 17200 3335 17250 3365
rect 17200 3315 17215 3335
rect 17235 3315 17250 3335
rect 17200 3285 17250 3315
rect 17200 3265 17215 3285
rect 17235 3265 17250 3285
rect 17200 3235 17250 3265
rect 17200 3215 17215 3235
rect 17235 3215 17250 3235
rect 17200 3185 17250 3215
rect 17200 3165 17215 3185
rect 17235 3165 17250 3185
rect 17200 3135 17250 3165
rect 17200 3115 17215 3135
rect 17235 3115 17250 3135
rect 17200 3085 17250 3115
rect 17200 3065 17215 3085
rect 17235 3065 17250 3085
rect 17200 3050 17250 3065
rect 17350 3535 17400 3550
rect 17350 3515 17365 3535
rect 17385 3515 17400 3535
rect 17350 3485 17400 3515
rect 17350 3465 17365 3485
rect 17385 3465 17400 3485
rect 17350 3435 17400 3465
rect 17350 3415 17365 3435
rect 17385 3415 17400 3435
rect 17350 3385 17400 3415
rect 17350 3365 17365 3385
rect 17385 3365 17400 3385
rect 17350 3335 17400 3365
rect 17350 3315 17365 3335
rect 17385 3315 17400 3335
rect 17350 3285 17400 3315
rect 17350 3265 17365 3285
rect 17385 3265 17400 3285
rect 17350 3235 17400 3265
rect 17350 3215 17365 3235
rect 17385 3215 17400 3235
rect 17350 3185 17400 3215
rect 17350 3165 17365 3185
rect 17385 3165 17400 3185
rect 17350 3135 17400 3165
rect 17350 3115 17365 3135
rect 17385 3115 17400 3135
rect 17350 3085 17400 3115
rect 17350 3065 17365 3085
rect 17385 3065 17400 3085
rect 17350 3050 17400 3065
rect 17500 3050 17550 3550
rect 17650 3050 17700 3550
rect 17800 3050 17850 3550
rect 17950 3535 18000 3550
rect 17950 3515 17965 3535
rect 17985 3515 18000 3535
rect 17950 3485 18000 3515
rect 17950 3465 17965 3485
rect 17985 3465 18000 3485
rect 17950 3435 18000 3465
rect 17950 3415 17965 3435
rect 17985 3415 18000 3435
rect 17950 3385 18000 3415
rect 17950 3365 17965 3385
rect 17985 3365 18000 3385
rect 17950 3335 18000 3365
rect 17950 3315 17965 3335
rect 17985 3315 18000 3335
rect 17950 3285 18000 3315
rect 17950 3265 17965 3285
rect 17985 3265 18000 3285
rect 17950 3235 18000 3265
rect 17950 3215 17965 3235
rect 17985 3215 18000 3235
rect 17950 3185 18000 3215
rect 17950 3165 17965 3185
rect 17985 3165 18000 3185
rect 17950 3135 18000 3165
rect 17950 3115 17965 3135
rect 17985 3115 18000 3135
rect 17950 3085 18000 3115
rect 17950 3065 17965 3085
rect 17985 3065 18000 3085
rect 17950 3050 18000 3065
rect 18100 3050 18150 3550
rect 18250 3050 18300 3550
rect 18400 3050 18450 3550
rect 18550 3535 18600 3550
rect 18550 3515 18565 3535
rect 18585 3515 18600 3535
rect 18550 3485 18600 3515
rect 18550 3465 18565 3485
rect 18585 3465 18600 3485
rect 18550 3435 18600 3465
rect 18550 3415 18565 3435
rect 18585 3415 18600 3435
rect 18550 3385 18600 3415
rect 18550 3365 18565 3385
rect 18585 3365 18600 3385
rect 18550 3335 18600 3365
rect 18550 3315 18565 3335
rect 18585 3315 18600 3335
rect 18550 3285 18600 3315
rect 18550 3265 18565 3285
rect 18585 3265 18600 3285
rect 18550 3235 18600 3265
rect 18550 3215 18565 3235
rect 18585 3215 18600 3235
rect 18550 3185 18600 3215
rect 18550 3165 18565 3185
rect 18585 3165 18600 3185
rect 18550 3135 18600 3165
rect 18550 3115 18565 3135
rect 18585 3115 18600 3135
rect 18550 3085 18600 3115
rect 18550 3065 18565 3085
rect 18585 3065 18600 3085
rect 18550 3050 18600 3065
rect 18700 3535 18750 3550
rect 18700 3515 18715 3535
rect 18735 3515 18750 3535
rect 18700 3485 18750 3515
rect 18700 3465 18715 3485
rect 18735 3465 18750 3485
rect 18700 3435 18750 3465
rect 18700 3415 18715 3435
rect 18735 3415 18750 3435
rect 18700 3385 18750 3415
rect 18700 3365 18715 3385
rect 18735 3365 18750 3385
rect 18700 3335 18750 3365
rect 18700 3315 18715 3335
rect 18735 3315 18750 3335
rect 18700 3285 18750 3315
rect 18700 3265 18715 3285
rect 18735 3265 18750 3285
rect 18700 3235 18750 3265
rect 18700 3215 18715 3235
rect 18735 3215 18750 3235
rect 18700 3185 18750 3215
rect 18700 3165 18715 3185
rect 18735 3165 18750 3185
rect 18700 3135 18750 3165
rect 18700 3115 18715 3135
rect 18735 3115 18750 3135
rect 18700 3085 18750 3115
rect 18700 3065 18715 3085
rect 18735 3065 18750 3085
rect 18700 3050 18750 3065
rect 18850 3535 18900 3550
rect 18850 3515 18865 3535
rect 18885 3515 18900 3535
rect 18850 3485 18900 3515
rect 18850 3465 18865 3485
rect 18885 3465 18900 3485
rect 18850 3435 18900 3465
rect 18850 3415 18865 3435
rect 18885 3415 18900 3435
rect 18850 3385 18900 3415
rect 18850 3365 18865 3385
rect 18885 3365 18900 3385
rect 18850 3335 18900 3365
rect 18850 3315 18865 3335
rect 18885 3315 18900 3335
rect 18850 3285 18900 3315
rect 18850 3265 18865 3285
rect 18885 3265 18900 3285
rect 18850 3235 18900 3265
rect 18850 3215 18865 3235
rect 18885 3215 18900 3235
rect 18850 3185 18900 3215
rect 18850 3165 18865 3185
rect 18885 3165 18900 3185
rect 18850 3135 18900 3165
rect 18850 3115 18865 3135
rect 18885 3115 18900 3135
rect 18850 3085 18900 3115
rect 18850 3065 18865 3085
rect 18885 3065 18900 3085
rect 18850 3050 18900 3065
rect 19000 3535 19050 3550
rect 19000 3515 19015 3535
rect 19035 3515 19050 3535
rect 19000 3485 19050 3515
rect 19000 3465 19015 3485
rect 19035 3465 19050 3485
rect 19000 3435 19050 3465
rect 19000 3415 19015 3435
rect 19035 3415 19050 3435
rect 19000 3385 19050 3415
rect 19000 3365 19015 3385
rect 19035 3365 19050 3385
rect 19000 3335 19050 3365
rect 19000 3315 19015 3335
rect 19035 3315 19050 3335
rect 19000 3285 19050 3315
rect 19000 3265 19015 3285
rect 19035 3265 19050 3285
rect 19000 3235 19050 3265
rect 19000 3215 19015 3235
rect 19035 3215 19050 3235
rect 19000 3185 19050 3215
rect 19000 3165 19015 3185
rect 19035 3165 19050 3185
rect 19000 3135 19050 3165
rect 19000 3115 19015 3135
rect 19035 3115 19050 3135
rect 19000 3085 19050 3115
rect 19000 3065 19015 3085
rect 19035 3065 19050 3085
rect 19000 3050 19050 3065
rect 19150 3535 19200 3550
rect 19150 3515 19165 3535
rect 19185 3515 19200 3535
rect 19150 3485 19200 3515
rect 19150 3465 19165 3485
rect 19185 3465 19200 3485
rect 19150 3435 19200 3465
rect 19150 3415 19165 3435
rect 19185 3415 19200 3435
rect 19150 3385 19200 3415
rect 19150 3365 19165 3385
rect 19185 3365 19200 3385
rect 19150 3335 19200 3365
rect 19150 3315 19165 3335
rect 19185 3315 19200 3335
rect 19150 3285 19200 3315
rect 19150 3265 19165 3285
rect 19185 3265 19200 3285
rect 19150 3235 19200 3265
rect 19150 3215 19165 3235
rect 19185 3215 19200 3235
rect 19150 3185 19200 3215
rect 19150 3165 19165 3185
rect 19185 3165 19200 3185
rect 19150 3135 19200 3165
rect 19150 3115 19165 3135
rect 19185 3115 19200 3135
rect 19150 3085 19200 3115
rect 19150 3065 19165 3085
rect 19185 3065 19200 3085
rect 19150 3050 19200 3065
rect 19300 3535 19350 3550
rect 19300 3515 19315 3535
rect 19335 3515 19350 3535
rect 19300 3485 19350 3515
rect 19300 3465 19315 3485
rect 19335 3465 19350 3485
rect 19300 3435 19350 3465
rect 19300 3415 19315 3435
rect 19335 3415 19350 3435
rect 19300 3385 19350 3415
rect 19300 3365 19315 3385
rect 19335 3365 19350 3385
rect 19300 3335 19350 3365
rect 19300 3315 19315 3335
rect 19335 3315 19350 3335
rect 19300 3285 19350 3315
rect 19300 3265 19315 3285
rect 19335 3265 19350 3285
rect 19300 3235 19350 3265
rect 19300 3215 19315 3235
rect 19335 3215 19350 3235
rect 19300 3185 19350 3215
rect 19300 3165 19315 3185
rect 19335 3165 19350 3185
rect 19300 3135 19350 3165
rect 19300 3115 19315 3135
rect 19335 3115 19350 3135
rect 19300 3085 19350 3115
rect 19300 3065 19315 3085
rect 19335 3065 19350 3085
rect 19300 3050 19350 3065
rect 19450 3535 19500 3550
rect 19450 3515 19465 3535
rect 19485 3515 19500 3535
rect 19450 3485 19500 3515
rect 19450 3465 19465 3485
rect 19485 3465 19500 3485
rect 19450 3435 19500 3465
rect 19450 3415 19465 3435
rect 19485 3415 19500 3435
rect 19450 3385 19500 3415
rect 19450 3365 19465 3385
rect 19485 3365 19500 3385
rect 19450 3335 19500 3365
rect 19450 3315 19465 3335
rect 19485 3315 19500 3335
rect 19450 3285 19500 3315
rect 19450 3265 19465 3285
rect 19485 3265 19500 3285
rect 19450 3235 19500 3265
rect 19450 3215 19465 3235
rect 19485 3215 19500 3235
rect 19450 3185 19500 3215
rect 19450 3165 19465 3185
rect 19485 3165 19500 3185
rect 19450 3135 19500 3165
rect 19450 3115 19465 3135
rect 19485 3115 19500 3135
rect 19450 3085 19500 3115
rect 19450 3065 19465 3085
rect 19485 3065 19500 3085
rect 19450 3050 19500 3065
rect 19600 3535 19650 3550
rect 19600 3515 19615 3535
rect 19635 3515 19650 3535
rect 19600 3485 19650 3515
rect 19600 3465 19615 3485
rect 19635 3465 19650 3485
rect 19600 3435 19650 3465
rect 19600 3415 19615 3435
rect 19635 3415 19650 3435
rect 19600 3385 19650 3415
rect 19600 3365 19615 3385
rect 19635 3365 19650 3385
rect 19600 3335 19650 3365
rect 19600 3315 19615 3335
rect 19635 3315 19650 3335
rect 19600 3285 19650 3315
rect 19600 3265 19615 3285
rect 19635 3265 19650 3285
rect 19600 3235 19650 3265
rect 19600 3215 19615 3235
rect 19635 3215 19650 3235
rect 19600 3185 19650 3215
rect 19600 3165 19615 3185
rect 19635 3165 19650 3185
rect 19600 3135 19650 3165
rect 19600 3115 19615 3135
rect 19635 3115 19650 3135
rect 19600 3085 19650 3115
rect 19600 3065 19615 3085
rect 19635 3065 19650 3085
rect 19600 3050 19650 3065
rect 19750 3535 19800 3550
rect 19750 3515 19765 3535
rect 19785 3515 19800 3535
rect 19750 3485 19800 3515
rect 19750 3465 19765 3485
rect 19785 3465 19800 3485
rect 19750 3435 19800 3465
rect 19750 3415 19765 3435
rect 19785 3415 19800 3435
rect 19750 3385 19800 3415
rect 19750 3365 19765 3385
rect 19785 3365 19800 3385
rect 19750 3335 19800 3365
rect 19750 3315 19765 3335
rect 19785 3315 19800 3335
rect 19750 3285 19800 3315
rect 19750 3265 19765 3285
rect 19785 3265 19800 3285
rect 19750 3235 19800 3265
rect 19750 3215 19765 3235
rect 19785 3215 19800 3235
rect 19750 3185 19800 3215
rect 19750 3165 19765 3185
rect 19785 3165 19800 3185
rect 19750 3135 19800 3165
rect 19750 3115 19765 3135
rect 19785 3115 19800 3135
rect 19750 3085 19800 3115
rect 19750 3065 19765 3085
rect 19785 3065 19800 3085
rect 19750 3050 19800 3065
rect 19900 3050 19950 3550
rect 20050 3050 20100 3550
rect 20200 3050 20250 3550
rect 20350 3535 20400 3550
rect 20350 3515 20365 3535
rect 20385 3515 20400 3535
rect 20350 3485 20400 3515
rect 20350 3465 20365 3485
rect 20385 3465 20400 3485
rect 20350 3435 20400 3465
rect 20350 3415 20365 3435
rect 20385 3415 20400 3435
rect 20350 3385 20400 3415
rect 20350 3365 20365 3385
rect 20385 3365 20400 3385
rect 20350 3335 20400 3365
rect 20350 3315 20365 3335
rect 20385 3315 20400 3335
rect 20350 3285 20400 3315
rect 20350 3265 20365 3285
rect 20385 3265 20400 3285
rect 20350 3235 20400 3265
rect 20350 3215 20365 3235
rect 20385 3215 20400 3235
rect 20350 3185 20400 3215
rect 20350 3165 20365 3185
rect 20385 3165 20400 3185
rect 20350 3135 20400 3165
rect 20350 3115 20365 3135
rect 20385 3115 20400 3135
rect 20350 3085 20400 3115
rect 20350 3065 20365 3085
rect 20385 3065 20400 3085
rect 20350 3050 20400 3065
rect 20500 3050 20550 3550
rect 20650 3050 20700 3550
rect 20800 3050 20850 3550
rect 20950 3535 21000 3550
rect 20950 3515 20965 3535
rect 20985 3515 21000 3535
rect 20950 3485 21000 3515
rect 20950 3465 20965 3485
rect 20985 3465 21000 3485
rect 20950 3435 21000 3465
rect 20950 3415 20965 3435
rect 20985 3415 21000 3435
rect 20950 3385 21000 3415
rect 20950 3365 20965 3385
rect 20985 3365 21000 3385
rect 20950 3335 21000 3365
rect 20950 3315 20965 3335
rect 20985 3315 21000 3335
rect 20950 3285 21000 3315
rect 20950 3265 20965 3285
rect 20985 3265 21000 3285
rect 20950 3235 21000 3265
rect 20950 3215 20965 3235
rect 20985 3215 21000 3235
rect 20950 3185 21000 3215
rect 20950 3165 20965 3185
rect 20985 3165 21000 3185
rect 20950 3135 21000 3165
rect 20950 3115 20965 3135
rect 20985 3115 21000 3135
rect 20950 3085 21000 3115
rect 20950 3065 20965 3085
rect 20985 3065 21000 3085
rect 20950 3050 21000 3065
rect 21100 3050 21150 3550
rect 21250 3050 21300 3550
rect 21400 3535 21450 3550
rect 21400 3515 21415 3535
rect 21435 3515 21450 3535
rect 21400 3485 21450 3515
rect 21400 3465 21415 3485
rect 21435 3465 21450 3485
rect 21400 3435 21450 3465
rect 21400 3415 21415 3435
rect 21435 3415 21450 3435
rect 21400 3385 21450 3415
rect 21400 3365 21415 3385
rect 21435 3365 21450 3385
rect 21400 3335 21450 3365
rect 21400 3315 21415 3335
rect 21435 3315 21450 3335
rect 21400 3285 21450 3315
rect 21400 3265 21415 3285
rect 21435 3265 21450 3285
rect 21400 3235 21450 3265
rect 21400 3215 21415 3235
rect 21435 3215 21450 3235
rect 21400 3185 21450 3215
rect 21400 3165 21415 3185
rect 21435 3165 21450 3185
rect 21400 3135 21450 3165
rect 21400 3115 21415 3135
rect 21435 3115 21450 3135
rect 21400 3085 21450 3115
rect 21400 3065 21415 3085
rect 21435 3065 21450 3085
rect 21400 3050 21450 3065
rect 21550 3050 21600 3550
rect 21700 3050 21750 3550
rect 21850 3535 21900 3550
rect 21850 3515 21865 3535
rect 21885 3515 21900 3535
rect 21850 3485 21900 3515
rect 21850 3465 21865 3485
rect 21885 3465 21900 3485
rect 21850 3435 21900 3465
rect 21850 3415 21865 3435
rect 21885 3415 21900 3435
rect 21850 3385 21900 3415
rect 21850 3365 21865 3385
rect 21885 3365 21900 3385
rect 21850 3335 21900 3365
rect 21850 3315 21865 3335
rect 21885 3315 21900 3335
rect 21850 3285 21900 3315
rect 21850 3265 21865 3285
rect 21885 3265 21900 3285
rect 21850 3235 21900 3265
rect 21850 3215 21865 3235
rect 21885 3215 21900 3235
rect 21850 3185 21900 3215
rect 21850 3165 21865 3185
rect 21885 3165 21900 3185
rect 21850 3135 21900 3165
rect 21850 3115 21865 3135
rect 21885 3115 21900 3135
rect 21850 3085 21900 3115
rect 21850 3065 21865 3085
rect 21885 3065 21900 3085
rect 21850 3050 21900 3065
rect 22000 3050 22050 3550
rect 22150 3050 22200 3550
rect 22300 3050 22350 3550
rect 22450 3535 22500 3550
rect 22450 3515 22465 3535
rect 22485 3515 22500 3535
rect 22450 3485 22500 3515
rect 22450 3465 22465 3485
rect 22485 3465 22500 3485
rect 22450 3435 22500 3465
rect 22450 3415 22465 3435
rect 22485 3415 22500 3435
rect 22450 3385 22500 3415
rect 22450 3365 22465 3385
rect 22485 3365 22500 3385
rect 22450 3335 22500 3365
rect 22450 3315 22465 3335
rect 22485 3315 22500 3335
rect 22450 3285 22500 3315
rect 22450 3265 22465 3285
rect 22485 3265 22500 3285
rect 22450 3235 22500 3265
rect 22450 3215 22465 3235
rect 22485 3215 22500 3235
rect 22450 3185 22500 3215
rect 22450 3165 22465 3185
rect 22485 3165 22500 3185
rect 22450 3135 22500 3165
rect 22450 3115 22465 3135
rect 22485 3115 22500 3135
rect 22450 3085 22500 3115
rect 22450 3065 22465 3085
rect 22485 3065 22500 3085
rect 22450 3050 22500 3065
rect 22600 3050 22650 3550
rect 22750 3050 22800 3550
rect 22900 3050 22950 3550
rect 23050 3535 23100 3550
rect 23050 3515 23065 3535
rect 23085 3515 23100 3535
rect 23050 3485 23100 3515
rect 23050 3465 23065 3485
rect 23085 3465 23100 3485
rect 23050 3435 23100 3465
rect 23050 3415 23065 3435
rect 23085 3415 23100 3435
rect 23050 3385 23100 3415
rect 23050 3365 23065 3385
rect 23085 3365 23100 3385
rect 23050 3335 23100 3365
rect 23050 3315 23065 3335
rect 23085 3315 23100 3335
rect 23050 3285 23100 3315
rect 23050 3265 23065 3285
rect 23085 3265 23100 3285
rect 23050 3235 23100 3265
rect 23050 3215 23065 3235
rect 23085 3215 23100 3235
rect 23050 3185 23100 3215
rect 23050 3165 23065 3185
rect 23085 3165 23100 3185
rect 23050 3135 23100 3165
rect 23050 3115 23065 3135
rect 23085 3115 23100 3135
rect 23050 3085 23100 3115
rect 23050 3065 23065 3085
rect 23085 3065 23100 3085
rect 23050 3050 23100 3065
rect 23200 3050 23250 3550
rect 23350 3050 23400 3550
rect 23500 3535 23550 3550
rect 23500 3515 23515 3535
rect 23535 3515 23550 3535
rect 23500 3485 23550 3515
rect 23500 3465 23515 3485
rect 23535 3465 23550 3485
rect 23500 3435 23550 3465
rect 23500 3415 23515 3435
rect 23535 3415 23550 3435
rect 23500 3385 23550 3415
rect 23500 3365 23515 3385
rect 23535 3365 23550 3385
rect 23500 3335 23550 3365
rect 23500 3315 23515 3335
rect 23535 3315 23550 3335
rect 23500 3285 23550 3315
rect 23500 3265 23515 3285
rect 23535 3265 23550 3285
rect 23500 3235 23550 3265
rect 23500 3215 23515 3235
rect 23535 3215 23550 3235
rect 23500 3185 23550 3215
rect 23500 3165 23515 3185
rect 23535 3165 23550 3185
rect 23500 3135 23550 3165
rect 23500 3115 23515 3135
rect 23535 3115 23550 3135
rect 23500 3085 23550 3115
rect 23500 3065 23515 3085
rect 23535 3065 23550 3085
rect 23500 3050 23550 3065
rect 23650 3050 23700 3550
rect 23800 3050 23850 3550
rect 23950 3535 24000 3550
rect 23950 3515 23965 3535
rect 23985 3515 24000 3535
rect 23950 3485 24000 3515
rect 23950 3465 23965 3485
rect 23985 3465 24000 3485
rect 23950 3435 24000 3465
rect 23950 3415 23965 3435
rect 23985 3415 24000 3435
rect 23950 3385 24000 3415
rect 23950 3365 23965 3385
rect 23985 3365 24000 3385
rect 23950 3335 24000 3365
rect 23950 3315 23965 3335
rect 23985 3315 24000 3335
rect 23950 3285 24000 3315
rect 23950 3265 23965 3285
rect 23985 3265 24000 3285
rect 23950 3235 24000 3265
rect 23950 3215 23965 3235
rect 23985 3215 24000 3235
rect 23950 3185 24000 3215
rect 23950 3165 23965 3185
rect 23985 3165 24000 3185
rect 23950 3135 24000 3165
rect 23950 3115 23965 3135
rect 23985 3115 24000 3135
rect 23950 3085 24000 3115
rect 23950 3065 23965 3085
rect 23985 3065 24000 3085
rect 23950 3050 24000 3065
rect 24100 3050 24150 3550
rect 24250 3050 24300 3550
rect 24400 3050 24450 3550
rect 24550 3535 24600 3550
rect 24550 3515 24565 3535
rect 24585 3515 24600 3535
rect 24550 3485 24600 3515
rect 24550 3465 24565 3485
rect 24585 3465 24600 3485
rect 24550 3435 24600 3465
rect 24550 3415 24565 3435
rect 24585 3415 24600 3435
rect 24550 3385 24600 3415
rect 24550 3365 24565 3385
rect 24585 3365 24600 3385
rect 24550 3335 24600 3365
rect 24550 3315 24565 3335
rect 24585 3315 24600 3335
rect 24550 3285 24600 3315
rect 24550 3265 24565 3285
rect 24585 3265 24600 3285
rect 24550 3235 24600 3265
rect 24550 3215 24565 3235
rect 24585 3215 24600 3235
rect 24550 3185 24600 3215
rect 24550 3165 24565 3185
rect 24585 3165 24600 3185
rect 24550 3135 24600 3165
rect 24550 3115 24565 3135
rect 24585 3115 24600 3135
rect 24550 3085 24600 3115
rect 24550 3065 24565 3085
rect 24585 3065 24600 3085
rect 24550 3050 24600 3065
rect 24700 3050 24750 3550
rect 24850 3050 24900 3550
rect 25000 3050 25050 3550
rect 25150 3535 25200 3550
rect 25150 3515 25165 3535
rect 25185 3515 25200 3535
rect 25150 3485 25200 3515
rect 25150 3465 25165 3485
rect 25185 3465 25200 3485
rect 25150 3435 25200 3465
rect 25150 3415 25165 3435
rect 25185 3415 25200 3435
rect 25150 3385 25200 3415
rect 25150 3365 25165 3385
rect 25185 3365 25200 3385
rect 25150 3335 25200 3365
rect 25150 3315 25165 3335
rect 25185 3315 25200 3335
rect 25150 3285 25200 3315
rect 25150 3265 25165 3285
rect 25185 3265 25200 3285
rect 25150 3235 25200 3265
rect 25150 3215 25165 3235
rect 25185 3215 25200 3235
rect 25150 3185 25200 3215
rect 25150 3165 25165 3185
rect 25185 3165 25200 3185
rect 25150 3135 25200 3165
rect 25150 3115 25165 3135
rect 25185 3115 25200 3135
rect 25150 3085 25200 3115
rect 25150 3065 25165 3085
rect 25185 3065 25200 3085
rect 25150 3050 25200 3065
rect 25300 3050 25350 3550
rect 25450 3050 25500 3550
rect 25600 3535 25650 3550
rect 25600 3515 25615 3535
rect 25635 3515 25650 3535
rect 25600 3485 25650 3515
rect 25600 3465 25615 3485
rect 25635 3465 25650 3485
rect 25600 3435 25650 3465
rect 25600 3415 25615 3435
rect 25635 3415 25650 3435
rect 25600 3385 25650 3415
rect 25600 3365 25615 3385
rect 25635 3365 25650 3385
rect 25600 3335 25650 3365
rect 25600 3315 25615 3335
rect 25635 3315 25650 3335
rect 25600 3285 25650 3315
rect 25600 3265 25615 3285
rect 25635 3265 25650 3285
rect 25600 3235 25650 3265
rect 25600 3215 25615 3235
rect 25635 3215 25650 3235
rect 25600 3185 25650 3215
rect 25600 3165 25615 3185
rect 25635 3165 25650 3185
rect 25600 3135 25650 3165
rect 25600 3115 25615 3135
rect 25635 3115 25650 3135
rect 25600 3085 25650 3115
rect 25600 3065 25615 3085
rect 25635 3065 25650 3085
rect 25600 3050 25650 3065
rect 25750 3050 25800 3550
rect 25900 3050 25950 3550
rect 26050 3535 26100 3550
rect 26050 3515 26065 3535
rect 26085 3515 26100 3535
rect 26050 3485 26100 3515
rect 26050 3465 26065 3485
rect 26085 3465 26100 3485
rect 26050 3435 26100 3465
rect 26050 3415 26065 3435
rect 26085 3415 26100 3435
rect 26050 3385 26100 3415
rect 26050 3365 26065 3385
rect 26085 3365 26100 3385
rect 26050 3335 26100 3365
rect 26050 3315 26065 3335
rect 26085 3315 26100 3335
rect 26050 3285 26100 3315
rect 26050 3265 26065 3285
rect 26085 3265 26100 3285
rect 26050 3235 26100 3265
rect 26050 3215 26065 3235
rect 26085 3215 26100 3235
rect 26050 3185 26100 3215
rect 26050 3165 26065 3185
rect 26085 3165 26100 3185
rect 26050 3135 26100 3165
rect 26050 3115 26065 3135
rect 26085 3115 26100 3135
rect 26050 3085 26100 3115
rect 26050 3065 26065 3085
rect 26085 3065 26100 3085
rect 26050 3050 26100 3065
rect 26200 3050 26250 3550
rect 26350 3050 26400 3550
rect 26500 3050 26550 3550
rect 26650 3535 26700 3550
rect 26650 3515 26665 3535
rect 26685 3515 26700 3535
rect 26650 3485 26700 3515
rect 26650 3465 26665 3485
rect 26685 3465 26700 3485
rect 26650 3435 26700 3465
rect 26650 3415 26665 3435
rect 26685 3415 26700 3435
rect 26650 3385 26700 3415
rect 26650 3365 26665 3385
rect 26685 3365 26700 3385
rect 26650 3335 26700 3365
rect 26650 3315 26665 3335
rect 26685 3315 26700 3335
rect 26650 3285 26700 3315
rect 26650 3265 26665 3285
rect 26685 3265 26700 3285
rect 26650 3235 26700 3265
rect 26650 3215 26665 3235
rect 26685 3215 26700 3235
rect 26650 3185 26700 3215
rect 26650 3165 26665 3185
rect 26685 3165 26700 3185
rect 26650 3135 26700 3165
rect 26650 3115 26665 3135
rect 26685 3115 26700 3135
rect 26650 3085 26700 3115
rect 26650 3065 26665 3085
rect 26685 3065 26700 3085
rect 26650 3050 26700 3065
rect 26800 3050 26850 3550
rect 26950 3050 27000 3550
rect 27100 3050 27150 3550
rect 27250 3535 27300 3550
rect 27250 3515 27265 3535
rect 27285 3515 27300 3535
rect 27250 3485 27300 3515
rect 27250 3465 27265 3485
rect 27285 3465 27300 3485
rect 27250 3435 27300 3465
rect 27250 3415 27265 3435
rect 27285 3415 27300 3435
rect 27250 3385 27300 3415
rect 27250 3365 27265 3385
rect 27285 3365 27300 3385
rect 27250 3335 27300 3365
rect 27250 3315 27265 3335
rect 27285 3315 27300 3335
rect 27250 3285 27300 3315
rect 27250 3265 27265 3285
rect 27285 3265 27300 3285
rect 27250 3235 27300 3265
rect 27250 3215 27265 3235
rect 27285 3215 27300 3235
rect 27250 3185 27300 3215
rect 27250 3165 27265 3185
rect 27285 3165 27300 3185
rect 27250 3135 27300 3165
rect 27250 3115 27265 3135
rect 27285 3115 27300 3135
rect 27250 3085 27300 3115
rect 27250 3065 27265 3085
rect 27285 3065 27300 3085
rect 27250 3050 27300 3065
rect 27400 3050 27450 3550
rect 27550 3050 27600 3550
rect 27700 3535 27750 3550
rect 27700 3515 27715 3535
rect 27735 3515 27750 3535
rect 27700 3485 27750 3515
rect 27700 3465 27715 3485
rect 27735 3465 27750 3485
rect 27700 3435 27750 3465
rect 27700 3415 27715 3435
rect 27735 3415 27750 3435
rect 27700 3385 27750 3415
rect 27700 3365 27715 3385
rect 27735 3365 27750 3385
rect 27700 3335 27750 3365
rect 27700 3315 27715 3335
rect 27735 3315 27750 3335
rect 27700 3285 27750 3315
rect 27700 3265 27715 3285
rect 27735 3265 27750 3285
rect 27700 3235 27750 3265
rect 27700 3215 27715 3235
rect 27735 3215 27750 3235
rect 27700 3185 27750 3215
rect 27700 3165 27715 3185
rect 27735 3165 27750 3185
rect 27700 3135 27750 3165
rect 27700 3115 27715 3135
rect 27735 3115 27750 3135
rect 27700 3085 27750 3115
rect 27700 3065 27715 3085
rect 27735 3065 27750 3085
rect 27700 3050 27750 3065
rect 27850 3050 27900 3550
rect 28000 3050 28050 3550
rect 28150 3535 28200 3550
rect 28150 3515 28165 3535
rect 28185 3515 28200 3535
rect 28150 3485 28200 3515
rect 28150 3465 28165 3485
rect 28185 3465 28200 3485
rect 28150 3435 28200 3465
rect 28150 3415 28165 3435
rect 28185 3415 28200 3435
rect 28150 3385 28200 3415
rect 28150 3365 28165 3385
rect 28185 3365 28200 3385
rect 28150 3335 28200 3365
rect 28150 3315 28165 3335
rect 28185 3315 28200 3335
rect 28150 3285 28200 3315
rect 28150 3265 28165 3285
rect 28185 3265 28200 3285
rect 28150 3235 28200 3265
rect 28150 3215 28165 3235
rect 28185 3215 28200 3235
rect 28150 3185 28200 3215
rect 28150 3165 28165 3185
rect 28185 3165 28200 3185
rect 28150 3135 28200 3165
rect 28150 3115 28165 3135
rect 28185 3115 28200 3135
rect 28150 3085 28200 3115
rect 28150 3065 28165 3085
rect 28185 3065 28200 3085
rect 28150 3050 28200 3065
rect 28300 3050 28350 3550
rect 28450 3050 28500 3550
rect 28600 3050 28650 3550
rect 28750 3535 28800 3550
rect 28750 3515 28765 3535
rect 28785 3515 28800 3535
rect 28750 3485 28800 3515
rect 28750 3465 28765 3485
rect 28785 3465 28800 3485
rect 28750 3435 28800 3465
rect 28750 3415 28765 3435
rect 28785 3415 28800 3435
rect 28750 3385 28800 3415
rect 28750 3365 28765 3385
rect 28785 3365 28800 3385
rect 28750 3335 28800 3365
rect 28750 3315 28765 3335
rect 28785 3315 28800 3335
rect 28750 3285 28800 3315
rect 28750 3265 28765 3285
rect 28785 3265 28800 3285
rect 28750 3235 28800 3265
rect 28750 3215 28765 3235
rect 28785 3215 28800 3235
rect 28750 3185 28800 3215
rect 28750 3165 28765 3185
rect 28785 3165 28800 3185
rect 28750 3135 28800 3165
rect 28750 3115 28765 3135
rect 28785 3115 28800 3135
rect 28750 3085 28800 3115
rect 28750 3065 28765 3085
rect 28785 3065 28800 3085
rect 28750 3050 28800 3065
rect 28900 3050 28950 3550
rect 29050 3050 29100 3550
rect 29200 3050 29250 3550
rect 29350 3535 29400 3550
rect 29350 3515 29365 3535
rect 29385 3515 29400 3535
rect 29350 3485 29400 3515
rect 29350 3465 29365 3485
rect 29385 3465 29400 3485
rect 29350 3435 29400 3465
rect 29350 3415 29365 3435
rect 29385 3415 29400 3435
rect 29350 3385 29400 3415
rect 29350 3365 29365 3385
rect 29385 3365 29400 3385
rect 29350 3335 29400 3365
rect 29350 3315 29365 3335
rect 29385 3315 29400 3335
rect 29350 3285 29400 3315
rect 29350 3265 29365 3285
rect 29385 3265 29400 3285
rect 29350 3235 29400 3265
rect 29350 3215 29365 3235
rect 29385 3215 29400 3235
rect 29350 3185 29400 3215
rect 29350 3165 29365 3185
rect 29385 3165 29400 3185
rect 29350 3135 29400 3165
rect 29350 3115 29365 3135
rect 29385 3115 29400 3135
rect 29350 3085 29400 3115
rect 29350 3065 29365 3085
rect 29385 3065 29400 3085
rect 29350 3050 29400 3065
rect 29500 3535 29550 3550
rect 29500 3515 29515 3535
rect 29535 3515 29550 3535
rect 29500 3485 29550 3515
rect 29500 3465 29515 3485
rect 29535 3465 29550 3485
rect 29500 3435 29550 3465
rect 29500 3415 29515 3435
rect 29535 3415 29550 3435
rect 29500 3385 29550 3415
rect 29500 3365 29515 3385
rect 29535 3365 29550 3385
rect 29500 3335 29550 3365
rect 29500 3315 29515 3335
rect 29535 3315 29550 3335
rect 29500 3285 29550 3315
rect 29500 3265 29515 3285
rect 29535 3265 29550 3285
rect 29500 3235 29550 3265
rect 29500 3215 29515 3235
rect 29535 3215 29550 3235
rect 29500 3185 29550 3215
rect 29500 3165 29515 3185
rect 29535 3165 29550 3185
rect 29500 3135 29550 3165
rect 29500 3115 29515 3135
rect 29535 3115 29550 3135
rect 29500 3085 29550 3115
rect 29500 3065 29515 3085
rect 29535 3065 29550 3085
rect 29500 3050 29550 3065
rect 29650 3535 29700 3550
rect 29650 3515 29665 3535
rect 29685 3515 29700 3535
rect 29650 3485 29700 3515
rect 29650 3465 29665 3485
rect 29685 3465 29700 3485
rect 29650 3435 29700 3465
rect 29650 3415 29665 3435
rect 29685 3415 29700 3435
rect 29650 3385 29700 3415
rect 29650 3365 29665 3385
rect 29685 3365 29700 3385
rect 29650 3335 29700 3365
rect 29650 3315 29665 3335
rect 29685 3315 29700 3335
rect 29650 3285 29700 3315
rect 29650 3265 29665 3285
rect 29685 3265 29700 3285
rect 29650 3235 29700 3265
rect 29650 3215 29665 3235
rect 29685 3215 29700 3235
rect 29650 3185 29700 3215
rect 29650 3165 29665 3185
rect 29685 3165 29700 3185
rect 29650 3135 29700 3165
rect 29650 3115 29665 3135
rect 29685 3115 29700 3135
rect 29650 3085 29700 3115
rect 29650 3065 29665 3085
rect 29685 3065 29700 3085
rect 29650 3050 29700 3065
rect 29800 3535 29850 3550
rect 29800 3515 29815 3535
rect 29835 3515 29850 3535
rect 29800 3485 29850 3515
rect 29800 3465 29815 3485
rect 29835 3465 29850 3485
rect 29800 3435 29850 3465
rect 29800 3415 29815 3435
rect 29835 3415 29850 3435
rect 29800 3385 29850 3415
rect 29800 3365 29815 3385
rect 29835 3365 29850 3385
rect 29800 3335 29850 3365
rect 29800 3315 29815 3335
rect 29835 3315 29850 3335
rect 29800 3285 29850 3315
rect 29800 3265 29815 3285
rect 29835 3265 29850 3285
rect 29800 3235 29850 3265
rect 29800 3215 29815 3235
rect 29835 3215 29850 3235
rect 29800 3185 29850 3215
rect 29800 3165 29815 3185
rect 29835 3165 29850 3185
rect 29800 3135 29850 3165
rect 29800 3115 29815 3135
rect 29835 3115 29850 3135
rect 29800 3085 29850 3115
rect 29800 3065 29815 3085
rect 29835 3065 29850 3085
rect 29800 3050 29850 3065
rect 29950 3535 30000 3550
rect 29950 3515 29965 3535
rect 29985 3515 30000 3535
rect 29950 3485 30000 3515
rect 29950 3465 29965 3485
rect 29985 3465 30000 3485
rect 29950 3435 30000 3465
rect 29950 3415 29965 3435
rect 29985 3415 30000 3435
rect 29950 3385 30000 3415
rect 29950 3365 29965 3385
rect 29985 3365 30000 3385
rect 29950 3335 30000 3365
rect 29950 3315 29965 3335
rect 29985 3315 30000 3335
rect 29950 3285 30000 3315
rect 29950 3265 29965 3285
rect 29985 3265 30000 3285
rect 29950 3235 30000 3265
rect 29950 3215 29965 3235
rect 29985 3215 30000 3235
rect 29950 3185 30000 3215
rect 29950 3165 29965 3185
rect 29985 3165 30000 3185
rect 29950 3135 30000 3165
rect 29950 3115 29965 3135
rect 29985 3115 30000 3135
rect 29950 3085 30000 3115
rect 29950 3065 29965 3085
rect 29985 3065 30000 3085
rect 29950 3050 30000 3065
rect 30100 3535 30150 3550
rect 30100 3515 30115 3535
rect 30135 3515 30150 3535
rect 30100 3485 30150 3515
rect 30100 3465 30115 3485
rect 30135 3465 30150 3485
rect 30100 3435 30150 3465
rect 30100 3415 30115 3435
rect 30135 3415 30150 3435
rect 30100 3385 30150 3415
rect 30100 3365 30115 3385
rect 30135 3365 30150 3385
rect 30100 3335 30150 3365
rect 30100 3315 30115 3335
rect 30135 3315 30150 3335
rect 30100 3285 30150 3315
rect 30100 3265 30115 3285
rect 30135 3265 30150 3285
rect 30100 3235 30150 3265
rect 30100 3215 30115 3235
rect 30135 3215 30150 3235
rect 30100 3185 30150 3215
rect 30100 3165 30115 3185
rect 30135 3165 30150 3185
rect 30100 3135 30150 3165
rect 30100 3115 30115 3135
rect 30135 3115 30150 3135
rect 30100 3085 30150 3115
rect 30100 3065 30115 3085
rect 30135 3065 30150 3085
rect 30100 3050 30150 3065
rect 30250 3535 30300 3550
rect 30250 3515 30265 3535
rect 30285 3515 30300 3535
rect 30250 3485 30300 3515
rect 30250 3465 30265 3485
rect 30285 3465 30300 3485
rect 30250 3435 30300 3465
rect 30250 3415 30265 3435
rect 30285 3415 30300 3435
rect 30250 3385 30300 3415
rect 30250 3365 30265 3385
rect 30285 3365 30300 3385
rect 30250 3335 30300 3365
rect 30250 3315 30265 3335
rect 30285 3315 30300 3335
rect 30250 3285 30300 3315
rect 30250 3265 30265 3285
rect 30285 3265 30300 3285
rect 30250 3235 30300 3265
rect 30250 3215 30265 3235
rect 30285 3215 30300 3235
rect 30250 3185 30300 3215
rect 30250 3165 30265 3185
rect 30285 3165 30300 3185
rect 30250 3135 30300 3165
rect 30250 3115 30265 3135
rect 30285 3115 30300 3135
rect 30250 3085 30300 3115
rect 30250 3065 30265 3085
rect 30285 3065 30300 3085
rect 30250 3050 30300 3065
rect 30400 3535 30450 3550
rect 30400 3515 30415 3535
rect 30435 3515 30450 3535
rect 30400 3485 30450 3515
rect 30400 3465 30415 3485
rect 30435 3465 30450 3485
rect 30400 3435 30450 3465
rect 30400 3415 30415 3435
rect 30435 3415 30450 3435
rect 30400 3385 30450 3415
rect 30400 3365 30415 3385
rect 30435 3365 30450 3385
rect 30400 3335 30450 3365
rect 30400 3315 30415 3335
rect 30435 3315 30450 3335
rect 30400 3285 30450 3315
rect 30400 3265 30415 3285
rect 30435 3265 30450 3285
rect 30400 3235 30450 3265
rect 30400 3215 30415 3235
rect 30435 3215 30450 3235
rect 30400 3185 30450 3215
rect 30400 3165 30415 3185
rect 30435 3165 30450 3185
rect 30400 3135 30450 3165
rect 30400 3115 30415 3135
rect 30435 3115 30450 3135
rect 30400 3085 30450 3115
rect 30400 3065 30415 3085
rect 30435 3065 30450 3085
rect 30400 3050 30450 3065
rect 30550 3535 30600 3550
rect 30550 3515 30565 3535
rect 30585 3515 30600 3535
rect 30550 3485 30600 3515
rect 30550 3465 30565 3485
rect 30585 3465 30600 3485
rect 30550 3435 30600 3465
rect 30550 3415 30565 3435
rect 30585 3415 30600 3435
rect 30550 3385 30600 3415
rect 30550 3365 30565 3385
rect 30585 3365 30600 3385
rect 30550 3335 30600 3365
rect 30550 3315 30565 3335
rect 30585 3315 30600 3335
rect 30550 3285 30600 3315
rect 30550 3265 30565 3285
rect 30585 3265 30600 3285
rect 30550 3235 30600 3265
rect 30550 3215 30565 3235
rect 30585 3215 30600 3235
rect 30550 3185 30600 3215
rect 30550 3165 30565 3185
rect 30585 3165 30600 3185
rect 30550 3135 30600 3165
rect 30550 3115 30565 3135
rect 30585 3115 30600 3135
rect 30550 3085 30600 3115
rect 30550 3065 30565 3085
rect 30585 3065 30600 3085
rect 30550 3050 30600 3065
rect 30700 3535 30750 3550
rect 30700 3515 30715 3535
rect 30735 3515 30750 3535
rect 30700 3485 30750 3515
rect 30700 3465 30715 3485
rect 30735 3465 30750 3485
rect 30700 3435 30750 3465
rect 30700 3415 30715 3435
rect 30735 3415 30750 3435
rect 30700 3385 30750 3415
rect 30700 3365 30715 3385
rect 30735 3365 30750 3385
rect 30700 3335 30750 3365
rect 30700 3315 30715 3335
rect 30735 3315 30750 3335
rect 30700 3285 30750 3315
rect 30700 3265 30715 3285
rect 30735 3265 30750 3285
rect 30700 3235 30750 3265
rect 30700 3215 30715 3235
rect 30735 3215 30750 3235
rect 30700 3185 30750 3215
rect 30700 3165 30715 3185
rect 30735 3165 30750 3185
rect 30700 3135 30750 3165
rect 30700 3115 30715 3135
rect 30735 3115 30750 3135
rect 30700 3085 30750 3115
rect 30700 3065 30715 3085
rect 30735 3065 30750 3085
rect 30700 3050 30750 3065
rect 30850 3535 30900 3550
rect 30850 3515 30865 3535
rect 30885 3515 30900 3535
rect 30850 3485 30900 3515
rect 30850 3465 30865 3485
rect 30885 3465 30900 3485
rect 30850 3435 30900 3465
rect 30850 3415 30865 3435
rect 30885 3415 30900 3435
rect 30850 3385 30900 3415
rect 30850 3365 30865 3385
rect 30885 3365 30900 3385
rect 30850 3335 30900 3365
rect 30850 3315 30865 3335
rect 30885 3315 30900 3335
rect 30850 3285 30900 3315
rect 30850 3265 30865 3285
rect 30885 3265 30900 3285
rect 30850 3235 30900 3265
rect 30850 3215 30865 3235
rect 30885 3215 30900 3235
rect 30850 3185 30900 3215
rect 30850 3165 30865 3185
rect 30885 3165 30900 3185
rect 30850 3135 30900 3165
rect 30850 3115 30865 3135
rect 30885 3115 30900 3135
rect 30850 3085 30900 3115
rect 30850 3065 30865 3085
rect 30885 3065 30900 3085
rect 30850 3050 30900 3065
rect 31000 3535 31050 3550
rect 31000 3515 31015 3535
rect 31035 3515 31050 3535
rect 31000 3485 31050 3515
rect 31000 3465 31015 3485
rect 31035 3465 31050 3485
rect 31000 3435 31050 3465
rect 31000 3415 31015 3435
rect 31035 3415 31050 3435
rect 31000 3385 31050 3415
rect 31000 3365 31015 3385
rect 31035 3365 31050 3385
rect 31000 3335 31050 3365
rect 31000 3315 31015 3335
rect 31035 3315 31050 3335
rect 31000 3285 31050 3315
rect 31000 3265 31015 3285
rect 31035 3265 31050 3285
rect 31000 3235 31050 3265
rect 31000 3215 31015 3235
rect 31035 3215 31050 3235
rect 31000 3185 31050 3215
rect 31000 3165 31015 3185
rect 31035 3165 31050 3185
rect 31000 3135 31050 3165
rect 31000 3115 31015 3135
rect 31035 3115 31050 3135
rect 31000 3085 31050 3115
rect 31000 3065 31015 3085
rect 31035 3065 31050 3085
rect 31000 3050 31050 3065
rect 31150 3535 31200 3550
rect 31150 3515 31165 3535
rect 31185 3515 31200 3535
rect 31150 3485 31200 3515
rect 31150 3465 31165 3485
rect 31185 3465 31200 3485
rect 31150 3435 31200 3465
rect 31150 3415 31165 3435
rect 31185 3415 31200 3435
rect 31150 3385 31200 3415
rect 31150 3365 31165 3385
rect 31185 3365 31200 3385
rect 31150 3335 31200 3365
rect 31150 3315 31165 3335
rect 31185 3315 31200 3335
rect 31150 3285 31200 3315
rect 31150 3265 31165 3285
rect 31185 3265 31200 3285
rect 31150 3235 31200 3265
rect 31150 3215 31165 3235
rect 31185 3215 31200 3235
rect 31150 3185 31200 3215
rect 31150 3165 31165 3185
rect 31185 3165 31200 3185
rect 31150 3135 31200 3165
rect 31150 3115 31165 3135
rect 31185 3115 31200 3135
rect 31150 3085 31200 3115
rect 31150 3065 31165 3085
rect 31185 3065 31200 3085
rect 31150 3050 31200 3065
rect 31300 3535 31350 3550
rect 31300 3515 31315 3535
rect 31335 3515 31350 3535
rect 31300 3485 31350 3515
rect 31300 3465 31315 3485
rect 31335 3465 31350 3485
rect 31300 3435 31350 3465
rect 31300 3415 31315 3435
rect 31335 3415 31350 3435
rect 31300 3385 31350 3415
rect 31300 3365 31315 3385
rect 31335 3365 31350 3385
rect 31300 3335 31350 3365
rect 31300 3315 31315 3335
rect 31335 3315 31350 3335
rect 31300 3285 31350 3315
rect 31300 3265 31315 3285
rect 31335 3265 31350 3285
rect 31300 3235 31350 3265
rect 31300 3215 31315 3235
rect 31335 3215 31350 3235
rect 31300 3185 31350 3215
rect 31300 3165 31315 3185
rect 31335 3165 31350 3185
rect 31300 3135 31350 3165
rect 31300 3115 31315 3135
rect 31335 3115 31350 3135
rect 31300 3085 31350 3115
rect 31300 3065 31315 3085
rect 31335 3065 31350 3085
rect 31300 3050 31350 3065
rect 31450 3535 31500 3550
rect 31450 3515 31465 3535
rect 31485 3515 31500 3535
rect 31450 3485 31500 3515
rect 31450 3465 31465 3485
rect 31485 3465 31500 3485
rect 31450 3435 31500 3465
rect 31450 3415 31465 3435
rect 31485 3415 31500 3435
rect 31450 3385 31500 3415
rect 31450 3365 31465 3385
rect 31485 3365 31500 3385
rect 31450 3335 31500 3365
rect 31450 3315 31465 3335
rect 31485 3315 31500 3335
rect 31450 3285 31500 3315
rect 31450 3265 31465 3285
rect 31485 3265 31500 3285
rect 31450 3235 31500 3265
rect 31450 3215 31465 3235
rect 31485 3215 31500 3235
rect 31450 3185 31500 3215
rect 31450 3165 31465 3185
rect 31485 3165 31500 3185
rect 31450 3135 31500 3165
rect 31450 3115 31465 3135
rect 31485 3115 31500 3135
rect 31450 3085 31500 3115
rect 31450 3065 31465 3085
rect 31485 3065 31500 3085
rect 31450 3050 31500 3065
rect 31600 3050 31650 3550
rect 31750 3050 31800 3550
rect 31900 3050 31950 3550
rect 32050 3535 32100 3550
rect 32050 3515 32065 3535
rect 32085 3515 32100 3535
rect 32050 3485 32100 3515
rect 32050 3465 32065 3485
rect 32085 3465 32100 3485
rect 32050 3435 32100 3465
rect 32050 3415 32065 3435
rect 32085 3415 32100 3435
rect 32050 3385 32100 3415
rect 32050 3365 32065 3385
rect 32085 3365 32100 3385
rect 32050 3335 32100 3365
rect 32050 3315 32065 3335
rect 32085 3315 32100 3335
rect 32050 3285 32100 3315
rect 32050 3265 32065 3285
rect 32085 3265 32100 3285
rect 32050 3235 32100 3265
rect 32050 3215 32065 3235
rect 32085 3215 32100 3235
rect 32050 3185 32100 3215
rect 32050 3165 32065 3185
rect 32085 3165 32100 3185
rect 32050 3135 32100 3165
rect 32050 3115 32065 3135
rect 32085 3115 32100 3135
rect 32050 3085 32100 3115
rect 32050 3065 32065 3085
rect 32085 3065 32100 3085
rect 32050 3050 32100 3065
<< mvndiffc >>
rect -635 1565 -615 1585
rect -635 1515 -615 1535
rect -635 1465 -615 1485
rect -635 1415 -615 1435
rect -635 1365 -615 1385
rect -635 1315 -615 1335
rect -635 1265 -615 1285
rect -635 1215 -615 1235
rect -635 1165 -615 1185
rect -635 1115 -615 1135
rect -635 1065 -615 1085
rect -635 1015 -615 1035
rect -635 965 -615 985
rect -635 915 -615 935
rect -485 1565 -465 1585
rect -485 1515 -465 1535
rect -485 1465 -465 1485
rect -485 1415 -465 1435
rect -485 1365 -465 1385
rect -485 1315 -465 1335
rect -485 1265 -465 1285
rect -485 1215 -465 1235
rect -485 1165 -465 1185
rect -485 1115 -465 1135
rect -485 1065 -465 1085
rect -485 1015 -465 1035
rect -485 965 -465 985
rect -485 915 -465 935
rect -335 1565 -315 1585
rect -335 1515 -315 1535
rect -335 1465 -315 1485
rect -335 1415 -315 1435
rect -335 1365 -315 1385
rect -335 1315 -315 1335
rect -335 1265 -315 1285
rect -335 1215 -315 1235
rect -335 1165 -315 1185
rect -335 1115 -315 1135
rect -335 1065 -315 1085
rect -335 1015 -315 1035
rect -335 965 -315 985
rect -335 915 -315 935
rect -185 1565 -165 1585
rect -185 1515 -165 1535
rect -185 1465 -165 1485
rect -185 1415 -165 1435
rect -185 1365 -165 1385
rect -185 1315 -165 1335
rect -185 1265 -165 1285
rect -185 1215 -165 1235
rect -185 1165 -165 1185
rect -185 1115 -165 1135
rect -185 1065 -165 1085
rect -185 1015 -165 1035
rect -185 965 -165 985
rect -185 915 -165 935
rect -35 1565 -15 1585
rect -35 1515 -15 1535
rect -35 1465 -15 1485
rect -35 1415 -15 1435
rect -35 1365 -15 1385
rect -35 1315 -15 1335
rect -35 1265 -15 1285
rect -35 1215 -15 1235
rect -35 1165 -15 1185
rect -35 1115 -15 1135
rect -35 1065 -15 1085
rect -35 1015 -15 1035
rect -35 965 -15 985
rect -35 915 -15 935
rect 1165 1565 1185 1585
rect 1165 1515 1185 1535
rect 1165 1465 1185 1485
rect 1165 1415 1185 1435
rect 1165 1365 1185 1385
rect 1165 1315 1185 1335
rect 1165 1265 1185 1285
rect 1165 1215 1185 1235
rect 1165 1165 1185 1185
rect 1165 1115 1185 1135
rect 1165 1065 1185 1085
rect 1165 1015 1185 1035
rect 1165 965 1185 985
rect 1165 915 1185 935
rect 1465 1565 1485 1585
rect 1465 1515 1485 1535
rect 1465 1465 1485 1485
rect 1465 1415 1485 1435
rect 1465 1365 1485 1385
rect 1465 1315 1485 1335
rect 1465 1265 1485 1285
rect 1465 1215 1485 1235
rect 1465 1165 1485 1185
rect 1465 1115 1485 1135
rect 1465 1065 1485 1085
rect 1465 1015 1485 1035
rect 1465 965 1485 985
rect 1465 915 1485 935
rect 1765 1565 1785 1585
rect 1765 1515 1785 1535
rect 1765 1465 1785 1485
rect 1765 1415 1785 1435
rect 1765 1365 1785 1385
rect 1765 1315 1785 1335
rect 1765 1265 1785 1285
rect 1765 1215 1785 1235
rect 1765 1165 1785 1185
rect 1765 1115 1785 1135
rect 1765 1065 1785 1085
rect 1765 1015 1785 1035
rect 1765 965 1785 985
rect 1765 915 1785 935
rect 2065 1565 2085 1585
rect 2065 1515 2085 1535
rect 2065 1465 2085 1485
rect 2065 1415 2085 1435
rect 2065 1365 2085 1385
rect 2065 1315 2085 1335
rect 2065 1265 2085 1285
rect 2065 1215 2085 1235
rect 2065 1165 2085 1185
rect 2065 1115 2085 1135
rect 2065 1065 2085 1085
rect 2065 1015 2085 1035
rect 2065 965 2085 985
rect 2065 915 2085 935
rect 2365 1565 2385 1585
rect 2365 1515 2385 1535
rect 2365 1465 2385 1485
rect 2365 1415 2385 1435
rect 2365 1365 2385 1385
rect 2365 1315 2385 1335
rect 2365 1265 2385 1285
rect 2365 1215 2385 1235
rect 2365 1165 2385 1185
rect 2365 1115 2385 1135
rect 2365 1065 2385 1085
rect 2365 1015 2385 1035
rect 2365 965 2385 985
rect 2365 915 2385 935
rect 2665 1565 2685 1585
rect 2665 1515 2685 1535
rect 2665 1465 2685 1485
rect 2665 1415 2685 1435
rect 2665 1365 2685 1385
rect 2665 1315 2685 1335
rect 2665 1265 2685 1285
rect 2665 1215 2685 1235
rect 2665 1165 2685 1185
rect 2665 1115 2685 1135
rect 2665 1065 2685 1085
rect 2665 1015 2685 1035
rect 2665 965 2685 985
rect 2665 915 2685 935
rect 2965 1565 2985 1585
rect 2965 1515 2985 1535
rect 2965 1465 2985 1485
rect 2965 1415 2985 1435
rect 2965 1365 2985 1385
rect 2965 1315 2985 1335
rect 2965 1265 2985 1285
rect 2965 1215 2985 1235
rect 2965 1165 2985 1185
rect 2965 1115 2985 1135
rect 2965 1065 2985 1085
rect 2965 1015 2985 1035
rect 2965 965 2985 985
rect 2965 915 2985 935
rect 3265 1565 3285 1585
rect 3265 1515 3285 1535
rect 3265 1465 3285 1485
rect 3265 1415 3285 1435
rect 3265 1365 3285 1385
rect 3265 1315 3285 1335
rect 3265 1265 3285 1285
rect 3265 1215 3285 1235
rect 3265 1165 3285 1185
rect 3265 1115 3285 1135
rect 3265 1065 3285 1085
rect 3265 1015 3285 1035
rect 3265 965 3285 985
rect 3265 915 3285 935
rect 3565 1565 3585 1585
rect 3565 1515 3585 1535
rect 3565 1465 3585 1485
rect 3565 1415 3585 1435
rect 3565 1365 3585 1385
rect 3565 1315 3585 1335
rect 3565 1265 3585 1285
rect 3565 1215 3585 1235
rect 3565 1165 3585 1185
rect 3565 1115 3585 1135
rect 3565 1065 3585 1085
rect 3565 1015 3585 1035
rect 3565 965 3585 985
rect 3565 915 3585 935
rect 3715 1565 3735 1585
rect 3715 1515 3735 1535
rect 3715 1465 3735 1485
rect 3715 1415 3735 1435
rect 3715 1365 3735 1385
rect 3715 1315 3735 1335
rect 3715 1265 3735 1285
rect 3715 1215 3735 1235
rect 3715 1165 3735 1185
rect 3715 1115 3735 1135
rect 3715 1065 3735 1085
rect 3715 1015 3735 1035
rect 3715 965 3735 985
rect 3715 915 3735 935
rect 3865 1565 3885 1585
rect 3865 1515 3885 1535
rect 3865 1465 3885 1485
rect 3865 1415 3885 1435
rect 3865 1365 3885 1385
rect 3865 1315 3885 1335
rect 3865 1265 3885 1285
rect 3865 1215 3885 1235
rect 3865 1165 3885 1185
rect 3865 1115 3885 1135
rect 3865 1065 3885 1085
rect 3865 1015 3885 1035
rect 3865 965 3885 985
rect 3865 915 3885 935
rect 4015 1565 4035 1585
rect 4015 1515 4035 1535
rect 4015 1465 4035 1485
rect 4015 1415 4035 1435
rect 4015 1365 4035 1385
rect 4015 1315 4035 1335
rect 4015 1265 4035 1285
rect 4015 1215 4035 1235
rect 4015 1165 4035 1185
rect 4015 1115 4035 1135
rect 4015 1065 4035 1085
rect 4015 1015 4035 1035
rect 4015 965 4035 985
rect 4015 915 4035 935
rect 4165 1565 4185 1585
rect 4165 1515 4185 1535
rect 4165 1465 4185 1485
rect 4165 1415 4185 1435
rect 4165 1365 4185 1385
rect 4165 1315 4185 1335
rect 4165 1265 4185 1285
rect 4165 1215 4185 1235
rect 4165 1165 4185 1185
rect 4165 1115 4185 1135
rect 4165 1065 4185 1085
rect 4165 1015 4185 1035
rect 4165 965 4185 985
rect 4165 915 4185 935
rect 4315 1565 4335 1585
rect 4315 1515 4335 1535
rect 4315 1465 4335 1485
rect 4315 1415 4335 1435
rect 4315 1365 4335 1385
rect 4315 1315 4335 1335
rect 4315 1265 4335 1285
rect 4315 1215 4335 1235
rect 4315 1165 4335 1185
rect 4315 1115 4335 1135
rect 4315 1065 4335 1085
rect 4315 1015 4335 1035
rect 4315 965 4335 985
rect 4315 915 4335 935
rect 4465 1565 4485 1585
rect 4465 1515 4485 1535
rect 4465 1465 4485 1485
rect 4465 1415 4485 1435
rect 4465 1365 4485 1385
rect 4465 1315 4485 1335
rect 4465 1265 4485 1285
rect 4465 1215 4485 1235
rect 4465 1165 4485 1185
rect 4465 1115 4485 1135
rect 4465 1065 4485 1085
rect 4465 1015 4485 1035
rect 4465 965 4485 985
rect 4465 915 4485 935
rect 4615 1565 4635 1585
rect 4615 1515 4635 1535
rect 4615 1465 4635 1485
rect 4615 1415 4635 1435
rect 4615 1365 4635 1385
rect 4615 1315 4635 1335
rect 4615 1265 4635 1285
rect 4615 1215 4635 1235
rect 4615 1165 4635 1185
rect 4615 1115 4635 1135
rect 4615 1065 4635 1085
rect 4615 1015 4635 1035
rect 4615 965 4635 985
rect 4615 915 4635 935
rect 4765 1565 4785 1585
rect 4765 1515 4785 1535
rect 4765 1465 4785 1485
rect 4765 1415 4785 1435
rect 4765 1365 4785 1385
rect 4765 1315 4785 1335
rect 4765 1265 4785 1285
rect 4765 1215 4785 1235
rect 4765 1165 4785 1185
rect 4765 1115 4785 1135
rect 4765 1065 4785 1085
rect 4765 1015 4785 1035
rect 4765 965 4785 985
rect 4765 915 4785 935
rect 5065 1565 5085 1585
rect 5065 1515 5085 1535
rect 5065 1465 5085 1485
rect 5065 1415 5085 1435
rect 5065 1365 5085 1385
rect 5065 1315 5085 1335
rect 5065 1265 5085 1285
rect 5065 1215 5085 1235
rect 5065 1165 5085 1185
rect 5065 1115 5085 1135
rect 5065 1065 5085 1085
rect 5065 1015 5085 1035
rect 5065 965 5085 985
rect 5065 915 5085 935
rect 5365 1565 5385 1585
rect 5365 1515 5385 1535
rect 5365 1465 5385 1485
rect 5365 1415 5385 1435
rect 5365 1365 5385 1385
rect 5365 1315 5385 1335
rect 5365 1265 5385 1285
rect 5365 1215 5385 1235
rect 5365 1165 5385 1185
rect 5365 1115 5385 1135
rect 5365 1065 5385 1085
rect 5365 1015 5385 1035
rect 5365 965 5385 985
rect 5365 915 5385 935
rect 5665 1565 5685 1585
rect 5665 1515 5685 1535
rect 5665 1465 5685 1485
rect 5665 1415 5685 1435
rect 5665 1365 5685 1385
rect 5665 1315 5685 1335
rect 5665 1265 5685 1285
rect 5665 1215 5685 1235
rect 5665 1165 5685 1185
rect 5665 1115 5685 1135
rect 5665 1065 5685 1085
rect 5665 1015 5685 1035
rect 5665 965 5685 985
rect 5665 915 5685 935
rect 5965 1565 5985 1585
rect 5965 1515 5985 1535
rect 5965 1465 5985 1485
rect 5965 1415 5985 1435
rect 5965 1365 5985 1385
rect 5965 1315 5985 1335
rect 5965 1265 5985 1285
rect 5965 1215 5985 1235
rect 5965 1165 5985 1185
rect 5965 1115 5985 1135
rect 5965 1065 5985 1085
rect 5965 1015 5985 1035
rect 5965 965 5985 985
rect 5965 915 5985 935
rect 6265 1565 6285 1585
rect 6265 1515 6285 1535
rect 6265 1465 6285 1485
rect 6265 1415 6285 1435
rect 6265 1365 6285 1385
rect 6265 1315 6285 1335
rect 6265 1265 6285 1285
rect 6265 1215 6285 1235
rect 6265 1165 6285 1185
rect 6265 1115 6285 1135
rect 6265 1065 6285 1085
rect 6265 1015 6285 1035
rect 6265 965 6285 985
rect 6265 915 6285 935
rect 6565 1565 6585 1585
rect 6565 1515 6585 1535
rect 6565 1465 6585 1485
rect 6565 1415 6585 1435
rect 6565 1365 6585 1385
rect 6565 1315 6585 1335
rect 6565 1265 6585 1285
rect 6565 1215 6585 1235
rect 6565 1165 6585 1185
rect 6565 1115 6585 1135
rect 6565 1065 6585 1085
rect 6565 1015 6585 1035
rect 6565 965 6585 985
rect 6565 915 6585 935
rect 6865 1565 6885 1585
rect 6865 1515 6885 1535
rect 6865 1465 6885 1485
rect 6865 1415 6885 1435
rect 6865 1365 6885 1385
rect 6865 1315 6885 1335
rect 6865 1265 6885 1285
rect 6865 1215 6885 1235
rect 6865 1165 6885 1185
rect 6865 1115 6885 1135
rect 6865 1065 6885 1085
rect 6865 1015 6885 1035
rect 6865 965 6885 985
rect 6865 915 6885 935
rect 7165 1565 7185 1585
rect 7165 1515 7185 1535
rect 7165 1465 7185 1485
rect 7165 1415 7185 1435
rect 7165 1365 7185 1385
rect 7165 1315 7185 1335
rect 7165 1265 7185 1285
rect 7165 1215 7185 1235
rect 7165 1165 7185 1185
rect 7165 1115 7185 1135
rect 7165 1065 7185 1085
rect 7165 1015 7185 1035
rect 7165 965 7185 985
rect 7165 915 7185 935
rect 8365 1565 8385 1585
rect 8365 1515 8385 1535
rect 8365 1465 8385 1485
rect 8365 1415 8385 1435
rect 8365 1365 8385 1385
rect 8365 1315 8385 1335
rect 8365 1265 8385 1285
rect 8365 1215 8385 1235
rect 8365 1165 8385 1185
rect 8365 1115 8385 1135
rect 8365 1065 8385 1085
rect 8365 1015 8385 1035
rect 8365 965 8385 985
rect 8365 915 8385 935
rect 9565 1565 9585 1585
rect 9565 1515 9585 1535
rect 9565 1465 9585 1485
rect 9565 1415 9585 1435
rect 9565 1365 9585 1385
rect 9565 1315 9585 1335
rect 9565 1265 9585 1285
rect 9565 1215 9585 1235
rect 9565 1165 9585 1185
rect 9565 1115 9585 1135
rect 9565 1065 9585 1085
rect 9565 1015 9585 1035
rect 9565 965 9585 985
rect 9565 915 9585 935
rect 10765 1565 10785 1585
rect 10765 1515 10785 1535
rect 10765 1465 10785 1485
rect 10765 1415 10785 1435
rect 10765 1365 10785 1385
rect 10765 1315 10785 1335
rect 10765 1265 10785 1285
rect 10765 1215 10785 1235
rect 10765 1165 10785 1185
rect 10765 1115 10785 1135
rect 10765 1065 10785 1085
rect 10765 1015 10785 1035
rect 10765 965 10785 985
rect 10765 915 10785 935
rect 11965 1565 11985 1585
rect 11965 1515 11985 1535
rect 11965 1465 11985 1485
rect 11965 1415 11985 1435
rect 11965 1365 11985 1385
rect 11965 1315 11985 1335
rect 11965 1265 11985 1285
rect 11965 1215 11985 1235
rect 11965 1165 11985 1185
rect 11965 1115 11985 1135
rect 11965 1065 11985 1085
rect 11965 1015 11985 1035
rect 11965 965 11985 985
rect 11965 915 11985 935
rect 12265 1565 12285 1585
rect 12265 1515 12285 1535
rect 12265 1465 12285 1485
rect 12265 1415 12285 1435
rect 12265 1365 12285 1385
rect 12265 1315 12285 1335
rect 12265 1265 12285 1285
rect 12265 1215 12285 1235
rect 12265 1165 12285 1185
rect 12265 1115 12285 1135
rect 12265 1065 12285 1085
rect 12265 1015 12285 1035
rect 12265 965 12285 985
rect 12265 915 12285 935
rect 12565 1565 12585 1585
rect 12565 1515 12585 1535
rect 12565 1465 12585 1485
rect 12565 1415 12585 1435
rect 12565 1365 12585 1385
rect 12565 1315 12585 1335
rect 12565 1265 12585 1285
rect 12565 1215 12585 1235
rect 12565 1165 12585 1185
rect 12565 1115 12585 1135
rect 12565 1065 12585 1085
rect 12565 1015 12585 1035
rect 12565 965 12585 985
rect 12565 915 12585 935
rect 12865 1565 12885 1585
rect 12865 1515 12885 1535
rect 12865 1465 12885 1485
rect 12865 1415 12885 1435
rect 12865 1365 12885 1385
rect 12865 1315 12885 1335
rect 12865 1265 12885 1285
rect 12865 1215 12885 1235
rect 12865 1165 12885 1185
rect 12865 1115 12885 1135
rect 12865 1065 12885 1085
rect 12865 1015 12885 1035
rect 12865 965 12885 985
rect 12865 915 12885 935
rect 13165 1565 13185 1585
rect 13165 1515 13185 1535
rect 13165 1465 13185 1485
rect 13165 1415 13185 1435
rect 13165 1365 13185 1385
rect 13165 1315 13185 1335
rect 13165 1265 13185 1285
rect 13165 1215 13185 1235
rect 13165 1165 13185 1185
rect 13165 1115 13185 1135
rect 13165 1065 13185 1085
rect 13165 1015 13185 1035
rect 13165 965 13185 985
rect 13165 915 13185 935
rect 13465 1565 13485 1585
rect 13465 1515 13485 1535
rect 13465 1465 13485 1485
rect 13465 1415 13485 1435
rect 13465 1365 13485 1385
rect 13465 1315 13485 1335
rect 13465 1265 13485 1285
rect 13465 1215 13485 1235
rect 13465 1165 13485 1185
rect 13465 1115 13485 1135
rect 13465 1065 13485 1085
rect 13465 1015 13485 1035
rect 13465 965 13485 985
rect 13465 915 13485 935
rect 13765 1565 13785 1585
rect 13765 1515 13785 1535
rect 13765 1465 13785 1485
rect 13765 1415 13785 1435
rect 13765 1365 13785 1385
rect 13765 1315 13785 1335
rect 13765 1265 13785 1285
rect 13765 1215 13785 1235
rect 13765 1165 13785 1185
rect 13765 1115 13785 1135
rect 13765 1065 13785 1085
rect 13765 1015 13785 1035
rect 13765 965 13785 985
rect 13765 915 13785 935
rect 14065 1565 14085 1585
rect 14065 1515 14085 1535
rect 14065 1465 14085 1485
rect 14065 1415 14085 1435
rect 14065 1365 14085 1385
rect 14065 1315 14085 1335
rect 14065 1265 14085 1285
rect 14065 1215 14085 1235
rect 14065 1165 14085 1185
rect 14065 1115 14085 1135
rect 14065 1065 14085 1085
rect 14065 1015 14085 1035
rect 14065 965 14085 985
rect 14065 915 14085 935
rect 14365 1565 14385 1585
rect 14365 1515 14385 1535
rect 14365 1465 14385 1485
rect 14365 1415 14385 1435
rect 14365 1365 14385 1385
rect 14365 1315 14385 1335
rect 14365 1265 14385 1285
rect 14365 1215 14385 1235
rect 14365 1165 14385 1185
rect 14365 1115 14385 1135
rect 14365 1065 14385 1085
rect 14365 1015 14385 1035
rect 14365 965 14385 985
rect 14365 915 14385 935
rect 15565 1565 15585 1585
rect 15565 1515 15585 1535
rect 15565 1465 15585 1485
rect 15565 1415 15585 1435
rect 15565 1365 15585 1385
rect 15565 1315 15585 1335
rect 15565 1265 15585 1285
rect 15565 1215 15585 1235
rect 15565 1165 15585 1185
rect 15565 1115 15585 1135
rect 15565 1065 15585 1085
rect 15565 1015 15585 1035
rect 15565 965 15585 985
rect 15565 915 15585 935
rect 16765 1565 16785 1585
rect 16765 1515 16785 1535
rect 16765 1465 16785 1485
rect 16765 1415 16785 1435
rect 16765 1365 16785 1385
rect 16765 1315 16785 1335
rect 16765 1265 16785 1285
rect 16765 1215 16785 1235
rect 16765 1165 16785 1185
rect 16765 1115 16785 1135
rect 16765 1065 16785 1085
rect 16765 1015 16785 1035
rect 16765 965 16785 985
rect 16765 915 16785 935
rect 17965 1565 17985 1585
rect 17965 1515 17985 1535
rect 17965 1465 17985 1485
rect 17965 1415 17985 1435
rect 17965 1365 17985 1385
rect 17965 1315 17985 1335
rect 17965 1265 17985 1285
rect 17965 1215 17985 1235
rect 17965 1165 17985 1185
rect 17965 1115 17985 1135
rect 17965 1065 17985 1085
rect 17965 1015 17985 1035
rect 17965 965 17985 985
rect 17965 915 17985 935
rect 19165 1565 19185 1585
rect 19165 1515 19185 1535
rect 19165 1465 19185 1485
rect 19165 1415 19185 1435
rect 19165 1365 19185 1385
rect 19165 1315 19185 1335
rect 19165 1265 19185 1285
rect 19165 1215 19185 1235
rect 19165 1165 19185 1185
rect 19165 1115 19185 1135
rect 19165 1065 19185 1085
rect 19165 1015 19185 1035
rect 19165 965 19185 985
rect 19165 915 19185 935
rect 20365 1565 20385 1585
rect 20365 1515 20385 1535
rect 20365 1465 20385 1485
rect 20365 1415 20385 1435
rect 20365 1365 20385 1385
rect 20365 1315 20385 1335
rect 20365 1265 20385 1285
rect 20365 1215 20385 1235
rect 20365 1165 20385 1185
rect 20365 1115 20385 1135
rect 20365 1065 20385 1085
rect 20365 1015 20385 1035
rect 20365 965 20385 985
rect 20365 915 20385 935
rect 21565 1565 21585 1585
rect 21565 1515 21585 1535
rect 21565 1465 21585 1485
rect 21565 1415 21585 1435
rect 21565 1365 21585 1385
rect 21565 1315 21585 1335
rect 21565 1265 21585 1285
rect 21565 1215 21585 1235
rect 21565 1165 21585 1185
rect 21565 1115 21585 1135
rect 21565 1065 21585 1085
rect 21565 1015 21585 1035
rect 21565 965 21585 985
rect 21565 915 21585 935
rect 22465 1565 22485 1585
rect 22465 1515 22485 1535
rect 22465 1465 22485 1485
rect 22465 1415 22485 1435
rect 22465 1365 22485 1385
rect 22465 1315 22485 1335
rect 22465 1265 22485 1285
rect 22465 1215 22485 1235
rect 22465 1165 22485 1185
rect 22465 1115 22485 1135
rect 22465 1065 22485 1085
rect 22465 1015 22485 1035
rect 22465 965 22485 985
rect 22465 915 22485 935
rect 23365 1565 23385 1585
rect 23365 1515 23385 1535
rect 23365 1465 23385 1485
rect 23365 1415 23385 1435
rect 23365 1365 23385 1385
rect 23365 1315 23385 1335
rect 23365 1265 23385 1285
rect 23365 1215 23385 1235
rect 23365 1165 23385 1185
rect 23365 1115 23385 1135
rect 23365 1065 23385 1085
rect 23365 1015 23385 1035
rect 23365 965 23385 985
rect 23365 915 23385 935
rect 24565 1565 24585 1585
rect 24565 1515 24585 1535
rect 24565 1465 24585 1485
rect 24565 1415 24585 1435
rect 24565 1365 24585 1385
rect 24565 1315 24585 1335
rect 24565 1265 24585 1285
rect 24565 1215 24585 1235
rect 24565 1165 24585 1185
rect 24565 1115 24585 1135
rect 24565 1065 24585 1085
rect 24565 1015 24585 1035
rect 24565 965 24585 985
rect 24565 915 24585 935
rect 25765 1565 25785 1585
rect 25765 1515 25785 1535
rect 25765 1465 25785 1485
rect 25765 1415 25785 1435
rect 25765 1365 25785 1385
rect 25765 1315 25785 1335
rect 25765 1265 25785 1285
rect 25765 1215 25785 1235
rect 25765 1165 25785 1185
rect 25765 1115 25785 1135
rect 25765 1065 25785 1085
rect 25765 1015 25785 1035
rect 25765 965 25785 985
rect 25765 915 25785 935
rect 26665 1565 26685 1585
rect 26665 1515 26685 1535
rect 26665 1465 26685 1485
rect 26665 1415 26685 1435
rect 26665 1365 26685 1385
rect 26665 1315 26685 1335
rect 26665 1265 26685 1285
rect 26665 1215 26685 1235
rect 26665 1165 26685 1185
rect 26665 1115 26685 1135
rect 26665 1065 26685 1085
rect 26665 1015 26685 1035
rect 26665 965 26685 985
rect 26665 915 26685 935
rect 27565 1565 27585 1585
rect 27565 1515 27585 1535
rect 27565 1465 27585 1485
rect 27565 1415 27585 1435
rect 27565 1365 27585 1385
rect 27565 1315 27585 1335
rect 27565 1265 27585 1285
rect 27565 1215 27585 1235
rect 27565 1165 27585 1185
rect 27565 1115 27585 1135
rect 27565 1065 27585 1085
rect 27565 1015 27585 1035
rect 27565 965 27585 985
rect 27565 915 27585 935
rect 28765 1565 28785 1585
rect 28765 1515 28785 1535
rect 28765 1465 28785 1485
rect 28765 1415 28785 1435
rect 28765 1365 28785 1385
rect 28765 1315 28785 1335
rect 28765 1265 28785 1285
rect 28765 1215 28785 1235
rect 28765 1165 28785 1185
rect 28765 1115 28785 1135
rect 28765 1065 28785 1085
rect 28765 1015 28785 1035
rect 28765 965 28785 985
rect 28765 915 28785 935
rect -635 715 -615 735
rect -635 665 -615 685
rect -635 615 -615 635
rect -635 565 -615 585
rect -635 515 -615 535
rect -635 465 -615 485
rect -635 415 -615 435
rect -635 365 -615 385
rect -635 315 -615 335
rect -635 265 -615 285
rect -635 215 -615 235
rect -635 165 -615 185
rect -635 115 -615 135
rect -635 65 -615 85
rect -485 715 -465 735
rect -485 665 -465 685
rect -485 615 -465 635
rect -485 565 -465 585
rect -485 515 -465 535
rect -485 465 -465 485
rect -485 415 -465 435
rect -485 365 -465 385
rect -485 315 -465 335
rect -485 265 -465 285
rect -485 215 -465 235
rect -485 165 -465 185
rect -485 115 -465 135
rect -485 65 -465 85
rect -335 715 -315 735
rect -335 665 -315 685
rect -335 615 -315 635
rect -335 565 -315 585
rect -335 515 -315 535
rect -335 465 -315 485
rect -335 415 -315 435
rect -335 365 -315 385
rect -335 315 -315 335
rect -335 265 -315 285
rect -335 215 -315 235
rect -335 165 -315 185
rect -335 115 -315 135
rect -335 65 -315 85
rect -185 715 -165 735
rect -185 665 -165 685
rect -185 615 -165 635
rect -185 565 -165 585
rect -185 515 -165 535
rect -185 465 -165 485
rect -185 415 -165 435
rect -185 365 -165 385
rect -185 315 -165 335
rect -185 265 -165 285
rect -185 215 -165 235
rect -185 165 -165 185
rect -185 115 -165 135
rect -185 65 -165 85
rect -35 715 -15 735
rect -35 665 -15 685
rect -35 615 -15 635
rect -35 565 -15 585
rect -35 515 -15 535
rect -35 465 -15 485
rect -35 415 -15 435
rect -35 365 -15 385
rect -35 315 -15 335
rect -35 265 -15 285
rect -35 215 -15 235
rect -35 165 -15 185
rect -35 115 -15 135
rect -35 65 -15 85
rect 1165 715 1185 735
rect 1165 665 1185 685
rect 1165 615 1185 635
rect 1165 565 1185 585
rect 1165 515 1185 535
rect 1165 465 1185 485
rect 1165 415 1185 435
rect 1165 365 1185 385
rect 1165 315 1185 335
rect 1165 265 1185 285
rect 1165 215 1185 235
rect 1165 165 1185 185
rect 1165 115 1185 135
rect 1165 65 1185 85
rect 1465 715 1485 735
rect 1465 665 1485 685
rect 1465 615 1485 635
rect 1465 565 1485 585
rect 1465 515 1485 535
rect 1465 465 1485 485
rect 1465 415 1485 435
rect 1465 365 1485 385
rect 1465 315 1485 335
rect 1465 265 1485 285
rect 1465 215 1485 235
rect 1465 165 1485 185
rect 1465 115 1485 135
rect 1465 65 1485 85
rect 1765 715 1785 735
rect 1765 665 1785 685
rect 1765 615 1785 635
rect 1765 565 1785 585
rect 1765 515 1785 535
rect 1765 465 1785 485
rect 1765 415 1785 435
rect 1765 365 1785 385
rect 1765 315 1785 335
rect 1765 265 1785 285
rect 1765 215 1785 235
rect 1765 165 1785 185
rect 1765 115 1785 135
rect 1765 65 1785 85
rect 2065 715 2085 735
rect 2065 665 2085 685
rect 2065 615 2085 635
rect 2065 565 2085 585
rect 2065 515 2085 535
rect 2065 465 2085 485
rect 2065 415 2085 435
rect 2065 365 2085 385
rect 2065 315 2085 335
rect 2065 265 2085 285
rect 2065 215 2085 235
rect 2065 165 2085 185
rect 2065 115 2085 135
rect 2065 65 2085 85
rect 2365 715 2385 735
rect 2365 665 2385 685
rect 2365 615 2385 635
rect 2365 565 2385 585
rect 2365 515 2385 535
rect 2365 465 2385 485
rect 2365 415 2385 435
rect 2365 365 2385 385
rect 2365 315 2385 335
rect 2365 265 2385 285
rect 2365 215 2385 235
rect 2365 165 2385 185
rect 2365 115 2385 135
rect 2365 65 2385 85
rect 2665 715 2685 735
rect 2665 665 2685 685
rect 2665 615 2685 635
rect 2665 565 2685 585
rect 2665 515 2685 535
rect 2665 465 2685 485
rect 2665 415 2685 435
rect 2665 365 2685 385
rect 2665 315 2685 335
rect 2665 265 2685 285
rect 2665 215 2685 235
rect 2665 165 2685 185
rect 2665 115 2685 135
rect 2665 65 2685 85
rect 2965 715 2985 735
rect 2965 665 2985 685
rect 2965 615 2985 635
rect 2965 565 2985 585
rect 2965 515 2985 535
rect 2965 465 2985 485
rect 2965 415 2985 435
rect 2965 365 2985 385
rect 2965 315 2985 335
rect 2965 265 2985 285
rect 2965 215 2985 235
rect 2965 165 2985 185
rect 2965 115 2985 135
rect 2965 65 2985 85
rect 3265 715 3285 735
rect 3265 665 3285 685
rect 3265 615 3285 635
rect 3265 565 3285 585
rect 3265 515 3285 535
rect 3265 465 3285 485
rect 3265 415 3285 435
rect 3265 365 3285 385
rect 3265 315 3285 335
rect 3265 265 3285 285
rect 3265 215 3285 235
rect 3265 165 3285 185
rect 3265 115 3285 135
rect 3265 65 3285 85
rect 3565 715 3585 735
rect 3565 665 3585 685
rect 3565 615 3585 635
rect 3565 565 3585 585
rect 3565 515 3585 535
rect 3565 465 3585 485
rect 3565 415 3585 435
rect 3565 365 3585 385
rect 3565 315 3585 335
rect 3565 265 3585 285
rect 3565 215 3585 235
rect 3565 165 3585 185
rect 3565 115 3585 135
rect 3565 65 3585 85
rect 3715 715 3735 735
rect 3715 665 3735 685
rect 3715 615 3735 635
rect 3715 565 3735 585
rect 3715 515 3735 535
rect 3715 465 3735 485
rect 3715 415 3735 435
rect 3715 365 3735 385
rect 3715 315 3735 335
rect 3715 265 3735 285
rect 3715 215 3735 235
rect 3715 165 3735 185
rect 3715 115 3735 135
rect 3715 65 3735 85
rect 3865 715 3885 735
rect 3865 665 3885 685
rect 3865 615 3885 635
rect 3865 565 3885 585
rect 3865 515 3885 535
rect 3865 465 3885 485
rect 3865 415 3885 435
rect 3865 365 3885 385
rect 3865 315 3885 335
rect 3865 265 3885 285
rect 3865 215 3885 235
rect 3865 165 3885 185
rect 3865 115 3885 135
rect 3865 65 3885 85
rect 4015 715 4035 735
rect 4015 665 4035 685
rect 4015 615 4035 635
rect 4015 565 4035 585
rect 4015 515 4035 535
rect 4015 465 4035 485
rect 4015 415 4035 435
rect 4015 365 4035 385
rect 4015 315 4035 335
rect 4015 265 4035 285
rect 4015 215 4035 235
rect 4015 165 4035 185
rect 4015 115 4035 135
rect 4015 65 4035 85
rect 4165 715 4185 735
rect 4165 665 4185 685
rect 4165 615 4185 635
rect 4165 565 4185 585
rect 4165 515 4185 535
rect 4165 465 4185 485
rect 4165 415 4185 435
rect 4165 365 4185 385
rect 4165 315 4185 335
rect 4165 265 4185 285
rect 4165 215 4185 235
rect 4165 165 4185 185
rect 4165 115 4185 135
rect 4165 65 4185 85
rect 4315 715 4335 735
rect 4315 665 4335 685
rect 4315 615 4335 635
rect 4315 565 4335 585
rect 4315 515 4335 535
rect 4315 465 4335 485
rect 4315 415 4335 435
rect 4315 365 4335 385
rect 4315 315 4335 335
rect 4315 265 4335 285
rect 4315 215 4335 235
rect 4315 165 4335 185
rect 4315 115 4335 135
rect 4315 65 4335 85
rect 4465 715 4485 735
rect 4465 665 4485 685
rect 4465 615 4485 635
rect 4465 565 4485 585
rect 4465 515 4485 535
rect 4465 465 4485 485
rect 4465 415 4485 435
rect 4465 365 4485 385
rect 4465 315 4485 335
rect 4465 265 4485 285
rect 4465 215 4485 235
rect 4465 165 4485 185
rect 4465 115 4485 135
rect 4465 65 4485 85
rect 4615 715 4635 735
rect 4615 665 4635 685
rect 4615 615 4635 635
rect 4615 565 4635 585
rect 4615 515 4635 535
rect 4615 465 4635 485
rect 4615 415 4635 435
rect 4615 365 4635 385
rect 4615 315 4635 335
rect 4615 265 4635 285
rect 4615 215 4635 235
rect 4615 165 4635 185
rect 4615 115 4635 135
rect 4615 65 4635 85
rect 4765 715 4785 735
rect 4765 665 4785 685
rect 4765 615 4785 635
rect 4765 565 4785 585
rect 4765 515 4785 535
rect 4765 465 4785 485
rect 4765 415 4785 435
rect 4765 365 4785 385
rect 4765 315 4785 335
rect 4765 265 4785 285
rect 4765 215 4785 235
rect 4765 165 4785 185
rect 4765 115 4785 135
rect 4765 65 4785 85
rect 5065 715 5085 735
rect 5065 665 5085 685
rect 5065 615 5085 635
rect 5065 565 5085 585
rect 5065 515 5085 535
rect 5065 465 5085 485
rect 5065 415 5085 435
rect 5065 365 5085 385
rect 5065 315 5085 335
rect 5065 265 5085 285
rect 5065 215 5085 235
rect 5065 165 5085 185
rect 5065 115 5085 135
rect 5065 65 5085 85
rect 5365 715 5385 735
rect 5365 665 5385 685
rect 5365 615 5385 635
rect 5365 565 5385 585
rect 5365 515 5385 535
rect 5365 465 5385 485
rect 5365 415 5385 435
rect 5365 365 5385 385
rect 5365 315 5385 335
rect 5365 265 5385 285
rect 5365 215 5385 235
rect 5365 165 5385 185
rect 5365 115 5385 135
rect 5365 65 5385 85
rect 5665 715 5685 735
rect 5665 665 5685 685
rect 5665 615 5685 635
rect 5665 565 5685 585
rect 5665 515 5685 535
rect 5665 465 5685 485
rect 5665 415 5685 435
rect 5665 365 5685 385
rect 5665 315 5685 335
rect 5665 265 5685 285
rect 5665 215 5685 235
rect 5665 165 5685 185
rect 5665 115 5685 135
rect 5665 65 5685 85
rect 5965 715 5985 735
rect 5965 665 5985 685
rect 5965 615 5985 635
rect 5965 565 5985 585
rect 5965 515 5985 535
rect 5965 465 5985 485
rect 5965 415 5985 435
rect 5965 365 5985 385
rect 5965 315 5985 335
rect 5965 265 5985 285
rect 5965 215 5985 235
rect 5965 165 5985 185
rect 5965 115 5985 135
rect 5965 65 5985 85
rect 6265 715 6285 735
rect 6265 665 6285 685
rect 6265 615 6285 635
rect 6265 565 6285 585
rect 6265 515 6285 535
rect 6265 465 6285 485
rect 6265 415 6285 435
rect 6265 365 6285 385
rect 6265 315 6285 335
rect 6265 265 6285 285
rect 6265 215 6285 235
rect 6265 165 6285 185
rect 6265 115 6285 135
rect 6265 65 6285 85
rect 6565 715 6585 735
rect 6565 665 6585 685
rect 6565 615 6585 635
rect 6565 565 6585 585
rect 6565 515 6585 535
rect 6565 465 6585 485
rect 6565 415 6585 435
rect 6565 365 6585 385
rect 6565 315 6585 335
rect 6565 265 6585 285
rect 6565 215 6585 235
rect 6565 165 6585 185
rect 6565 115 6585 135
rect 6565 65 6585 85
rect 6865 715 6885 735
rect 6865 665 6885 685
rect 6865 615 6885 635
rect 6865 565 6885 585
rect 6865 515 6885 535
rect 6865 465 6885 485
rect 6865 415 6885 435
rect 6865 365 6885 385
rect 6865 315 6885 335
rect 6865 265 6885 285
rect 6865 215 6885 235
rect 6865 165 6885 185
rect 6865 115 6885 135
rect 6865 65 6885 85
rect 7165 715 7185 735
rect 7165 665 7185 685
rect 7165 615 7185 635
rect 7165 565 7185 585
rect 7165 515 7185 535
rect 7165 465 7185 485
rect 7165 415 7185 435
rect 7165 365 7185 385
rect 7165 315 7185 335
rect 7165 265 7185 285
rect 7165 215 7185 235
rect 7165 165 7185 185
rect 7165 115 7185 135
rect 7165 65 7185 85
rect 8365 715 8385 735
rect 8365 665 8385 685
rect 8365 615 8385 635
rect 8365 565 8385 585
rect 8365 515 8385 535
rect 8365 465 8385 485
rect 8365 415 8385 435
rect 8365 365 8385 385
rect 8365 315 8385 335
rect 8365 265 8385 285
rect 8365 215 8385 235
rect 8365 165 8385 185
rect 8365 115 8385 135
rect 8365 65 8385 85
rect 9565 715 9585 735
rect 9565 665 9585 685
rect 9565 615 9585 635
rect 9565 565 9585 585
rect 9565 515 9585 535
rect 9565 465 9585 485
rect 9565 415 9585 435
rect 9565 365 9585 385
rect 9565 315 9585 335
rect 9565 265 9585 285
rect 9565 215 9585 235
rect 9565 165 9585 185
rect 9565 115 9585 135
rect 9565 65 9585 85
rect 10765 715 10785 735
rect 10765 665 10785 685
rect 10765 615 10785 635
rect 10765 565 10785 585
rect 10765 515 10785 535
rect 10765 465 10785 485
rect 10765 415 10785 435
rect 10765 365 10785 385
rect 10765 315 10785 335
rect 10765 265 10785 285
rect 10765 215 10785 235
rect 10765 165 10785 185
rect 10765 115 10785 135
rect 10765 65 10785 85
rect 11965 715 11985 735
rect 11965 665 11985 685
rect 11965 615 11985 635
rect 11965 565 11985 585
rect 11965 515 11985 535
rect 11965 465 11985 485
rect 11965 415 11985 435
rect 11965 365 11985 385
rect 11965 315 11985 335
rect 11965 265 11985 285
rect 11965 215 11985 235
rect 11965 165 11985 185
rect 11965 115 11985 135
rect 11965 65 11985 85
rect 12265 715 12285 735
rect 12265 665 12285 685
rect 12265 615 12285 635
rect 12265 565 12285 585
rect 12265 515 12285 535
rect 12265 465 12285 485
rect 12265 415 12285 435
rect 12265 365 12285 385
rect 12265 315 12285 335
rect 12265 265 12285 285
rect 12265 215 12285 235
rect 12265 165 12285 185
rect 12265 115 12285 135
rect 12265 65 12285 85
rect 12565 715 12585 735
rect 12565 665 12585 685
rect 12565 615 12585 635
rect 12565 565 12585 585
rect 12565 515 12585 535
rect 12565 465 12585 485
rect 12565 415 12585 435
rect 12565 365 12585 385
rect 12565 315 12585 335
rect 12565 265 12585 285
rect 12565 215 12585 235
rect 12565 165 12585 185
rect 12565 115 12585 135
rect 12565 65 12585 85
rect 12865 715 12885 735
rect 12865 665 12885 685
rect 12865 615 12885 635
rect 12865 565 12885 585
rect 12865 515 12885 535
rect 12865 465 12885 485
rect 12865 415 12885 435
rect 12865 365 12885 385
rect 12865 315 12885 335
rect 12865 265 12885 285
rect 12865 215 12885 235
rect 12865 165 12885 185
rect 12865 115 12885 135
rect 12865 65 12885 85
rect 13165 715 13185 735
rect 13165 665 13185 685
rect 13165 615 13185 635
rect 13165 565 13185 585
rect 13165 515 13185 535
rect 13165 465 13185 485
rect 13165 415 13185 435
rect 13165 365 13185 385
rect 13165 315 13185 335
rect 13165 265 13185 285
rect 13165 215 13185 235
rect 13165 165 13185 185
rect 13165 115 13185 135
rect 13165 65 13185 85
rect 13465 715 13485 735
rect 13465 665 13485 685
rect 13465 615 13485 635
rect 13465 565 13485 585
rect 13465 515 13485 535
rect 13465 465 13485 485
rect 13465 415 13485 435
rect 13465 365 13485 385
rect 13465 315 13485 335
rect 13465 265 13485 285
rect 13465 215 13485 235
rect 13465 165 13485 185
rect 13465 115 13485 135
rect 13465 65 13485 85
rect 13765 715 13785 735
rect 13765 665 13785 685
rect 13765 615 13785 635
rect 13765 565 13785 585
rect 13765 515 13785 535
rect 13765 465 13785 485
rect 13765 415 13785 435
rect 13765 365 13785 385
rect 13765 315 13785 335
rect 13765 265 13785 285
rect 13765 215 13785 235
rect 13765 165 13785 185
rect 13765 115 13785 135
rect 13765 65 13785 85
rect 14065 715 14085 735
rect 14065 665 14085 685
rect 14065 615 14085 635
rect 14065 565 14085 585
rect 14065 515 14085 535
rect 14065 465 14085 485
rect 14065 415 14085 435
rect 14065 365 14085 385
rect 14065 315 14085 335
rect 14065 265 14085 285
rect 14065 215 14085 235
rect 14065 165 14085 185
rect 14065 115 14085 135
rect 14065 65 14085 85
rect 14365 715 14385 735
rect 14365 665 14385 685
rect 14365 615 14385 635
rect 14365 565 14385 585
rect 14365 515 14385 535
rect 14365 465 14385 485
rect 14365 415 14385 435
rect 14365 365 14385 385
rect 14365 315 14385 335
rect 14365 265 14385 285
rect 14365 215 14385 235
rect 14365 165 14385 185
rect 14365 115 14385 135
rect 14365 65 14385 85
rect 15565 715 15585 735
rect 15565 665 15585 685
rect 15565 615 15585 635
rect 15565 565 15585 585
rect 15565 515 15585 535
rect 15565 465 15585 485
rect 15565 415 15585 435
rect 15565 365 15585 385
rect 15565 315 15585 335
rect 15565 265 15585 285
rect 15565 215 15585 235
rect 15565 165 15585 185
rect 15565 115 15585 135
rect 15565 65 15585 85
rect 16765 715 16785 735
rect 16765 665 16785 685
rect 16765 615 16785 635
rect 16765 565 16785 585
rect 16765 515 16785 535
rect 16765 465 16785 485
rect 16765 415 16785 435
rect 16765 365 16785 385
rect 16765 315 16785 335
rect 16765 265 16785 285
rect 16765 215 16785 235
rect 16765 165 16785 185
rect 16765 115 16785 135
rect 16765 65 16785 85
rect 17965 715 17985 735
rect 17965 665 17985 685
rect 17965 615 17985 635
rect 17965 565 17985 585
rect 17965 515 17985 535
rect 17965 465 17985 485
rect 17965 415 17985 435
rect 17965 365 17985 385
rect 17965 315 17985 335
rect 17965 265 17985 285
rect 17965 215 17985 235
rect 17965 165 17985 185
rect 17965 115 17985 135
rect 17965 65 17985 85
rect 19165 715 19185 735
rect 19165 665 19185 685
rect 19165 615 19185 635
rect 19165 565 19185 585
rect 19165 515 19185 535
rect 19165 465 19185 485
rect 19165 415 19185 435
rect 19165 365 19185 385
rect 19165 315 19185 335
rect 19165 265 19185 285
rect 19165 215 19185 235
rect 19165 165 19185 185
rect 19165 115 19185 135
rect 19165 65 19185 85
rect 20365 715 20385 735
rect 20365 665 20385 685
rect 20365 615 20385 635
rect 20365 565 20385 585
rect 20365 515 20385 535
rect 20365 465 20385 485
rect 20365 415 20385 435
rect 20365 365 20385 385
rect 20365 315 20385 335
rect 20365 265 20385 285
rect 20365 215 20385 235
rect 20365 165 20385 185
rect 20365 115 20385 135
rect 20365 65 20385 85
rect 21565 715 21585 735
rect 21565 665 21585 685
rect 21565 615 21585 635
rect 21565 565 21585 585
rect 21565 515 21585 535
rect 21565 465 21585 485
rect 21565 415 21585 435
rect 21565 365 21585 385
rect 21565 315 21585 335
rect 21565 265 21585 285
rect 21565 215 21585 235
rect 21565 165 21585 185
rect 21565 115 21585 135
rect 21565 65 21585 85
rect 22465 715 22485 735
rect 22465 665 22485 685
rect 22465 615 22485 635
rect 22465 565 22485 585
rect 22465 515 22485 535
rect 22465 465 22485 485
rect 22465 415 22485 435
rect 22465 365 22485 385
rect 22465 315 22485 335
rect 22465 265 22485 285
rect 22465 215 22485 235
rect 22465 165 22485 185
rect 22465 115 22485 135
rect 22465 65 22485 85
rect 23365 715 23385 735
rect 23365 665 23385 685
rect 23365 615 23385 635
rect 23365 565 23385 585
rect 23365 515 23385 535
rect 23365 465 23385 485
rect 23365 415 23385 435
rect 23365 365 23385 385
rect 23365 315 23385 335
rect 23365 265 23385 285
rect 23365 215 23385 235
rect 23365 165 23385 185
rect 23365 115 23385 135
rect 23365 65 23385 85
rect 24565 715 24585 735
rect 24565 665 24585 685
rect 24565 615 24585 635
rect 24565 565 24585 585
rect 24565 515 24585 535
rect 24565 465 24585 485
rect 24565 415 24585 435
rect 24565 365 24585 385
rect 24565 315 24585 335
rect 24565 265 24585 285
rect 24565 215 24585 235
rect 24565 165 24585 185
rect 24565 115 24585 135
rect 24565 65 24585 85
rect 25765 715 25785 735
rect 25765 665 25785 685
rect 25765 615 25785 635
rect 25765 565 25785 585
rect 25765 515 25785 535
rect 25765 465 25785 485
rect 25765 415 25785 435
rect 25765 365 25785 385
rect 25765 315 25785 335
rect 25765 265 25785 285
rect 25765 215 25785 235
rect 25765 165 25785 185
rect 25765 115 25785 135
rect 25765 65 25785 85
rect 26665 715 26685 735
rect 26665 665 26685 685
rect 26665 615 26685 635
rect 26665 565 26685 585
rect 26665 515 26685 535
rect 26665 465 26685 485
rect 26665 415 26685 435
rect 26665 365 26685 385
rect 26665 315 26685 335
rect 26665 265 26685 285
rect 26665 215 26685 235
rect 26665 165 26685 185
rect 26665 115 26685 135
rect 26665 65 26685 85
rect 27565 715 27585 735
rect 27565 665 27585 685
rect 27565 615 27585 635
rect 27565 565 27585 585
rect 27565 515 27585 535
rect 27565 465 27585 485
rect 27565 415 27585 435
rect 27565 365 27585 385
rect 27565 315 27585 335
rect 27565 265 27585 285
rect 27565 215 27585 235
rect 27565 165 27585 185
rect 27565 115 27585 135
rect 27565 65 27585 85
rect 28765 715 28785 735
rect 28765 665 28785 685
rect 28765 615 28785 635
rect 28765 565 28785 585
rect 28765 515 28785 535
rect 28765 465 28785 485
rect 28765 415 28785 435
rect 28765 365 28785 385
rect 28765 315 28785 335
rect 28765 265 28785 285
rect 28765 215 28785 235
rect 28765 165 28785 185
rect 28765 115 28785 135
rect 28765 65 28785 85
rect -635 -135 -615 -115
rect -635 -185 -615 -165
rect -635 -235 -615 -215
rect -635 -285 -615 -265
rect -635 -335 -615 -315
rect -635 -385 -615 -365
rect -635 -435 -615 -415
rect -635 -485 -615 -465
rect -635 -535 -615 -515
rect -635 -585 -615 -565
rect -635 -635 -615 -615
rect -635 -685 -615 -665
rect -635 -735 -615 -715
rect -635 -785 -615 -765
rect -485 -135 -465 -115
rect -485 -185 -465 -165
rect -485 -235 -465 -215
rect -485 -285 -465 -265
rect -485 -335 -465 -315
rect -485 -385 -465 -365
rect -485 -435 -465 -415
rect -485 -485 -465 -465
rect -485 -535 -465 -515
rect -485 -585 -465 -565
rect -485 -635 -465 -615
rect -485 -685 -465 -665
rect -485 -735 -465 -715
rect -485 -785 -465 -765
rect -335 -135 -315 -115
rect -335 -185 -315 -165
rect -335 -235 -315 -215
rect -335 -285 -315 -265
rect -335 -335 -315 -315
rect -335 -385 -315 -365
rect -335 -435 -315 -415
rect -335 -485 -315 -465
rect -335 -535 -315 -515
rect -335 -585 -315 -565
rect -335 -635 -315 -615
rect -335 -685 -315 -665
rect -335 -735 -315 -715
rect -335 -785 -315 -765
rect -185 -135 -165 -115
rect -185 -185 -165 -165
rect -185 -235 -165 -215
rect -185 -285 -165 -265
rect -185 -335 -165 -315
rect -185 -385 -165 -365
rect -185 -435 -165 -415
rect -185 -485 -165 -465
rect -185 -535 -165 -515
rect -185 -585 -165 -565
rect -185 -635 -165 -615
rect -185 -685 -165 -665
rect -185 -735 -165 -715
rect -185 -785 -165 -765
rect -35 -135 -15 -115
rect -35 -185 -15 -165
rect -35 -235 -15 -215
rect -35 -285 -15 -265
rect -35 -335 -15 -315
rect -35 -385 -15 -365
rect -35 -435 -15 -415
rect -35 -485 -15 -465
rect -35 -535 -15 -515
rect -35 -585 -15 -565
rect -35 -635 -15 -615
rect -35 -685 -15 -665
rect -35 -735 -15 -715
rect -35 -785 -15 -765
rect 1165 -135 1185 -115
rect 1165 -185 1185 -165
rect 1165 -235 1185 -215
rect 1165 -285 1185 -265
rect 1165 -335 1185 -315
rect 1165 -385 1185 -365
rect 1165 -435 1185 -415
rect 1165 -485 1185 -465
rect 1165 -535 1185 -515
rect 1165 -585 1185 -565
rect 1165 -635 1185 -615
rect 1165 -685 1185 -665
rect 1165 -735 1185 -715
rect 1165 -785 1185 -765
rect 1465 -135 1485 -115
rect 1465 -185 1485 -165
rect 1465 -235 1485 -215
rect 1465 -285 1485 -265
rect 1465 -335 1485 -315
rect 1465 -385 1485 -365
rect 1465 -435 1485 -415
rect 1465 -485 1485 -465
rect 1465 -535 1485 -515
rect 1465 -585 1485 -565
rect 1465 -635 1485 -615
rect 1465 -685 1485 -665
rect 1465 -735 1485 -715
rect 1465 -785 1485 -765
rect 1765 -135 1785 -115
rect 1765 -185 1785 -165
rect 1765 -235 1785 -215
rect 1765 -285 1785 -265
rect 1765 -335 1785 -315
rect 1765 -385 1785 -365
rect 1765 -435 1785 -415
rect 1765 -485 1785 -465
rect 1765 -535 1785 -515
rect 1765 -585 1785 -565
rect 1765 -635 1785 -615
rect 1765 -685 1785 -665
rect 1765 -735 1785 -715
rect 1765 -785 1785 -765
rect 2065 -135 2085 -115
rect 2065 -185 2085 -165
rect 2065 -235 2085 -215
rect 2065 -285 2085 -265
rect 2065 -335 2085 -315
rect 2065 -385 2085 -365
rect 2065 -435 2085 -415
rect 2065 -485 2085 -465
rect 2065 -535 2085 -515
rect 2065 -585 2085 -565
rect 2065 -635 2085 -615
rect 2065 -685 2085 -665
rect 2065 -735 2085 -715
rect 2065 -785 2085 -765
rect 2365 -135 2385 -115
rect 2365 -185 2385 -165
rect 2365 -235 2385 -215
rect 2365 -285 2385 -265
rect 2365 -335 2385 -315
rect 2365 -385 2385 -365
rect 2365 -435 2385 -415
rect 2365 -485 2385 -465
rect 2365 -535 2385 -515
rect 2365 -585 2385 -565
rect 2365 -635 2385 -615
rect 2365 -685 2385 -665
rect 2365 -735 2385 -715
rect 2365 -785 2385 -765
rect 2665 -135 2685 -115
rect 2665 -185 2685 -165
rect 2665 -235 2685 -215
rect 2665 -285 2685 -265
rect 2665 -335 2685 -315
rect 2665 -385 2685 -365
rect 2665 -435 2685 -415
rect 2665 -485 2685 -465
rect 2665 -535 2685 -515
rect 2665 -585 2685 -565
rect 2665 -635 2685 -615
rect 2665 -685 2685 -665
rect 2665 -735 2685 -715
rect 2665 -785 2685 -765
rect 2965 -135 2985 -115
rect 2965 -185 2985 -165
rect 2965 -235 2985 -215
rect 2965 -285 2985 -265
rect 2965 -335 2985 -315
rect 2965 -385 2985 -365
rect 2965 -435 2985 -415
rect 2965 -485 2985 -465
rect 2965 -535 2985 -515
rect 2965 -585 2985 -565
rect 2965 -635 2985 -615
rect 2965 -685 2985 -665
rect 2965 -735 2985 -715
rect 2965 -785 2985 -765
rect 3265 -135 3285 -115
rect 3265 -185 3285 -165
rect 3265 -235 3285 -215
rect 3265 -285 3285 -265
rect 3265 -335 3285 -315
rect 3265 -385 3285 -365
rect 3265 -435 3285 -415
rect 3265 -485 3285 -465
rect 3265 -535 3285 -515
rect 3265 -585 3285 -565
rect 3265 -635 3285 -615
rect 3265 -685 3285 -665
rect 3265 -735 3285 -715
rect 3265 -785 3285 -765
rect 3565 -135 3585 -115
rect 3565 -185 3585 -165
rect 3565 -235 3585 -215
rect 3565 -285 3585 -265
rect 3565 -335 3585 -315
rect 3565 -385 3585 -365
rect 3565 -435 3585 -415
rect 3565 -485 3585 -465
rect 3565 -535 3585 -515
rect 3565 -585 3585 -565
rect 3565 -635 3585 -615
rect 3565 -685 3585 -665
rect 3565 -735 3585 -715
rect 3565 -785 3585 -765
rect 3715 -135 3735 -115
rect 3715 -185 3735 -165
rect 3715 -235 3735 -215
rect 3715 -285 3735 -265
rect 3715 -335 3735 -315
rect 3715 -385 3735 -365
rect 3715 -435 3735 -415
rect 3715 -485 3735 -465
rect 3715 -535 3735 -515
rect 3715 -585 3735 -565
rect 3715 -635 3735 -615
rect 3715 -685 3735 -665
rect 3715 -735 3735 -715
rect 3715 -785 3735 -765
rect 3865 -135 3885 -115
rect 3865 -185 3885 -165
rect 3865 -235 3885 -215
rect 3865 -285 3885 -265
rect 3865 -335 3885 -315
rect 3865 -385 3885 -365
rect 3865 -435 3885 -415
rect 3865 -485 3885 -465
rect 3865 -535 3885 -515
rect 3865 -585 3885 -565
rect 3865 -635 3885 -615
rect 3865 -685 3885 -665
rect 3865 -735 3885 -715
rect 3865 -785 3885 -765
rect 4015 -135 4035 -115
rect 4015 -185 4035 -165
rect 4015 -235 4035 -215
rect 4015 -285 4035 -265
rect 4015 -335 4035 -315
rect 4015 -385 4035 -365
rect 4015 -435 4035 -415
rect 4015 -485 4035 -465
rect 4015 -535 4035 -515
rect 4015 -585 4035 -565
rect 4015 -635 4035 -615
rect 4015 -685 4035 -665
rect 4015 -735 4035 -715
rect 4015 -785 4035 -765
rect 4165 -135 4185 -115
rect 4165 -185 4185 -165
rect 4165 -235 4185 -215
rect 4165 -285 4185 -265
rect 4165 -335 4185 -315
rect 4165 -385 4185 -365
rect 4165 -435 4185 -415
rect 4165 -485 4185 -465
rect 4165 -535 4185 -515
rect 4165 -585 4185 -565
rect 4165 -635 4185 -615
rect 4165 -685 4185 -665
rect 4165 -735 4185 -715
rect 4165 -785 4185 -765
rect 4315 -135 4335 -115
rect 4315 -185 4335 -165
rect 4315 -235 4335 -215
rect 4315 -285 4335 -265
rect 4315 -335 4335 -315
rect 4315 -385 4335 -365
rect 4315 -435 4335 -415
rect 4315 -485 4335 -465
rect 4315 -535 4335 -515
rect 4315 -585 4335 -565
rect 4315 -635 4335 -615
rect 4315 -685 4335 -665
rect 4315 -735 4335 -715
rect 4315 -785 4335 -765
rect 4465 -135 4485 -115
rect 4465 -185 4485 -165
rect 4465 -235 4485 -215
rect 4465 -285 4485 -265
rect 4465 -335 4485 -315
rect 4465 -385 4485 -365
rect 4465 -435 4485 -415
rect 4465 -485 4485 -465
rect 4465 -535 4485 -515
rect 4465 -585 4485 -565
rect 4465 -635 4485 -615
rect 4465 -685 4485 -665
rect 4465 -735 4485 -715
rect 4465 -785 4485 -765
rect 4615 -135 4635 -115
rect 4615 -185 4635 -165
rect 4615 -235 4635 -215
rect 4615 -285 4635 -265
rect 4615 -335 4635 -315
rect 4615 -385 4635 -365
rect 4615 -435 4635 -415
rect 4615 -485 4635 -465
rect 4615 -535 4635 -515
rect 4615 -585 4635 -565
rect 4615 -635 4635 -615
rect 4615 -685 4635 -665
rect 4615 -735 4635 -715
rect 4615 -785 4635 -765
rect 4765 -135 4785 -115
rect 4765 -185 4785 -165
rect 4765 -235 4785 -215
rect 4765 -285 4785 -265
rect 4765 -335 4785 -315
rect 4765 -385 4785 -365
rect 4765 -435 4785 -415
rect 4765 -485 4785 -465
rect 4765 -535 4785 -515
rect 4765 -585 4785 -565
rect 4765 -635 4785 -615
rect 4765 -685 4785 -665
rect 4765 -735 4785 -715
rect 4765 -785 4785 -765
rect 5065 -135 5085 -115
rect 5065 -185 5085 -165
rect 5065 -235 5085 -215
rect 5065 -285 5085 -265
rect 5065 -335 5085 -315
rect 5065 -385 5085 -365
rect 5065 -435 5085 -415
rect 5065 -485 5085 -465
rect 5065 -535 5085 -515
rect 5065 -585 5085 -565
rect 5065 -635 5085 -615
rect 5065 -685 5085 -665
rect 5065 -735 5085 -715
rect 5065 -785 5085 -765
rect 5365 -135 5385 -115
rect 5365 -185 5385 -165
rect 5365 -235 5385 -215
rect 5365 -285 5385 -265
rect 5365 -335 5385 -315
rect 5365 -385 5385 -365
rect 5365 -435 5385 -415
rect 5365 -485 5385 -465
rect 5365 -535 5385 -515
rect 5365 -585 5385 -565
rect 5365 -635 5385 -615
rect 5365 -685 5385 -665
rect 5365 -735 5385 -715
rect 5365 -785 5385 -765
rect 5665 -135 5685 -115
rect 5665 -185 5685 -165
rect 5665 -235 5685 -215
rect 5665 -285 5685 -265
rect 5665 -335 5685 -315
rect 5665 -385 5685 -365
rect 5665 -435 5685 -415
rect 5665 -485 5685 -465
rect 5665 -535 5685 -515
rect 5665 -585 5685 -565
rect 5665 -635 5685 -615
rect 5665 -685 5685 -665
rect 5665 -735 5685 -715
rect 5665 -785 5685 -765
rect 5965 -135 5985 -115
rect 5965 -185 5985 -165
rect 5965 -235 5985 -215
rect 5965 -285 5985 -265
rect 5965 -335 5985 -315
rect 5965 -385 5985 -365
rect 5965 -435 5985 -415
rect 5965 -485 5985 -465
rect 5965 -535 5985 -515
rect 5965 -585 5985 -565
rect 5965 -635 5985 -615
rect 5965 -685 5985 -665
rect 5965 -735 5985 -715
rect 5965 -785 5985 -765
rect 6265 -135 6285 -115
rect 6265 -185 6285 -165
rect 6265 -235 6285 -215
rect 6265 -285 6285 -265
rect 6265 -335 6285 -315
rect 6265 -385 6285 -365
rect 6265 -435 6285 -415
rect 6265 -485 6285 -465
rect 6265 -535 6285 -515
rect 6265 -585 6285 -565
rect 6265 -635 6285 -615
rect 6265 -685 6285 -665
rect 6265 -735 6285 -715
rect 6265 -785 6285 -765
rect 6565 -135 6585 -115
rect 6565 -185 6585 -165
rect 6565 -235 6585 -215
rect 6565 -285 6585 -265
rect 6565 -335 6585 -315
rect 6565 -385 6585 -365
rect 6565 -435 6585 -415
rect 6565 -485 6585 -465
rect 6565 -535 6585 -515
rect 6565 -585 6585 -565
rect 6565 -635 6585 -615
rect 6565 -685 6585 -665
rect 6565 -735 6585 -715
rect 6565 -785 6585 -765
rect 6865 -135 6885 -115
rect 6865 -185 6885 -165
rect 6865 -235 6885 -215
rect 6865 -285 6885 -265
rect 6865 -335 6885 -315
rect 6865 -385 6885 -365
rect 6865 -435 6885 -415
rect 6865 -485 6885 -465
rect 6865 -535 6885 -515
rect 6865 -585 6885 -565
rect 6865 -635 6885 -615
rect 6865 -685 6885 -665
rect 6865 -735 6885 -715
rect 6865 -785 6885 -765
rect 7165 -135 7185 -115
rect 7165 -185 7185 -165
rect 7165 -235 7185 -215
rect 7165 -285 7185 -265
rect 7165 -335 7185 -315
rect 7165 -385 7185 -365
rect 7165 -435 7185 -415
rect 7165 -485 7185 -465
rect 7165 -535 7185 -515
rect 7165 -585 7185 -565
rect 7165 -635 7185 -615
rect 7165 -685 7185 -665
rect 7165 -735 7185 -715
rect 7165 -785 7185 -765
rect 8365 -135 8385 -115
rect 8365 -185 8385 -165
rect 8365 -235 8385 -215
rect 8365 -285 8385 -265
rect 8365 -335 8385 -315
rect 8365 -385 8385 -365
rect 8365 -435 8385 -415
rect 8365 -485 8385 -465
rect 8365 -535 8385 -515
rect 8365 -585 8385 -565
rect 8365 -635 8385 -615
rect 8365 -685 8385 -665
rect 8365 -735 8385 -715
rect 8365 -785 8385 -765
rect 9565 -135 9585 -115
rect 9565 -185 9585 -165
rect 9565 -235 9585 -215
rect 9565 -285 9585 -265
rect 9565 -335 9585 -315
rect 9565 -385 9585 -365
rect 9565 -435 9585 -415
rect 9565 -485 9585 -465
rect 9565 -535 9585 -515
rect 9565 -585 9585 -565
rect 9565 -635 9585 -615
rect 9565 -685 9585 -665
rect 9565 -735 9585 -715
rect 9565 -785 9585 -765
rect 10765 -135 10785 -115
rect 10765 -185 10785 -165
rect 10765 -235 10785 -215
rect 10765 -285 10785 -265
rect 10765 -335 10785 -315
rect 10765 -385 10785 -365
rect 10765 -435 10785 -415
rect 10765 -485 10785 -465
rect 10765 -535 10785 -515
rect 10765 -585 10785 -565
rect 10765 -635 10785 -615
rect 10765 -685 10785 -665
rect 10765 -735 10785 -715
rect 10765 -785 10785 -765
rect 11965 -135 11985 -115
rect 11965 -185 11985 -165
rect 11965 -235 11985 -215
rect 11965 -285 11985 -265
rect 11965 -335 11985 -315
rect 11965 -385 11985 -365
rect 11965 -435 11985 -415
rect 11965 -485 11985 -465
rect 11965 -535 11985 -515
rect 11965 -585 11985 -565
rect 11965 -635 11985 -615
rect 11965 -685 11985 -665
rect 11965 -735 11985 -715
rect 11965 -785 11985 -765
rect 12265 -135 12285 -115
rect 12265 -185 12285 -165
rect 12265 -235 12285 -215
rect 12265 -285 12285 -265
rect 12265 -335 12285 -315
rect 12265 -385 12285 -365
rect 12265 -435 12285 -415
rect 12265 -485 12285 -465
rect 12265 -535 12285 -515
rect 12265 -585 12285 -565
rect 12265 -635 12285 -615
rect 12265 -685 12285 -665
rect 12265 -735 12285 -715
rect 12265 -785 12285 -765
rect 12565 -135 12585 -115
rect 12565 -185 12585 -165
rect 12565 -235 12585 -215
rect 12565 -285 12585 -265
rect 12565 -335 12585 -315
rect 12565 -385 12585 -365
rect 12565 -435 12585 -415
rect 12565 -485 12585 -465
rect 12565 -535 12585 -515
rect 12565 -585 12585 -565
rect 12565 -635 12585 -615
rect 12565 -685 12585 -665
rect 12565 -735 12585 -715
rect 12565 -785 12585 -765
rect 12865 -135 12885 -115
rect 12865 -185 12885 -165
rect 12865 -235 12885 -215
rect 12865 -285 12885 -265
rect 12865 -335 12885 -315
rect 12865 -385 12885 -365
rect 12865 -435 12885 -415
rect 12865 -485 12885 -465
rect 12865 -535 12885 -515
rect 12865 -585 12885 -565
rect 12865 -635 12885 -615
rect 12865 -685 12885 -665
rect 12865 -735 12885 -715
rect 12865 -785 12885 -765
rect 13165 -135 13185 -115
rect 13165 -185 13185 -165
rect 13165 -235 13185 -215
rect 13165 -285 13185 -265
rect 13165 -335 13185 -315
rect 13165 -385 13185 -365
rect 13165 -435 13185 -415
rect 13165 -485 13185 -465
rect 13165 -535 13185 -515
rect 13165 -585 13185 -565
rect 13165 -635 13185 -615
rect 13165 -685 13185 -665
rect 13165 -735 13185 -715
rect 13165 -785 13185 -765
rect 13465 -135 13485 -115
rect 13465 -185 13485 -165
rect 13465 -235 13485 -215
rect 13465 -285 13485 -265
rect 13465 -335 13485 -315
rect 13465 -385 13485 -365
rect 13465 -435 13485 -415
rect 13465 -485 13485 -465
rect 13465 -535 13485 -515
rect 13465 -585 13485 -565
rect 13465 -635 13485 -615
rect 13465 -685 13485 -665
rect 13465 -735 13485 -715
rect 13465 -785 13485 -765
rect 13765 -135 13785 -115
rect 13765 -185 13785 -165
rect 13765 -235 13785 -215
rect 13765 -285 13785 -265
rect 13765 -335 13785 -315
rect 13765 -385 13785 -365
rect 13765 -435 13785 -415
rect 13765 -485 13785 -465
rect 13765 -535 13785 -515
rect 13765 -585 13785 -565
rect 13765 -635 13785 -615
rect 13765 -685 13785 -665
rect 13765 -735 13785 -715
rect 13765 -785 13785 -765
rect 14065 -135 14085 -115
rect 14065 -185 14085 -165
rect 14065 -235 14085 -215
rect 14065 -285 14085 -265
rect 14065 -335 14085 -315
rect 14065 -385 14085 -365
rect 14065 -435 14085 -415
rect 14065 -485 14085 -465
rect 14065 -535 14085 -515
rect 14065 -585 14085 -565
rect 14065 -635 14085 -615
rect 14065 -685 14085 -665
rect 14065 -735 14085 -715
rect 14065 -785 14085 -765
rect 14365 -135 14385 -115
rect 14365 -185 14385 -165
rect 14365 -235 14385 -215
rect 14365 -285 14385 -265
rect 14365 -335 14385 -315
rect 14365 -385 14385 -365
rect 14365 -435 14385 -415
rect 14365 -485 14385 -465
rect 14365 -535 14385 -515
rect 14365 -585 14385 -565
rect 14365 -635 14385 -615
rect 14365 -685 14385 -665
rect 14365 -735 14385 -715
rect 14365 -785 14385 -765
rect 15565 -135 15585 -115
rect 15565 -185 15585 -165
rect 15565 -235 15585 -215
rect 15565 -285 15585 -265
rect 15565 -335 15585 -315
rect 15565 -385 15585 -365
rect 15565 -435 15585 -415
rect 15565 -485 15585 -465
rect 15565 -535 15585 -515
rect 15565 -585 15585 -565
rect 15565 -635 15585 -615
rect 15565 -685 15585 -665
rect 15565 -735 15585 -715
rect 15565 -785 15585 -765
rect 16765 -135 16785 -115
rect 16765 -185 16785 -165
rect 16765 -235 16785 -215
rect 16765 -285 16785 -265
rect 16765 -335 16785 -315
rect 16765 -385 16785 -365
rect 16765 -435 16785 -415
rect 16765 -485 16785 -465
rect 16765 -535 16785 -515
rect 16765 -585 16785 -565
rect 16765 -635 16785 -615
rect 16765 -685 16785 -665
rect 16765 -735 16785 -715
rect 16765 -785 16785 -765
rect 17965 -135 17985 -115
rect 17965 -185 17985 -165
rect 17965 -235 17985 -215
rect 17965 -285 17985 -265
rect 17965 -335 17985 -315
rect 17965 -385 17985 -365
rect 17965 -435 17985 -415
rect 17965 -485 17985 -465
rect 17965 -535 17985 -515
rect 17965 -585 17985 -565
rect 17965 -635 17985 -615
rect 17965 -685 17985 -665
rect 17965 -735 17985 -715
rect 17965 -785 17985 -765
rect 19165 -135 19185 -115
rect 19165 -185 19185 -165
rect 19165 -235 19185 -215
rect 19165 -285 19185 -265
rect 19165 -335 19185 -315
rect 19165 -385 19185 -365
rect 19165 -435 19185 -415
rect 19165 -485 19185 -465
rect 19165 -535 19185 -515
rect 19165 -585 19185 -565
rect 19165 -635 19185 -615
rect 19165 -685 19185 -665
rect 19165 -735 19185 -715
rect 19165 -785 19185 -765
rect 20365 -135 20385 -115
rect 20365 -185 20385 -165
rect 20365 -235 20385 -215
rect 20365 -285 20385 -265
rect 20365 -335 20385 -315
rect 20365 -385 20385 -365
rect 20365 -435 20385 -415
rect 20365 -485 20385 -465
rect 20365 -535 20385 -515
rect 20365 -585 20385 -565
rect 20365 -635 20385 -615
rect 20365 -685 20385 -665
rect 20365 -735 20385 -715
rect 20365 -785 20385 -765
rect 21565 -135 21585 -115
rect 21565 -185 21585 -165
rect 21565 -235 21585 -215
rect 21565 -285 21585 -265
rect 21565 -335 21585 -315
rect 21565 -385 21585 -365
rect 21565 -435 21585 -415
rect 21565 -485 21585 -465
rect 21565 -535 21585 -515
rect 21565 -585 21585 -565
rect 21565 -635 21585 -615
rect 21565 -685 21585 -665
rect 21565 -735 21585 -715
rect 21565 -785 21585 -765
rect 22465 -135 22485 -115
rect 22465 -185 22485 -165
rect 22465 -235 22485 -215
rect 22465 -285 22485 -265
rect 22465 -335 22485 -315
rect 22465 -385 22485 -365
rect 22465 -435 22485 -415
rect 22465 -485 22485 -465
rect 22465 -535 22485 -515
rect 22465 -585 22485 -565
rect 22465 -635 22485 -615
rect 22465 -685 22485 -665
rect 22465 -735 22485 -715
rect 22465 -785 22485 -765
rect 23365 -135 23385 -115
rect 23365 -185 23385 -165
rect 23365 -235 23385 -215
rect 23365 -285 23385 -265
rect 23365 -335 23385 -315
rect 23365 -385 23385 -365
rect 23365 -435 23385 -415
rect 23365 -485 23385 -465
rect 23365 -535 23385 -515
rect 23365 -585 23385 -565
rect 23365 -635 23385 -615
rect 23365 -685 23385 -665
rect 23365 -735 23385 -715
rect 23365 -785 23385 -765
rect 24565 -135 24585 -115
rect 24565 -185 24585 -165
rect 24565 -235 24585 -215
rect 24565 -285 24585 -265
rect 24565 -335 24585 -315
rect 24565 -385 24585 -365
rect 24565 -435 24585 -415
rect 24565 -485 24585 -465
rect 24565 -535 24585 -515
rect 24565 -585 24585 -565
rect 24565 -635 24585 -615
rect 24565 -685 24585 -665
rect 24565 -735 24585 -715
rect 24565 -785 24585 -765
rect 25765 -135 25785 -115
rect 25765 -185 25785 -165
rect 25765 -235 25785 -215
rect 25765 -285 25785 -265
rect 25765 -335 25785 -315
rect 25765 -385 25785 -365
rect 25765 -435 25785 -415
rect 25765 -485 25785 -465
rect 25765 -535 25785 -515
rect 25765 -585 25785 -565
rect 25765 -635 25785 -615
rect 25765 -685 25785 -665
rect 25765 -735 25785 -715
rect 25765 -785 25785 -765
rect 26665 -135 26685 -115
rect 26665 -185 26685 -165
rect 26665 -235 26685 -215
rect 26665 -285 26685 -265
rect 26665 -335 26685 -315
rect 26665 -385 26685 -365
rect 26665 -435 26685 -415
rect 26665 -485 26685 -465
rect 26665 -535 26685 -515
rect 26665 -585 26685 -565
rect 26665 -635 26685 -615
rect 26665 -685 26685 -665
rect 26665 -735 26685 -715
rect 26665 -785 26685 -765
rect 27565 -135 27585 -115
rect 27565 -185 27585 -165
rect 27565 -235 27585 -215
rect 27565 -285 27585 -265
rect 27565 -335 27585 -315
rect 27565 -385 27585 -365
rect 27565 -435 27585 -415
rect 27565 -485 27585 -465
rect 27565 -535 27585 -515
rect 27565 -585 27585 -565
rect 27565 -635 27585 -615
rect 27565 -685 27585 -665
rect 27565 -735 27585 -715
rect 27565 -785 27585 -765
rect 28765 -135 28785 -115
rect 28765 -185 28785 -165
rect 28765 -235 28785 -215
rect 28765 -285 28785 -265
rect 28765 -335 28785 -315
rect 28765 -385 28785 -365
rect 28765 -435 28785 -415
rect 28765 -485 28785 -465
rect 28765 -535 28785 -515
rect 28765 -585 28785 -565
rect 28765 -635 28785 -615
rect 28765 -685 28785 -665
rect 28765 -735 28785 -715
rect 28765 -785 28785 -765
rect -635 -985 -615 -965
rect -635 -1035 -615 -1015
rect -635 -1085 -615 -1065
rect -635 -1135 -615 -1115
rect -635 -1185 -615 -1165
rect -635 -1235 -615 -1215
rect -635 -1285 -615 -1265
rect -635 -1335 -615 -1315
rect -635 -1385 -615 -1365
rect -635 -1435 -615 -1415
rect -635 -1485 -615 -1465
rect -635 -1535 -615 -1515
rect -635 -1585 -615 -1565
rect -635 -1635 -615 -1615
rect -485 -985 -465 -965
rect -485 -1035 -465 -1015
rect -485 -1085 -465 -1065
rect -485 -1135 -465 -1115
rect -485 -1185 -465 -1165
rect -485 -1235 -465 -1215
rect -485 -1285 -465 -1265
rect -485 -1335 -465 -1315
rect -485 -1385 -465 -1365
rect -485 -1435 -465 -1415
rect -485 -1485 -465 -1465
rect -485 -1535 -465 -1515
rect -485 -1585 -465 -1565
rect -485 -1635 -465 -1615
rect -335 -985 -315 -965
rect -335 -1035 -315 -1015
rect -335 -1085 -315 -1065
rect -335 -1135 -315 -1115
rect -335 -1185 -315 -1165
rect -335 -1235 -315 -1215
rect -335 -1285 -315 -1265
rect -335 -1335 -315 -1315
rect -335 -1385 -315 -1365
rect -335 -1435 -315 -1415
rect -335 -1485 -315 -1465
rect -335 -1535 -315 -1515
rect -335 -1585 -315 -1565
rect -335 -1635 -315 -1615
rect -185 -985 -165 -965
rect -185 -1035 -165 -1015
rect -185 -1085 -165 -1065
rect -185 -1135 -165 -1115
rect -185 -1185 -165 -1165
rect -185 -1235 -165 -1215
rect -185 -1285 -165 -1265
rect -185 -1335 -165 -1315
rect -185 -1385 -165 -1365
rect -185 -1435 -165 -1415
rect -185 -1485 -165 -1465
rect -185 -1535 -165 -1515
rect -185 -1585 -165 -1565
rect -185 -1635 -165 -1615
rect -35 -985 -15 -965
rect -35 -1035 -15 -1015
rect -35 -1085 -15 -1065
rect -35 -1135 -15 -1115
rect -35 -1185 -15 -1165
rect -35 -1235 -15 -1215
rect -35 -1285 -15 -1265
rect -35 -1335 -15 -1315
rect -35 -1385 -15 -1365
rect -35 -1435 -15 -1415
rect -35 -1485 -15 -1465
rect -35 -1535 -15 -1515
rect -35 -1585 -15 -1565
rect -35 -1635 -15 -1615
rect 1165 -985 1185 -965
rect 1165 -1035 1185 -1015
rect 1165 -1085 1185 -1065
rect 1165 -1135 1185 -1115
rect 1165 -1185 1185 -1165
rect 1165 -1235 1185 -1215
rect 1165 -1285 1185 -1265
rect 1165 -1335 1185 -1315
rect 1165 -1385 1185 -1365
rect 1165 -1435 1185 -1415
rect 1165 -1485 1185 -1465
rect 1165 -1535 1185 -1515
rect 1165 -1585 1185 -1565
rect 1165 -1635 1185 -1615
rect 1465 -985 1485 -965
rect 1465 -1035 1485 -1015
rect 1465 -1085 1485 -1065
rect 1465 -1135 1485 -1115
rect 1465 -1185 1485 -1165
rect 1465 -1235 1485 -1215
rect 1465 -1285 1485 -1265
rect 1465 -1335 1485 -1315
rect 1465 -1385 1485 -1365
rect 1465 -1435 1485 -1415
rect 1465 -1485 1485 -1465
rect 1465 -1535 1485 -1515
rect 1465 -1585 1485 -1565
rect 1465 -1635 1485 -1615
rect 1765 -985 1785 -965
rect 1765 -1035 1785 -1015
rect 1765 -1085 1785 -1065
rect 1765 -1135 1785 -1115
rect 1765 -1185 1785 -1165
rect 1765 -1235 1785 -1215
rect 1765 -1285 1785 -1265
rect 1765 -1335 1785 -1315
rect 1765 -1385 1785 -1365
rect 1765 -1435 1785 -1415
rect 1765 -1485 1785 -1465
rect 1765 -1535 1785 -1515
rect 1765 -1585 1785 -1565
rect 1765 -1635 1785 -1615
rect 2065 -985 2085 -965
rect 2065 -1035 2085 -1015
rect 2065 -1085 2085 -1065
rect 2065 -1135 2085 -1115
rect 2065 -1185 2085 -1165
rect 2065 -1235 2085 -1215
rect 2065 -1285 2085 -1265
rect 2065 -1335 2085 -1315
rect 2065 -1385 2085 -1365
rect 2065 -1435 2085 -1415
rect 2065 -1485 2085 -1465
rect 2065 -1535 2085 -1515
rect 2065 -1585 2085 -1565
rect 2065 -1635 2085 -1615
rect 2365 -985 2385 -965
rect 2365 -1035 2385 -1015
rect 2365 -1085 2385 -1065
rect 2365 -1135 2385 -1115
rect 2365 -1185 2385 -1165
rect 2365 -1235 2385 -1215
rect 2365 -1285 2385 -1265
rect 2365 -1335 2385 -1315
rect 2365 -1385 2385 -1365
rect 2365 -1435 2385 -1415
rect 2365 -1485 2385 -1465
rect 2365 -1535 2385 -1515
rect 2365 -1585 2385 -1565
rect 2365 -1635 2385 -1615
rect 2665 -985 2685 -965
rect 2665 -1035 2685 -1015
rect 2665 -1085 2685 -1065
rect 2665 -1135 2685 -1115
rect 2665 -1185 2685 -1165
rect 2665 -1235 2685 -1215
rect 2665 -1285 2685 -1265
rect 2665 -1335 2685 -1315
rect 2665 -1385 2685 -1365
rect 2665 -1435 2685 -1415
rect 2665 -1485 2685 -1465
rect 2665 -1535 2685 -1515
rect 2665 -1585 2685 -1565
rect 2665 -1635 2685 -1615
rect 2965 -985 2985 -965
rect 2965 -1035 2985 -1015
rect 2965 -1085 2985 -1065
rect 2965 -1135 2985 -1115
rect 2965 -1185 2985 -1165
rect 2965 -1235 2985 -1215
rect 2965 -1285 2985 -1265
rect 2965 -1335 2985 -1315
rect 2965 -1385 2985 -1365
rect 2965 -1435 2985 -1415
rect 2965 -1485 2985 -1465
rect 2965 -1535 2985 -1515
rect 2965 -1585 2985 -1565
rect 2965 -1635 2985 -1615
rect 3265 -985 3285 -965
rect 3265 -1035 3285 -1015
rect 3265 -1085 3285 -1065
rect 3265 -1135 3285 -1115
rect 3265 -1185 3285 -1165
rect 3265 -1235 3285 -1215
rect 3265 -1285 3285 -1265
rect 3265 -1335 3285 -1315
rect 3265 -1385 3285 -1365
rect 3265 -1435 3285 -1415
rect 3265 -1485 3285 -1465
rect 3265 -1535 3285 -1515
rect 3265 -1585 3285 -1565
rect 3265 -1635 3285 -1615
rect 3565 -985 3585 -965
rect 3565 -1035 3585 -1015
rect 3565 -1085 3585 -1065
rect 3565 -1135 3585 -1115
rect 3565 -1185 3585 -1165
rect 3565 -1235 3585 -1215
rect 3565 -1285 3585 -1265
rect 3565 -1335 3585 -1315
rect 3565 -1385 3585 -1365
rect 3565 -1435 3585 -1415
rect 3565 -1485 3585 -1465
rect 3565 -1535 3585 -1515
rect 3565 -1585 3585 -1565
rect 3565 -1635 3585 -1615
rect 3715 -985 3735 -965
rect 3715 -1035 3735 -1015
rect 3715 -1085 3735 -1065
rect 3715 -1135 3735 -1115
rect 3715 -1185 3735 -1165
rect 3715 -1235 3735 -1215
rect 3715 -1285 3735 -1265
rect 3715 -1335 3735 -1315
rect 3715 -1385 3735 -1365
rect 3715 -1435 3735 -1415
rect 3715 -1485 3735 -1465
rect 3715 -1535 3735 -1515
rect 3715 -1585 3735 -1565
rect 3715 -1635 3735 -1615
rect 3865 -985 3885 -965
rect 3865 -1035 3885 -1015
rect 3865 -1085 3885 -1065
rect 3865 -1135 3885 -1115
rect 3865 -1185 3885 -1165
rect 3865 -1235 3885 -1215
rect 3865 -1285 3885 -1265
rect 3865 -1335 3885 -1315
rect 3865 -1385 3885 -1365
rect 3865 -1435 3885 -1415
rect 3865 -1485 3885 -1465
rect 3865 -1535 3885 -1515
rect 3865 -1585 3885 -1565
rect 3865 -1635 3885 -1615
rect 4015 -985 4035 -965
rect 4015 -1035 4035 -1015
rect 4015 -1085 4035 -1065
rect 4015 -1135 4035 -1115
rect 4015 -1185 4035 -1165
rect 4015 -1235 4035 -1215
rect 4015 -1285 4035 -1265
rect 4015 -1335 4035 -1315
rect 4015 -1385 4035 -1365
rect 4015 -1435 4035 -1415
rect 4015 -1485 4035 -1465
rect 4015 -1535 4035 -1515
rect 4015 -1585 4035 -1565
rect 4015 -1635 4035 -1615
rect 4165 -985 4185 -965
rect 4165 -1035 4185 -1015
rect 4165 -1085 4185 -1065
rect 4165 -1135 4185 -1115
rect 4165 -1185 4185 -1165
rect 4165 -1235 4185 -1215
rect 4165 -1285 4185 -1265
rect 4165 -1335 4185 -1315
rect 4165 -1385 4185 -1365
rect 4165 -1435 4185 -1415
rect 4165 -1485 4185 -1465
rect 4165 -1535 4185 -1515
rect 4165 -1585 4185 -1565
rect 4165 -1635 4185 -1615
rect 4315 -985 4335 -965
rect 4315 -1035 4335 -1015
rect 4315 -1085 4335 -1065
rect 4315 -1135 4335 -1115
rect 4315 -1185 4335 -1165
rect 4315 -1235 4335 -1215
rect 4315 -1285 4335 -1265
rect 4315 -1335 4335 -1315
rect 4315 -1385 4335 -1365
rect 4315 -1435 4335 -1415
rect 4315 -1485 4335 -1465
rect 4315 -1535 4335 -1515
rect 4315 -1585 4335 -1565
rect 4315 -1635 4335 -1615
rect 4465 -985 4485 -965
rect 4465 -1035 4485 -1015
rect 4465 -1085 4485 -1065
rect 4465 -1135 4485 -1115
rect 4465 -1185 4485 -1165
rect 4465 -1235 4485 -1215
rect 4465 -1285 4485 -1265
rect 4465 -1335 4485 -1315
rect 4465 -1385 4485 -1365
rect 4465 -1435 4485 -1415
rect 4465 -1485 4485 -1465
rect 4465 -1535 4485 -1515
rect 4465 -1585 4485 -1565
rect 4465 -1635 4485 -1615
rect 4615 -985 4635 -965
rect 4615 -1035 4635 -1015
rect 4615 -1085 4635 -1065
rect 4615 -1135 4635 -1115
rect 4615 -1185 4635 -1165
rect 4615 -1235 4635 -1215
rect 4615 -1285 4635 -1265
rect 4615 -1335 4635 -1315
rect 4615 -1385 4635 -1365
rect 4615 -1435 4635 -1415
rect 4615 -1485 4635 -1465
rect 4615 -1535 4635 -1515
rect 4615 -1585 4635 -1565
rect 4615 -1635 4635 -1615
rect 4765 -985 4785 -965
rect 4765 -1035 4785 -1015
rect 4765 -1085 4785 -1065
rect 4765 -1135 4785 -1115
rect 4765 -1185 4785 -1165
rect 4765 -1235 4785 -1215
rect 4765 -1285 4785 -1265
rect 4765 -1335 4785 -1315
rect 4765 -1385 4785 -1365
rect 4765 -1435 4785 -1415
rect 4765 -1485 4785 -1465
rect 4765 -1535 4785 -1515
rect 4765 -1585 4785 -1565
rect 4765 -1635 4785 -1615
rect 5065 -985 5085 -965
rect 5065 -1035 5085 -1015
rect 5065 -1085 5085 -1065
rect 5065 -1135 5085 -1115
rect 5065 -1185 5085 -1165
rect 5065 -1235 5085 -1215
rect 5065 -1285 5085 -1265
rect 5065 -1335 5085 -1315
rect 5065 -1385 5085 -1365
rect 5065 -1435 5085 -1415
rect 5065 -1485 5085 -1465
rect 5065 -1535 5085 -1515
rect 5065 -1585 5085 -1565
rect 5065 -1635 5085 -1615
rect 5365 -985 5385 -965
rect 5365 -1035 5385 -1015
rect 5365 -1085 5385 -1065
rect 5365 -1135 5385 -1115
rect 5365 -1185 5385 -1165
rect 5365 -1235 5385 -1215
rect 5365 -1285 5385 -1265
rect 5365 -1335 5385 -1315
rect 5365 -1385 5385 -1365
rect 5365 -1435 5385 -1415
rect 5365 -1485 5385 -1465
rect 5365 -1535 5385 -1515
rect 5365 -1585 5385 -1565
rect 5365 -1635 5385 -1615
rect 5665 -985 5685 -965
rect 5665 -1035 5685 -1015
rect 5665 -1085 5685 -1065
rect 5665 -1135 5685 -1115
rect 5665 -1185 5685 -1165
rect 5665 -1235 5685 -1215
rect 5665 -1285 5685 -1265
rect 5665 -1335 5685 -1315
rect 5665 -1385 5685 -1365
rect 5665 -1435 5685 -1415
rect 5665 -1485 5685 -1465
rect 5665 -1535 5685 -1515
rect 5665 -1585 5685 -1565
rect 5665 -1635 5685 -1615
rect 5965 -985 5985 -965
rect 5965 -1035 5985 -1015
rect 5965 -1085 5985 -1065
rect 5965 -1135 5985 -1115
rect 5965 -1185 5985 -1165
rect 5965 -1235 5985 -1215
rect 5965 -1285 5985 -1265
rect 5965 -1335 5985 -1315
rect 5965 -1385 5985 -1365
rect 5965 -1435 5985 -1415
rect 5965 -1485 5985 -1465
rect 5965 -1535 5985 -1515
rect 5965 -1585 5985 -1565
rect 5965 -1635 5985 -1615
rect 6265 -985 6285 -965
rect 6265 -1035 6285 -1015
rect 6265 -1085 6285 -1065
rect 6265 -1135 6285 -1115
rect 6265 -1185 6285 -1165
rect 6265 -1235 6285 -1215
rect 6265 -1285 6285 -1265
rect 6265 -1335 6285 -1315
rect 6265 -1385 6285 -1365
rect 6265 -1435 6285 -1415
rect 6265 -1485 6285 -1465
rect 6265 -1535 6285 -1515
rect 6265 -1585 6285 -1565
rect 6265 -1635 6285 -1615
rect 6565 -985 6585 -965
rect 6565 -1035 6585 -1015
rect 6565 -1085 6585 -1065
rect 6565 -1135 6585 -1115
rect 6565 -1185 6585 -1165
rect 6565 -1235 6585 -1215
rect 6565 -1285 6585 -1265
rect 6565 -1335 6585 -1315
rect 6565 -1385 6585 -1365
rect 6565 -1435 6585 -1415
rect 6565 -1485 6585 -1465
rect 6565 -1535 6585 -1515
rect 6565 -1585 6585 -1565
rect 6565 -1635 6585 -1615
rect 6865 -985 6885 -965
rect 6865 -1035 6885 -1015
rect 6865 -1085 6885 -1065
rect 6865 -1135 6885 -1115
rect 6865 -1185 6885 -1165
rect 6865 -1235 6885 -1215
rect 6865 -1285 6885 -1265
rect 6865 -1335 6885 -1315
rect 6865 -1385 6885 -1365
rect 6865 -1435 6885 -1415
rect 6865 -1485 6885 -1465
rect 6865 -1535 6885 -1515
rect 6865 -1585 6885 -1565
rect 6865 -1635 6885 -1615
rect 7165 -985 7185 -965
rect 7165 -1035 7185 -1015
rect 7165 -1085 7185 -1065
rect 7165 -1135 7185 -1115
rect 7165 -1185 7185 -1165
rect 7165 -1235 7185 -1215
rect 7165 -1285 7185 -1265
rect 7165 -1335 7185 -1315
rect 7165 -1385 7185 -1365
rect 7165 -1435 7185 -1415
rect 7165 -1485 7185 -1465
rect 7165 -1535 7185 -1515
rect 7165 -1585 7185 -1565
rect 7165 -1635 7185 -1615
rect 8365 -985 8385 -965
rect 8365 -1035 8385 -1015
rect 8365 -1085 8385 -1065
rect 8365 -1135 8385 -1115
rect 8365 -1185 8385 -1165
rect 8365 -1235 8385 -1215
rect 8365 -1285 8385 -1265
rect 8365 -1335 8385 -1315
rect 8365 -1385 8385 -1365
rect 8365 -1435 8385 -1415
rect 8365 -1485 8385 -1465
rect 8365 -1535 8385 -1515
rect 8365 -1585 8385 -1565
rect 8365 -1635 8385 -1615
rect 9565 -985 9585 -965
rect 9565 -1035 9585 -1015
rect 9565 -1085 9585 -1065
rect 9565 -1135 9585 -1115
rect 9565 -1185 9585 -1165
rect 9565 -1235 9585 -1215
rect 9565 -1285 9585 -1265
rect 9565 -1335 9585 -1315
rect 9565 -1385 9585 -1365
rect 9565 -1435 9585 -1415
rect 9565 -1485 9585 -1465
rect 9565 -1535 9585 -1515
rect 9565 -1585 9585 -1565
rect 9565 -1635 9585 -1615
rect 10765 -985 10785 -965
rect 10765 -1035 10785 -1015
rect 10765 -1085 10785 -1065
rect 10765 -1135 10785 -1115
rect 10765 -1185 10785 -1165
rect 10765 -1235 10785 -1215
rect 10765 -1285 10785 -1265
rect 10765 -1335 10785 -1315
rect 10765 -1385 10785 -1365
rect 10765 -1435 10785 -1415
rect 10765 -1485 10785 -1465
rect 10765 -1535 10785 -1515
rect 10765 -1585 10785 -1565
rect 10765 -1635 10785 -1615
rect 11965 -985 11985 -965
rect 11965 -1035 11985 -1015
rect 11965 -1085 11985 -1065
rect 11965 -1135 11985 -1115
rect 11965 -1185 11985 -1165
rect 11965 -1235 11985 -1215
rect 11965 -1285 11985 -1265
rect 11965 -1335 11985 -1315
rect 11965 -1385 11985 -1365
rect 11965 -1435 11985 -1415
rect 11965 -1485 11985 -1465
rect 11965 -1535 11985 -1515
rect 11965 -1585 11985 -1565
rect 11965 -1635 11985 -1615
rect 12265 -985 12285 -965
rect 12265 -1035 12285 -1015
rect 12265 -1085 12285 -1065
rect 12265 -1135 12285 -1115
rect 12265 -1185 12285 -1165
rect 12265 -1235 12285 -1215
rect 12265 -1285 12285 -1265
rect 12265 -1335 12285 -1315
rect 12265 -1385 12285 -1365
rect 12265 -1435 12285 -1415
rect 12265 -1485 12285 -1465
rect 12265 -1535 12285 -1515
rect 12265 -1585 12285 -1565
rect 12265 -1635 12285 -1615
rect 12565 -985 12585 -965
rect 12565 -1035 12585 -1015
rect 12565 -1085 12585 -1065
rect 12565 -1135 12585 -1115
rect 12565 -1185 12585 -1165
rect 12565 -1235 12585 -1215
rect 12565 -1285 12585 -1265
rect 12565 -1335 12585 -1315
rect 12565 -1385 12585 -1365
rect 12565 -1435 12585 -1415
rect 12565 -1485 12585 -1465
rect 12565 -1535 12585 -1515
rect 12565 -1585 12585 -1565
rect 12565 -1635 12585 -1615
rect 12865 -985 12885 -965
rect 12865 -1035 12885 -1015
rect 12865 -1085 12885 -1065
rect 12865 -1135 12885 -1115
rect 12865 -1185 12885 -1165
rect 12865 -1235 12885 -1215
rect 12865 -1285 12885 -1265
rect 12865 -1335 12885 -1315
rect 12865 -1385 12885 -1365
rect 12865 -1435 12885 -1415
rect 12865 -1485 12885 -1465
rect 12865 -1535 12885 -1515
rect 12865 -1585 12885 -1565
rect 12865 -1635 12885 -1615
rect 13165 -985 13185 -965
rect 13165 -1035 13185 -1015
rect 13165 -1085 13185 -1065
rect 13165 -1135 13185 -1115
rect 13165 -1185 13185 -1165
rect 13165 -1235 13185 -1215
rect 13165 -1285 13185 -1265
rect 13165 -1335 13185 -1315
rect 13165 -1385 13185 -1365
rect 13165 -1435 13185 -1415
rect 13165 -1485 13185 -1465
rect 13165 -1535 13185 -1515
rect 13165 -1585 13185 -1565
rect 13165 -1635 13185 -1615
rect 13465 -985 13485 -965
rect 13465 -1035 13485 -1015
rect 13465 -1085 13485 -1065
rect 13465 -1135 13485 -1115
rect 13465 -1185 13485 -1165
rect 13465 -1235 13485 -1215
rect 13465 -1285 13485 -1265
rect 13465 -1335 13485 -1315
rect 13465 -1385 13485 -1365
rect 13465 -1435 13485 -1415
rect 13465 -1485 13485 -1465
rect 13465 -1535 13485 -1515
rect 13465 -1585 13485 -1565
rect 13465 -1635 13485 -1615
rect 13765 -985 13785 -965
rect 13765 -1035 13785 -1015
rect 13765 -1085 13785 -1065
rect 13765 -1135 13785 -1115
rect 13765 -1185 13785 -1165
rect 13765 -1235 13785 -1215
rect 13765 -1285 13785 -1265
rect 13765 -1335 13785 -1315
rect 13765 -1385 13785 -1365
rect 13765 -1435 13785 -1415
rect 13765 -1485 13785 -1465
rect 13765 -1535 13785 -1515
rect 13765 -1585 13785 -1565
rect 13765 -1635 13785 -1615
rect 14065 -985 14085 -965
rect 14065 -1035 14085 -1015
rect 14065 -1085 14085 -1065
rect 14065 -1135 14085 -1115
rect 14065 -1185 14085 -1165
rect 14065 -1235 14085 -1215
rect 14065 -1285 14085 -1265
rect 14065 -1335 14085 -1315
rect 14065 -1385 14085 -1365
rect 14065 -1435 14085 -1415
rect 14065 -1485 14085 -1465
rect 14065 -1535 14085 -1515
rect 14065 -1585 14085 -1565
rect 14065 -1635 14085 -1615
rect 14365 -985 14385 -965
rect 14365 -1035 14385 -1015
rect 14365 -1085 14385 -1065
rect 14365 -1135 14385 -1115
rect 14365 -1185 14385 -1165
rect 14365 -1235 14385 -1215
rect 14365 -1285 14385 -1265
rect 14365 -1335 14385 -1315
rect 14365 -1385 14385 -1365
rect 14365 -1435 14385 -1415
rect 14365 -1485 14385 -1465
rect 14365 -1535 14385 -1515
rect 14365 -1585 14385 -1565
rect 14365 -1635 14385 -1615
rect 15565 -985 15585 -965
rect 15565 -1035 15585 -1015
rect 15565 -1085 15585 -1065
rect 15565 -1135 15585 -1115
rect 15565 -1185 15585 -1165
rect 15565 -1235 15585 -1215
rect 15565 -1285 15585 -1265
rect 15565 -1335 15585 -1315
rect 15565 -1385 15585 -1365
rect 15565 -1435 15585 -1415
rect 15565 -1485 15585 -1465
rect 15565 -1535 15585 -1515
rect 15565 -1585 15585 -1565
rect 15565 -1635 15585 -1615
rect 16765 -985 16785 -965
rect 16765 -1035 16785 -1015
rect 16765 -1085 16785 -1065
rect 16765 -1135 16785 -1115
rect 16765 -1185 16785 -1165
rect 16765 -1235 16785 -1215
rect 16765 -1285 16785 -1265
rect 16765 -1335 16785 -1315
rect 16765 -1385 16785 -1365
rect 16765 -1435 16785 -1415
rect 16765 -1485 16785 -1465
rect 16765 -1535 16785 -1515
rect 16765 -1585 16785 -1565
rect 16765 -1635 16785 -1615
rect 17965 -985 17985 -965
rect 17965 -1035 17985 -1015
rect 17965 -1085 17985 -1065
rect 17965 -1135 17985 -1115
rect 17965 -1185 17985 -1165
rect 17965 -1235 17985 -1215
rect 17965 -1285 17985 -1265
rect 17965 -1335 17985 -1315
rect 17965 -1385 17985 -1365
rect 17965 -1435 17985 -1415
rect 17965 -1485 17985 -1465
rect 17965 -1535 17985 -1515
rect 17965 -1585 17985 -1565
rect 17965 -1635 17985 -1615
rect 19165 -985 19185 -965
rect 19165 -1035 19185 -1015
rect 19165 -1085 19185 -1065
rect 19165 -1135 19185 -1115
rect 19165 -1185 19185 -1165
rect 19165 -1235 19185 -1215
rect 19165 -1285 19185 -1265
rect 19165 -1335 19185 -1315
rect 19165 -1385 19185 -1365
rect 19165 -1435 19185 -1415
rect 19165 -1485 19185 -1465
rect 19165 -1535 19185 -1515
rect 19165 -1585 19185 -1565
rect 19165 -1635 19185 -1615
rect 20365 -985 20385 -965
rect 20365 -1035 20385 -1015
rect 20365 -1085 20385 -1065
rect 20365 -1135 20385 -1115
rect 20365 -1185 20385 -1165
rect 20365 -1235 20385 -1215
rect 20365 -1285 20385 -1265
rect 20365 -1335 20385 -1315
rect 20365 -1385 20385 -1365
rect 20365 -1435 20385 -1415
rect 20365 -1485 20385 -1465
rect 20365 -1535 20385 -1515
rect 20365 -1585 20385 -1565
rect 20365 -1635 20385 -1615
rect 21565 -985 21585 -965
rect 21565 -1035 21585 -1015
rect 21565 -1085 21585 -1065
rect 21565 -1135 21585 -1115
rect 21565 -1185 21585 -1165
rect 21565 -1235 21585 -1215
rect 21565 -1285 21585 -1265
rect 21565 -1335 21585 -1315
rect 21565 -1385 21585 -1365
rect 21565 -1435 21585 -1415
rect 21565 -1485 21585 -1465
rect 21565 -1535 21585 -1515
rect 21565 -1585 21585 -1565
rect 21565 -1635 21585 -1615
rect 22465 -985 22485 -965
rect 22465 -1035 22485 -1015
rect 22465 -1085 22485 -1065
rect 22465 -1135 22485 -1115
rect 22465 -1185 22485 -1165
rect 22465 -1235 22485 -1215
rect 22465 -1285 22485 -1265
rect 22465 -1335 22485 -1315
rect 22465 -1385 22485 -1365
rect 22465 -1435 22485 -1415
rect 22465 -1485 22485 -1465
rect 22465 -1535 22485 -1515
rect 22465 -1585 22485 -1565
rect 22465 -1635 22485 -1615
rect 23365 -985 23385 -965
rect 23365 -1035 23385 -1015
rect 23365 -1085 23385 -1065
rect 23365 -1135 23385 -1115
rect 23365 -1185 23385 -1165
rect 23365 -1235 23385 -1215
rect 23365 -1285 23385 -1265
rect 23365 -1335 23385 -1315
rect 23365 -1385 23385 -1365
rect 23365 -1435 23385 -1415
rect 23365 -1485 23385 -1465
rect 23365 -1535 23385 -1515
rect 23365 -1585 23385 -1565
rect 23365 -1635 23385 -1615
rect 24565 -985 24585 -965
rect 24565 -1035 24585 -1015
rect 24565 -1085 24585 -1065
rect 24565 -1135 24585 -1115
rect 24565 -1185 24585 -1165
rect 24565 -1235 24585 -1215
rect 24565 -1285 24585 -1265
rect 24565 -1335 24585 -1315
rect 24565 -1385 24585 -1365
rect 24565 -1435 24585 -1415
rect 24565 -1485 24585 -1465
rect 24565 -1535 24585 -1515
rect 24565 -1585 24585 -1565
rect 24565 -1635 24585 -1615
rect 25765 -985 25785 -965
rect 25765 -1035 25785 -1015
rect 25765 -1085 25785 -1065
rect 25765 -1135 25785 -1115
rect 25765 -1185 25785 -1165
rect 25765 -1235 25785 -1215
rect 25765 -1285 25785 -1265
rect 25765 -1335 25785 -1315
rect 25765 -1385 25785 -1365
rect 25765 -1435 25785 -1415
rect 25765 -1485 25785 -1465
rect 25765 -1535 25785 -1515
rect 25765 -1585 25785 -1565
rect 25765 -1635 25785 -1615
rect 26665 -985 26685 -965
rect 26665 -1035 26685 -1015
rect 26665 -1085 26685 -1065
rect 26665 -1135 26685 -1115
rect 26665 -1185 26685 -1165
rect 26665 -1235 26685 -1215
rect 26665 -1285 26685 -1265
rect 26665 -1335 26685 -1315
rect 26665 -1385 26685 -1365
rect 26665 -1435 26685 -1415
rect 26665 -1485 26685 -1465
rect 26665 -1535 26685 -1515
rect 26665 -1585 26685 -1565
rect 26665 -1635 26685 -1615
rect 27565 -985 27585 -965
rect 27565 -1035 27585 -1015
rect 27565 -1085 27585 -1065
rect 27565 -1135 27585 -1115
rect 27565 -1185 27585 -1165
rect 27565 -1235 27585 -1215
rect 27565 -1285 27585 -1265
rect 27565 -1335 27585 -1315
rect 27565 -1385 27585 -1365
rect 27565 -1435 27585 -1415
rect 27565 -1485 27585 -1465
rect 27565 -1535 27585 -1515
rect 27565 -1585 27585 -1565
rect 27565 -1635 27585 -1615
rect 28765 -985 28785 -965
rect 28765 -1035 28785 -1015
rect 28765 -1085 28785 -1065
rect 28765 -1135 28785 -1115
rect 28765 -1185 28785 -1165
rect 28765 -1235 28785 -1215
rect 28765 -1285 28785 -1265
rect 28765 -1335 28785 -1315
rect 28765 -1385 28785 -1365
rect 28765 -1435 28785 -1415
rect 28765 -1485 28785 -1465
rect 28765 -1535 28785 -1515
rect 28765 -1585 28785 -1565
rect 28765 -1635 28785 -1615
<< mvpdiffc >>
rect -635 5465 -615 5485
rect -635 5415 -615 5435
rect -635 5365 -615 5385
rect -635 5315 -615 5335
rect -635 5265 -615 5285
rect -635 5215 -615 5235
rect -635 5165 -615 5185
rect -635 5115 -615 5135
rect -635 5065 -615 5085
rect -635 5015 -615 5035
rect -485 5465 -465 5485
rect -485 5415 -465 5435
rect -485 5365 -465 5385
rect -485 5315 -465 5335
rect -485 5265 -465 5285
rect -485 5215 -465 5235
rect -485 5165 -465 5185
rect -485 5115 -465 5135
rect -485 5065 -465 5085
rect -485 5015 -465 5035
rect -335 5465 -315 5485
rect -335 5415 -315 5435
rect -335 5365 -315 5385
rect -335 5315 -315 5335
rect -335 5265 -315 5285
rect -335 5215 -315 5235
rect -335 5165 -315 5185
rect -335 5115 -315 5135
rect -335 5065 -315 5085
rect -335 5015 -315 5035
rect -185 5465 -165 5485
rect -185 5415 -165 5435
rect -185 5365 -165 5385
rect -185 5315 -165 5335
rect -185 5265 -165 5285
rect -185 5215 -165 5235
rect -185 5165 -165 5185
rect -185 5115 -165 5135
rect -185 5065 -165 5085
rect -185 5015 -165 5035
rect -35 5465 -15 5485
rect -35 5415 -15 5435
rect -35 5365 -15 5385
rect -35 5315 -15 5335
rect -35 5265 -15 5285
rect -35 5215 -15 5235
rect -35 5165 -15 5185
rect -35 5115 -15 5135
rect -35 5065 -15 5085
rect -35 5015 -15 5035
rect 565 5465 585 5485
rect 565 5415 585 5435
rect 565 5365 585 5385
rect 565 5315 585 5335
rect 565 5265 585 5285
rect 565 5215 585 5235
rect 565 5165 585 5185
rect 565 5115 585 5135
rect 565 5065 585 5085
rect 565 5015 585 5035
rect 715 5465 735 5485
rect 715 5415 735 5435
rect 715 5365 735 5385
rect 715 5315 735 5335
rect 715 5265 735 5285
rect 715 5215 735 5235
rect 715 5165 735 5185
rect 715 5115 735 5135
rect 715 5065 735 5085
rect 715 5015 735 5035
rect 865 5465 885 5485
rect 865 5415 885 5435
rect 865 5365 885 5385
rect 865 5315 885 5335
rect 865 5265 885 5285
rect 865 5215 885 5235
rect 865 5165 885 5185
rect 865 5115 885 5135
rect 865 5065 885 5085
rect 865 5015 885 5035
rect 1015 5465 1035 5485
rect 1015 5415 1035 5435
rect 1015 5365 1035 5385
rect 1015 5315 1035 5335
rect 1015 5265 1035 5285
rect 1015 5215 1035 5235
rect 1015 5165 1035 5185
rect 1015 5115 1035 5135
rect 1015 5065 1035 5085
rect 1015 5015 1035 5035
rect 1165 5465 1185 5485
rect 1165 5415 1185 5435
rect 1165 5365 1185 5385
rect 1165 5315 1185 5335
rect 1165 5265 1185 5285
rect 1165 5215 1185 5235
rect 1165 5165 1185 5185
rect 1165 5115 1185 5135
rect 1165 5065 1185 5085
rect 1165 5015 1185 5035
rect 1315 5465 1335 5485
rect 1315 5415 1335 5435
rect 1315 5365 1335 5385
rect 1315 5315 1335 5335
rect 1315 5265 1335 5285
rect 1315 5215 1335 5235
rect 1315 5165 1335 5185
rect 1315 5115 1335 5135
rect 1315 5065 1335 5085
rect 1315 5015 1335 5035
rect 1465 5465 1485 5485
rect 1465 5415 1485 5435
rect 1465 5365 1485 5385
rect 1465 5315 1485 5335
rect 1465 5265 1485 5285
rect 1465 5215 1485 5235
rect 1465 5165 1485 5185
rect 1465 5115 1485 5135
rect 1465 5065 1485 5085
rect 1465 5015 1485 5035
rect 1615 5465 1635 5485
rect 1615 5415 1635 5435
rect 1615 5365 1635 5385
rect 1615 5315 1635 5335
rect 1615 5265 1635 5285
rect 1615 5215 1635 5235
rect 1615 5165 1635 5185
rect 1615 5115 1635 5135
rect 1615 5065 1635 5085
rect 1615 5015 1635 5035
rect 1765 5465 1785 5485
rect 1765 5415 1785 5435
rect 1765 5365 1785 5385
rect 1765 5315 1785 5335
rect 1765 5265 1785 5285
rect 1765 5215 1785 5235
rect 1765 5165 1785 5185
rect 1765 5115 1785 5135
rect 1765 5065 1785 5085
rect 1765 5015 1785 5035
rect 1915 5465 1935 5485
rect 1915 5415 1935 5435
rect 1915 5365 1935 5385
rect 1915 5315 1935 5335
rect 1915 5265 1935 5285
rect 1915 5215 1935 5235
rect 1915 5165 1935 5185
rect 1915 5115 1935 5135
rect 1915 5065 1935 5085
rect 1915 5015 1935 5035
rect 2065 5465 2085 5485
rect 2065 5415 2085 5435
rect 2065 5365 2085 5385
rect 2065 5315 2085 5335
rect 2065 5265 2085 5285
rect 2065 5215 2085 5235
rect 2065 5165 2085 5185
rect 2065 5115 2085 5135
rect 2065 5065 2085 5085
rect 2065 5015 2085 5035
rect 2215 5465 2235 5485
rect 2215 5415 2235 5435
rect 2215 5365 2235 5385
rect 2215 5315 2235 5335
rect 2215 5265 2235 5285
rect 2215 5215 2235 5235
rect 2215 5165 2235 5185
rect 2215 5115 2235 5135
rect 2215 5065 2235 5085
rect 2215 5015 2235 5035
rect 2365 5465 2385 5485
rect 2365 5415 2385 5435
rect 2365 5365 2385 5385
rect 2365 5315 2385 5335
rect 2365 5265 2385 5285
rect 2365 5215 2385 5235
rect 2365 5165 2385 5185
rect 2365 5115 2385 5135
rect 2365 5065 2385 5085
rect 2365 5015 2385 5035
rect 2515 5465 2535 5485
rect 2515 5415 2535 5435
rect 2515 5365 2535 5385
rect 2515 5315 2535 5335
rect 2515 5265 2535 5285
rect 2515 5215 2535 5235
rect 2515 5165 2535 5185
rect 2515 5115 2535 5135
rect 2515 5065 2535 5085
rect 2515 5015 2535 5035
rect 2665 5465 2685 5485
rect 2665 5415 2685 5435
rect 2665 5365 2685 5385
rect 2665 5315 2685 5335
rect 2665 5265 2685 5285
rect 2665 5215 2685 5235
rect 2665 5165 2685 5185
rect 2665 5115 2685 5135
rect 2665 5065 2685 5085
rect 2665 5015 2685 5035
rect 2815 5465 2835 5485
rect 2815 5415 2835 5435
rect 2815 5365 2835 5385
rect 2815 5315 2835 5335
rect 2815 5265 2835 5285
rect 2815 5215 2835 5235
rect 2815 5165 2835 5185
rect 2815 5115 2835 5135
rect 2815 5065 2835 5085
rect 2815 5015 2835 5035
rect 2965 5465 2985 5485
rect 2965 5415 2985 5435
rect 2965 5365 2985 5385
rect 2965 5315 2985 5335
rect 2965 5265 2985 5285
rect 2965 5215 2985 5235
rect 2965 5165 2985 5185
rect 2965 5115 2985 5135
rect 2965 5065 2985 5085
rect 2965 5015 2985 5035
rect 3115 5465 3135 5485
rect 3115 5415 3135 5435
rect 3115 5365 3135 5385
rect 3115 5315 3135 5335
rect 3115 5265 3135 5285
rect 3115 5215 3135 5235
rect 3115 5165 3135 5185
rect 3115 5115 3135 5135
rect 3115 5065 3135 5085
rect 3115 5015 3135 5035
rect 3265 5465 3285 5485
rect 3265 5415 3285 5435
rect 3265 5365 3285 5385
rect 3265 5315 3285 5335
rect 3265 5265 3285 5285
rect 3265 5215 3285 5235
rect 3265 5165 3285 5185
rect 3265 5115 3285 5135
rect 3265 5065 3285 5085
rect 3265 5015 3285 5035
rect 3415 5465 3435 5485
rect 3415 5415 3435 5435
rect 3415 5365 3435 5385
rect 3415 5315 3435 5335
rect 3415 5265 3435 5285
rect 3415 5215 3435 5235
rect 3415 5165 3435 5185
rect 3415 5115 3435 5135
rect 3415 5065 3435 5085
rect 3415 5015 3435 5035
rect 3565 5465 3585 5485
rect 3565 5415 3585 5435
rect 3565 5365 3585 5385
rect 3565 5315 3585 5335
rect 3565 5265 3585 5285
rect 3565 5215 3585 5235
rect 3565 5165 3585 5185
rect 3565 5115 3585 5135
rect 3565 5065 3585 5085
rect 3565 5015 3585 5035
rect 4165 5465 4185 5485
rect 4165 5415 4185 5435
rect 4165 5365 4185 5385
rect 4165 5315 4185 5335
rect 4165 5265 4185 5285
rect 4165 5215 4185 5235
rect 4165 5165 4185 5185
rect 4165 5115 4185 5135
rect 4165 5065 4185 5085
rect 4165 5015 4185 5035
rect 4765 5465 4785 5485
rect 4765 5415 4785 5435
rect 4765 5365 4785 5385
rect 4765 5315 4785 5335
rect 4765 5265 4785 5285
rect 4765 5215 4785 5235
rect 4765 5165 4785 5185
rect 4765 5115 4785 5135
rect 4765 5065 4785 5085
rect 4765 5015 4785 5035
rect 4915 5465 4935 5485
rect 4915 5415 4935 5435
rect 4915 5365 4935 5385
rect 4915 5315 4935 5335
rect 4915 5265 4935 5285
rect 4915 5215 4935 5235
rect 4915 5165 4935 5185
rect 4915 5115 4935 5135
rect 4915 5065 4935 5085
rect 4915 5015 4935 5035
rect 5065 5465 5085 5485
rect 5065 5415 5085 5435
rect 5065 5365 5085 5385
rect 5065 5315 5085 5335
rect 5065 5265 5085 5285
rect 5065 5215 5085 5235
rect 5065 5165 5085 5185
rect 5065 5115 5085 5135
rect 5065 5065 5085 5085
rect 5065 5015 5085 5035
rect 5215 5465 5235 5485
rect 5215 5415 5235 5435
rect 5215 5365 5235 5385
rect 5215 5315 5235 5335
rect 5215 5265 5235 5285
rect 5215 5215 5235 5235
rect 5215 5165 5235 5185
rect 5215 5115 5235 5135
rect 5215 5065 5235 5085
rect 5215 5015 5235 5035
rect 5365 5465 5385 5485
rect 5365 5415 5385 5435
rect 5365 5365 5385 5385
rect 5365 5315 5385 5335
rect 5365 5265 5385 5285
rect 5365 5215 5385 5235
rect 5365 5165 5385 5185
rect 5365 5115 5385 5135
rect 5365 5065 5385 5085
rect 5365 5015 5385 5035
rect 5515 5465 5535 5485
rect 5515 5415 5535 5435
rect 5515 5365 5535 5385
rect 5515 5315 5535 5335
rect 5515 5265 5535 5285
rect 5515 5215 5535 5235
rect 5515 5165 5535 5185
rect 5515 5115 5535 5135
rect 5515 5065 5535 5085
rect 5515 5015 5535 5035
rect 5665 5465 5685 5485
rect 5665 5415 5685 5435
rect 5665 5365 5685 5385
rect 5665 5315 5685 5335
rect 5665 5265 5685 5285
rect 5665 5215 5685 5235
rect 5665 5165 5685 5185
rect 5665 5115 5685 5135
rect 5665 5065 5685 5085
rect 5665 5015 5685 5035
rect 5815 5465 5835 5485
rect 5815 5415 5835 5435
rect 5815 5365 5835 5385
rect 5815 5315 5835 5335
rect 5815 5265 5835 5285
rect 5815 5215 5835 5235
rect 5815 5165 5835 5185
rect 5815 5115 5835 5135
rect 5815 5065 5835 5085
rect 5815 5015 5835 5035
rect 5965 5465 5985 5485
rect 5965 5415 5985 5435
rect 5965 5365 5985 5385
rect 5965 5315 5985 5335
rect 5965 5265 5985 5285
rect 5965 5215 5985 5235
rect 5965 5165 5985 5185
rect 5965 5115 5985 5135
rect 5965 5065 5985 5085
rect 5965 5015 5985 5035
rect 6115 5465 6135 5485
rect 6115 5415 6135 5435
rect 6115 5365 6135 5385
rect 6115 5315 6135 5335
rect 6115 5265 6135 5285
rect 6115 5215 6135 5235
rect 6115 5165 6135 5185
rect 6115 5115 6135 5135
rect 6115 5065 6135 5085
rect 6115 5015 6135 5035
rect 6265 5465 6285 5485
rect 6265 5415 6285 5435
rect 6265 5365 6285 5385
rect 6265 5315 6285 5335
rect 6265 5265 6285 5285
rect 6265 5215 6285 5235
rect 6265 5165 6285 5185
rect 6265 5115 6285 5135
rect 6265 5065 6285 5085
rect 6265 5015 6285 5035
rect 6415 5465 6435 5485
rect 6415 5415 6435 5435
rect 6415 5365 6435 5385
rect 6415 5315 6435 5335
rect 6415 5265 6435 5285
rect 6415 5215 6435 5235
rect 6415 5165 6435 5185
rect 6415 5115 6435 5135
rect 6415 5065 6435 5085
rect 6415 5015 6435 5035
rect 6565 5465 6585 5485
rect 6565 5415 6585 5435
rect 6565 5365 6585 5385
rect 6565 5315 6585 5335
rect 6565 5265 6585 5285
rect 6565 5215 6585 5235
rect 6565 5165 6585 5185
rect 6565 5115 6585 5135
rect 6565 5065 6585 5085
rect 6565 5015 6585 5035
rect 6715 5465 6735 5485
rect 6715 5415 6735 5435
rect 6715 5365 6735 5385
rect 6715 5315 6735 5335
rect 6715 5265 6735 5285
rect 6715 5215 6735 5235
rect 6715 5165 6735 5185
rect 6715 5115 6735 5135
rect 6715 5065 6735 5085
rect 6715 5015 6735 5035
rect 6865 5465 6885 5485
rect 6865 5415 6885 5435
rect 6865 5365 6885 5385
rect 6865 5315 6885 5335
rect 6865 5265 6885 5285
rect 6865 5215 6885 5235
rect 6865 5165 6885 5185
rect 6865 5115 6885 5135
rect 6865 5065 6885 5085
rect 6865 5015 6885 5035
rect 7015 5465 7035 5485
rect 7015 5415 7035 5435
rect 7015 5365 7035 5385
rect 7015 5315 7035 5335
rect 7015 5265 7035 5285
rect 7015 5215 7035 5235
rect 7015 5165 7035 5185
rect 7015 5115 7035 5135
rect 7015 5065 7035 5085
rect 7015 5015 7035 5035
rect 7165 5465 7185 5485
rect 7165 5415 7185 5435
rect 7165 5365 7185 5385
rect 7165 5315 7185 5335
rect 7165 5265 7185 5285
rect 7165 5215 7185 5235
rect 7165 5165 7185 5185
rect 7165 5115 7185 5135
rect 7165 5065 7185 5085
rect 7165 5015 7185 5035
rect 7315 5465 7335 5485
rect 7315 5415 7335 5435
rect 7315 5365 7335 5385
rect 7315 5315 7335 5335
rect 7315 5265 7335 5285
rect 7315 5215 7335 5235
rect 7315 5165 7335 5185
rect 7315 5115 7335 5135
rect 7315 5065 7335 5085
rect 7315 5015 7335 5035
rect 7465 5465 7485 5485
rect 7465 5415 7485 5435
rect 7465 5365 7485 5385
rect 7465 5315 7485 5335
rect 7465 5265 7485 5285
rect 7465 5215 7485 5235
rect 7465 5165 7485 5185
rect 7465 5115 7485 5135
rect 7465 5065 7485 5085
rect 7465 5015 7485 5035
rect 7615 5465 7635 5485
rect 7615 5415 7635 5435
rect 7615 5365 7635 5385
rect 7615 5315 7635 5335
rect 7615 5265 7635 5285
rect 7615 5215 7635 5235
rect 7615 5165 7635 5185
rect 7615 5115 7635 5135
rect 7615 5065 7635 5085
rect 7615 5015 7635 5035
rect 7765 5465 7785 5485
rect 7765 5415 7785 5435
rect 7765 5365 7785 5385
rect 7765 5315 7785 5335
rect 7765 5265 7785 5285
rect 7765 5215 7785 5235
rect 7765 5165 7785 5185
rect 7765 5115 7785 5135
rect 7765 5065 7785 5085
rect 7765 5015 7785 5035
rect 8365 5465 8385 5485
rect 8365 5415 8385 5435
rect 8365 5365 8385 5385
rect 8365 5315 8385 5335
rect 8365 5265 8385 5285
rect 8365 5215 8385 5235
rect 8365 5165 8385 5185
rect 8365 5115 8385 5135
rect 8365 5065 8385 5085
rect 8365 5015 8385 5035
rect 8515 5465 8535 5485
rect 8515 5415 8535 5435
rect 8515 5365 8535 5385
rect 8515 5315 8535 5335
rect 8515 5265 8535 5285
rect 8515 5215 8535 5235
rect 8515 5165 8535 5185
rect 8515 5115 8535 5135
rect 8515 5065 8535 5085
rect 8515 5015 8535 5035
rect 8665 5465 8685 5485
rect 8665 5415 8685 5435
rect 8665 5365 8685 5385
rect 8665 5315 8685 5335
rect 8665 5265 8685 5285
rect 8665 5215 8685 5235
rect 8665 5165 8685 5185
rect 8665 5115 8685 5135
rect 8665 5065 8685 5085
rect 8665 5015 8685 5035
rect 8815 5465 8835 5485
rect 8815 5415 8835 5435
rect 8815 5365 8835 5385
rect 8815 5315 8835 5335
rect 8815 5265 8835 5285
rect 8815 5215 8835 5235
rect 8815 5165 8835 5185
rect 8815 5115 8835 5135
rect 8815 5065 8835 5085
rect 8815 5015 8835 5035
rect 8965 5465 8985 5485
rect 8965 5415 8985 5435
rect 8965 5365 8985 5385
rect 8965 5315 8985 5335
rect 8965 5265 8985 5285
rect 8965 5215 8985 5235
rect 8965 5165 8985 5185
rect 8965 5115 8985 5135
rect 8965 5065 8985 5085
rect 8965 5015 8985 5035
rect 9115 5465 9135 5485
rect 9115 5415 9135 5435
rect 9115 5365 9135 5385
rect 9115 5315 9135 5335
rect 9115 5265 9135 5285
rect 9115 5215 9135 5235
rect 9115 5165 9135 5185
rect 9115 5115 9135 5135
rect 9115 5065 9135 5085
rect 9115 5015 9135 5035
rect 9265 5465 9285 5485
rect 9265 5415 9285 5435
rect 9265 5365 9285 5385
rect 9265 5315 9285 5335
rect 9265 5265 9285 5285
rect 9265 5215 9285 5235
rect 9265 5165 9285 5185
rect 9265 5115 9285 5135
rect 9265 5065 9285 5085
rect 9265 5015 9285 5035
rect 9415 5465 9435 5485
rect 9415 5415 9435 5435
rect 9415 5365 9435 5385
rect 9415 5315 9435 5335
rect 9415 5265 9435 5285
rect 9415 5215 9435 5235
rect 9415 5165 9435 5185
rect 9415 5115 9435 5135
rect 9415 5065 9435 5085
rect 9415 5015 9435 5035
rect 9565 5465 9585 5485
rect 9565 5415 9585 5435
rect 9565 5365 9585 5385
rect 9565 5315 9585 5335
rect 9565 5265 9585 5285
rect 9565 5215 9585 5235
rect 9565 5165 9585 5185
rect 9565 5115 9585 5135
rect 9565 5065 9585 5085
rect 9565 5015 9585 5035
rect 9715 5465 9735 5485
rect 9715 5415 9735 5435
rect 9715 5365 9735 5385
rect 9715 5315 9735 5335
rect 9715 5265 9735 5285
rect 9715 5215 9735 5235
rect 9715 5165 9735 5185
rect 9715 5115 9735 5135
rect 9715 5065 9735 5085
rect 9715 5015 9735 5035
rect 9865 5465 9885 5485
rect 9865 5415 9885 5435
rect 9865 5365 9885 5385
rect 9865 5315 9885 5335
rect 9865 5265 9885 5285
rect 9865 5215 9885 5235
rect 9865 5165 9885 5185
rect 9865 5115 9885 5135
rect 9865 5065 9885 5085
rect 9865 5015 9885 5035
rect 10015 5465 10035 5485
rect 10015 5415 10035 5435
rect 10015 5365 10035 5385
rect 10015 5315 10035 5335
rect 10015 5265 10035 5285
rect 10015 5215 10035 5235
rect 10015 5165 10035 5185
rect 10015 5115 10035 5135
rect 10015 5065 10035 5085
rect 10015 5015 10035 5035
rect 10165 5465 10185 5485
rect 10165 5415 10185 5435
rect 10165 5365 10185 5385
rect 10165 5315 10185 5335
rect 10165 5265 10185 5285
rect 10165 5215 10185 5235
rect 10165 5165 10185 5185
rect 10165 5115 10185 5135
rect 10165 5065 10185 5085
rect 10165 5015 10185 5035
rect 10315 5465 10335 5485
rect 10315 5415 10335 5435
rect 10315 5365 10335 5385
rect 10315 5315 10335 5335
rect 10315 5265 10335 5285
rect 10315 5215 10335 5235
rect 10315 5165 10335 5185
rect 10315 5115 10335 5135
rect 10315 5065 10335 5085
rect 10315 5015 10335 5035
rect 10465 5465 10485 5485
rect 10465 5415 10485 5435
rect 10465 5365 10485 5385
rect 10465 5315 10485 5335
rect 10465 5265 10485 5285
rect 10465 5215 10485 5235
rect 10465 5165 10485 5185
rect 10465 5115 10485 5135
rect 10465 5065 10485 5085
rect 10465 5015 10485 5035
rect 10615 5465 10635 5485
rect 10615 5415 10635 5435
rect 10615 5365 10635 5385
rect 10615 5315 10635 5335
rect 10615 5265 10635 5285
rect 10615 5215 10635 5235
rect 10615 5165 10635 5185
rect 10615 5115 10635 5135
rect 10615 5065 10635 5085
rect 10615 5015 10635 5035
rect 10765 5465 10785 5485
rect 10765 5415 10785 5435
rect 10765 5365 10785 5385
rect 10765 5315 10785 5335
rect 10765 5265 10785 5285
rect 10765 5215 10785 5235
rect 10765 5165 10785 5185
rect 10765 5115 10785 5135
rect 10765 5065 10785 5085
rect 10765 5015 10785 5035
rect 11365 5465 11385 5485
rect 11365 5415 11385 5435
rect 11365 5365 11385 5385
rect 11365 5315 11385 5335
rect 11365 5265 11385 5285
rect 11365 5215 11385 5235
rect 11365 5165 11385 5185
rect 11365 5115 11385 5135
rect 11365 5065 11385 5085
rect 11365 5015 11385 5035
rect 11965 5465 11985 5485
rect 11965 5415 11985 5435
rect 11965 5365 11985 5385
rect 11965 5315 11985 5335
rect 11965 5265 11985 5285
rect 11965 5215 11985 5235
rect 11965 5165 11985 5185
rect 11965 5115 11985 5135
rect 11965 5065 11985 5085
rect 11965 5015 11985 5035
rect 12565 5465 12585 5485
rect 12565 5415 12585 5435
rect 12565 5365 12585 5385
rect 12565 5315 12585 5335
rect 12565 5265 12585 5285
rect 12565 5215 12585 5235
rect 12565 5165 12585 5185
rect 12565 5115 12585 5135
rect 12565 5065 12585 5085
rect 12565 5015 12585 5035
rect 13165 5465 13185 5485
rect 13165 5415 13185 5435
rect 13165 5365 13185 5385
rect 13165 5315 13185 5335
rect 13165 5265 13185 5285
rect 13165 5215 13185 5235
rect 13165 5165 13185 5185
rect 13165 5115 13185 5135
rect 13165 5065 13185 5085
rect 13165 5015 13185 5035
rect 13765 5465 13785 5485
rect 13765 5415 13785 5435
rect 13765 5365 13785 5385
rect 13765 5315 13785 5335
rect 13765 5265 13785 5285
rect 13765 5215 13785 5235
rect 13765 5165 13785 5185
rect 13765 5115 13785 5135
rect 13765 5065 13785 5085
rect 13765 5015 13785 5035
rect 14365 5465 14385 5485
rect 14365 5415 14385 5435
rect 14365 5365 14385 5385
rect 14365 5315 14385 5335
rect 14365 5265 14385 5285
rect 14365 5215 14385 5235
rect 14365 5165 14385 5185
rect 14365 5115 14385 5135
rect 14365 5065 14385 5085
rect 14365 5015 14385 5035
rect 14965 5465 14985 5485
rect 14965 5415 14985 5435
rect 14965 5365 14985 5385
rect 14965 5315 14985 5335
rect 14965 5265 14985 5285
rect 14965 5215 14985 5235
rect 14965 5165 14985 5185
rect 14965 5115 14985 5135
rect 14965 5065 14985 5085
rect 14965 5015 14985 5035
rect 15565 5465 15585 5485
rect 15565 5415 15585 5435
rect 15565 5365 15585 5385
rect 15565 5315 15585 5335
rect 15565 5265 15585 5285
rect 15565 5215 15585 5235
rect 15565 5165 15585 5185
rect 15565 5115 15585 5135
rect 15565 5065 15585 5085
rect 15565 5015 15585 5035
rect 16165 5465 16185 5485
rect 16165 5415 16185 5435
rect 16165 5365 16185 5385
rect 16165 5315 16185 5335
rect 16165 5265 16185 5285
rect 16165 5215 16185 5235
rect 16165 5165 16185 5185
rect 16165 5115 16185 5135
rect 16165 5065 16185 5085
rect 16165 5015 16185 5035
rect 16315 5465 16335 5485
rect 16315 5415 16335 5435
rect 16315 5365 16335 5385
rect 16315 5315 16335 5335
rect 16315 5265 16335 5285
rect 16315 5215 16335 5235
rect 16315 5165 16335 5185
rect 16315 5115 16335 5135
rect 16315 5065 16335 5085
rect 16315 5015 16335 5035
rect 16465 5465 16485 5485
rect 16465 5415 16485 5435
rect 16465 5365 16485 5385
rect 16465 5315 16485 5335
rect 16465 5265 16485 5285
rect 16465 5215 16485 5235
rect 16465 5165 16485 5185
rect 16465 5115 16485 5135
rect 16465 5065 16485 5085
rect 16465 5015 16485 5035
rect 16615 5465 16635 5485
rect 16615 5415 16635 5435
rect 16615 5365 16635 5385
rect 16615 5315 16635 5335
rect 16615 5265 16635 5285
rect 16615 5215 16635 5235
rect 16615 5165 16635 5185
rect 16615 5115 16635 5135
rect 16615 5065 16635 5085
rect 16615 5015 16635 5035
rect 16765 5465 16785 5485
rect 16765 5415 16785 5435
rect 16765 5365 16785 5385
rect 16765 5315 16785 5335
rect 16765 5265 16785 5285
rect 16765 5215 16785 5235
rect 16765 5165 16785 5185
rect 16765 5115 16785 5135
rect 16765 5065 16785 5085
rect 16765 5015 16785 5035
rect 16915 5465 16935 5485
rect 16915 5415 16935 5435
rect 16915 5365 16935 5385
rect 16915 5315 16935 5335
rect 16915 5265 16935 5285
rect 16915 5215 16935 5235
rect 16915 5165 16935 5185
rect 16915 5115 16935 5135
rect 16915 5065 16935 5085
rect 16915 5015 16935 5035
rect 17065 5465 17085 5485
rect 17065 5415 17085 5435
rect 17065 5365 17085 5385
rect 17065 5315 17085 5335
rect 17065 5265 17085 5285
rect 17065 5215 17085 5235
rect 17065 5165 17085 5185
rect 17065 5115 17085 5135
rect 17065 5065 17085 5085
rect 17065 5015 17085 5035
rect 17215 5465 17235 5485
rect 17215 5415 17235 5435
rect 17215 5365 17235 5385
rect 17215 5315 17235 5335
rect 17215 5265 17235 5285
rect 17215 5215 17235 5235
rect 17215 5165 17235 5185
rect 17215 5115 17235 5135
rect 17215 5065 17235 5085
rect 17215 5015 17235 5035
rect 17365 5465 17385 5485
rect 17365 5415 17385 5435
rect 17365 5365 17385 5385
rect 17365 5315 17385 5335
rect 17365 5265 17385 5285
rect 17365 5215 17385 5235
rect 17365 5165 17385 5185
rect 17365 5115 17385 5135
rect 17365 5065 17385 5085
rect 17365 5015 17385 5035
rect 17965 5465 17985 5485
rect 17965 5415 17985 5435
rect 17965 5365 17985 5385
rect 17965 5315 17985 5335
rect 17965 5265 17985 5285
rect 17965 5215 17985 5235
rect 17965 5165 17985 5185
rect 17965 5115 17985 5135
rect 17965 5065 17985 5085
rect 17965 5015 17985 5035
rect 18565 5465 18585 5485
rect 18565 5415 18585 5435
rect 18565 5365 18585 5385
rect 18565 5315 18585 5335
rect 18565 5265 18585 5285
rect 18565 5215 18585 5235
rect 18565 5165 18585 5185
rect 18565 5115 18585 5135
rect 18565 5065 18585 5085
rect 18565 5015 18585 5035
rect 18715 5465 18735 5485
rect 18715 5415 18735 5435
rect 18715 5365 18735 5385
rect 18715 5315 18735 5335
rect 18715 5265 18735 5285
rect 18715 5215 18735 5235
rect 18715 5165 18735 5185
rect 18715 5115 18735 5135
rect 18715 5065 18735 5085
rect 18715 5015 18735 5035
rect 18865 5465 18885 5485
rect 18865 5415 18885 5435
rect 18865 5365 18885 5385
rect 18865 5315 18885 5335
rect 18865 5265 18885 5285
rect 18865 5215 18885 5235
rect 18865 5165 18885 5185
rect 18865 5115 18885 5135
rect 18865 5065 18885 5085
rect 18865 5015 18885 5035
rect 19015 5465 19035 5485
rect 19015 5415 19035 5435
rect 19015 5365 19035 5385
rect 19015 5315 19035 5335
rect 19015 5265 19035 5285
rect 19015 5215 19035 5235
rect 19015 5165 19035 5185
rect 19015 5115 19035 5135
rect 19015 5065 19035 5085
rect 19015 5015 19035 5035
rect 19165 5465 19185 5485
rect 19165 5415 19185 5435
rect 19165 5365 19185 5385
rect 19165 5315 19185 5335
rect 19165 5265 19185 5285
rect 19165 5215 19185 5235
rect 19165 5165 19185 5185
rect 19165 5115 19185 5135
rect 19165 5065 19185 5085
rect 19165 5015 19185 5035
rect 19315 5465 19335 5485
rect 19315 5415 19335 5435
rect 19315 5365 19335 5385
rect 19315 5315 19335 5335
rect 19315 5265 19335 5285
rect 19315 5215 19335 5235
rect 19315 5165 19335 5185
rect 19315 5115 19335 5135
rect 19315 5065 19335 5085
rect 19315 5015 19335 5035
rect 19465 5465 19485 5485
rect 19465 5415 19485 5435
rect 19465 5365 19485 5385
rect 19465 5315 19485 5335
rect 19465 5265 19485 5285
rect 19465 5215 19485 5235
rect 19465 5165 19485 5185
rect 19465 5115 19485 5135
rect 19465 5065 19485 5085
rect 19465 5015 19485 5035
rect 19615 5465 19635 5485
rect 19615 5415 19635 5435
rect 19615 5365 19635 5385
rect 19615 5315 19635 5335
rect 19615 5265 19635 5285
rect 19615 5215 19635 5235
rect 19615 5165 19635 5185
rect 19615 5115 19635 5135
rect 19615 5065 19635 5085
rect 19615 5015 19635 5035
rect 19765 5465 19785 5485
rect 19765 5415 19785 5435
rect 19765 5365 19785 5385
rect 19765 5315 19785 5335
rect 19765 5265 19785 5285
rect 19765 5215 19785 5235
rect 19765 5165 19785 5185
rect 19765 5115 19785 5135
rect 19765 5065 19785 5085
rect 19765 5015 19785 5035
rect 20365 5465 20385 5485
rect 20365 5415 20385 5435
rect 20365 5365 20385 5385
rect 20365 5315 20385 5335
rect 20365 5265 20385 5285
rect 20365 5215 20385 5235
rect 20365 5165 20385 5185
rect 20365 5115 20385 5135
rect 20365 5065 20385 5085
rect 20365 5015 20385 5035
rect 20965 5465 20985 5485
rect 20965 5415 20985 5435
rect 20965 5365 20985 5385
rect 20965 5315 20985 5335
rect 20965 5265 20985 5285
rect 20965 5215 20985 5235
rect 20965 5165 20985 5185
rect 20965 5115 20985 5135
rect 20965 5065 20985 5085
rect 20965 5015 20985 5035
rect 21415 5465 21435 5485
rect 21415 5415 21435 5435
rect 21415 5365 21435 5385
rect 21415 5315 21435 5335
rect 21415 5265 21435 5285
rect 21415 5215 21435 5235
rect 21415 5165 21435 5185
rect 21415 5115 21435 5135
rect 21415 5065 21435 5085
rect 21415 5015 21435 5035
rect 21865 5465 21885 5485
rect 21865 5415 21885 5435
rect 21865 5365 21885 5385
rect 21865 5315 21885 5335
rect 21865 5265 21885 5285
rect 21865 5215 21885 5235
rect 21865 5165 21885 5185
rect 21865 5115 21885 5135
rect 21865 5065 21885 5085
rect 21865 5015 21885 5035
rect 22465 5465 22485 5485
rect 22465 5415 22485 5435
rect 22465 5365 22485 5385
rect 22465 5315 22485 5335
rect 22465 5265 22485 5285
rect 22465 5215 22485 5235
rect 22465 5165 22485 5185
rect 22465 5115 22485 5135
rect 22465 5065 22485 5085
rect 22465 5015 22485 5035
rect 23065 5465 23085 5485
rect 23065 5415 23085 5435
rect 23065 5365 23085 5385
rect 23065 5315 23085 5335
rect 23065 5265 23085 5285
rect 23065 5215 23085 5235
rect 23065 5165 23085 5185
rect 23065 5115 23085 5135
rect 23065 5065 23085 5085
rect 23065 5015 23085 5035
rect 23515 5465 23535 5485
rect 23515 5415 23535 5435
rect 23515 5365 23535 5385
rect 23515 5315 23535 5335
rect 23515 5265 23535 5285
rect 23515 5215 23535 5235
rect 23515 5165 23535 5185
rect 23515 5115 23535 5135
rect 23515 5065 23535 5085
rect 23515 5015 23535 5035
rect 23965 5465 23985 5485
rect 23965 5415 23985 5435
rect 23965 5365 23985 5385
rect 23965 5315 23985 5335
rect 23965 5265 23985 5285
rect 23965 5215 23985 5235
rect 23965 5165 23985 5185
rect 23965 5115 23985 5135
rect 23965 5065 23985 5085
rect 23965 5015 23985 5035
rect 24565 5465 24585 5485
rect 24565 5415 24585 5435
rect 24565 5365 24585 5385
rect 24565 5315 24585 5335
rect 24565 5265 24585 5285
rect 24565 5215 24585 5235
rect 24565 5165 24585 5185
rect 24565 5115 24585 5135
rect 24565 5065 24585 5085
rect 24565 5015 24585 5035
rect 25165 5465 25185 5485
rect 25165 5415 25185 5435
rect 25165 5365 25185 5385
rect 25165 5315 25185 5335
rect 25165 5265 25185 5285
rect 25165 5215 25185 5235
rect 25165 5165 25185 5185
rect 25165 5115 25185 5135
rect 25165 5065 25185 5085
rect 25165 5015 25185 5035
rect 25615 5465 25635 5485
rect 25615 5415 25635 5435
rect 25615 5365 25635 5385
rect 25615 5315 25635 5335
rect 25615 5265 25635 5285
rect 25615 5215 25635 5235
rect 25615 5165 25635 5185
rect 25615 5115 25635 5135
rect 25615 5065 25635 5085
rect 25615 5015 25635 5035
rect 26065 5465 26085 5485
rect 26065 5415 26085 5435
rect 26065 5365 26085 5385
rect 26065 5315 26085 5335
rect 26065 5265 26085 5285
rect 26065 5215 26085 5235
rect 26065 5165 26085 5185
rect 26065 5115 26085 5135
rect 26065 5065 26085 5085
rect 26065 5015 26085 5035
rect 26665 5465 26685 5485
rect 26665 5415 26685 5435
rect 26665 5365 26685 5385
rect 26665 5315 26685 5335
rect 26665 5265 26685 5285
rect 26665 5215 26685 5235
rect 26665 5165 26685 5185
rect 26665 5115 26685 5135
rect 26665 5065 26685 5085
rect 26665 5015 26685 5035
rect 27265 5465 27285 5485
rect 27265 5415 27285 5435
rect 27265 5365 27285 5385
rect 27265 5315 27285 5335
rect 27265 5265 27285 5285
rect 27265 5215 27285 5235
rect 27265 5165 27285 5185
rect 27265 5115 27285 5135
rect 27265 5065 27285 5085
rect 27265 5015 27285 5035
rect 27715 5465 27735 5485
rect 27715 5415 27735 5435
rect 27715 5365 27735 5385
rect 27715 5315 27735 5335
rect 27715 5265 27735 5285
rect 27715 5215 27735 5235
rect 27715 5165 27735 5185
rect 27715 5115 27735 5135
rect 27715 5065 27735 5085
rect 27715 5015 27735 5035
rect 28165 5465 28185 5485
rect 28165 5415 28185 5435
rect 28165 5365 28185 5385
rect 28165 5315 28185 5335
rect 28165 5265 28185 5285
rect 28165 5215 28185 5235
rect 28165 5165 28185 5185
rect 28165 5115 28185 5135
rect 28165 5065 28185 5085
rect 28165 5015 28185 5035
rect 28765 5465 28785 5485
rect 28765 5415 28785 5435
rect 28765 5365 28785 5385
rect 28765 5315 28785 5335
rect 28765 5265 28785 5285
rect 28765 5215 28785 5235
rect 28765 5165 28785 5185
rect 28765 5115 28785 5135
rect 28765 5065 28785 5085
rect 28765 5015 28785 5035
rect 29365 5465 29385 5485
rect 29365 5415 29385 5435
rect 29365 5365 29385 5385
rect 29365 5315 29385 5335
rect 29365 5265 29385 5285
rect 29365 5215 29385 5235
rect 29365 5165 29385 5185
rect 29365 5115 29385 5135
rect 29365 5065 29385 5085
rect 29365 5015 29385 5035
rect 29515 5465 29535 5485
rect 29515 5415 29535 5435
rect 29515 5365 29535 5385
rect 29515 5315 29535 5335
rect 29515 5265 29535 5285
rect 29515 5215 29535 5235
rect 29515 5165 29535 5185
rect 29515 5115 29535 5135
rect 29515 5065 29535 5085
rect 29515 5015 29535 5035
rect 29665 5465 29685 5485
rect 29665 5415 29685 5435
rect 29665 5365 29685 5385
rect 29665 5315 29685 5335
rect 29665 5265 29685 5285
rect 29665 5215 29685 5235
rect 29665 5165 29685 5185
rect 29665 5115 29685 5135
rect 29665 5065 29685 5085
rect 29665 5015 29685 5035
rect 29815 5465 29835 5485
rect 29815 5415 29835 5435
rect 29815 5365 29835 5385
rect 29815 5315 29835 5335
rect 29815 5265 29835 5285
rect 29815 5215 29835 5235
rect 29815 5165 29835 5185
rect 29815 5115 29835 5135
rect 29815 5065 29835 5085
rect 29815 5015 29835 5035
rect 29965 5465 29985 5485
rect 29965 5415 29985 5435
rect 29965 5365 29985 5385
rect 29965 5315 29985 5335
rect 29965 5265 29985 5285
rect 29965 5215 29985 5235
rect 29965 5165 29985 5185
rect 29965 5115 29985 5135
rect 29965 5065 29985 5085
rect 29965 5015 29985 5035
rect 30115 5465 30135 5485
rect 30115 5415 30135 5435
rect 30115 5365 30135 5385
rect 30115 5315 30135 5335
rect 30115 5265 30135 5285
rect 30115 5215 30135 5235
rect 30115 5165 30135 5185
rect 30115 5115 30135 5135
rect 30115 5065 30135 5085
rect 30115 5015 30135 5035
rect 30265 5465 30285 5485
rect 30265 5415 30285 5435
rect 30265 5365 30285 5385
rect 30265 5315 30285 5335
rect 30265 5265 30285 5285
rect 30265 5215 30285 5235
rect 30265 5165 30285 5185
rect 30265 5115 30285 5135
rect 30265 5065 30285 5085
rect 30265 5015 30285 5035
rect 30415 5465 30435 5485
rect 30415 5415 30435 5435
rect 30415 5365 30435 5385
rect 30415 5315 30435 5335
rect 30415 5265 30435 5285
rect 30415 5215 30435 5235
rect 30415 5165 30435 5185
rect 30415 5115 30435 5135
rect 30415 5065 30435 5085
rect 30415 5015 30435 5035
rect 30565 5465 30585 5485
rect 30565 5415 30585 5435
rect 30565 5365 30585 5385
rect 30565 5315 30585 5335
rect 30565 5265 30585 5285
rect 30565 5215 30585 5235
rect 30565 5165 30585 5185
rect 30565 5115 30585 5135
rect 30565 5065 30585 5085
rect 30565 5015 30585 5035
rect 30715 5465 30735 5485
rect 30715 5415 30735 5435
rect 30715 5365 30735 5385
rect 30715 5315 30735 5335
rect 30715 5265 30735 5285
rect 30715 5215 30735 5235
rect 30715 5165 30735 5185
rect 30715 5115 30735 5135
rect 30715 5065 30735 5085
rect 30715 5015 30735 5035
rect 30865 5465 30885 5485
rect 30865 5415 30885 5435
rect 30865 5365 30885 5385
rect 30865 5315 30885 5335
rect 30865 5265 30885 5285
rect 30865 5215 30885 5235
rect 30865 5165 30885 5185
rect 30865 5115 30885 5135
rect 30865 5065 30885 5085
rect 30865 5015 30885 5035
rect 31015 5465 31035 5485
rect 31015 5415 31035 5435
rect 31015 5365 31035 5385
rect 31015 5315 31035 5335
rect 31015 5265 31035 5285
rect 31015 5215 31035 5235
rect 31015 5165 31035 5185
rect 31015 5115 31035 5135
rect 31015 5065 31035 5085
rect 31015 5015 31035 5035
rect 31165 5465 31185 5485
rect 31165 5415 31185 5435
rect 31165 5365 31185 5385
rect 31165 5315 31185 5335
rect 31165 5265 31185 5285
rect 31165 5215 31185 5235
rect 31165 5165 31185 5185
rect 31165 5115 31185 5135
rect 31165 5065 31185 5085
rect 31165 5015 31185 5035
rect 31315 5465 31335 5485
rect 31315 5415 31335 5435
rect 31315 5365 31335 5385
rect 31315 5315 31335 5335
rect 31315 5265 31335 5285
rect 31315 5215 31335 5235
rect 31315 5165 31335 5185
rect 31315 5115 31335 5135
rect 31315 5065 31335 5085
rect 31315 5015 31335 5035
rect 31465 5465 31485 5485
rect 31465 5415 31485 5435
rect 31465 5365 31485 5385
rect 31465 5315 31485 5335
rect 31465 5265 31485 5285
rect 31465 5215 31485 5235
rect 31465 5165 31485 5185
rect 31465 5115 31485 5135
rect 31465 5065 31485 5085
rect 31465 5015 31485 5035
rect 32065 5465 32085 5485
rect 32065 5415 32085 5435
rect 32065 5365 32085 5385
rect 32065 5315 32085 5335
rect 32065 5265 32085 5285
rect 32065 5215 32085 5235
rect 32065 5165 32085 5185
rect 32065 5115 32085 5135
rect 32065 5065 32085 5085
rect 32065 5015 32085 5035
rect -635 4815 -615 4835
rect -635 4765 -615 4785
rect -635 4715 -615 4735
rect -635 4665 -615 4685
rect -635 4615 -615 4635
rect -635 4565 -615 4585
rect -635 4515 -615 4535
rect -635 4465 -615 4485
rect -635 4415 -615 4435
rect -635 4365 -615 4385
rect -485 4815 -465 4835
rect -485 4765 -465 4785
rect -485 4715 -465 4735
rect -485 4665 -465 4685
rect -485 4615 -465 4635
rect -485 4565 -465 4585
rect -485 4515 -465 4535
rect -485 4465 -465 4485
rect -485 4415 -465 4435
rect -485 4365 -465 4385
rect -335 4815 -315 4835
rect -335 4765 -315 4785
rect -335 4715 -315 4735
rect -335 4665 -315 4685
rect -335 4615 -315 4635
rect -335 4565 -315 4585
rect -335 4515 -315 4535
rect -335 4465 -315 4485
rect -335 4415 -315 4435
rect -335 4365 -315 4385
rect -185 4815 -165 4835
rect -185 4765 -165 4785
rect -185 4715 -165 4735
rect -185 4665 -165 4685
rect -185 4615 -165 4635
rect -185 4565 -165 4585
rect -185 4515 -165 4535
rect -185 4465 -165 4485
rect -185 4415 -165 4435
rect -185 4365 -165 4385
rect -35 4815 -15 4835
rect -35 4765 -15 4785
rect -35 4715 -15 4735
rect -35 4665 -15 4685
rect -35 4615 -15 4635
rect -35 4565 -15 4585
rect -35 4515 -15 4535
rect -35 4465 -15 4485
rect -35 4415 -15 4435
rect -35 4365 -15 4385
rect 565 4815 585 4835
rect 565 4765 585 4785
rect 565 4715 585 4735
rect 565 4665 585 4685
rect 565 4615 585 4635
rect 565 4565 585 4585
rect 565 4515 585 4535
rect 565 4465 585 4485
rect 565 4415 585 4435
rect 565 4365 585 4385
rect 715 4815 735 4835
rect 715 4765 735 4785
rect 715 4715 735 4735
rect 715 4665 735 4685
rect 715 4615 735 4635
rect 715 4565 735 4585
rect 715 4515 735 4535
rect 715 4465 735 4485
rect 715 4415 735 4435
rect 715 4365 735 4385
rect 865 4815 885 4835
rect 865 4765 885 4785
rect 865 4715 885 4735
rect 865 4665 885 4685
rect 865 4615 885 4635
rect 865 4565 885 4585
rect 865 4515 885 4535
rect 865 4465 885 4485
rect 865 4415 885 4435
rect 865 4365 885 4385
rect 1015 4815 1035 4835
rect 1015 4765 1035 4785
rect 1015 4715 1035 4735
rect 1015 4665 1035 4685
rect 1015 4615 1035 4635
rect 1015 4565 1035 4585
rect 1015 4515 1035 4535
rect 1015 4465 1035 4485
rect 1015 4415 1035 4435
rect 1015 4365 1035 4385
rect 1165 4815 1185 4835
rect 1165 4765 1185 4785
rect 1165 4715 1185 4735
rect 1165 4665 1185 4685
rect 1165 4615 1185 4635
rect 1165 4565 1185 4585
rect 1165 4515 1185 4535
rect 1165 4465 1185 4485
rect 1165 4415 1185 4435
rect 1165 4365 1185 4385
rect 1315 4815 1335 4835
rect 1315 4765 1335 4785
rect 1315 4715 1335 4735
rect 1315 4665 1335 4685
rect 1315 4615 1335 4635
rect 1315 4565 1335 4585
rect 1315 4515 1335 4535
rect 1315 4465 1335 4485
rect 1315 4415 1335 4435
rect 1315 4365 1335 4385
rect 1465 4815 1485 4835
rect 1465 4765 1485 4785
rect 1465 4715 1485 4735
rect 1465 4665 1485 4685
rect 1465 4615 1485 4635
rect 1465 4565 1485 4585
rect 1465 4515 1485 4535
rect 1465 4465 1485 4485
rect 1465 4415 1485 4435
rect 1465 4365 1485 4385
rect 1615 4815 1635 4835
rect 1615 4765 1635 4785
rect 1615 4715 1635 4735
rect 1615 4665 1635 4685
rect 1615 4615 1635 4635
rect 1615 4565 1635 4585
rect 1615 4515 1635 4535
rect 1615 4465 1635 4485
rect 1615 4415 1635 4435
rect 1615 4365 1635 4385
rect 1765 4815 1785 4835
rect 1765 4765 1785 4785
rect 1765 4715 1785 4735
rect 1765 4665 1785 4685
rect 1765 4615 1785 4635
rect 1765 4565 1785 4585
rect 1765 4515 1785 4535
rect 1765 4465 1785 4485
rect 1765 4415 1785 4435
rect 1765 4365 1785 4385
rect 1915 4815 1935 4835
rect 1915 4765 1935 4785
rect 1915 4715 1935 4735
rect 1915 4665 1935 4685
rect 1915 4615 1935 4635
rect 1915 4565 1935 4585
rect 1915 4515 1935 4535
rect 1915 4465 1935 4485
rect 1915 4415 1935 4435
rect 1915 4365 1935 4385
rect 2065 4815 2085 4835
rect 2065 4765 2085 4785
rect 2065 4715 2085 4735
rect 2065 4665 2085 4685
rect 2065 4615 2085 4635
rect 2065 4565 2085 4585
rect 2065 4515 2085 4535
rect 2065 4465 2085 4485
rect 2065 4415 2085 4435
rect 2065 4365 2085 4385
rect 2215 4815 2235 4835
rect 2215 4765 2235 4785
rect 2215 4715 2235 4735
rect 2215 4665 2235 4685
rect 2215 4615 2235 4635
rect 2215 4565 2235 4585
rect 2215 4515 2235 4535
rect 2215 4465 2235 4485
rect 2215 4415 2235 4435
rect 2215 4365 2235 4385
rect 2365 4815 2385 4835
rect 2365 4765 2385 4785
rect 2365 4715 2385 4735
rect 2365 4665 2385 4685
rect 2365 4615 2385 4635
rect 2365 4565 2385 4585
rect 2365 4515 2385 4535
rect 2365 4465 2385 4485
rect 2365 4415 2385 4435
rect 2365 4365 2385 4385
rect 2515 4815 2535 4835
rect 2515 4765 2535 4785
rect 2515 4715 2535 4735
rect 2515 4665 2535 4685
rect 2515 4615 2535 4635
rect 2515 4565 2535 4585
rect 2515 4515 2535 4535
rect 2515 4465 2535 4485
rect 2515 4415 2535 4435
rect 2515 4365 2535 4385
rect 2665 4815 2685 4835
rect 2665 4765 2685 4785
rect 2665 4715 2685 4735
rect 2665 4665 2685 4685
rect 2665 4615 2685 4635
rect 2665 4565 2685 4585
rect 2665 4515 2685 4535
rect 2665 4465 2685 4485
rect 2665 4415 2685 4435
rect 2665 4365 2685 4385
rect 2815 4815 2835 4835
rect 2815 4765 2835 4785
rect 2815 4715 2835 4735
rect 2815 4665 2835 4685
rect 2815 4615 2835 4635
rect 2815 4565 2835 4585
rect 2815 4515 2835 4535
rect 2815 4465 2835 4485
rect 2815 4415 2835 4435
rect 2815 4365 2835 4385
rect 2965 4815 2985 4835
rect 2965 4765 2985 4785
rect 2965 4715 2985 4735
rect 2965 4665 2985 4685
rect 2965 4615 2985 4635
rect 2965 4565 2985 4585
rect 2965 4515 2985 4535
rect 2965 4465 2985 4485
rect 2965 4415 2985 4435
rect 2965 4365 2985 4385
rect 3115 4815 3135 4835
rect 3115 4765 3135 4785
rect 3115 4715 3135 4735
rect 3115 4665 3135 4685
rect 3115 4615 3135 4635
rect 3115 4565 3135 4585
rect 3115 4515 3135 4535
rect 3115 4465 3135 4485
rect 3115 4415 3135 4435
rect 3115 4365 3135 4385
rect 3265 4815 3285 4835
rect 3265 4765 3285 4785
rect 3265 4715 3285 4735
rect 3265 4665 3285 4685
rect 3265 4615 3285 4635
rect 3265 4565 3285 4585
rect 3265 4515 3285 4535
rect 3265 4465 3285 4485
rect 3265 4415 3285 4435
rect 3265 4365 3285 4385
rect 3415 4815 3435 4835
rect 3415 4765 3435 4785
rect 3415 4715 3435 4735
rect 3415 4665 3435 4685
rect 3415 4615 3435 4635
rect 3415 4565 3435 4585
rect 3415 4515 3435 4535
rect 3415 4465 3435 4485
rect 3415 4415 3435 4435
rect 3415 4365 3435 4385
rect 3565 4815 3585 4835
rect 3565 4765 3585 4785
rect 3565 4715 3585 4735
rect 3565 4665 3585 4685
rect 3565 4615 3585 4635
rect 3565 4565 3585 4585
rect 3565 4515 3585 4535
rect 3565 4465 3585 4485
rect 3565 4415 3585 4435
rect 3565 4365 3585 4385
rect 4165 4815 4185 4835
rect 4165 4765 4185 4785
rect 4165 4715 4185 4735
rect 4165 4665 4185 4685
rect 4165 4615 4185 4635
rect 4165 4565 4185 4585
rect 4165 4515 4185 4535
rect 4165 4465 4185 4485
rect 4165 4415 4185 4435
rect 4165 4365 4185 4385
rect 4765 4815 4785 4835
rect 4765 4765 4785 4785
rect 4765 4715 4785 4735
rect 4765 4665 4785 4685
rect 4765 4615 4785 4635
rect 4765 4565 4785 4585
rect 4765 4515 4785 4535
rect 4765 4465 4785 4485
rect 4765 4415 4785 4435
rect 4765 4365 4785 4385
rect 4915 4815 4935 4835
rect 4915 4765 4935 4785
rect 4915 4715 4935 4735
rect 4915 4665 4935 4685
rect 4915 4615 4935 4635
rect 4915 4565 4935 4585
rect 4915 4515 4935 4535
rect 4915 4465 4935 4485
rect 4915 4415 4935 4435
rect 4915 4365 4935 4385
rect 5065 4815 5085 4835
rect 5065 4765 5085 4785
rect 5065 4715 5085 4735
rect 5065 4665 5085 4685
rect 5065 4615 5085 4635
rect 5065 4565 5085 4585
rect 5065 4515 5085 4535
rect 5065 4465 5085 4485
rect 5065 4415 5085 4435
rect 5065 4365 5085 4385
rect 5215 4815 5235 4835
rect 5215 4765 5235 4785
rect 5215 4715 5235 4735
rect 5215 4665 5235 4685
rect 5215 4615 5235 4635
rect 5215 4565 5235 4585
rect 5215 4515 5235 4535
rect 5215 4465 5235 4485
rect 5215 4415 5235 4435
rect 5215 4365 5235 4385
rect 5365 4815 5385 4835
rect 5365 4765 5385 4785
rect 5365 4715 5385 4735
rect 5365 4665 5385 4685
rect 5365 4615 5385 4635
rect 5365 4565 5385 4585
rect 5365 4515 5385 4535
rect 5365 4465 5385 4485
rect 5365 4415 5385 4435
rect 5365 4365 5385 4385
rect 5515 4815 5535 4835
rect 5515 4765 5535 4785
rect 5515 4715 5535 4735
rect 5515 4665 5535 4685
rect 5515 4615 5535 4635
rect 5515 4565 5535 4585
rect 5515 4515 5535 4535
rect 5515 4465 5535 4485
rect 5515 4415 5535 4435
rect 5515 4365 5535 4385
rect 5665 4815 5685 4835
rect 5665 4765 5685 4785
rect 5665 4715 5685 4735
rect 5665 4665 5685 4685
rect 5665 4615 5685 4635
rect 5665 4565 5685 4585
rect 5665 4515 5685 4535
rect 5665 4465 5685 4485
rect 5665 4415 5685 4435
rect 5665 4365 5685 4385
rect 5815 4815 5835 4835
rect 5815 4765 5835 4785
rect 5815 4715 5835 4735
rect 5815 4665 5835 4685
rect 5815 4615 5835 4635
rect 5815 4565 5835 4585
rect 5815 4515 5835 4535
rect 5815 4465 5835 4485
rect 5815 4415 5835 4435
rect 5815 4365 5835 4385
rect 5965 4815 5985 4835
rect 5965 4765 5985 4785
rect 5965 4715 5985 4735
rect 5965 4665 5985 4685
rect 5965 4615 5985 4635
rect 5965 4565 5985 4585
rect 5965 4515 5985 4535
rect 5965 4465 5985 4485
rect 5965 4415 5985 4435
rect 5965 4365 5985 4385
rect 6115 4815 6135 4835
rect 6115 4765 6135 4785
rect 6115 4715 6135 4735
rect 6115 4665 6135 4685
rect 6115 4615 6135 4635
rect 6115 4565 6135 4585
rect 6115 4515 6135 4535
rect 6115 4465 6135 4485
rect 6115 4415 6135 4435
rect 6115 4365 6135 4385
rect 6265 4815 6285 4835
rect 6265 4765 6285 4785
rect 6265 4715 6285 4735
rect 6265 4665 6285 4685
rect 6265 4615 6285 4635
rect 6265 4565 6285 4585
rect 6265 4515 6285 4535
rect 6265 4465 6285 4485
rect 6265 4415 6285 4435
rect 6265 4365 6285 4385
rect 6415 4815 6435 4835
rect 6415 4765 6435 4785
rect 6415 4715 6435 4735
rect 6415 4665 6435 4685
rect 6415 4615 6435 4635
rect 6415 4565 6435 4585
rect 6415 4515 6435 4535
rect 6415 4465 6435 4485
rect 6415 4415 6435 4435
rect 6415 4365 6435 4385
rect 6565 4815 6585 4835
rect 6565 4765 6585 4785
rect 6565 4715 6585 4735
rect 6565 4665 6585 4685
rect 6565 4615 6585 4635
rect 6565 4565 6585 4585
rect 6565 4515 6585 4535
rect 6565 4465 6585 4485
rect 6565 4415 6585 4435
rect 6565 4365 6585 4385
rect 6715 4815 6735 4835
rect 6715 4765 6735 4785
rect 6715 4715 6735 4735
rect 6715 4665 6735 4685
rect 6715 4615 6735 4635
rect 6715 4565 6735 4585
rect 6715 4515 6735 4535
rect 6715 4465 6735 4485
rect 6715 4415 6735 4435
rect 6715 4365 6735 4385
rect 6865 4815 6885 4835
rect 6865 4765 6885 4785
rect 6865 4715 6885 4735
rect 6865 4665 6885 4685
rect 6865 4615 6885 4635
rect 6865 4565 6885 4585
rect 6865 4515 6885 4535
rect 6865 4465 6885 4485
rect 6865 4415 6885 4435
rect 6865 4365 6885 4385
rect 7015 4815 7035 4835
rect 7015 4765 7035 4785
rect 7015 4715 7035 4735
rect 7015 4665 7035 4685
rect 7015 4615 7035 4635
rect 7015 4565 7035 4585
rect 7015 4515 7035 4535
rect 7015 4465 7035 4485
rect 7015 4415 7035 4435
rect 7015 4365 7035 4385
rect 7165 4815 7185 4835
rect 7165 4765 7185 4785
rect 7165 4715 7185 4735
rect 7165 4665 7185 4685
rect 7165 4615 7185 4635
rect 7165 4565 7185 4585
rect 7165 4515 7185 4535
rect 7165 4465 7185 4485
rect 7165 4415 7185 4435
rect 7165 4365 7185 4385
rect 7315 4815 7335 4835
rect 7315 4765 7335 4785
rect 7315 4715 7335 4735
rect 7315 4665 7335 4685
rect 7315 4615 7335 4635
rect 7315 4565 7335 4585
rect 7315 4515 7335 4535
rect 7315 4465 7335 4485
rect 7315 4415 7335 4435
rect 7315 4365 7335 4385
rect 7465 4815 7485 4835
rect 7465 4765 7485 4785
rect 7465 4715 7485 4735
rect 7465 4665 7485 4685
rect 7465 4615 7485 4635
rect 7465 4565 7485 4585
rect 7465 4515 7485 4535
rect 7465 4465 7485 4485
rect 7465 4415 7485 4435
rect 7465 4365 7485 4385
rect 7615 4815 7635 4835
rect 7615 4765 7635 4785
rect 7615 4715 7635 4735
rect 7615 4665 7635 4685
rect 7615 4615 7635 4635
rect 7615 4565 7635 4585
rect 7615 4515 7635 4535
rect 7615 4465 7635 4485
rect 7615 4415 7635 4435
rect 7615 4365 7635 4385
rect 7765 4815 7785 4835
rect 7765 4765 7785 4785
rect 7765 4715 7785 4735
rect 7765 4665 7785 4685
rect 7765 4615 7785 4635
rect 7765 4565 7785 4585
rect 7765 4515 7785 4535
rect 7765 4465 7785 4485
rect 7765 4415 7785 4435
rect 7765 4365 7785 4385
rect 8365 4815 8385 4835
rect 8365 4765 8385 4785
rect 8365 4715 8385 4735
rect 8365 4665 8385 4685
rect 8365 4615 8385 4635
rect 8365 4565 8385 4585
rect 8365 4515 8385 4535
rect 8365 4465 8385 4485
rect 8365 4415 8385 4435
rect 8365 4365 8385 4385
rect 8515 4815 8535 4835
rect 8515 4765 8535 4785
rect 8515 4715 8535 4735
rect 8515 4665 8535 4685
rect 8515 4615 8535 4635
rect 8515 4565 8535 4585
rect 8515 4515 8535 4535
rect 8515 4465 8535 4485
rect 8515 4415 8535 4435
rect 8515 4365 8535 4385
rect 8665 4815 8685 4835
rect 8665 4765 8685 4785
rect 8665 4715 8685 4735
rect 8665 4665 8685 4685
rect 8665 4615 8685 4635
rect 8665 4565 8685 4585
rect 8665 4515 8685 4535
rect 8665 4465 8685 4485
rect 8665 4415 8685 4435
rect 8665 4365 8685 4385
rect 8815 4815 8835 4835
rect 8815 4765 8835 4785
rect 8815 4715 8835 4735
rect 8815 4665 8835 4685
rect 8815 4615 8835 4635
rect 8815 4565 8835 4585
rect 8815 4515 8835 4535
rect 8815 4465 8835 4485
rect 8815 4415 8835 4435
rect 8815 4365 8835 4385
rect 8965 4815 8985 4835
rect 8965 4765 8985 4785
rect 8965 4715 8985 4735
rect 8965 4665 8985 4685
rect 8965 4615 8985 4635
rect 8965 4565 8985 4585
rect 8965 4515 8985 4535
rect 8965 4465 8985 4485
rect 8965 4415 8985 4435
rect 8965 4365 8985 4385
rect 9115 4815 9135 4835
rect 9115 4765 9135 4785
rect 9115 4715 9135 4735
rect 9115 4665 9135 4685
rect 9115 4615 9135 4635
rect 9115 4565 9135 4585
rect 9115 4515 9135 4535
rect 9115 4465 9135 4485
rect 9115 4415 9135 4435
rect 9115 4365 9135 4385
rect 9265 4815 9285 4835
rect 9265 4765 9285 4785
rect 9265 4715 9285 4735
rect 9265 4665 9285 4685
rect 9265 4615 9285 4635
rect 9265 4565 9285 4585
rect 9265 4515 9285 4535
rect 9265 4465 9285 4485
rect 9265 4415 9285 4435
rect 9265 4365 9285 4385
rect 9415 4815 9435 4835
rect 9415 4765 9435 4785
rect 9415 4715 9435 4735
rect 9415 4665 9435 4685
rect 9415 4615 9435 4635
rect 9415 4565 9435 4585
rect 9415 4515 9435 4535
rect 9415 4465 9435 4485
rect 9415 4415 9435 4435
rect 9415 4365 9435 4385
rect 9565 4815 9585 4835
rect 9565 4765 9585 4785
rect 9565 4715 9585 4735
rect 9565 4665 9585 4685
rect 9565 4615 9585 4635
rect 9565 4565 9585 4585
rect 9565 4515 9585 4535
rect 9565 4465 9585 4485
rect 9565 4415 9585 4435
rect 9565 4365 9585 4385
rect 9715 4815 9735 4835
rect 9715 4765 9735 4785
rect 9715 4715 9735 4735
rect 9715 4665 9735 4685
rect 9715 4615 9735 4635
rect 9715 4565 9735 4585
rect 9715 4515 9735 4535
rect 9715 4465 9735 4485
rect 9715 4415 9735 4435
rect 9715 4365 9735 4385
rect 9865 4815 9885 4835
rect 9865 4765 9885 4785
rect 9865 4715 9885 4735
rect 9865 4665 9885 4685
rect 9865 4615 9885 4635
rect 9865 4565 9885 4585
rect 9865 4515 9885 4535
rect 9865 4465 9885 4485
rect 9865 4415 9885 4435
rect 9865 4365 9885 4385
rect 10015 4815 10035 4835
rect 10015 4765 10035 4785
rect 10015 4715 10035 4735
rect 10015 4665 10035 4685
rect 10015 4615 10035 4635
rect 10015 4565 10035 4585
rect 10015 4515 10035 4535
rect 10015 4465 10035 4485
rect 10015 4415 10035 4435
rect 10015 4365 10035 4385
rect 10165 4815 10185 4835
rect 10165 4765 10185 4785
rect 10165 4715 10185 4735
rect 10165 4665 10185 4685
rect 10165 4615 10185 4635
rect 10165 4565 10185 4585
rect 10165 4515 10185 4535
rect 10165 4465 10185 4485
rect 10165 4415 10185 4435
rect 10165 4365 10185 4385
rect 10315 4815 10335 4835
rect 10315 4765 10335 4785
rect 10315 4715 10335 4735
rect 10315 4665 10335 4685
rect 10315 4615 10335 4635
rect 10315 4565 10335 4585
rect 10315 4515 10335 4535
rect 10315 4465 10335 4485
rect 10315 4415 10335 4435
rect 10315 4365 10335 4385
rect 10465 4815 10485 4835
rect 10465 4765 10485 4785
rect 10465 4715 10485 4735
rect 10465 4665 10485 4685
rect 10465 4615 10485 4635
rect 10465 4565 10485 4585
rect 10465 4515 10485 4535
rect 10465 4465 10485 4485
rect 10465 4415 10485 4435
rect 10465 4365 10485 4385
rect 10615 4815 10635 4835
rect 10615 4765 10635 4785
rect 10615 4715 10635 4735
rect 10615 4665 10635 4685
rect 10615 4615 10635 4635
rect 10615 4565 10635 4585
rect 10615 4515 10635 4535
rect 10615 4465 10635 4485
rect 10615 4415 10635 4435
rect 10615 4365 10635 4385
rect 10765 4815 10785 4835
rect 10765 4765 10785 4785
rect 10765 4715 10785 4735
rect 10765 4665 10785 4685
rect 10765 4615 10785 4635
rect 10765 4565 10785 4585
rect 10765 4515 10785 4535
rect 10765 4465 10785 4485
rect 10765 4415 10785 4435
rect 10765 4365 10785 4385
rect 11365 4815 11385 4835
rect 11365 4765 11385 4785
rect 11365 4715 11385 4735
rect 11365 4665 11385 4685
rect 11365 4615 11385 4635
rect 11365 4565 11385 4585
rect 11365 4515 11385 4535
rect 11365 4465 11385 4485
rect 11365 4415 11385 4435
rect 11365 4365 11385 4385
rect 11965 4815 11985 4835
rect 11965 4765 11985 4785
rect 11965 4715 11985 4735
rect 11965 4665 11985 4685
rect 11965 4615 11985 4635
rect 11965 4565 11985 4585
rect 11965 4515 11985 4535
rect 11965 4465 11985 4485
rect 11965 4415 11985 4435
rect 11965 4365 11985 4385
rect 12565 4815 12585 4835
rect 12565 4765 12585 4785
rect 12565 4715 12585 4735
rect 12565 4665 12585 4685
rect 12565 4615 12585 4635
rect 12565 4565 12585 4585
rect 12565 4515 12585 4535
rect 12565 4465 12585 4485
rect 12565 4415 12585 4435
rect 12565 4365 12585 4385
rect 13165 4815 13185 4835
rect 13165 4765 13185 4785
rect 13165 4715 13185 4735
rect 13165 4665 13185 4685
rect 13165 4615 13185 4635
rect 13165 4565 13185 4585
rect 13165 4515 13185 4535
rect 13165 4465 13185 4485
rect 13165 4415 13185 4435
rect 13165 4365 13185 4385
rect 13765 4815 13785 4835
rect 13765 4765 13785 4785
rect 13765 4715 13785 4735
rect 13765 4665 13785 4685
rect 13765 4615 13785 4635
rect 13765 4565 13785 4585
rect 13765 4515 13785 4535
rect 13765 4465 13785 4485
rect 13765 4415 13785 4435
rect 13765 4365 13785 4385
rect 14365 4815 14385 4835
rect 14365 4765 14385 4785
rect 14365 4715 14385 4735
rect 14365 4665 14385 4685
rect 14365 4615 14385 4635
rect 14365 4565 14385 4585
rect 14365 4515 14385 4535
rect 14365 4465 14385 4485
rect 14365 4415 14385 4435
rect 14365 4365 14385 4385
rect 14965 4815 14985 4835
rect 14965 4765 14985 4785
rect 14965 4715 14985 4735
rect 14965 4665 14985 4685
rect 14965 4615 14985 4635
rect 14965 4565 14985 4585
rect 14965 4515 14985 4535
rect 14965 4465 14985 4485
rect 14965 4415 14985 4435
rect 14965 4365 14985 4385
rect 15565 4815 15585 4835
rect 15565 4765 15585 4785
rect 15565 4715 15585 4735
rect 15565 4665 15585 4685
rect 15565 4615 15585 4635
rect 15565 4565 15585 4585
rect 15565 4515 15585 4535
rect 15565 4465 15585 4485
rect 15565 4415 15585 4435
rect 15565 4365 15585 4385
rect 16165 4815 16185 4835
rect 16165 4765 16185 4785
rect 16165 4715 16185 4735
rect 16165 4665 16185 4685
rect 16165 4615 16185 4635
rect 16165 4565 16185 4585
rect 16165 4515 16185 4535
rect 16165 4465 16185 4485
rect 16165 4415 16185 4435
rect 16165 4365 16185 4385
rect 16315 4815 16335 4835
rect 16315 4765 16335 4785
rect 16315 4715 16335 4735
rect 16315 4665 16335 4685
rect 16315 4615 16335 4635
rect 16315 4565 16335 4585
rect 16315 4515 16335 4535
rect 16315 4465 16335 4485
rect 16315 4415 16335 4435
rect 16315 4365 16335 4385
rect 16465 4815 16485 4835
rect 16465 4765 16485 4785
rect 16465 4715 16485 4735
rect 16465 4665 16485 4685
rect 16465 4615 16485 4635
rect 16465 4565 16485 4585
rect 16465 4515 16485 4535
rect 16465 4465 16485 4485
rect 16465 4415 16485 4435
rect 16465 4365 16485 4385
rect 16615 4815 16635 4835
rect 16615 4765 16635 4785
rect 16615 4715 16635 4735
rect 16615 4665 16635 4685
rect 16615 4615 16635 4635
rect 16615 4565 16635 4585
rect 16615 4515 16635 4535
rect 16615 4465 16635 4485
rect 16615 4415 16635 4435
rect 16615 4365 16635 4385
rect 16765 4815 16785 4835
rect 16765 4765 16785 4785
rect 16765 4715 16785 4735
rect 16765 4665 16785 4685
rect 16765 4615 16785 4635
rect 16765 4565 16785 4585
rect 16765 4515 16785 4535
rect 16765 4465 16785 4485
rect 16765 4415 16785 4435
rect 16765 4365 16785 4385
rect 16915 4815 16935 4835
rect 16915 4765 16935 4785
rect 16915 4715 16935 4735
rect 16915 4665 16935 4685
rect 16915 4615 16935 4635
rect 16915 4565 16935 4585
rect 16915 4515 16935 4535
rect 16915 4465 16935 4485
rect 16915 4415 16935 4435
rect 16915 4365 16935 4385
rect 17065 4815 17085 4835
rect 17065 4765 17085 4785
rect 17065 4715 17085 4735
rect 17065 4665 17085 4685
rect 17065 4615 17085 4635
rect 17065 4565 17085 4585
rect 17065 4515 17085 4535
rect 17065 4465 17085 4485
rect 17065 4415 17085 4435
rect 17065 4365 17085 4385
rect 17215 4815 17235 4835
rect 17215 4765 17235 4785
rect 17215 4715 17235 4735
rect 17215 4665 17235 4685
rect 17215 4615 17235 4635
rect 17215 4565 17235 4585
rect 17215 4515 17235 4535
rect 17215 4465 17235 4485
rect 17215 4415 17235 4435
rect 17215 4365 17235 4385
rect 17365 4815 17385 4835
rect 17365 4765 17385 4785
rect 17365 4715 17385 4735
rect 17365 4665 17385 4685
rect 17365 4615 17385 4635
rect 17365 4565 17385 4585
rect 17365 4515 17385 4535
rect 17365 4465 17385 4485
rect 17365 4415 17385 4435
rect 17365 4365 17385 4385
rect 17965 4815 17985 4835
rect 17965 4765 17985 4785
rect 17965 4715 17985 4735
rect 17965 4665 17985 4685
rect 17965 4615 17985 4635
rect 17965 4565 17985 4585
rect 17965 4515 17985 4535
rect 17965 4465 17985 4485
rect 17965 4415 17985 4435
rect 17965 4365 17985 4385
rect 18565 4815 18585 4835
rect 18565 4765 18585 4785
rect 18565 4715 18585 4735
rect 18565 4665 18585 4685
rect 18565 4615 18585 4635
rect 18565 4565 18585 4585
rect 18565 4515 18585 4535
rect 18565 4465 18585 4485
rect 18565 4415 18585 4435
rect 18565 4365 18585 4385
rect 18715 4815 18735 4835
rect 18715 4765 18735 4785
rect 18715 4715 18735 4735
rect 18715 4665 18735 4685
rect 18715 4615 18735 4635
rect 18715 4565 18735 4585
rect 18715 4515 18735 4535
rect 18715 4465 18735 4485
rect 18715 4415 18735 4435
rect 18715 4365 18735 4385
rect 18865 4815 18885 4835
rect 18865 4765 18885 4785
rect 18865 4715 18885 4735
rect 18865 4665 18885 4685
rect 18865 4615 18885 4635
rect 18865 4565 18885 4585
rect 18865 4515 18885 4535
rect 18865 4465 18885 4485
rect 18865 4415 18885 4435
rect 18865 4365 18885 4385
rect 19015 4815 19035 4835
rect 19015 4765 19035 4785
rect 19015 4715 19035 4735
rect 19015 4665 19035 4685
rect 19015 4615 19035 4635
rect 19015 4565 19035 4585
rect 19015 4515 19035 4535
rect 19015 4465 19035 4485
rect 19015 4415 19035 4435
rect 19015 4365 19035 4385
rect 19165 4815 19185 4835
rect 19165 4765 19185 4785
rect 19165 4715 19185 4735
rect 19165 4665 19185 4685
rect 19165 4615 19185 4635
rect 19165 4565 19185 4585
rect 19165 4515 19185 4535
rect 19165 4465 19185 4485
rect 19165 4415 19185 4435
rect 19165 4365 19185 4385
rect 19315 4815 19335 4835
rect 19315 4765 19335 4785
rect 19315 4715 19335 4735
rect 19315 4665 19335 4685
rect 19315 4615 19335 4635
rect 19315 4565 19335 4585
rect 19315 4515 19335 4535
rect 19315 4465 19335 4485
rect 19315 4415 19335 4435
rect 19315 4365 19335 4385
rect 19465 4815 19485 4835
rect 19465 4765 19485 4785
rect 19465 4715 19485 4735
rect 19465 4665 19485 4685
rect 19465 4615 19485 4635
rect 19465 4565 19485 4585
rect 19465 4515 19485 4535
rect 19465 4465 19485 4485
rect 19465 4415 19485 4435
rect 19465 4365 19485 4385
rect 19615 4815 19635 4835
rect 19615 4765 19635 4785
rect 19615 4715 19635 4735
rect 19615 4665 19635 4685
rect 19615 4615 19635 4635
rect 19615 4565 19635 4585
rect 19615 4515 19635 4535
rect 19615 4465 19635 4485
rect 19615 4415 19635 4435
rect 19615 4365 19635 4385
rect 19765 4815 19785 4835
rect 19765 4765 19785 4785
rect 19765 4715 19785 4735
rect 19765 4665 19785 4685
rect 19765 4615 19785 4635
rect 19765 4565 19785 4585
rect 19765 4515 19785 4535
rect 19765 4465 19785 4485
rect 19765 4415 19785 4435
rect 19765 4365 19785 4385
rect 20365 4815 20385 4835
rect 20365 4765 20385 4785
rect 20365 4715 20385 4735
rect 20365 4665 20385 4685
rect 20365 4615 20385 4635
rect 20365 4565 20385 4585
rect 20365 4515 20385 4535
rect 20365 4465 20385 4485
rect 20365 4415 20385 4435
rect 20365 4365 20385 4385
rect 20965 4815 20985 4835
rect 20965 4765 20985 4785
rect 20965 4715 20985 4735
rect 20965 4665 20985 4685
rect 20965 4615 20985 4635
rect 20965 4565 20985 4585
rect 20965 4515 20985 4535
rect 20965 4465 20985 4485
rect 20965 4415 20985 4435
rect 20965 4365 20985 4385
rect 21415 4815 21435 4835
rect 21415 4765 21435 4785
rect 21415 4715 21435 4735
rect 21415 4665 21435 4685
rect 21415 4615 21435 4635
rect 21415 4565 21435 4585
rect 21415 4515 21435 4535
rect 21415 4465 21435 4485
rect 21415 4415 21435 4435
rect 21415 4365 21435 4385
rect 21865 4815 21885 4835
rect 21865 4765 21885 4785
rect 21865 4715 21885 4735
rect 21865 4665 21885 4685
rect 21865 4615 21885 4635
rect 21865 4565 21885 4585
rect 21865 4515 21885 4535
rect 21865 4465 21885 4485
rect 21865 4415 21885 4435
rect 21865 4365 21885 4385
rect 22465 4815 22485 4835
rect 22465 4765 22485 4785
rect 22465 4715 22485 4735
rect 22465 4665 22485 4685
rect 22465 4615 22485 4635
rect 22465 4565 22485 4585
rect 22465 4515 22485 4535
rect 22465 4465 22485 4485
rect 22465 4415 22485 4435
rect 22465 4365 22485 4385
rect 23065 4815 23085 4835
rect 23065 4765 23085 4785
rect 23065 4715 23085 4735
rect 23065 4665 23085 4685
rect 23065 4615 23085 4635
rect 23065 4565 23085 4585
rect 23065 4515 23085 4535
rect 23065 4465 23085 4485
rect 23065 4415 23085 4435
rect 23065 4365 23085 4385
rect 23515 4815 23535 4835
rect 23515 4765 23535 4785
rect 23515 4715 23535 4735
rect 23515 4665 23535 4685
rect 23515 4615 23535 4635
rect 23515 4565 23535 4585
rect 23515 4515 23535 4535
rect 23515 4465 23535 4485
rect 23515 4415 23535 4435
rect 23515 4365 23535 4385
rect 23965 4815 23985 4835
rect 23965 4765 23985 4785
rect 23965 4715 23985 4735
rect 23965 4665 23985 4685
rect 23965 4615 23985 4635
rect 23965 4565 23985 4585
rect 23965 4515 23985 4535
rect 23965 4465 23985 4485
rect 23965 4415 23985 4435
rect 23965 4365 23985 4385
rect 24565 4815 24585 4835
rect 24565 4765 24585 4785
rect 24565 4715 24585 4735
rect 24565 4665 24585 4685
rect 24565 4615 24585 4635
rect 24565 4565 24585 4585
rect 24565 4515 24585 4535
rect 24565 4465 24585 4485
rect 24565 4415 24585 4435
rect 24565 4365 24585 4385
rect 25165 4815 25185 4835
rect 25165 4765 25185 4785
rect 25165 4715 25185 4735
rect 25165 4665 25185 4685
rect 25165 4615 25185 4635
rect 25165 4565 25185 4585
rect 25165 4515 25185 4535
rect 25165 4465 25185 4485
rect 25165 4415 25185 4435
rect 25165 4365 25185 4385
rect 25615 4815 25635 4835
rect 25615 4765 25635 4785
rect 25615 4715 25635 4735
rect 25615 4665 25635 4685
rect 25615 4615 25635 4635
rect 25615 4565 25635 4585
rect 25615 4515 25635 4535
rect 25615 4465 25635 4485
rect 25615 4415 25635 4435
rect 25615 4365 25635 4385
rect 26065 4815 26085 4835
rect 26065 4765 26085 4785
rect 26065 4715 26085 4735
rect 26065 4665 26085 4685
rect 26065 4615 26085 4635
rect 26065 4565 26085 4585
rect 26065 4515 26085 4535
rect 26065 4465 26085 4485
rect 26065 4415 26085 4435
rect 26065 4365 26085 4385
rect 26665 4815 26685 4835
rect 26665 4765 26685 4785
rect 26665 4715 26685 4735
rect 26665 4665 26685 4685
rect 26665 4615 26685 4635
rect 26665 4565 26685 4585
rect 26665 4515 26685 4535
rect 26665 4465 26685 4485
rect 26665 4415 26685 4435
rect 26665 4365 26685 4385
rect 27265 4815 27285 4835
rect 27265 4765 27285 4785
rect 27265 4715 27285 4735
rect 27265 4665 27285 4685
rect 27265 4615 27285 4635
rect 27265 4565 27285 4585
rect 27265 4515 27285 4535
rect 27265 4465 27285 4485
rect 27265 4415 27285 4435
rect 27265 4365 27285 4385
rect 27715 4815 27735 4835
rect 27715 4765 27735 4785
rect 27715 4715 27735 4735
rect 27715 4665 27735 4685
rect 27715 4615 27735 4635
rect 27715 4565 27735 4585
rect 27715 4515 27735 4535
rect 27715 4465 27735 4485
rect 27715 4415 27735 4435
rect 27715 4365 27735 4385
rect 28165 4815 28185 4835
rect 28165 4765 28185 4785
rect 28165 4715 28185 4735
rect 28165 4665 28185 4685
rect 28165 4615 28185 4635
rect 28165 4565 28185 4585
rect 28165 4515 28185 4535
rect 28165 4465 28185 4485
rect 28165 4415 28185 4435
rect 28165 4365 28185 4385
rect 28765 4815 28785 4835
rect 28765 4765 28785 4785
rect 28765 4715 28785 4735
rect 28765 4665 28785 4685
rect 28765 4615 28785 4635
rect 28765 4565 28785 4585
rect 28765 4515 28785 4535
rect 28765 4465 28785 4485
rect 28765 4415 28785 4435
rect 28765 4365 28785 4385
rect 29365 4815 29385 4835
rect 29365 4765 29385 4785
rect 29365 4715 29385 4735
rect 29365 4665 29385 4685
rect 29365 4615 29385 4635
rect 29365 4565 29385 4585
rect 29365 4515 29385 4535
rect 29365 4465 29385 4485
rect 29365 4415 29385 4435
rect 29365 4365 29385 4385
rect 29515 4815 29535 4835
rect 29515 4765 29535 4785
rect 29515 4715 29535 4735
rect 29515 4665 29535 4685
rect 29515 4615 29535 4635
rect 29515 4565 29535 4585
rect 29515 4515 29535 4535
rect 29515 4465 29535 4485
rect 29515 4415 29535 4435
rect 29515 4365 29535 4385
rect 29665 4815 29685 4835
rect 29665 4765 29685 4785
rect 29665 4715 29685 4735
rect 29665 4665 29685 4685
rect 29665 4615 29685 4635
rect 29665 4565 29685 4585
rect 29665 4515 29685 4535
rect 29665 4465 29685 4485
rect 29665 4415 29685 4435
rect 29665 4365 29685 4385
rect 29815 4815 29835 4835
rect 29815 4765 29835 4785
rect 29815 4715 29835 4735
rect 29815 4665 29835 4685
rect 29815 4615 29835 4635
rect 29815 4565 29835 4585
rect 29815 4515 29835 4535
rect 29815 4465 29835 4485
rect 29815 4415 29835 4435
rect 29815 4365 29835 4385
rect 29965 4815 29985 4835
rect 29965 4765 29985 4785
rect 29965 4715 29985 4735
rect 29965 4665 29985 4685
rect 29965 4615 29985 4635
rect 29965 4565 29985 4585
rect 29965 4515 29985 4535
rect 29965 4465 29985 4485
rect 29965 4415 29985 4435
rect 29965 4365 29985 4385
rect 30115 4815 30135 4835
rect 30115 4765 30135 4785
rect 30115 4715 30135 4735
rect 30115 4665 30135 4685
rect 30115 4615 30135 4635
rect 30115 4565 30135 4585
rect 30115 4515 30135 4535
rect 30115 4465 30135 4485
rect 30115 4415 30135 4435
rect 30115 4365 30135 4385
rect 30265 4815 30285 4835
rect 30265 4765 30285 4785
rect 30265 4715 30285 4735
rect 30265 4665 30285 4685
rect 30265 4615 30285 4635
rect 30265 4565 30285 4585
rect 30265 4515 30285 4535
rect 30265 4465 30285 4485
rect 30265 4415 30285 4435
rect 30265 4365 30285 4385
rect 30415 4815 30435 4835
rect 30415 4765 30435 4785
rect 30415 4715 30435 4735
rect 30415 4665 30435 4685
rect 30415 4615 30435 4635
rect 30415 4565 30435 4585
rect 30415 4515 30435 4535
rect 30415 4465 30435 4485
rect 30415 4415 30435 4435
rect 30415 4365 30435 4385
rect 30565 4815 30585 4835
rect 30565 4765 30585 4785
rect 30565 4715 30585 4735
rect 30565 4665 30585 4685
rect 30565 4615 30585 4635
rect 30565 4565 30585 4585
rect 30565 4515 30585 4535
rect 30565 4465 30585 4485
rect 30565 4415 30585 4435
rect 30565 4365 30585 4385
rect 30715 4815 30735 4835
rect 30715 4765 30735 4785
rect 30715 4715 30735 4735
rect 30715 4665 30735 4685
rect 30715 4615 30735 4635
rect 30715 4565 30735 4585
rect 30715 4515 30735 4535
rect 30715 4465 30735 4485
rect 30715 4415 30735 4435
rect 30715 4365 30735 4385
rect 30865 4815 30885 4835
rect 30865 4765 30885 4785
rect 30865 4715 30885 4735
rect 30865 4665 30885 4685
rect 30865 4615 30885 4635
rect 30865 4565 30885 4585
rect 30865 4515 30885 4535
rect 30865 4465 30885 4485
rect 30865 4415 30885 4435
rect 30865 4365 30885 4385
rect 31015 4815 31035 4835
rect 31015 4765 31035 4785
rect 31015 4715 31035 4735
rect 31015 4665 31035 4685
rect 31015 4615 31035 4635
rect 31015 4565 31035 4585
rect 31015 4515 31035 4535
rect 31015 4465 31035 4485
rect 31015 4415 31035 4435
rect 31015 4365 31035 4385
rect 31165 4815 31185 4835
rect 31165 4765 31185 4785
rect 31165 4715 31185 4735
rect 31165 4665 31185 4685
rect 31165 4615 31185 4635
rect 31165 4565 31185 4585
rect 31165 4515 31185 4535
rect 31165 4465 31185 4485
rect 31165 4415 31185 4435
rect 31165 4365 31185 4385
rect 31315 4815 31335 4835
rect 31315 4765 31335 4785
rect 31315 4715 31335 4735
rect 31315 4665 31335 4685
rect 31315 4615 31335 4635
rect 31315 4565 31335 4585
rect 31315 4515 31335 4535
rect 31315 4465 31335 4485
rect 31315 4415 31335 4435
rect 31315 4365 31335 4385
rect 31465 4815 31485 4835
rect 31465 4765 31485 4785
rect 31465 4715 31485 4735
rect 31465 4665 31485 4685
rect 31465 4615 31485 4635
rect 31465 4565 31485 4585
rect 31465 4515 31485 4535
rect 31465 4465 31485 4485
rect 31465 4415 31485 4435
rect 31465 4365 31485 4385
rect 32065 4815 32085 4835
rect 32065 4765 32085 4785
rect 32065 4715 32085 4735
rect 32065 4665 32085 4685
rect 32065 4615 32085 4635
rect 32065 4565 32085 4585
rect 32065 4515 32085 4535
rect 32065 4465 32085 4485
rect 32065 4415 32085 4435
rect 32065 4365 32085 4385
rect -635 4165 -615 4185
rect -635 4115 -615 4135
rect -635 4065 -615 4085
rect -635 4015 -615 4035
rect -635 3965 -615 3985
rect -635 3915 -615 3935
rect -635 3865 -615 3885
rect -635 3815 -615 3835
rect -635 3765 -615 3785
rect -635 3715 -615 3735
rect -485 4165 -465 4185
rect -485 4115 -465 4135
rect -485 4065 -465 4085
rect -485 4015 -465 4035
rect -485 3965 -465 3985
rect -485 3915 -465 3935
rect -485 3865 -465 3885
rect -485 3815 -465 3835
rect -485 3765 -465 3785
rect -485 3715 -465 3735
rect -335 4165 -315 4185
rect -335 4115 -315 4135
rect -335 4065 -315 4085
rect -335 4015 -315 4035
rect -335 3965 -315 3985
rect -335 3915 -315 3935
rect -335 3865 -315 3885
rect -335 3815 -315 3835
rect -335 3765 -315 3785
rect -335 3715 -315 3735
rect -185 4165 -165 4185
rect -185 4115 -165 4135
rect -185 4065 -165 4085
rect -185 4015 -165 4035
rect -185 3965 -165 3985
rect -185 3915 -165 3935
rect -185 3865 -165 3885
rect -185 3815 -165 3835
rect -185 3765 -165 3785
rect -185 3715 -165 3735
rect -35 4165 -15 4185
rect -35 4115 -15 4135
rect -35 4065 -15 4085
rect -35 4015 -15 4035
rect -35 3965 -15 3985
rect -35 3915 -15 3935
rect -35 3865 -15 3885
rect -35 3815 -15 3835
rect -35 3765 -15 3785
rect -35 3715 -15 3735
rect 565 4165 585 4185
rect 565 4115 585 4135
rect 565 4065 585 4085
rect 565 4015 585 4035
rect 565 3965 585 3985
rect 565 3915 585 3935
rect 565 3865 585 3885
rect 565 3815 585 3835
rect 565 3765 585 3785
rect 565 3715 585 3735
rect 715 4165 735 4185
rect 715 4115 735 4135
rect 715 4065 735 4085
rect 715 4015 735 4035
rect 715 3965 735 3985
rect 715 3915 735 3935
rect 715 3865 735 3885
rect 715 3815 735 3835
rect 715 3765 735 3785
rect 715 3715 735 3735
rect 865 4165 885 4185
rect 865 4115 885 4135
rect 865 4065 885 4085
rect 865 4015 885 4035
rect 865 3965 885 3985
rect 865 3915 885 3935
rect 865 3865 885 3885
rect 865 3815 885 3835
rect 865 3765 885 3785
rect 865 3715 885 3735
rect 1015 4165 1035 4185
rect 1015 4115 1035 4135
rect 1015 4065 1035 4085
rect 1015 4015 1035 4035
rect 1015 3965 1035 3985
rect 1015 3915 1035 3935
rect 1015 3865 1035 3885
rect 1015 3815 1035 3835
rect 1015 3765 1035 3785
rect 1015 3715 1035 3735
rect 1165 4165 1185 4185
rect 1165 4115 1185 4135
rect 1165 4065 1185 4085
rect 1165 4015 1185 4035
rect 1165 3965 1185 3985
rect 1165 3915 1185 3935
rect 1165 3865 1185 3885
rect 1165 3815 1185 3835
rect 1165 3765 1185 3785
rect 1165 3715 1185 3735
rect 1315 4165 1335 4185
rect 1315 4115 1335 4135
rect 1315 4065 1335 4085
rect 1315 4015 1335 4035
rect 1315 3965 1335 3985
rect 1315 3915 1335 3935
rect 1315 3865 1335 3885
rect 1315 3815 1335 3835
rect 1315 3765 1335 3785
rect 1315 3715 1335 3735
rect 1465 4165 1485 4185
rect 1465 4115 1485 4135
rect 1465 4065 1485 4085
rect 1465 4015 1485 4035
rect 1465 3965 1485 3985
rect 1465 3915 1485 3935
rect 1465 3865 1485 3885
rect 1465 3815 1485 3835
rect 1465 3765 1485 3785
rect 1465 3715 1485 3735
rect 1615 4165 1635 4185
rect 1615 4115 1635 4135
rect 1615 4065 1635 4085
rect 1615 4015 1635 4035
rect 1615 3965 1635 3985
rect 1615 3915 1635 3935
rect 1615 3865 1635 3885
rect 1615 3815 1635 3835
rect 1615 3765 1635 3785
rect 1615 3715 1635 3735
rect 1765 4165 1785 4185
rect 1765 4115 1785 4135
rect 1765 4065 1785 4085
rect 1765 4015 1785 4035
rect 1765 3965 1785 3985
rect 1765 3915 1785 3935
rect 1765 3865 1785 3885
rect 1765 3815 1785 3835
rect 1765 3765 1785 3785
rect 1765 3715 1785 3735
rect 1915 4165 1935 4185
rect 1915 4115 1935 4135
rect 1915 4065 1935 4085
rect 1915 4015 1935 4035
rect 1915 3965 1935 3985
rect 1915 3915 1935 3935
rect 1915 3865 1935 3885
rect 1915 3815 1935 3835
rect 1915 3765 1935 3785
rect 1915 3715 1935 3735
rect 2065 4165 2085 4185
rect 2065 4115 2085 4135
rect 2065 4065 2085 4085
rect 2065 4015 2085 4035
rect 2065 3965 2085 3985
rect 2065 3915 2085 3935
rect 2065 3865 2085 3885
rect 2065 3815 2085 3835
rect 2065 3765 2085 3785
rect 2065 3715 2085 3735
rect 2215 4165 2235 4185
rect 2215 4115 2235 4135
rect 2215 4065 2235 4085
rect 2215 4015 2235 4035
rect 2215 3965 2235 3985
rect 2215 3915 2235 3935
rect 2215 3865 2235 3885
rect 2215 3815 2235 3835
rect 2215 3765 2235 3785
rect 2215 3715 2235 3735
rect 2365 4165 2385 4185
rect 2365 4115 2385 4135
rect 2365 4065 2385 4085
rect 2365 4015 2385 4035
rect 2365 3965 2385 3985
rect 2365 3915 2385 3935
rect 2365 3865 2385 3885
rect 2365 3815 2385 3835
rect 2365 3765 2385 3785
rect 2365 3715 2385 3735
rect 2515 4165 2535 4185
rect 2515 4115 2535 4135
rect 2515 4065 2535 4085
rect 2515 4015 2535 4035
rect 2515 3965 2535 3985
rect 2515 3915 2535 3935
rect 2515 3865 2535 3885
rect 2515 3815 2535 3835
rect 2515 3765 2535 3785
rect 2515 3715 2535 3735
rect 2665 4165 2685 4185
rect 2665 4115 2685 4135
rect 2665 4065 2685 4085
rect 2665 4015 2685 4035
rect 2665 3965 2685 3985
rect 2665 3915 2685 3935
rect 2665 3865 2685 3885
rect 2665 3815 2685 3835
rect 2665 3765 2685 3785
rect 2665 3715 2685 3735
rect 2815 4165 2835 4185
rect 2815 4115 2835 4135
rect 2815 4065 2835 4085
rect 2815 4015 2835 4035
rect 2815 3965 2835 3985
rect 2815 3915 2835 3935
rect 2815 3865 2835 3885
rect 2815 3815 2835 3835
rect 2815 3765 2835 3785
rect 2815 3715 2835 3735
rect 2965 4165 2985 4185
rect 2965 4115 2985 4135
rect 2965 4065 2985 4085
rect 2965 4015 2985 4035
rect 2965 3965 2985 3985
rect 2965 3915 2985 3935
rect 2965 3865 2985 3885
rect 2965 3815 2985 3835
rect 2965 3765 2985 3785
rect 2965 3715 2985 3735
rect 3115 4165 3135 4185
rect 3115 4115 3135 4135
rect 3115 4065 3135 4085
rect 3115 4015 3135 4035
rect 3115 3965 3135 3985
rect 3115 3915 3135 3935
rect 3115 3865 3135 3885
rect 3115 3815 3135 3835
rect 3115 3765 3135 3785
rect 3115 3715 3135 3735
rect 3265 4165 3285 4185
rect 3265 4115 3285 4135
rect 3265 4065 3285 4085
rect 3265 4015 3285 4035
rect 3265 3965 3285 3985
rect 3265 3915 3285 3935
rect 3265 3865 3285 3885
rect 3265 3815 3285 3835
rect 3265 3765 3285 3785
rect 3265 3715 3285 3735
rect 3415 4165 3435 4185
rect 3415 4115 3435 4135
rect 3415 4065 3435 4085
rect 3415 4015 3435 4035
rect 3415 3965 3435 3985
rect 3415 3915 3435 3935
rect 3415 3865 3435 3885
rect 3415 3815 3435 3835
rect 3415 3765 3435 3785
rect 3415 3715 3435 3735
rect 3565 4165 3585 4185
rect 3565 4115 3585 4135
rect 3565 4065 3585 4085
rect 3565 4015 3585 4035
rect 3565 3965 3585 3985
rect 3565 3915 3585 3935
rect 3565 3865 3585 3885
rect 3565 3815 3585 3835
rect 3565 3765 3585 3785
rect 3565 3715 3585 3735
rect 4165 4165 4185 4185
rect 4165 4115 4185 4135
rect 4165 4065 4185 4085
rect 4165 4015 4185 4035
rect 4165 3965 4185 3985
rect 4165 3915 4185 3935
rect 4165 3865 4185 3885
rect 4165 3815 4185 3835
rect 4165 3765 4185 3785
rect 4165 3715 4185 3735
rect 4765 4165 4785 4185
rect 4765 4115 4785 4135
rect 4765 4065 4785 4085
rect 4765 4015 4785 4035
rect 4765 3965 4785 3985
rect 4765 3915 4785 3935
rect 4765 3865 4785 3885
rect 4765 3815 4785 3835
rect 4765 3765 4785 3785
rect 4765 3715 4785 3735
rect 4915 4165 4935 4185
rect 4915 4115 4935 4135
rect 4915 4065 4935 4085
rect 4915 4015 4935 4035
rect 4915 3965 4935 3985
rect 4915 3915 4935 3935
rect 4915 3865 4935 3885
rect 4915 3815 4935 3835
rect 4915 3765 4935 3785
rect 4915 3715 4935 3735
rect 5065 4165 5085 4185
rect 5065 4115 5085 4135
rect 5065 4065 5085 4085
rect 5065 4015 5085 4035
rect 5065 3965 5085 3985
rect 5065 3915 5085 3935
rect 5065 3865 5085 3885
rect 5065 3815 5085 3835
rect 5065 3765 5085 3785
rect 5065 3715 5085 3735
rect 5215 4165 5235 4185
rect 5215 4115 5235 4135
rect 5215 4065 5235 4085
rect 5215 4015 5235 4035
rect 5215 3965 5235 3985
rect 5215 3915 5235 3935
rect 5215 3865 5235 3885
rect 5215 3815 5235 3835
rect 5215 3765 5235 3785
rect 5215 3715 5235 3735
rect 5365 4165 5385 4185
rect 5365 4115 5385 4135
rect 5365 4065 5385 4085
rect 5365 4015 5385 4035
rect 5365 3965 5385 3985
rect 5365 3915 5385 3935
rect 5365 3865 5385 3885
rect 5365 3815 5385 3835
rect 5365 3765 5385 3785
rect 5365 3715 5385 3735
rect 5515 4165 5535 4185
rect 5515 4115 5535 4135
rect 5515 4065 5535 4085
rect 5515 4015 5535 4035
rect 5515 3965 5535 3985
rect 5515 3915 5535 3935
rect 5515 3865 5535 3885
rect 5515 3815 5535 3835
rect 5515 3765 5535 3785
rect 5515 3715 5535 3735
rect 5665 4165 5685 4185
rect 5665 4115 5685 4135
rect 5665 4065 5685 4085
rect 5665 4015 5685 4035
rect 5665 3965 5685 3985
rect 5665 3915 5685 3935
rect 5665 3865 5685 3885
rect 5665 3815 5685 3835
rect 5665 3765 5685 3785
rect 5665 3715 5685 3735
rect 5815 4165 5835 4185
rect 5815 4115 5835 4135
rect 5815 4065 5835 4085
rect 5815 4015 5835 4035
rect 5815 3965 5835 3985
rect 5815 3915 5835 3935
rect 5815 3865 5835 3885
rect 5815 3815 5835 3835
rect 5815 3765 5835 3785
rect 5815 3715 5835 3735
rect 5965 4165 5985 4185
rect 5965 4115 5985 4135
rect 5965 4065 5985 4085
rect 5965 4015 5985 4035
rect 5965 3965 5985 3985
rect 5965 3915 5985 3935
rect 5965 3865 5985 3885
rect 5965 3815 5985 3835
rect 5965 3765 5985 3785
rect 5965 3715 5985 3735
rect 6115 4165 6135 4185
rect 6115 4115 6135 4135
rect 6115 4065 6135 4085
rect 6115 4015 6135 4035
rect 6115 3965 6135 3985
rect 6115 3915 6135 3935
rect 6115 3865 6135 3885
rect 6115 3815 6135 3835
rect 6115 3765 6135 3785
rect 6115 3715 6135 3735
rect 6265 4165 6285 4185
rect 6265 4115 6285 4135
rect 6265 4065 6285 4085
rect 6265 4015 6285 4035
rect 6265 3965 6285 3985
rect 6265 3915 6285 3935
rect 6265 3865 6285 3885
rect 6265 3815 6285 3835
rect 6265 3765 6285 3785
rect 6265 3715 6285 3735
rect 6415 4165 6435 4185
rect 6415 4115 6435 4135
rect 6415 4065 6435 4085
rect 6415 4015 6435 4035
rect 6415 3965 6435 3985
rect 6415 3915 6435 3935
rect 6415 3865 6435 3885
rect 6415 3815 6435 3835
rect 6415 3765 6435 3785
rect 6415 3715 6435 3735
rect 6565 4165 6585 4185
rect 6565 4115 6585 4135
rect 6565 4065 6585 4085
rect 6565 4015 6585 4035
rect 6565 3965 6585 3985
rect 6565 3915 6585 3935
rect 6565 3865 6585 3885
rect 6565 3815 6585 3835
rect 6565 3765 6585 3785
rect 6565 3715 6585 3735
rect 6715 4165 6735 4185
rect 6715 4115 6735 4135
rect 6715 4065 6735 4085
rect 6715 4015 6735 4035
rect 6715 3965 6735 3985
rect 6715 3915 6735 3935
rect 6715 3865 6735 3885
rect 6715 3815 6735 3835
rect 6715 3765 6735 3785
rect 6715 3715 6735 3735
rect 6865 4165 6885 4185
rect 6865 4115 6885 4135
rect 6865 4065 6885 4085
rect 6865 4015 6885 4035
rect 6865 3965 6885 3985
rect 6865 3915 6885 3935
rect 6865 3865 6885 3885
rect 6865 3815 6885 3835
rect 6865 3765 6885 3785
rect 6865 3715 6885 3735
rect 7015 4165 7035 4185
rect 7015 4115 7035 4135
rect 7015 4065 7035 4085
rect 7015 4015 7035 4035
rect 7015 3965 7035 3985
rect 7015 3915 7035 3935
rect 7015 3865 7035 3885
rect 7015 3815 7035 3835
rect 7015 3765 7035 3785
rect 7015 3715 7035 3735
rect 7165 4165 7185 4185
rect 7165 4115 7185 4135
rect 7165 4065 7185 4085
rect 7165 4015 7185 4035
rect 7165 3965 7185 3985
rect 7165 3915 7185 3935
rect 7165 3865 7185 3885
rect 7165 3815 7185 3835
rect 7165 3765 7185 3785
rect 7165 3715 7185 3735
rect 7315 4165 7335 4185
rect 7315 4115 7335 4135
rect 7315 4065 7335 4085
rect 7315 4015 7335 4035
rect 7315 3965 7335 3985
rect 7315 3915 7335 3935
rect 7315 3865 7335 3885
rect 7315 3815 7335 3835
rect 7315 3765 7335 3785
rect 7315 3715 7335 3735
rect 7465 4165 7485 4185
rect 7465 4115 7485 4135
rect 7465 4065 7485 4085
rect 7465 4015 7485 4035
rect 7465 3965 7485 3985
rect 7465 3915 7485 3935
rect 7465 3865 7485 3885
rect 7465 3815 7485 3835
rect 7465 3765 7485 3785
rect 7465 3715 7485 3735
rect 7615 4165 7635 4185
rect 7615 4115 7635 4135
rect 7615 4065 7635 4085
rect 7615 4015 7635 4035
rect 7615 3965 7635 3985
rect 7615 3915 7635 3935
rect 7615 3865 7635 3885
rect 7615 3815 7635 3835
rect 7615 3765 7635 3785
rect 7615 3715 7635 3735
rect 7765 4165 7785 4185
rect 7765 4115 7785 4135
rect 7765 4065 7785 4085
rect 7765 4015 7785 4035
rect 7765 3965 7785 3985
rect 7765 3915 7785 3935
rect 7765 3865 7785 3885
rect 7765 3815 7785 3835
rect 7765 3765 7785 3785
rect 7765 3715 7785 3735
rect 8365 4165 8385 4185
rect 8365 4115 8385 4135
rect 8365 4065 8385 4085
rect 8365 4015 8385 4035
rect 8365 3965 8385 3985
rect 8365 3915 8385 3935
rect 8365 3865 8385 3885
rect 8365 3815 8385 3835
rect 8365 3765 8385 3785
rect 8365 3715 8385 3735
rect 8515 4165 8535 4185
rect 8515 4115 8535 4135
rect 8515 4065 8535 4085
rect 8515 4015 8535 4035
rect 8515 3965 8535 3985
rect 8515 3915 8535 3935
rect 8515 3865 8535 3885
rect 8515 3815 8535 3835
rect 8515 3765 8535 3785
rect 8515 3715 8535 3735
rect 8665 4165 8685 4185
rect 8665 4115 8685 4135
rect 8665 4065 8685 4085
rect 8665 4015 8685 4035
rect 8665 3965 8685 3985
rect 8665 3915 8685 3935
rect 8665 3865 8685 3885
rect 8665 3815 8685 3835
rect 8665 3765 8685 3785
rect 8665 3715 8685 3735
rect 8815 4165 8835 4185
rect 8815 4115 8835 4135
rect 8815 4065 8835 4085
rect 8815 4015 8835 4035
rect 8815 3965 8835 3985
rect 8815 3915 8835 3935
rect 8815 3865 8835 3885
rect 8815 3815 8835 3835
rect 8815 3765 8835 3785
rect 8815 3715 8835 3735
rect 8965 4165 8985 4185
rect 8965 4115 8985 4135
rect 8965 4065 8985 4085
rect 8965 4015 8985 4035
rect 8965 3965 8985 3985
rect 8965 3915 8985 3935
rect 8965 3865 8985 3885
rect 8965 3815 8985 3835
rect 8965 3765 8985 3785
rect 8965 3715 8985 3735
rect 9115 4165 9135 4185
rect 9115 4115 9135 4135
rect 9115 4065 9135 4085
rect 9115 4015 9135 4035
rect 9115 3965 9135 3985
rect 9115 3915 9135 3935
rect 9115 3865 9135 3885
rect 9115 3815 9135 3835
rect 9115 3765 9135 3785
rect 9115 3715 9135 3735
rect 9265 4165 9285 4185
rect 9265 4115 9285 4135
rect 9265 4065 9285 4085
rect 9265 4015 9285 4035
rect 9265 3965 9285 3985
rect 9265 3915 9285 3935
rect 9265 3865 9285 3885
rect 9265 3815 9285 3835
rect 9265 3765 9285 3785
rect 9265 3715 9285 3735
rect 9415 4165 9435 4185
rect 9415 4115 9435 4135
rect 9415 4065 9435 4085
rect 9415 4015 9435 4035
rect 9415 3965 9435 3985
rect 9415 3915 9435 3935
rect 9415 3865 9435 3885
rect 9415 3815 9435 3835
rect 9415 3765 9435 3785
rect 9415 3715 9435 3735
rect 9565 4165 9585 4185
rect 9565 4115 9585 4135
rect 9565 4065 9585 4085
rect 9565 4015 9585 4035
rect 9565 3965 9585 3985
rect 9565 3915 9585 3935
rect 9565 3865 9585 3885
rect 9565 3815 9585 3835
rect 9565 3765 9585 3785
rect 9565 3715 9585 3735
rect 9715 4165 9735 4185
rect 9715 4115 9735 4135
rect 9715 4065 9735 4085
rect 9715 4015 9735 4035
rect 9715 3965 9735 3985
rect 9715 3915 9735 3935
rect 9715 3865 9735 3885
rect 9715 3815 9735 3835
rect 9715 3765 9735 3785
rect 9715 3715 9735 3735
rect 9865 4165 9885 4185
rect 9865 4115 9885 4135
rect 9865 4065 9885 4085
rect 9865 4015 9885 4035
rect 9865 3965 9885 3985
rect 9865 3915 9885 3935
rect 9865 3865 9885 3885
rect 9865 3815 9885 3835
rect 9865 3765 9885 3785
rect 9865 3715 9885 3735
rect 10015 4165 10035 4185
rect 10015 4115 10035 4135
rect 10015 4065 10035 4085
rect 10015 4015 10035 4035
rect 10015 3965 10035 3985
rect 10015 3915 10035 3935
rect 10015 3865 10035 3885
rect 10015 3815 10035 3835
rect 10015 3765 10035 3785
rect 10015 3715 10035 3735
rect 10165 4165 10185 4185
rect 10165 4115 10185 4135
rect 10165 4065 10185 4085
rect 10165 4015 10185 4035
rect 10165 3965 10185 3985
rect 10165 3915 10185 3935
rect 10165 3865 10185 3885
rect 10165 3815 10185 3835
rect 10165 3765 10185 3785
rect 10165 3715 10185 3735
rect 10315 4165 10335 4185
rect 10315 4115 10335 4135
rect 10315 4065 10335 4085
rect 10315 4015 10335 4035
rect 10315 3965 10335 3985
rect 10315 3915 10335 3935
rect 10315 3865 10335 3885
rect 10315 3815 10335 3835
rect 10315 3765 10335 3785
rect 10315 3715 10335 3735
rect 10465 4165 10485 4185
rect 10465 4115 10485 4135
rect 10465 4065 10485 4085
rect 10465 4015 10485 4035
rect 10465 3965 10485 3985
rect 10465 3915 10485 3935
rect 10465 3865 10485 3885
rect 10465 3815 10485 3835
rect 10465 3765 10485 3785
rect 10465 3715 10485 3735
rect 10615 4165 10635 4185
rect 10615 4115 10635 4135
rect 10615 4065 10635 4085
rect 10615 4015 10635 4035
rect 10615 3965 10635 3985
rect 10615 3915 10635 3935
rect 10615 3865 10635 3885
rect 10615 3815 10635 3835
rect 10615 3765 10635 3785
rect 10615 3715 10635 3735
rect 10765 4165 10785 4185
rect 10765 4115 10785 4135
rect 10765 4065 10785 4085
rect 10765 4015 10785 4035
rect 10765 3965 10785 3985
rect 10765 3915 10785 3935
rect 10765 3865 10785 3885
rect 10765 3815 10785 3835
rect 10765 3765 10785 3785
rect 10765 3715 10785 3735
rect 11365 4165 11385 4185
rect 11365 4115 11385 4135
rect 11365 4065 11385 4085
rect 11365 4015 11385 4035
rect 11365 3965 11385 3985
rect 11365 3915 11385 3935
rect 11365 3865 11385 3885
rect 11365 3815 11385 3835
rect 11365 3765 11385 3785
rect 11365 3715 11385 3735
rect 11965 4165 11985 4185
rect 11965 4115 11985 4135
rect 11965 4065 11985 4085
rect 11965 4015 11985 4035
rect 11965 3965 11985 3985
rect 11965 3915 11985 3935
rect 11965 3865 11985 3885
rect 11965 3815 11985 3835
rect 11965 3765 11985 3785
rect 11965 3715 11985 3735
rect 12565 4165 12585 4185
rect 12565 4115 12585 4135
rect 12565 4065 12585 4085
rect 12565 4015 12585 4035
rect 12565 3965 12585 3985
rect 12565 3915 12585 3935
rect 12565 3865 12585 3885
rect 12565 3815 12585 3835
rect 12565 3765 12585 3785
rect 12565 3715 12585 3735
rect 13165 4165 13185 4185
rect 13165 4115 13185 4135
rect 13165 4065 13185 4085
rect 13165 4015 13185 4035
rect 13165 3965 13185 3985
rect 13165 3915 13185 3935
rect 13165 3865 13185 3885
rect 13165 3815 13185 3835
rect 13165 3765 13185 3785
rect 13165 3715 13185 3735
rect 13765 4165 13785 4185
rect 13765 4115 13785 4135
rect 13765 4065 13785 4085
rect 13765 4015 13785 4035
rect 13765 3965 13785 3985
rect 13765 3915 13785 3935
rect 13765 3865 13785 3885
rect 13765 3815 13785 3835
rect 13765 3765 13785 3785
rect 13765 3715 13785 3735
rect 14365 4165 14385 4185
rect 14365 4115 14385 4135
rect 14365 4065 14385 4085
rect 14365 4015 14385 4035
rect 14365 3965 14385 3985
rect 14365 3915 14385 3935
rect 14365 3865 14385 3885
rect 14365 3815 14385 3835
rect 14365 3765 14385 3785
rect 14365 3715 14385 3735
rect 14965 4165 14985 4185
rect 14965 4115 14985 4135
rect 14965 4065 14985 4085
rect 14965 4015 14985 4035
rect 14965 3965 14985 3985
rect 14965 3915 14985 3935
rect 14965 3865 14985 3885
rect 14965 3815 14985 3835
rect 14965 3765 14985 3785
rect 14965 3715 14985 3735
rect 15565 4165 15585 4185
rect 15565 4115 15585 4135
rect 15565 4065 15585 4085
rect 15565 4015 15585 4035
rect 15565 3965 15585 3985
rect 15565 3915 15585 3935
rect 15565 3865 15585 3885
rect 15565 3815 15585 3835
rect 15565 3765 15585 3785
rect 15565 3715 15585 3735
rect 16165 4165 16185 4185
rect 16165 4115 16185 4135
rect 16165 4065 16185 4085
rect 16165 4015 16185 4035
rect 16165 3965 16185 3985
rect 16165 3915 16185 3935
rect 16165 3865 16185 3885
rect 16165 3815 16185 3835
rect 16165 3765 16185 3785
rect 16165 3715 16185 3735
rect 16315 4165 16335 4185
rect 16315 4115 16335 4135
rect 16315 4065 16335 4085
rect 16315 4015 16335 4035
rect 16315 3965 16335 3985
rect 16315 3915 16335 3935
rect 16315 3865 16335 3885
rect 16315 3815 16335 3835
rect 16315 3765 16335 3785
rect 16315 3715 16335 3735
rect 16465 4165 16485 4185
rect 16465 4115 16485 4135
rect 16465 4065 16485 4085
rect 16465 4015 16485 4035
rect 16465 3965 16485 3985
rect 16465 3915 16485 3935
rect 16465 3865 16485 3885
rect 16465 3815 16485 3835
rect 16465 3765 16485 3785
rect 16465 3715 16485 3735
rect 16615 4165 16635 4185
rect 16615 4115 16635 4135
rect 16615 4065 16635 4085
rect 16615 4015 16635 4035
rect 16615 3965 16635 3985
rect 16615 3915 16635 3935
rect 16615 3865 16635 3885
rect 16615 3815 16635 3835
rect 16615 3765 16635 3785
rect 16615 3715 16635 3735
rect 16765 4165 16785 4185
rect 16765 4115 16785 4135
rect 16765 4065 16785 4085
rect 16765 4015 16785 4035
rect 16765 3965 16785 3985
rect 16765 3915 16785 3935
rect 16765 3865 16785 3885
rect 16765 3815 16785 3835
rect 16765 3765 16785 3785
rect 16765 3715 16785 3735
rect 16915 4165 16935 4185
rect 16915 4115 16935 4135
rect 16915 4065 16935 4085
rect 16915 4015 16935 4035
rect 16915 3965 16935 3985
rect 16915 3915 16935 3935
rect 16915 3865 16935 3885
rect 16915 3815 16935 3835
rect 16915 3765 16935 3785
rect 16915 3715 16935 3735
rect 17065 4165 17085 4185
rect 17065 4115 17085 4135
rect 17065 4065 17085 4085
rect 17065 4015 17085 4035
rect 17065 3965 17085 3985
rect 17065 3915 17085 3935
rect 17065 3865 17085 3885
rect 17065 3815 17085 3835
rect 17065 3765 17085 3785
rect 17065 3715 17085 3735
rect 17215 4165 17235 4185
rect 17215 4115 17235 4135
rect 17215 4065 17235 4085
rect 17215 4015 17235 4035
rect 17215 3965 17235 3985
rect 17215 3915 17235 3935
rect 17215 3865 17235 3885
rect 17215 3815 17235 3835
rect 17215 3765 17235 3785
rect 17215 3715 17235 3735
rect 17365 4165 17385 4185
rect 17365 4115 17385 4135
rect 17365 4065 17385 4085
rect 17365 4015 17385 4035
rect 17365 3965 17385 3985
rect 17365 3915 17385 3935
rect 17365 3865 17385 3885
rect 17365 3815 17385 3835
rect 17365 3765 17385 3785
rect 17365 3715 17385 3735
rect 17965 4165 17985 4185
rect 17965 4115 17985 4135
rect 17965 4065 17985 4085
rect 17965 4015 17985 4035
rect 17965 3965 17985 3985
rect 17965 3915 17985 3935
rect 17965 3865 17985 3885
rect 17965 3815 17985 3835
rect 17965 3765 17985 3785
rect 17965 3715 17985 3735
rect 18565 4165 18585 4185
rect 18565 4115 18585 4135
rect 18565 4065 18585 4085
rect 18565 4015 18585 4035
rect 18565 3965 18585 3985
rect 18565 3915 18585 3935
rect 18565 3865 18585 3885
rect 18565 3815 18585 3835
rect 18565 3765 18585 3785
rect 18565 3715 18585 3735
rect 18715 4165 18735 4185
rect 18715 4115 18735 4135
rect 18715 4065 18735 4085
rect 18715 4015 18735 4035
rect 18715 3965 18735 3985
rect 18715 3915 18735 3935
rect 18715 3865 18735 3885
rect 18715 3815 18735 3835
rect 18715 3765 18735 3785
rect 18715 3715 18735 3735
rect 18865 4165 18885 4185
rect 18865 4115 18885 4135
rect 18865 4065 18885 4085
rect 18865 4015 18885 4035
rect 18865 3965 18885 3985
rect 18865 3915 18885 3935
rect 18865 3865 18885 3885
rect 18865 3815 18885 3835
rect 18865 3765 18885 3785
rect 18865 3715 18885 3735
rect 19015 4165 19035 4185
rect 19015 4115 19035 4135
rect 19015 4065 19035 4085
rect 19015 4015 19035 4035
rect 19015 3965 19035 3985
rect 19015 3915 19035 3935
rect 19015 3865 19035 3885
rect 19015 3815 19035 3835
rect 19015 3765 19035 3785
rect 19015 3715 19035 3735
rect 19165 4165 19185 4185
rect 19165 4115 19185 4135
rect 19165 4065 19185 4085
rect 19165 4015 19185 4035
rect 19165 3965 19185 3985
rect 19165 3915 19185 3935
rect 19165 3865 19185 3885
rect 19165 3815 19185 3835
rect 19165 3765 19185 3785
rect 19165 3715 19185 3735
rect 19315 4165 19335 4185
rect 19315 4115 19335 4135
rect 19315 4065 19335 4085
rect 19315 4015 19335 4035
rect 19315 3965 19335 3985
rect 19315 3915 19335 3935
rect 19315 3865 19335 3885
rect 19315 3815 19335 3835
rect 19315 3765 19335 3785
rect 19315 3715 19335 3735
rect 19465 4165 19485 4185
rect 19465 4115 19485 4135
rect 19465 4065 19485 4085
rect 19465 4015 19485 4035
rect 19465 3965 19485 3985
rect 19465 3915 19485 3935
rect 19465 3865 19485 3885
rect 19465 3815 19485 3835
rect 19465 3765 19485 3785
rect 19465 3715 19485 3735
rect 19615 4165 19635 4185
rect 19615 4115 19635 4135
rect 19615 4065 19635 4085
rect 19615 4015 19635 4035
rect 19615 3965 19635 3985
rect 19615 3915 19635 3935
rect 19615 3865 19635 3885
rect 19615 3815 19635 3835
rect 19615 3765 19635 3785
rect 19615 3715 19635 3735
rect 19765 4165 19785 4185
rect 19765 4115 19785 4135
rect 19765 4065 19785 4085
rect 19765 4015 19785 4035
rect 19765 3965 19785 3985
rect 19765 3915 19785 3935
rect 19765 3865 19785 3885
rect 19765 3815 19785 3835
rect 19765 3765 19785 3785
rect 19765 3715 19785 3735
rect 20365 4165 20385 4185
rect 20365 4115 20385 4135
rect 20365 4065 20385 4085
rect 20365 4015 20385 4035
rect 20365 3965 20385 3985
rect 20365 3915 20385 3935
rect 20365 3865 20385 3885
rect 20365 3815 20385 3835
rect 20365 3765 20385 3785
rect 20365 3715 20385 3735
rect 20965 4165 20985 4185
rect 20965 4115 20985 4135
rect 20965 4065 20985 4085
rect 20965 4015 20985 4035
rect 20965 3965 20985 3985
rect 20965 3915 20985 3935
rect 20965 3865 20985 3885
rect 20965 3815 20985 3835
rect 20965 3765 20985 3785
rect 20965 3715 20985 3735
rect 21415 4165 21435 4185
rect 21415 4115 21435 4135
rect 21415 4065 21435 4085
rect 21415 4015 21435 4035
rect 21415 3965 21435 3985
rect 21415 3915 21435 3935
rect 21415 3865 21435 3885
rect 21415 3815 21435 3835
rect 21415 3765 21435 3785
rect 21415 3715 21435 3735
rect 21865 4165 21885 4185
rect 21865 4115 21885 4135
rect 21865 4065 21885 4085
rect 21865 4015 21885 4035
rect 21865 3965 21885 3985
rect 21865 3915 21885 3935
rect 21865 3865 21885 3885
rect 21865 3815 21885 3835
rect 21865 3765 21885 3785
rect 21865 3715 21885 3735
rect 22465 4165 22485 4185
rect 22465 4115 22485 4135
rect 22465 4065 22485 4085
rect 22465 4015 22485 4035
rect 22465 3965 22485 3985
rect 22465 3915 22485 3935
rect 22465 3865 22485 3885
rect 22465 3815 22485 3835
rect 22465 3765 22485 3785
rect 22465 3715 22485 3735
rect 23065 4165 23085 4185
rect 23065 4115 23085 4135
rect 23065 4065 23085 4085
rect 23065 4015 23085 4035
rect 23065 3965 23085 3985
rect 23065 3915 23085 3935
rect 23065 3865 23085 3885
rect 23065 3815 23085 3835
rect 23065 3765 23085 3785
rect 23065 3715 23085 3735
rect 23515 4165 23535 4185
rect 23515 4115 23535 4135
rect 23515 4065 23535 4085
rect 23515 4015 23535 4035
rect 23515 3965 23535 3985
rect 23515 3915 23535 3935
rect 23515 3865 23535 3885
rect 23515 3815 23535 3835
rect 23515 3765 23535 3785
rect 23515 3715 23535 3735
rect 23965 4165 23985 4185
rect 23965 4115 23985 4135
rect 23965 4065 23985 4085
rect 23965 4015 23985 4035
rect 23965 3965 23985 3985
rect 23965 3915 23985 3935
rect 23965 3865 23985 3885
rect 23965 3815 23985 3835
rect 23965 3765 23985 3785
rect 23965 3715 23985 3735
rect 24565 4165 24585 4185
rect 24565 4115 24585 4135
rect 24565 4065 24585 4085
rect 24565 4015 24585 4035
rect 24565 3965 24585 3985
rect 24565 3915 24585 3935
rect 24565 3865 24585 3885
rect 24565 3815 24585 3835
rect 24565 3765 24585 3785
rect 24565 3715 24585 3735
rect 25165 4165 25185 4185
rect 25165 4115 25185 4135
rect 25165 4065 25185 4085
rect 25165 4015 25185 4035
rect 25165 3965 25185 3985
rect 25165 3915 25185 3935
rect 25165 3865 25185 3885
rect 25165 3815 25185 3835
rect 25165 3765 25185 3785
rect 25165 3715 25185 3735
rect 25615 4165 25635 4185
rect 25615 4115 25635 4135
rect 25615 4065 25635 4085
rect 25615 4015 25635 4035
rect 25615 3965 25635 3985
rect 25615 3915 25635 3935
rect 25615 3865 25635 3885
rect 25615 3815 25635 3835
rect 25615 3765 25635 3785
rect 25615 3715 25635 3735
rect 26065 4165 26085 4185
rect 26065 4115 26085 4135
rect 26065 4065 26085 4085
rect 26065 4015 26085 4035
rect 26065 3965 26085 3985
rect 26065 3915 26085 3935
rect 26065 3865 26085 3885
rect 26065 3815 26085 3835
rect 26065 3765 26085 3785
rect 26065 3715 26085 3735
rect 26665 4165 26685 4185
rect 26665 4115 26685 4135
rect 26665 4065 26685 4085
rect 26665 4015 26685 4035
rect 26665 3965 26685 3985
rect 26665 3915 26685 3935
rect 26665 3865 26685 3885
rect 26665 3815 26685 3835
rect 26665 3765 26685 3785
rect 26665 3715 26685 3735
rect 27265 4165 27285 4185
rect 27265 4115 27285 4135
rect 27265 4065 27285 4085
rect 27265 4015 27285 4035
rect 27265 3965 27285 3985
rect 27265 3915 27285 3935
rect 27265 3865 27285 3885
rect 27265 3815 27285 3835
rect 27265 3765 27285 3785
rect 27265 3715 27285 3735
rect 27715 4165 27735 4185
rect 27715 4115 27735 4135
rect 27715 4065 27735 4085
rect 27715 4015 27735 4035
rect 27715 3965 27735 3985
rect 27715 3915 27735 3935
rect 27715 3865 27735 3885
rect 27715 3815 27735 3835
rect 27715 3765 27735 3785
rect 27715 3715 27735 3735
rect 28165 4165 28185 4185
rect 28165 4115 28185 4135
rect 28165 4065 28185 4085
rect 28165 4015 28185 4035
rect 28165 3965 28185 3985
rect 28165 3915 28185 3935
rect 28165 3865 28185 3885
rect 28165 3815 28185 3835
rect 28165 3765 28185 3785
rect 28165 3715 28185 3735
rect 28765 4165 28785 4185
rect 28765 4115 28785 4135
rect 28765 4065 28785 4085
rect 28765 4015 28785 4035
rect 28765 3965 28785 3985
rect 28765 3915 28785 3935
rect 28765 3865 28785 3885
rect 28765 3815 28785 3835
rect 28765 3765 28785 3785
rect 28765 3715 28785 3735
rect 29365 4165 29385 4185
rect 29365 4115 29385 4135
rect 29365 4065 29385 4085
rect 29365 4015 29385 4035
rect 29365 3965 29385 3985
rect 29365 3915 29385 3935
rect 29365 3865 29385 3885
rect 29365 3815 29385 3835
rect 29365 3765 29385 3785
rect 29365 3715 29385 3735
rect 29515 4165 29535 4185
rect 29515 4115 29535 4135
rect 29515 4065 29535 4085
rect 29515 4015 29535 4035
rect 29515 3965 29535 3985
rect 29515 3915 29535 3935
rect 29515 3865 29535 3885
rect 29515 3815 29535 3835
rect 29515 3765 29535 3785
rect 29515 3715 29535 3735
rect 29665 4165 29685 4185
rect 29665 4115 29685 4135
rect 29665 4065 29685 4085
rect 29665 4015 29685 4035
rect 29665 3965 29685 3985
rect 29665 3915 29685 3935
rect 29665 3865 29685 3885
rect 29665 3815 29685 3835
rect 29665 3765 29685 3785
rect 29665 3715 29685 3735
rect 29815 4165 29835 4185
rect 29815 4115 29835 4135
rect 29815 4065 29835 4085
rect 29815 4015 29835 4035
rect 29815 3965 29835 3985
rect 29815 3915 29835 3935
rect 29815 3865 29835 3885
rect 29815 3815 29835 3835
rect 29815 3765 29835 3785
rect 29815 3715 29835 3735
rect 29965 4165 29985 4185
rect 29965 4115 29985 4135
rect 29965 4065 29985 4085
rect 29965 4015 29985 4035
rect 29965 3965 29985 3985
rect 29965 3915 29985 3935
rect 29965 3865 29985 3885
rect 29965 3815 29985 3835
rect 29965 3765 29985 3785
rect 29965 3715 29985 3735
rect 30115 4165 30135 4185
rect 30115 4115 30135 4135
rect 30115 4065 30135 4085
rect 30115 4015 30135 4035
rect 30115 3965 30135 3985
rect 30115 3915 30135 3935
rect 30115 3865 30135 3885
rect 30115 3815 30135 3835
rect 30115 3765 30135 3785
rect 30115 3715 30135 3735
rect 30265 4165 30285 4185
rect 30265 4115 30285 4135
rect 30265 4065 30285 4085
rect 30265 4015 30285 4035
rect 30265 3965 30285 3985
rect 30265 3915 30285 3935
rect 30265 3865 30285 3885
rect 30265 3815 30285 3835
rect 30265 3765 30285 3785
rect 30265 3715 30285 3735
rect 30415 4165 30435 4185
rect 30415 4115 30435 4135
rect 30415 4065 30435 4085
rect 30415 4015 30435 4035
rect 30415 3965 30435 3985
rect 30415 3915 30435 3935
rect 30415 3865 30435 3885
rect 30415 3815 30435 3835
rect 30415 3765 30435 3785
rect 30415 3715 30435 3735
rect 30565 4165 30585 4185
rect 30565 4115 30585 4135
rect 30565 4065 30585 4085
rect 30565 4015 30585 4035
rect 30565 3965 30585 3985
rect 30565 3915 30585 3935
rect 30565 3865 30585 3885
rect 30565 3815 30585 3835
rect 30565 3765 30585 3785
rect 30565 3715 30585 3735
rect 30715 4165 30735 4185
rect 30715 4115 30735 4135
rect 30715 4065 30735 4085
rect 30715 4015 30735 4035
rect 30715 3965 30735 3985
rect 30715 3915 30735 3935
rect 30715 3865 30735 3885
rect 30715 3815 30735 3835
rect 30715 3765 30735 3785
rect 30715 3715 30735 3735
rect 30865 4165 30885 4185
rect 30865 4115 30885 4135
rect 30865 4065 30885 4085
rect 30865 4015 30885 4035
rect 30865 3965 30885 3985
rect 30865 3915 30885 3935
rect 30865 3865 30885 3885
rect 30865 3815 30885 3835
rect 30865 3765 30885 3785
rect 30865 3715 30885 3735
rect 31015 4165 31035 4185
rect 31015 4115 31035 4135
rect 31015 4065 31035 4085
rect 31015 4015 31035 4035
rect 31015 3965 31035 3985
rect 31015 3915 31035 3935
rect 31015 3865 31035 3885
rect 31015 3815 31035 3835
rect 31015 3765 31035 3785
rect 31015 3715 31035 3735
rect 31165 4165 31185 4185
rect 31165 4115 31185 4135
rect 31165 4065 31185 4085
rect 31165 4015 31185 4035
rect 31165 3965 31185 3985
rect 31165 3915 31185 3935
rect 31165 3865 31185 3885
rect 31165 3815 31185 3835
rect 31165 3765 31185 3785
rect 31165 3715 31185 3735
rect 31315 4165 31335 4185
rect 31315 4115 31335 4135
rect 31315 4065 31335 4085
rect 31315 4015 31335 4035
rect 31315 3965 31335 3985
rect 31315 3915 31335 3935
rect 31315 3865 31335 3885
rect 31315 3815 31335 3835
rect 31315 3765 31335 3785
rect 31315 3715 31335 3735
rect 31465 4165 31485 4185
rect 31465 4115 31485 4135
rect 31465 4065 31485 4085
rect 31465 4015 31485 4035
rect 31465 3965 31485 3985
rect 31465 3915 31485 3935
rect 31465 3865 31485 3885
rect 31465 3815 31485 3835
rect 31465 3765 31485 3785
rect 31465 3715 31485 3735
rect 32065 4165 32085 4185
rect 32065 4115 32085 4135
rect 32065 4065 32085 4085
rect 32065 4015 32085 4035
rect 32065 3965 32085 3985
rect 32065 3915 32085 3935
rect 32065 3865 32085 3885
rect 32065 3815 32085 3835
rect 32065 3765 32085 3785
rect 32065 3715 32085 3735
rect -635 3515 -615 3535
rect -635 3465 -615 3485
rect -635 3415 -615 3435
rect -635 3365 -615 3385
rect -635 3315 -615 3335
rect -635 3265 -615 3285
rect -635 3215 -615 3235
rect -635 3165 -615 3185
rect -635 3115 -615 3135
rect -635 3065 -615 3085
rect -485 3515 -465 3535
rect -485 3465 -465 3485
rect -485 3415 -465 3435
rect -485 3365 -465 3385
rect -485 3315 -465 3335
rect -485 3265 -465 3285
rect -485 3215 -465 3235
rect -485 3165 -465 3185
rect -485 3115 -465 3135
rect -485 3065 -465 3085
rect -335 3515 -315 3535
rect -335 3465 -315 3485
rect -335 3415 -315 3435
rect -335 3365 -315 3385
rect -335 3315 -315 3335
rect -335 3265 -315 3285
rect -335 3215 -315 3235
rect -335 3165 -315 3185
rect -335 3115 -315 3135
rect -335 3065 -315 3085
rect -185 3515 -165 3535
rect -185 3465 -165 3485
rect -185 3415 -165 3435
rect -185 3365 -165 3385
rect -185 3315 -165 3335
rect -185 3265 -165 3285
rect -185 3215 -165 3235
rect -185 3165 -165 3185
rect -185 3115 -165 3135
rect -185 3065 -165 3085
rect -35 3515 -15 3535
rect -35 3465 -15 3485
rect -35 3415 -15 3435
rect -35 3365 -15 3385
rect -35 3315 -15 3335
rect -35 3265 -15 3285
rect -35 3215 -15 3235
rect -35 3165 -15 3185
rect -35 3115 -15 3135
rect -35 3065 -15 3085
rect 565 3515 585 3535
rect 565 3465 585 3485
rect 565 3415 585 3435
rect 565 3365 585 3385
rect 565 3315 585 3335
rect 565 3265 585 3285
rect 565 3215 585 3235
rect 565 3165 585 3185
rect 565 3115 585 3135
rect 565 3065 585 3085
rect 715 3515 735 3535
rect 715 3465 735 3485
rect 715 3415 735 3435
rect 715 3365 735 3385
rect 715 3315 735 3335
rect 715 3265 735 3285
rect 715 3215 735 3235
rect 715 3165 735 3185
rect 715 3115 735 3135
rect 715 3065 735 3085
rect 865 3515 885 3535
rect 865 3465 885 3485
rect 865 3415 885 3435
rect 865 3365 885 3385
rect 865 3315 885 3335
rect 865 3265 885 3285
rect 865 3215 885 3235
rect 865 3165 885 3185
rect 865 3115 885 3135
rect 865 3065 885 3085
rect 1015 3515 1035 3535
rect 1015 3465 1035 3485
rect 1015 3415 1035 3435
rect 1015 3365 1035 3385
rect 1015 3315 1035 3335
rect 1015 3265 1035 3285
rect 1015 3215 1035 3235
rect 1015 3165 1035 3185
rect 1015 3115 1035 3135
rect 1015 3065 1035 3085
rect 1165 3515 1185 3535
rect 1165 3465 1185 3485
rect 1165 3415 1185 3435
rect 1165 3365 1185 3385
rect 1165 3315 1185 3335
rect 1165 3265 1185 3285
rect 1165 3215 1185 3235
rect 1165 3165 1185 3185
rect 1165 3115 1185 3135
rect 1165 3065 1185 3085
rect 1315 3515 1335 3535
rect 1315 3465 1335 3485
rect 1315 3415 1335 3435
rect 1315 3365 1335 3385
rect 1315 3315 1335 3335
rect 1315 3265 1335 3285
rect 1315 3215 1335 3235
rect 1315 3165 1335 3185
rect 1315 3115 1335 3135
rect 1315 3065 1335 3085
rect 1465 3515 1485 3535
rect 1465 3465 1485 3485
rect 1465 3415 1485 3435
rect 1465 3365 1485 3385
rect 1465 3315 1485 3335
rect 1465 3265 1485 3285
rect 1465 3215 1485 3235
rect 1465 3165 1485 3185
rect 1465 3115 1485 3135
rect 1465 3065 1485 3085
rect 1615 3515 1635 3535
rect 1615 3465 1635 3485
rect 1615 3415 1635 3435
rect 1615 3365 1635 3385
rect 1615 3315 1635 3335
rect 1615 3265 1635 3285
rect 1615 3215 1635 3235
rect 1615 3165 1635 3185
rect 1615 3115 1635 3135
rect 1615 3065 1635 3085
rect 1765 3515 1785 3535
rect 1765 3465 1785 3485
rect 1765 3415 1785 3435
rect 1765 3365 1785 3385
rect 1765 3315 1785 3335
rect 1765 3265 1785 3285
rect 1765 3215 1785 3235
rect 1765 3165 1785 3185
rect 1765 3115 1785 3135
rect 1765 3065 1785 3085
rect 1915 3515 1935 3535
rect 1915 3465 1935 3485
rect 1915 3415 1935 3435
rect 1915 3365 1935 3385
rect 1915 3315 1935 3335
rect 1915 3265 1935 3285
rect 1915 3215 1935 3235
rect 1915 3165 1935 3185
rect 1915 3115 1935 3135
rect 1915 3065 1935 3085
rect 2065 3515 2085 3535
rect 2065 3465 2085 3485
rect 2065 3415 2085 3435
rect 2065 3365 2085 3385
rect 2065 3315 2085 3335
rect 2065 3265 2085 3285
rect 2065 3215 2085 3235
rect 2065 3165 2085 3185
rect 2065 3115 2085 3135
rect 2065 3065 2085 3085
rect 2215 3515 2235 3535
rect 2215 3465 2235 3485
rect 2215 3415 2235 3435
rect 2215 3365 2235 3385
rect 2215 3315 2235 3335
rect 2215 3265 2235 3285
rect 2215 3215 2235 3235
rect 2215 3165 2235 3185
rect 2215 3115 2235 3135
rect 2215 3065 2235 3085
rect 2365 3515 2385 3535
rect 2365 3465 2385 3485
rect 2365 3415 2385 3435
rect 2365 3365 2385 3385
rect 2365 3315 2385 3335
rect 2365 3265 2385 3285
rect 2365 3215 2385 3235
rect 2365 3165 2385 3185
rect 2365 3115 2385 3135
rect 2365 3065 2385 3085
rect 2515 3515 2535 3535
rect 2515 3465 2535 3485
rect 2515 3415 2535 3435
rect 2515 3365 2535 3385
rect 2515 3315 2535 3335
rect 2515 3265 2535 3285
rect 2515 3215 2535 3235
rect 2515 3165 2535 3185
rect 2515 3115 2535 3135
rect 2515 3065 2535 3085
rect 2665 3515 2685 3535
rect 2665 3465 2685 3485
rect 2665 3415 2685 3435
rect 2665 3365 2685 3385
rect 2665 3315 2685 3335
rect 2665 3265 2685 3285
rect 2665 3215 2685 3235
rect 2665 3165 2685 3185
rect 2665 3115 2685 3135
rect 2665 3065 2685 3085
rect 2815 3515 2835 3535
rect 2815 3465 2835 3485
rect 2815 3415 2835 3435
rect 2815 3365 2835 3385
rect 2815 3315 2835 3335
rect 2815 3265 2835 3285
rect 2815 3215 2835 3235
rect 2815 3165 2835 3185
rect 2815 3115 2835 3135
rect 2815 3065 2835 3085
rect 2965 3515 2985 3535
rect 2965 3465 2985 3485
rect 2965 3415 2985 3435
rect 2965 3365 2985 3385
rect 2965 3315 2985 3335
rect 2965 3265 2985 3285
rect 2965 3215 2985 3235
rect 2965 3165 2985 3185
rect 2965 3115 2985 3135
rect 2965 3065 2985 3085
rect 3115 3515 3135 3535
rect 3115 3465 3135 3485
rect 3115 3415 3135 3435
rect 3115 3365 3135 3385
rect 3115 3315 3135 3335
rect 3115 3265 3135 3285
rect 3115 3215 3135 3235
rect 3115 3165 3135 3185
rect 3115 3115 3135 3135
rect 3115 3065 3135 3085
rect 3265 3515 3285 3535
rect 3265 3465 3285 3485
rect 3265 3415 3285 3435
rect 3265 3365 3285 3385
rect 3265 3315 3285 3335
rect 3265 3265 3285 3285
rect 3265 3215 3285 3235
rect 3265 3165 3285 3185
rect 3265 3115 3285 3135
rect 3265 3065 3285 3085
rect 3415 3515 3435 3535
rect 3415 3465 3435 3485
rect 3415 3415 3435 3435
rect 3415 3365 3435 3385
rect 3415 3315 3435 3335
rect 3415 3265 3435 3285
rect 3415 3215 3435 3235
rect 3415 3165 3435 3185
rect 3415 3115 3435 3135
rect 3415 3065 3435 3085
rect 3565 3515 3585 3535
rect 3565 3465 3585 3485
rect 3565 3415 3585 3435
rect 3565 3365 3585 3385
rect 3565 3315 3585 3335
rect 3565 3265 3585 3285
rect 3565 3215 3585 3235
rect 3565 3165 3585 3185
rect 3565 3115 3585 3135
rect 3565 3065 3585 3085
rect 4165 3515 4185 3535
rect 4165 3465 4185 3485
rect 4165 3415 4185 3435
rect 4165 3365 4185 3385
rect 4165 3315 4185 3335
rect 4165 3265 4185 3285
rect 4165 3215 4185 3235
rect 4165 3165 4185 3185
rect 4165 3115 4185 3135
rect 4165 3065 4185 3085
rect 4765 3515 4785 3535
rect 4765 3465 4785 3485
rect 4765 3415 4785 3435
rect 4765 3365 4785 3385
rect 4765 3315 4785 3335
rect 4765 3265 4785 3285
rect 4765 3215 4785 3235
rect 4765 3165 4785 3185
rect 4765 3115 4785 3135
rect 4765 3065 4785 3085
rect 4915 3515 4935 3535
rect 4915 3465 4935 3485
rect 4915 3415 4935 3435
rect 4915 3365 4935 3385
rect 4915 3315 4935 3335
rect 4915 3265 4935 3285
rect 4915 3215 4935 3235
rect 4915 3165 4935 3185
rect 4915 3115 4935 3135
rect 4915 3065 4935 3085
rect 5065 3515 5085 3535
rect 5065 3465 5085 3485
rect 5065 3415 5085 3435
rect 5065 3365 5085 3385
rect 5065 3315 5085 3335
rect 5065 3265 5085 3285
rect 5065 3215 5085 3235
rect 5065 3165 5085 3185
rect 5065 3115 5085 3135
rect 5065 3065 5085 3085
rect 5215 3515 5235 3535
rect 5215 3465 5235 3485
rect 5215 3415 5235 3435
rect 5215 3365 5235 3385
rect 5215 3315 5235 3335
rect 5215 3265 5235 3285
rect 5215 3215 5235 3235
rect 5215 3165 5235 3185
rect 5215 3115 5235 3135
rect 5215 3065 5235 3085
rect 5365 3515 5385 3535
rect 5365 3465 5385 3485
rect 5365 3415 5385 3435
rect 5365 3365 5385 3385
rect 5365 3315 5385 3335
rect 5365 3265 5385 3285
rect 5365 3215 5385 3235
rect 5365 3165 5385 3185
rect 5365 3115 5385 3135
rect 5365 3065 5385 3085
rect 5515 3515 5535 3535
rect 5515 3465 5535 3485
rect 5515 3415 5535 3435
rect 5515 3365 5535 3385
rect 5515 3315 5535 3335
rect 5515 3265 5535 3285
rect 5515 3215 5535 3235
rect 5515 3165 5535 3185
rect 5515 3115 5535 3135
rect 5515 3065 5535 3085
rect 5665 3515 5685 3535
rect 5665 3465 5685 3485
rect 5665 3415 5685 3435
rect 5665 3365 5685 3385
rect 5665 3315 5685 3335
rect 5665 3265 5685 3285
rect 5665 3215 5685 3235
rect 5665 3165 5685 3185
rect 5665 3115 5685 3135
rect 5665 3065 5685 3085
rect 5815 3515 5835 3535
rect 5815 3465 5835 3485
rect 5815 3415 5835 3435
rect 5815 3365 5835 3385
rect 5815 3315 5835 3335
rect 5815 3265 5835 3285
rect 5815 3215 5835 3235
rect 5815 3165 5835 3185
rect 5815 3115 5835 3135
rect 5815 3065 5835 3085
rect 5965 3515 5985 3535
rect 5965 3465 5985 3485
rect 5965 3415 5985 3435
rect 5965 3365 5985 3385
rect 5965 3315 5985 3335
rect 5965 3265 5985 3285
rect 5965 3215 5985 3235
rect 5965 3165 5985 3185
rect 5965 3115 5985 3135
rect 5965 3065 5985 3085
rect 6115 3515 6135 3535
rect 6115 3465 6135 3485
rect 6115 3415 6135 3435
rect 6115 3365 6135 3385
rect 6115 3315 6135 3335
rect 6115 3265 6135 3285
rect 6115 3215 6135 3235
rect 6115 3165 6135 3185
rect 6115 3115 6135 3135
rect 6115 3065 6135 3085
rect 6265 3515 6285 3535
rect 6265 3465 6285 3485
rect 6265 3415 6285 3435
rect 6265 3365 6285 3385
rect 6265 3315 6285 3335
rect 6265 3265 6285 3285
rect 6265 3215 6285 3235
rect 6265 3165 6285 3185
rect 6265 3115 6285 3135
rect 6265 3065 6285 3085
rect 6415 3515 6435 3535
rect 6415 3465 6435 3485
rect 6415 3415 6435 3435
rect 6415 3365 6435 3385
rect 6415 3315 6435 3335
rect 6415 3265 6435 3285
rect 6415 3215 6435 3235
rect 6415 3165 6435 3185
rect 6415 3115 6435 3135
rect 6415 3065 6435 3085
rect 6565 3515 6585 3535
rect 6565 3465 6585 3485
rect 6565 3415 6585 3435
rect 6565 3365 6585 3385
rect 6565 3315 6585 3335
rect 6565 3265 6585 3285
rect 6565 3215 6585 3235
rect 6565 3165 6585 3185
rect 6565 3115 6585 3135
rect 6565 3065 6585 3085
rect 6715 3515 6735 3535
rect 6715 3465 6735 3485
rect 6715 3415 6735 3435
rect 6715 3365 6735 3385
rect 6715 3315 6735 3335
rect 6715 3265 6735 3285
rect 6715 3215 6735 3235
rect 6715 3165 6735 3185
rect 6715 3115 6735 3135
rect 6715 3065 6735 3085
rect 6865 3515 6885 3535
rect 6865 3465 6885 3485
rect 6865 3415 6885 3435
rect 6865 3365 6885 3385
rect 6865 3315 6885 3335
rect 6865 3265 6885 3285
rect 6865 3215 6885 3235
rect 6865 3165 6885 3185
rect 6865 3115 6885 3135
rect 6865 3065 6885 3085
rect 7015 3515 7035 3535
rect 7015 3465 7035 3485
rect 7015 3415 7035 3435
rect 7015 3365 7035 3385
rect 7015 3315 7035 3335
rect 7015 3265 7035 3285
rect 7015 3215 7035 3235
rect 7015 3165 7035 3185
rect 7015 3115 7035 3135
rect 7015 3065 7035 3085
rect 7165 3515 7185 3535
rect 7165 3465 7185 3485
rect 7165 3415 7185 3435
rect 7165 3365 7185 3385
rect 7165 3315 7185 3335
rect 7165 3265 7185 3285
rect 7165 3215 7185 3235
rect 7165 3165 7185 3185
rect 7165 3115 7185 3135
rect 7165 3065 7185 3085
rect 7315 3515 7335 3535
rect 7315 3465 7335 3485
rect 7315 3415 7335 3435
rect 7315 3365 7335 3385
rect 7315 3315 7335 3335
rect 7315 3265 7335 3285
rect 7315 3215 7335 3235
rect 7315 3165 7335 3185
rect 7315 3115 7335 3135
rect 7315 3065 7335 3085
rect 7465 3515 7485 3535
rect 7465 3465 7485 3485
rect 7465 3415 7485 3435
rect 7465 3365 7485 3385
rect 7465 3315 7485 3335
rect 7465 3265 7485 3285
rect 7465 3215 7485 3235
rect 7465 3165 7485 3185
rect 7465 3115 7485 3135
rect 7465 3065 7485 3085
rect 7615 3515 7635 3535
rect 7615 3465 7635 3485
rect 7615 3415 7635 3435
rect 7615 3365 7635 3385
rect 7615 3315 7635 3335
rect 7615 3265 7635 3285
rect 7615 3215 7635 3235
rect 7615 3165 7635 3185
rect 7615 3115 7635 3135
rect 7615 3065 7635 3085
rect 7765 3515 7785 3535
rect 7765 3465 7785 3485
rect 7765 3415 7785 3435
rect 7765 3365 7785 3385
rect 7765 3315 7785 3335
rect 7765 3265 7785 3285
rect 7765 3215 7785 3235
rect 7765 3165 7785 3185
rect 7765 3115 7785 3135
rect 7765 3065 7785 3085
rect 8365 3515 8385 3535
rect 8365 3465 8385 3485
rect 8365 3415 8385 3435
rect 8365 3365 8385 3385
rect 8365 3315 8385 3335
rect 8365 3265 8385 3285
rect 8365 3215 8385 3235
rect 8365 3165 8385 3185
rect 8365 3115 8385 3135
rect 8365 3065 8385 3085
rect 8515 3515 8535 3535
rect 8515 3465 8535 3485
rect 8515 3415 8535 3435
rect 8515 3365 8535 3385
rect 8515 3315 8535 3335
rect 8515 3265 8535 3285
rect 8515 3215 8535 3235
rect 8515 3165 8535 3185
rect 8515 3115 8535 3135
rect 8515 3065 8535 3085
rect 8665 3515 8685 3535
rect 8665 3465 8685 3485
rect 8665 3415 8685 3435
rect 8665 3365 8685 3385
rect 8665 3315 8685 3335
rect 8665 3265 8685 3285
rect 8665 3215 8685 3235
rect 8665 3165 8685 3185
rect 8665 3115 8685 3135
rect 8665 3065 8685 3085
rect 8815 3515 8835 3535
rect 8815 3465 8835 3485
rect 8815 3415 8835 3435
rect 8815 3365 8835 3385
rect 8815 3315 8835 3335
rect 8815 3265 8835 3285
rect 8815 3215 8835 3235
rect 8815 3165 8835 3185
rect 8815 3115 8835 3135
rect 8815 3065 8835 3085
rect 8965 3515 8985 3535
rect 8965 3465 8985 3485
rect 8965 3415 8985 3435
rect 8965 3365 8985 3385
rect 8965 3315 8985 3335
rect 8965 3265 8985 3285
rect 8965 3215 8985 3235
rect 8965 3165 8985 3185
rect 8965 3115 8985 3135
rect 8965 3065 8985 3085
rect 9115 3515 9135 3535
rect 9115 3465 9135 3485
rect 9115 3415 9135 3435
rect 9115 3365 9135 3385
rect 9115 3315 9135 3335
rect 9115 3265 9135 3285
rect 9115 3215 9135 3235
rect 9115 3165 9135 3185
rect 9115 3115 9135 3135
rect 9115 3065 9135 3085
rect 9265 3515 9285 3535
rect 9265 3465 9285 3485
rect 9265 3415 9285 3435
rect 9265 3365 9285 3385
rect 9265 3315 9285 3335
rect 9265 3265 9285 3285
rect 9265 3215 9285 3235
rect 9265 3165 9285 3185
rect 9265 3115 9285 3135
rect 9265 3065 9285 3085
rect 9415 3515 9435 3535
rect 9415 3465 9435 3485
rect 9415 3415 9435 3435
rect 9415 3365 9435 3385
rect 9415 3315 9435 3335
rect 9415 3265 9435 3285
rect 9415 3215 9435 3235
rect 9415 3165 9435 3185
rect 9415 3115 9435 3135
rect 9415 3065 9435 3085
rect 9565 3515 9585 3535
rect 9565 3465 9585 3485
rect 9565 3415 9585 3435
rect 9565 3365 9585 3385
rect 9565 3315 9585 3335
rect 9565 3265 9585 3285
rect 9565 3215 9585 3235
rect 9565 3165 9585 3185
rect 9565 3115 9585 3135
rect 9565 3065 9585 3085
rect 9715 3515 9735 3535
rect 9715 3465 9735 3485
rect 9715 3415 9735 3435
rect 9715 3365 9735 3385
rect 9715 3315 9735 3335
rect 9715 3265 9735 3285
rect 9715 3215 9735 3235
rect 9715 3165 9735 3185
rect 9715 3115 9735 3135
rect 9715 3065 9735 3085
rect 9865 3515 9885 3535
rect 9865 3465 9885 3485
rect 9865 3415 9885 3435
rect 9865 3365 9885 3385
rect 9865 3315 9885 3335
rect 9865 3265 9885 3285
rect 9865 3215 9885 3235
rect 9865 3165 9885 3185
rect 9865 3115 9885 3135
rect 9865 3065 9885 3085
rect 10015 3515 10035 3535
rect 10015 3465 10035 3485
rect 10015 3415 10035 3435
rect 10015 3365 10035 3385
rect 10015 3315 10035 3335
rect 10015 3265 10035 3285
rect 10015 3215 10035 3235
rect 10015 3165 10035 3185
rect 10015 3115 10035 3135
rect 10015 3065 10035 3085
rect 10165 3515 10185 3535
rect 10165 3465 10185 3485
rect 10165 3415 10185 3435
rect 10165 3365 10185 3385
rect 10165 3315 10185 3335
rect 10165 3265 10185 3285
rect 10165 3215 10185 3235
rect 10165 3165 10185 3185
rect 10165 3115 10185 3135
rect 10165 3065 10185 3085
rect 10315 3515 10335 3535
rect 10315 3465 10335 3485
rect 10315 3415 10335 3435
rect 10315 3365 10335 3385
rect 10315 3315 10335 3335
rect 10315 3265 10335 3285
rect 10315 3215 10335 3235
rect 10315 3165 10335 3185
rect 10315 3115 10335 3135
rect 10315 3065 10335 3085
rect 10465 3515 10485 3535
rect 10465 3465 10485 3485
rect 10465 3415 10485 3435
rect 10465 3365 10485 3385
rect 10465 3315 10485 3335
rect 10465 3265 10485 3285
rect 10465 3215 10485 3235
rect 10465 3165 10485 3185
rect 10465 3115 10485 3135
rect 10465 3065 10485 3085
rect 10615 3515 10635 3535
rect 10615 3465 10635 3485
rect 10615 3415 10635 3435
rect 10615 3365 10635 3385
rect 10615 3315 10635 3335
rect 10615 3265 10635 3285
rect 10615 3215 10635 3235
rect 10615 3165 10635 3185
rect 10615 3115 10635 3135
rect 10615 3065 10635 3085
rect 10765 3515 10785 3535
rect 10765 3465 10785 3485
rect 10765 3415 10785 3435
rect 10765 3365 10785 3385
rect 10765 3315 10785 3335
rect 10765 3265 10785 3285
rect 10765 3215 10785 3235
rect 10765 3165 10785 3185
rect 10765 3115 10785 3135
rect 10765 3065 10785 3085
rect 11365 3515 11385 3535
rect 11365 3465 11385 3485
rect 11365 3415 11385 3435
rect 11365 3365 11385 3385
rect 11365 3315 11385 3335
rect 11365 3265 11385 3285
rect 11365 3215 11385 3235
rect 11365 3165 11385 3185
rect 11365 3115 11385 3135
rect 11365 3065 11385 3085
rect 11965 3515 11985 3535
rect 11965 3465 11985 3485
rect 11965 3415 11985 3435
rect 11965 3365 11985 3385
rect 11965 3315 11985 3335
rect 11965 3265 11985 3285
rect 11965 3215 11985 3235
rect 11965 3165 11985 3185
rect 11965 3115 11985 3135
rect 11965 3065 11985 3085
rect 12565 3515 12585 3535
rect 12565 3465 12585 3485
rect 12565 3415 12585 3435
rect 12565 3365 12585 3385
rect 12565 3315 12585 3335
rect 12565 3265 12585 3285
rect 12565 3215 12585 3235
rect 12565 3165 12585 3185
rect 12565 3115 12585 3135
rect 12565 3065 12585 3085
rect 13165 3515 13185 3535
rect 13165 3465 13185 3485
rect 13165 3415 13185 3435
rect 13165 3365 13185 3385
rect 13165 3315 13185 3335
rect 13165 3265 13185 3285
rect 13165 3215 13185 3235
rect 13165 3165 13185 3185
rect 13165 3115 13185 3135
rect 13165 3065 13185 3085
rect 13765 3515 13785 3535
rect 13765 3465 13785 3485
rect 13765 3415 13785 3435
rect 13765 3365 13785 3385
rect 13765 3315 13785 3335
rect 13765 3265 13785 3285
rect 13765 3215 13785 3235
rect 13765 3165 13785 3185
rect 13765 3115 13785 3135
rect 13765 3065 13785 3085
rect 14365 3515 14385 3535
rect 14365 3465 14385 3485
rect 14365 3415 14385 3435
rect 14365 3365 14385 3385
rect 14365 3315 14385 3335
rect 14365 3265 14385 3285
rect 14365 3215 14385 3235
rect 14365 3165 14385 3185
rect 14365 3115 14385 3135
rect 14365 3065 14385 3085
rect 14965 3515 14985 3535
rect 14965 3465 14985 3485
rect 14965 3415 14985 3435
rect 14965 3365 14985 3385
rect 14965 3315 14985 3335
rect 14965 3265 14985 3285
rect 14965 3215 14985 3235
rect 14965 3165 14985 3185
rect 14965 3115 14985 3135
rect 14965 3065 14985 3085
rect 15565 3515 15585 3535
rect 15565 3465 15585 3485
rect 15565 3415 15585 3435
rect 15565 3365 15585 3385
rect 15565 3315 15585 3335
rect 15565 3265 15585 3285
rect 15565 3215 15585 3235
rect 15565 3165 15585 3185
rect 15565 3115 15585 3135
rect 15565 3065 15585 3085
rect 16165 3515 16185 3535
rect 16165 3465 16185 3485
rect 16165 3415 16185 3435
rect 16165 3365 16185 3385
rect 16165 3315 16185 3335
rect 16165 3265 16185 3285
rect 16165 3215 16185 3235
rect 16165 3165 16185 3185
rect 16165 3115 16185 3135
rect 16165 3065 16185 3085
rect 16315 3515 16335 3535
rect 16315 3465 16335 3485
rect 16315 3415 16335 3435
rect 16315 3365 16335 3385
rect 16315 3315 16335 3335
rect 16315 3265 16335 3285
rect 16315 3215 16335 3235
rect 16315 3165 16335 3185
rect 16315 3115 16335 3135
rect 16315 3065 16335 3085
rect 16465 3515 16485 3535
rect 16465 3465 16485 3485
rect 16465 3415 16485 3435
rect 16465 3365 16485 3385
rect 16465 3315 16485 3335
rect 16465 3265 16485 3285
rect 16465 3215 16485 3235
rect 16465 3165 16485 3185
rect 16465 3115 16485 3135
rect 16465 3065 16485 3085
rect 16615 3515 16635 3535
rect 16615 3465 16635 3485
rect 16615 3415 16635 3435
rect 16615 3365 16635 3385
rect 16615 3315 16635 3335
rect 16615 3265 16635 3285
rect 16615 3215 16635 3235
rect 16615 3165 16635 3185
rect 16615 3115 16635 3135
rect 16615 3065 16635 3085
rect 16765 3515 16785 3535
rect 16765 3465 16785 3485
rect 16765 3415 16785 3435
rect 16765 3365 16785 3385
rect 16765 3315 16785 3335
rect 16765 3265 16785 3285
rect 16765 3215 16785 3235
rect 16765 3165 16785 3185
rect 16765 3115 16785 3135
rect 16765 3065 16785 3085
rect 16915 3515 16935 3535
rect 16915 3465 16935 3485
rect 16915 3415 16935 3435
rect 16915 3365 16935 3385
rect 16915 3315 16935 3335
rect 16915 3265 16935 3285
rect 16915 3215 16935 3235
rect 16915 3165 16935 3185
rect 16915 3115 16935 3135
rect 16915 3065 16935 3085
rect 17065 3515 17085 3535
rect 17065 3465 17085 3485
rect 17065 3415 17085 3435
rect 17065 3365 17085 3385
rect 17065 3315 17085 3335
rect 17065 3265 17085 3285
rect 17065 3215 17085 3235
rect 17065 3165 17085 3185
rect 17065 3115 17085 3135
rect 17065 3065 17085 3085
rect 17215 3515 17235 3535
rect 17215 3465 17235 3485
rect 17215 3415 17235 3435
rect 17215 3365 17235 3385
rect 17215 3315 17235 3335
rect 17215 3265 17235 3285
rect 17215 3215 17235 3235
rect 17215 3165 17235 3185
rect 17215 3115 17235 3135
rect 17215 3065 17235 3085
rect 17365 3515 17385 3535
rect 17365 3465 17385 3485
rect 17365 3415 17385 3435
rect 17365 3365 17385 3385
rect 17365 3315 17385 3335
rect 17365 3265 17385 3285
rect 17365 3215 17385 3235
rect 17365 3165 17385 3185
rect 17365 3115 17385 3135
rect 17365 3065 17385 3085
rect 17965 3515 17985 3535
rect 17965 3465 17985 3485
rect 17965 3415 17985 3435
rect 17965 3365 17985 3385
rect 17965 3315 17985 3335
rect 17965 3265 17985 3285
rect 17965 3215 17985 3235
rect 17965 3165 17985 3185
rect 17965 3115 17985 3135
rect 17965 3065 17985 3085
rect 18565 3515 18585 3535
rect 18565 3465 18585 3485
rect 18565 3415 18585 3435
rect 18565 3365 18585 3385
rect 18565 3315 18585 3335
rect 18565 3265 18585 3285
rect 18565 3215 18585 3235
rect 18565 3165 18585 3185
rect 18565 3115 18585 3135
rect 18565 3065 18585 3085
rect 18715 3515 18735 3535
rect 18715 3465 18735 3485
rect 18715 3415 18735 3435
rect 18715 3365 18735 3385
rect 18715 3315 18735 3335
rect 18715 3265 18735 3285
rect 18715 3215 18735 3235
rect 18715 3165 18735 3185
rect 18715 3115 18735 3135
rect 18715 3065 18735 3085
rect 18865 3515 18885 3535
rect 18865 3465 18885 3485
rect 18865 3415 18885 3435
rect 18865 3365 18885 3385
rect 18865 3315 18885 3335
rect 18865 3265 18885 3285
rect 18865 3215 18885 3235
rect 18865 3165 18885 3185
rect 18865 3115 18885 3135
rect 18865 3065 18885 3085
rect 19015 3515 19035 3535
rect 19015 3465 19035 3485
rect 19015 3415 19035 3435
rect 19015 3365 19035 3385
rect 19015 3315 19035 3335
rect 19015 3265 19035 3285
rect 19015 3215 19035 3235
rect 19015 3165 19035 3185
rect 19015 3115 19035 3135
rect 19015 3065 19035 3085
rect 19165 3515 19185 3535
rect 19165 3465 19185 3485
rect 19165 3415 19185 3435
rect 19165 3365 19185 3385
rect 19165 3315 19185 3335
rect 19165 3265 19185 3285
rect 19165 3215 19185 3235
rect 19165 3165 19185 3185
rect 19165 3115 19185 3135
rect 19165 3065 19185 3085
rect 19315 3515 19335 3535
rect 19315 3465 19335 3485
rect 19315 3415 19335 3435
rect 19315 3365 19335 3385
rect 19315 3315 19335 3335
rect 19315 3265 19335 3285
rect 19315 3215 19335 3235
rect 19315 3165 19335 3185
rect 19315 3115 19335 3135
rect 19315 3065 19335 3085
rect 19465 3515 19485 3535
rect 19465 3465 19485 3485
rect 19465 3415 19485 3435
rect 19465 3365 19485 3385
rect 19465 3315 19485 3335
rect 19465 3265 19485 3285
rect 19465 3215 19485 3235
rect 19465 3165 19485 3185
rect 19465 3115 19485 3135
rect 19465 3065 19485 3085
rect 19615 3515 19635 3535
rect 19615 3465 19635 3485
rect 19615 3415 19635 3435
rect 19615 3365 19635 3385
rect 19615 3315 19635 3335
rect 19615 3265 19635 3285
rect 19615 3215 19635 3235
rect 19615 3165 19635 3185
rect 19615 3115 19635 3135
rect 19615 3065 19635 3085
rect 19765 3515 19785 3535
rect 19765 3465 19785 3485
rect 19765 3415 19785 3435
rect 19765 3365 19785 3385
rect 19765 3315 19785 3335
rect 19765 3265 19785 3285
rect 19765 3215 19785 3235
rect 19765 3165 19785 3185
rect 19765 3115 19785 3135
rect 19765 3065 19785 3085
rect 20365 3515 20385 3535
rect 20365 3465 20385 3485
rect 20365 3415 20385 3435
rect 20365 3365 20385 3385
rect 20365 3315 20385 3335
rect 20365 3265 20385 3285
rect 20365 3215 20385 3235
rect 20365 3165 20385 3185
rect 20365 3115 20385 3135
rect 20365 3065 20385 3085
rect 20965 3515 20985 3535
rect 20965 3465 20985 3485
rect 20965 3415 20985 3435
rect 20965 3365 20985 3385
rect 20965 3315 20985 3335
rect 20965 3265 20985 3285
rect 20965 3215 20985 3235
rect 20965 3165 20985 3185
rect 20965 3115 20985 3135
rect 20965 3065 20985 3085
rect 21415 3515 21435 3535
rect 21415 3465 21435 3485
rect 21415 3415 21435 3435
rect 21415 3365 21435 3385
rect 21415 3315 21435 3335
rect 21415 3265 21435 3285
rect 21415 3215 21435 3235
rect 21415 3165 21435 3185
rect 21415 3115 21435 3135
rect 21415 3065 21435 3085
rect 21865 3515 21885 3535
rect 21865 3465 21885 3485
rect 21865 3415 21885 3435
rect 21865 3365 21885 3385
rect 21865 3315 21885 3335
rect 21865 3265 21885 3285
rect 21865 3215 21885 3235
rect 21865 3165 21885 3185
rect 21865 3115 21885 3135
rect 21865 3065 21885 3085
rect 22465 3515 22485 3535
rect 22465 3465 22485 3485
rect 22465 3415 22485 3435
rect 22465 3365 22485 3385
rect 22465 3315 22485 3335
rect 22465 3265 22485 3285
rect 22465 3215 22485 3235
rect 22465 3165 22485 3185
rect 22465 3115 22485 3135
rect 22465 3065 22485 3085
rect 23065 3515 23085 3535
rect 23065 3465 23085 3485
rect 23065 3415 23085 3435
rect 23065 3365 23085 3385
rect 23065 3315 23085 3335
rect 23065 3265 23085 3285
rect 23065 3215 23085 3235
rect 23065 3165 23085 3185
rect 23065 3115 23085 3135
rect 23065 3065 23085 3085
rect 23515 3515 23535 3535
rect 23515 3465 23535 3485
rect 23515 3415 23535 3435
rect 23515 3365 23535 3385
rect 23515 3315 23535 3335
rect 23515 3265 23535 3285
rect 23515 3215 23535 3235
rect 23515 3165 23535 3185
rect 23515 3115 23535 3135
rect 23515 3065 23535 3085
rect 23965 3515 23985 3535
rect 23965 3465 23985 3485
rect 23965 3415 23985 3435
rect 23965 3365 23985 3385
rect 23965 3315 23985 3335
rect 23965 3265 23985 3285
rect 23965 3215 23985 3235
rect 23965 3165 23985 3185
rect 23965 3115 23985 3135
rect 23965 3065 23985 3085
rect 24565 3515 24585 3535
rect 24565 3465 24585 3485
rect 24565 3415 24585 3435
rect 24565 3365 24585 3385
rect 24565 3315 24585 3335
rect 24565 3265 24585 3285
rect 24565 3215 24585 3235
rect 24565 3165 24585 3185
rect 24565 3115 24585 3135
rect 24565 3065 24585 3085
rect 25165 3515 25185 3535
rect 25165 3465 25185 3485
rect 25165 3415 25185 3435
rect 25165 3365 25185 3385
rect 25165 3315 25185 3335
rect 25165 3265 25185 3285
rect 25165 3215 25185 3235
rect 25165 3165 25185 3185
rect 25165 3115 25185 3135
rect 25165 3065 25185 3085
rect 25615 3515 25635 3535
rect 25615 3465 25635 3485
rect 25615 3415 25635 3435
rect 25615 3365 25635 3385
rect 25615 3315 25635 3335
rect 25615 3265 25635 3285
rect 25615 3215 25635 3235
rect 25615 3165 25635 3185
rect 25615 3115 25635 3135
rect 25615 3065 25635 3085
rect 26065 3515 26085 3535
rect 26065 3465 26085 3485
rect 26065 3415 26085 3435
rect 26065 3365 26085 3385
rect 26065 3315 26085 3335
rect 26065 3265 26085 3285
rect 26065 3215 26085 3235
rect 26065 3165 26085 3185
rect 26065 3115 26085 3135
rect 26065 3065 26085 3085
rect 26665 3515 26685 3535
rect 26665 3465 26685 3485
rect 26665 3415 26685 3435
rect 26665 3365 26685 3385
rect 26665 3315 26685 3335
rect 26665 3265 26685 3285
rect 26665 3215 26685 3235
rect 26665 3165 26685 3185
rect 26665 3115 26685 3135
rect 26665 3065 26685 3085
rect 27265 3515 27285 3535
rect 27265 3465 27285 3485
rect 27265 3415 27285 3435
rect 27265 3365 27285 3385
rect 27265 3315 27285 3335
rect 27265 3265 27285 3285
rect 27265 3215 27285 3235
rect 27265 3165 27285 3185
rect 27265 3115 27285 3135
rect 27265 3065 27285 3085
rect 27715 3515 27735 3535
rect 27715 3465 27735 3485
rect 27715 3415 27735 3435
rect 27715 3365 27735 3385
rect 27715 3315 27735 3335
rect 27715 3265 27735 3285
rect 27715 3215 27735 3235
rect 27715 3165 27735 3185
rect 27715 3115 27735 3135
rect 27715 3065 27735 3085
rect 28165 3515 28185 3535
rect 28165 3465 28185 3485
rect 28165 3415 28185 3435
rect 28165 3365 28185 3385
rect 28165 3315 28185 3335
rect 28165 3265 28185 3285
rect 28165 3215 28185 3235
rect 28165 3165 28185 3185
rect 28165 3115 28185 3135
rect 28165 3065 28185 3085
rect 28765 3515 28785 3535
rect 28765 3465 28785 3485
rect 28765 3415 28785 3435
rect 28765 3365 28785 3385
rect 28765 3315 28785 3335
rect 28765 3265 28785 3285
rect 28765 3215 28785 3235
rect 28765 3165 28785 3185
rect 28765 3115 28785 3135
rect 28765 3065 28785 3085
rect 29365 3515 29385 3535
rect 29365 3465 29385 3485
rect 29365 3415 29385 3435
rect 29365 3365 29385 3385
rect 29365 3315 29385 3335
rect 29365 3265 29385 3285
rect 29365 3215 29385 3235
rect 29365 3165 29385 3185
rect 29365 3115 29385 3135
rect 29365 3065 29385 3085
rect 29515 3515 29535 3535
rect 29515 3465 29535 3485
rect 29515 3415 29535 3435
rect 29515 3365 29535 3385
rect 29515 3315 29535 3335
rect 29515 3265 29535 3285
rect 29515 3215 29535 3235
rect 29515 3165 29535 3185
rect 29515 3115 29535 3135
rect 29515 3065 29535 3085
rect 29665 3515 29685 3535
rect 29665 3465 29685 3485
rect 29665 3415 29685 3435
rect 29665 3365 29685 3385
rect 29665 3315 29685 3335
rect 29665 3265 29685 3285
rect 29665 3215 29685 3235
rect 29665 3165 29685 3185
rect 29665 3115 29685 3135
rect 29665 3065 29685 3085
rect 29815 3515 29835 3535
rect 29815 3465 29835 3485
rect 29815 3415 29835 3435
rect 29815 3365 29835 3385
rect 29815 3315 29835 3335
rect 29815 3265 29835 3285
rect 29815 3215 29835 3235
rect 29815 3165 29835 3185
rect 29815 3115 29835 3135
rect 29815 3065 29835 3085
rect 29965 3515 29985 3535
rect 29965 3465 29985 3485
rect 29965 3415 29985 3435
rect 29965 3365 29985 3385
rect 29965 3315 29985 3335
rect 29965 3265 29985 3285
rect 29965 3215 29985 3235
rect 29965 3165 29985 3185
rect 29965 3115 29985 3135
rect 29965 3065 29985 3085
rect 30115 3515 30135 3535
rect 30115 3465 30135 3485
rect 30115 3415 30135 3435
rect 30115 3365 30135 3385
rect 30115 3315 30135 3335
rect 30115 3265 30135 3285
rect 30115 3215 30135 3235
rect 30115 3165 30135 3185
rect 30115 3115 30135 3135
rect 30115 3065 30135 3085
rect 30265 3515 30285 3535
rect 30265 3465 30285 3485
rect 30265 3415 30285 3435
rect 30265 3365 30285 3385
rect 30265 3315 30285 3335
rect 30265 3265 30285 3285
rect 30265 3215 30285 3235
rect 30265 3165 30285 3185
rect 30265 3115 30285 3135
rect 30265 3065 30285 3085
rect 30415 3515 30435 3535
rect 30415 3465 30435 3485
rect 30415 3415 30435 3435
rect 30415 3365 30435 3385
rect 30415 3315 30435 3335
rect 30415 3265 30435 3285
rect 30415 3215 30435 3235
rect 30415 3165 30435 3185
rect 30415 3115 30435 3135
rect 30415 3065 30435 3085
rect 30565 3515 30585 3535
rect 30565 3465 30585 3485
rect 30565 3415 30585 3435
rect 30565 3365 30585 3385
rect 30565 3315 30585 3335
rect 30565 3265 30585 3285
rect 30565 3215 30585 3235
rect 30565 3165 30585 3185
rect 30565 3115 30585 3135
rect 30565 3065 30585 3085
rect 30715 3515 30735 3535
rect 30715 3465 30735 3485
rect 30715 3415 30735 3435
rect 30715 3365 30735 3385
rect 30715 3315 30735 3335
rect 30715 3265 30735 3285
rect 30715 3215 30735 3235
rect 30715 3165 30735 3185
rect 30715 3115 30735 3135
rect 30715 3065 30735 3085
rect 30865 3515 30885 3535
rect 30865 3465 30885 3485
rect 30865 3415 30885 3435
rect 30865 3365 30885 3385
rect 30865 3315 30885 3335
rect 30865 3265 30885 3285
rect 30865 3215 30885 3235
rect 30865 3165 30885 3185
rect 30865 3115 30885 3135
rect 30865 3065 30885 3085
rect 31015 3515 31035 3535
rect 31015 3465 31035 3485
rect 31015 3415 31035 3435
rect 31015 3365 31035 3385
rect 31015 3315 31035 3335
rect 31015 3265 31035 3285
rect 31015 3215 31035 3235
rect 31015 3165 31035 3185
rect 31015 3115 31035 3135
rect 31015 3065 31035 3085
rect 31165 3515 31185 3535
rect 31165 3465 31185 3485
rect 31165 3415 31185 3435
rect 31165 3365 31185 3385
rect 31165 3315 31185 3335
rect 31165 3265 31185 3285
rect 31165 3215 31185 3235
rect 31165 3165 31185 3185
rect 31165 3115 31185 3135
rect 31165 3065 31185 3085
rect 31315 3515 31335 3535
rect 31315 3465 31335 3485
rect 31315 3415 31335 3435
rect 31315 3365 31335 3385
rect 31315 3315 31335 3335
rect 31315 3265 31335 3285
rect 31315 3215 31335 3235
rect 31315 3165 31335 3185
rect 31315 3115 31335 3135
rect 31315 3065 31335 3085
rect 31465 3515 31485 3535
rect 31465 3465 31485 3485
rect 31465 3415 31485 3435
rect 31465 3365 31485 3385
rect 31465 3315 31485 3335
rect 31465 3265 31485 3285
rect 31465 3215 31485 3235
rect 31465 3165 31485 3185
rect 31465 3115 31485 3135
rect 31465 3065 31485 3085
rect 32065 3515 32085 3535
rect 32065 3465 32085 3485
rect 32065 3415 32085 3435
rect 32065 3365 32085 3385
rect 32065 3315 32085 3335
rect 32065 3265 32085 3285
rect 32065 3215 32085 3235
rect 32065 3165 32085 3185
rect 32065 3115 32085 3135
rect 32065 3065 32085 3085
<< mvpsubdiff >>
rect -900 2835 32100 2850
rect -900 2815 -885 2835
rect -865 2815 -835 2835
rect -815 2815 -785 2835
rect -765 2815 -735 2835
rect -715 2815 -685 2835
rect -665 2815 -635 2835
rect -615 2815 -585 2835
rect -565 2815 -535 2835
rect -515 2815 -485 2835
rect -465 2815 -435 2835
rect -415 2815 -385 2835
rect -365 2815 -335 2835
rect -315 2815 -285 2835
rect -265 2815 -235 2835
rect -215 2815 -185 2835
rect -165 2815 -135 2835
rect -115 2815 -85 2835
rect -65 2815 -35 2835
rect -15 2815 15 2835
rect 35 2815 65 2835
rect 85 2815 115 2835
rect 135 2815 165 2835
rect 185 2815 215 2835
rect 235 2815 265 2835
rect 285 2815 315 2835
rect 335 2815 365 2835
rect 385 2815 415 2835
rect 435 2815 465 2835
rect 485 2815 515 2835
rect 535 2815 565 2835
rect 585 2815 615 2835
rect 635 2815 665 2835
rect 685 2815 715 2835
rect 735 2815 765 2835
rect 785 2815 815 2835
rect 835 2815 865 2835
rect 885 2815 915 2835
rect 935 2815 965 2835
rect 985 2815 1015 2835
rect 1035 2815 1065 2835
rect 1085 2815 1115 2835
rect 1135 2815 1165 2835
rect 1185 2815 1215 2835
rect 1235 2815 1265 2835
rect 1285 2815 1315 2835
rect 1335 2815 1365 2835
rect 1385 2815 1415 2835
rect 1435 2815 1465 2835
rect 1485 2815 1515 2835
rect 1535 2815 1565 2835
rect 1585 2815 1615 2835
rect 1635 2815 1665 2835
rect 1685 2815 1715 2835
rect 1735 2815 1765 2835
rect 1785 2815 1815 2835
rect 1835 2815 1865 2835
rect 1885 2815 1915 2835
rect 1935 2815 1965 2835
rect 1985 2815 2015 2835
rect 2035 2815 2065 2835
rect 2085 2815 2115 2835
rect 2135 2815 2165 2835
rect 2185 2815 2215 2835
rect 2235 2815 2265 2835
rect 2285 2815 2315 2835
rect 2335 2815 2365 2835
rect 2385 2815 2415 2835
rect 2435 2815 2465 2835
rect 2485 2815 2515 2835
rect 2535 2815 2565 2835
rect 2585 2815 2615 2835
rect 2635 2815 2665 2835
rect 2685 2815 2715 2835
rect 2735 2815 2765 2835
rect 2785 2815 2815 2835
rect 2835 2815 2865 2835
rect 2885 2815 2915 2835
rect 2935 2815 2965 2835
rect 2985 2815 3015 2835
rect 3035 2815 3065 2835
rect 3085 2815 3115 2835
rect 3135 2815 3165 2835
rect 3185 2815 3215 2835
rect 3235 2815 3265 2835
rect 3285 2815 3315 2835
rect 3335 2815 3365 2835
rect 3385 2815 3415 2835
rect 3435 2815 3465 2835
rect 3485 2815 3515 2835
rect 3535 2815 3565 2835
rect 3585 2815 3615 2835
rect 3635 2815 3665 2835
rect 3685 2815 3715 2835
rect 3735 2815 3765 2835
rect 3785 2815 3815 2835
rect 3835 2815 3865 2835
rect 3885 2815 3915 2835
rect 3935 2815 3965 2835
rect 3985 2815 4015 2835
rect 4035 2815 4065 2835
rect 4085 2815 4115 2835
rect 4135 2815 4165 2835
rect 4185 2815 4215 2835
rect 4235 2815 4265 2835
rect 4285 2815 4315 2835
rect 4335 2815 4365 2835
rect 4385 2815 4415 2835
rect 4435 2815 4465 2835
rect 4485 2815 4515 2835
rect 4535 2815 4565 2835
rect 4585 2815 4615 2835
rect 4635 2815 4665 2835
rect 4685 2815 4715 2835
rect 4735 2815 4765 2835
rect 4785 2815 4815 2835
rect 4835 2815 4865 2835
rect 4885 2815 4915 2835
rect 4935 2815 4965 2835
rect 4985 2815 5015 2835
rect 5035 2815 5065 2835
rect 5085 2815 5115 2835
rect 5135 2815 5165 2835
rect 5185 2815 5215 2835
rect 5235 2815 5265 2835
rect 5285 2815 5315 2835
rect 5335 2815 5365 2835
rect 5385 2815 5415 2835
rect 5435 2815 5465 2835
rect 5485 2815 5515 2835
rect 5535 2815 5565 2835
rect 5585 2815 5615 2835
rect 5635 2815 5665 2835
rect 5685 2815 5715 2835
rect 5735 2815 5765 2835
rect 5785 2815 5815 2835
rect 5835 2815 5865 2835
rect 5885 2815 5915 2835
rect 5935 2815 5965 2835
rect 5985 2815 6015 2835
rect 6035 2815 6065 2835
rect 6085 2815 6115 2835
rect 6135 2815 6165 2835
rect 6185 2815 6215 2835
rect 6235 2815 6265 2835
rect 6285 2815 6315 2835
rect 6335 2815 6365 2835
rect 6385 2815 6415 2835
rect 6435 2815 6465 2835
rect 6485 2815 6515 2835
rect 6535 2815 6565 2835
rect 6585 2815 6615 2835
rect 6635 2815 6665 2835
rect 6685 2815 6715 2835
rect 6735 2815 6765 2835
rect 6785 2815 6815 2835
rect 6835 2815 6865 2835
rect 6885 2815 6915 2835
rect 6935 2815 6965 2835
rect 6985 2815 7015 2835
rect 7035 2815 7065 2835
rect 7085 2815 7115 2835
rect 7135 2815 7165 2835
rect 7185 2815 7215 2835
rect 7235 2815 7265 2835
rect 7285 2815 7315 2835
rect 7335 2815 7365 2835
rect 7385 2815 7415 2835
rect 7435 2815 7465 2835
rect 7485 2815 7515 2835
rect 7535 2815 7565 2835
rect 7585 2815 7615 2835
rect 7635 2815 7665 2835
rect 7685 2815 7715 2835
rect 7735 2815 7765 2835
rect 7785 2815 7815 2835
rect 7835 2815 7865 2835
rect 7885 2815 7915 2835
rect 7935 2815 7965 2835
rect 7985 2815 8015 2835
rect 8035 2815 8065 2835
rect 8085 2815 8115 2835
rect 8135 2815 8165 2835
rect 8185 2815 8215 2835
rect 8235 2815 8265 2835
rect 8285 2815 8315 2835
rect 8335 2815 8365 2835
rect 8385 2815 8415 2835
rect 8435 2815 8465 2835
rect 8485 2815 8515 2835
rect 8535 2815 8565 2835
rect 8585 2815 8615 2835
rect 8635 2815 8665 2835
rect 8685 2815 8715 2835
rect 8735 2815 8765 2835
rect 8785 2815 8815 2835
rect 8835 2815 8865 2835
rect 8885 2815 8915 2835
rect 8935 2815 8965 2835
rect 8985 2815 9015 2835
rect 9035 2815 9065 2835
rect 9085 2815 9115 2835
rect 9135 2815 9165 2835
rect 9185 2815 9215 2835
rect 9235 2815 9265 2835
rect 9285 2815 9315 2835
rect 9335 2815 9365 2835
rect 9385 2815 9415 2835
rect 9435 2815 9465 2835
rect 9485 2815 9515 2835
rect 9535 2815 9565 2835
rect 9585 2815 9615 2835
rect 9635 2815 9665 2835
rect 9685 2815 9715 2835
rect 9735 2815 9765 2835
rect 9785 2815 9815 2835
rect 9835 2815 9865 2835
rect 9885 2815 9915 2835
rect 9935 2815 9965 2835
rect 9985 2815 10015 2835
rect 10035 2815 10065 2835
rect 10085 2815 10115 2835
rect 10135 2815 10165 2835
rect 10185 2815 10215 2835
rect 10235 2815 10265 2835
rect 10285 2815 10315 2835
rect 10335 2815 10365 2835
rect 10385 2815 10415 2835
rect 10435 2815 10465 2835
rect 10485 2815 10515 2835
rect 10535 2815 10565 2835
rect 10585 2815 10615 2835
rect 10635 2815 10665 2835
rect 10685 2815 10715 2835
rect 10735 2815 10765 2835
rect 10785 2815 10815 2835
rect 10835 2815 10865 2835
rect 10885 2815 10915 2835
rect 10935 2815 10965 2835
rect 10985 2815 11015 2835
rect 11035 2815 11065 2835
rect 11085 2815 11115 2835
rect 11135 2815 11165 2835
rect 11185 2815 11215 2835
rect 11235 2815 11265 2835
rect 11285 2815 11315 2835
rect 11335 2815 11365 2835
rect 11385 2815 11415 2835
rect 11435 2815 11465 2835
rect 11485 2815 11515 2835
rect 11535 2815 11565 2835
rect 11585 2815 11615 2835
rect 11635 2815 11665 2835
rect 11685 2815 11715 2835
rect 11735 2815 11765 2835
rect 11785 2815 11815 2835
rect 11835 2815 11865 2835
rect 11885 2815 11915 2835
rect 11935 2815 11965 2835
rect 11985 2815 12015 2835
rect 12035 2815 12065 2835
rect 12085 2815 12115 2835
rect 12135 2815 12165 2835
rect 12185 2815 12215 2835
rect 12235 2815 12265 2835
rect 12285 2815 12315 2835
rect 12335 2815 12365 2835
rect 12385 2815 12415 2835
rect 12435 2815 12465 2835
rect 12485 2815 12515 2835
rect 12535 2815 12565 2835
rect 12585 2815 12615 2835
rect 12635 2815 12665 2835
rect 12685 2815 12715 2835
rect 12735 2815 12765 2835
rect 12785 2815 12815 2835
rect 12835 2815 12865 2835
rect 12885 2815 12915 2835
rect 12935 2815 12965 2835
rect 12985 2815 13015 2835
rect 13035 2815 13065 2835
rect 13085 2815 13115 2835
rect 13135 2815 13165 2835
rect 13185 2815 13215 2835
rect 13235 2815 13265 2835
rect 13285 2815 13315 2835
rect 13335 2815 13365 2835
rect 13385 2815 13415 2835
rect 13435 2815 13465 2835
rect 13485 2815 13515 2835
rect 13535 2815 13565 2835
rect 13585 2815 13615 2835
rect 13635 2815 13665 2835
rect 13685 2815 13715 2835
rect 13735 2815 13765 2835
rect 13785 2815 13815 2835
rect 13835 2815 13865 2835
rect 13885 2815 13915 2835
rect 13935 2815 13965 2835
rect 13985 2815 14015 2835
rect 14035 2815 14065 2835
rect 14085 2815 14115 2835
rect 14135 2815 14165 2835
rect 14185 2815 14215 2835
rect 14235 2815 14265 2835
rect 14285 2815 14315 2835
rect 14335 2815 14365 2835
rect 14385 2815 14415 2835
rect 14435 2815 14465 2835
rect 14485 2815 14515 2835
rect 14535 2815 14565 2835
rect 14585 2815 14615 2835
rect 14635 2815 14665 2835
rect 14685 2815 14715 2835
rect 14735 2815 14765 2835
rect 14785 2815 14815 2835
rect 14835 2815 14865 2835
rect 14885 2815 14915 2835
rect 14935 2815 14965 2835
rect 14985 2815 15015 2835
rect 15035 2815 15065 2835
rect 15085 2815 15115 2835
rect 15135 2815 15165 2835
rect 15185 2815 15215 2835
rect 15235 2815 15265 2835
rect 15285 2815 15315 2835
rect 15335 2815 15365 2835
rect 15385 2815 15415 2835
rect 15435 2815 15465 2835
rect 15485 2815 15515 2835
rect 15535 2815 15565 2835
rect 15585 2815 15615 2835
rect 15635 2815 15665 2835
rect 15685 2815 15715 2835
rect 15735 2815 15765 2835
rect 15785 2815 15815 2835
rect 15835 2815 15865 2835
rect 15885 2815 15915 2835
rect 15935 2815 15965 2835
rect 15985 2815 16015 2835
rect 16035 2815 16065 2835
rect 16085 2815 16115 2835
rect 16135 2815 16165 2835
rect 16185 2815 16215 2835
rect 16235 2815 16265 2835
rect 16285 2815 16315 2835
rect 16335 2815 16365 2835
rect 16385 2815 16415 2835
rect 16435 2815 16465 2835
rect 16485 2815 16515 2835
rect 16535 2815 16565 2835
rect 16585 2815 16615 2835
rect 16635 2815 16665 2835
rect 16685 2815 16715 2835
rect 16735 2815 16765 2835
rect 16785 2815 16815 2835
rect 16835 2815 16865 2835
rect 16885 2815 16915 2835
rect 16935 2815 16965 2835
rect 16985 2815 17015 2835
rect 17035 2815 17065 2835
rect 17085 2815 17115 2835
rect 17135 2815 17165 2835
rect 17185 2815 17215 2835
rect 17235 2815 17265 2835
rect 17285 2815 17315 2835
rect 17335 2815 17365 2835
rect 17385 2815 17415 2835
rect 17435 2815 17465 2835
rect 17485 2815 17515 2835
rect 17535 2815 17565 2835
rect 17585 2815 17615 2835
rect 17635 2815 17665 2835
rect 17685 2815 17715 2835
rect 17735 2815 17765 2835
rect 17785 2815 17815 2835
rect 17835 2815 17865 2835
rect 17885 2815 17915 2835
rect 17935 2815 17965 2835
rect 17985 2815 18015 2835
rect 18035 2815 18065 2835
rect 18085 2815 18115 2835
rect 18135 2815 18165 2835
rect 18185 2815 18215 2835
rect 18235 2815 18265 2835
rect 18285 2815 18315 2835
rect 18335 2815 18365 2835
rect 18385 2815 18415 2835
rect 18435 2815 18465 2835
rect 18485 2815 18515 2835
rect 18535 2815 18565 2835
rect 18585 2815 18615 2835
rect 18635 2815 18665 2835
rect 18685 2815 18715 2835
rect 18735 2815 18765 2835
rect 18785 2815 18815 2835
rect 18835 2815 18865 2835
rect 18885 2815 18915 2835
rect 18935 2815 18965 2835
rect 18985 2815 19015 2835
rect 19035 2815 19065 2835
rect 19085 2815 19115 2835
rect 19135 2815 19165 2835
rect 19185 2815 19215 2835
rect 19235 2815 19265 2835
rect 19285 2815 19315 2835
rect 19335 2815 19365 2835
rect 19385 2815 19415 2835
rect 19435 2815 19465 2835
rect 19485 2815 19515 2835
rect 19535 2815 19565 2835
rect 19585 2815 19615 2835
rect 19635 2815 19665 2835
rect 19685 2815 19715 2835
rect 19735 2815 19765 2835
rect 19785 2815 19815 2835
rect 19835 2815 19865 2835
rect 19885 2815 19915 2835
rect 19935 2815 19965 2835
rect 19985 2815 20015 2835
rect 20035 2815 20065 2835
rect 20085 2815 20115 2835
rect 20135 2815 20165 2835
rect 20185 2815 20215 2835
rect 20235 2815 20265 2835
rect 20285 2815 20315 2835
rect 20335 2815 20365 2835
rect 20385 2815 20415 2835
rect 20435 2815 20465 2835
rect 20485 2815 20515 2835
rect 20535 2815 20565 2835
rect 20585 2815 20615 2835
rect 20635 2815 20665 2835
rect 20685 2815 20715 2835
rect 20735 2815 20765 2835
rect 20785 2815 20815 2835
rect 20835 2815 20865 2835
rect 20885 2815 20915 2835
rect 20935 2815 20965 2835
rect 20985 2815 21015 2835
rect 21035 2815 21065 2835
rect 21085 2815 21115 2835
rect 21135 2815 21165 2835
rect 21185 2815 21215 2835
rect 21235 2815 21265 2835
rect 21285 2815 21315 2835
rect 21335 2815 21365 2835
rect 21385 2815 21415 2835
rect 21435 2815 21465 2835
rect 21485 2815 21515 2835
rect 21535 2815 21565 2835
rect 21585 2815 21615 2835
rect 21635 2815 21665 2835
rect 21685 2815 21715 2835
rect 21735 2815 21765 2835
rect 21785 2815 21815 2835
rect 21835 2815 21865 2835
rect 21885 2815 21915 2835
rect 21935 2815 21965 2835
rect 21985 2815 22015 2835
rect 22035 2815 22065 2835
rect 22085 2815 22115 2835
rect 22135 2815 22165 2835
rect 22185 2815 22215 2835
rect 22235 2815 22265 2835
rect 22285 2815 22315 2835
rect 22335 2815 22365 2835
rect 22385 2815 22415 2835
rect 22435 2815 22465 2835
rect 22485 2815 22515 2835
rect 22535 2815 22565 2835
rect 22585 2815 22615 2835
rect 22635 2815 22665 2835
rect 22685 2815 22715 2835
rect 22735 2815 22765 2835
rect 22785 2815 22815 2835
rect 22835 2815 22865 2835
rect 22885 2815 22915 2835
rect 22935 2815 22965 2835
rect 22985 2815 23015 2835
rect 23035 2815 23065 2835
rect 23085 2815 23115 2835
rect 23135 2815 23165 2835
rect 23185 2815 23215 2835
rect 23235 2815 23265 2835
rect 23285 2815 23315 2835
rect 23335 2815 23365 2835
rect 23385 2815 23415 2835
rect 23435 2815 23465 2835
rect 23485 2815 23515 2835
rect 23535 2815 23565 2835
rect 23585 2815 23615 2835
rect 23635 2815 23665 2835
rect 23685 2815 23715 2835
rect 23735 2815 23765 2835
rect 23785 2815 23815 2835
rect 23835 2815 23865 2835
rect 23885 2815 23915 2835
rect 23935 2815 23965 2835
rect 23985 2815 24015 2835
rect 24035 2815 24065 2835
rect 24085 2815 24115 2835
rect 24135 2815 24165 2835
rect 24185 2815 24215 2835
rect 24235 2815 24265 2835
rect 24285 2815 24315 2835
rect 24335 2815 24365 2835
rect 24385 2815 24415 2835
rect 24435 2815 24465 2835
rect 24485 2815 24515 2835
rect 24535 2815 24565 2835
rect 24585 2815 24615 2835
rect 24635 2815 24665 2835
rect 24685 2815 24715 2835
rect 24735 2815 24765 2835
rect 24785 2815 24815 2835
rect 24835 2815 24865 2835
rect 24885 2815 24915 2835
rect 24935 2815 24965 2835
rect 24985 2815 25015 2835
rect 25035 2815 25065 2835
rect 25085 2815 25115 2835
rect 25135 2815 25165 2835
rect 25185 2815 25215 2835
rect 25235 2815 25265 2835
rect 25285 2815 25315 2835
rect 25335 2815 25365 2835
rect 25385 2815 25415 2835
rect 25435 2815 25465 2835
rect 25485 2815 25515 2835
rect 25535 2815 25565 2835
rect 25585 2815 25615 2835
rect 25635 2815 25665 2835
rect 25685 2815 25715 2835
rect 25735 2815 25765 2835
rect 25785 2815 25815 2835
rect 25835 2815 25865 2835
rect 25885 2815 25915 2835
rect 25935 2815 25965 2835
rect 25985 2815 26015 2835
rect 26035 2815 26065 2835
rect 26085 2815 26115 2835
rect 26135 2815 26165 2835
rect 26185 2815 26215 2835
rect 26235 2815 26265 2835
rect 26285 2815 26315 2835
rect 26335 2815 26365 2835
rect 26385 2815 26415 2835
rect 26435 2815 26465 2835
rect 26485 2815 26515 2835
rect 26535 2815 26565 2835
rect 26585 2815 26615 2835
rect 26635 2815 26665 2835
rect 26685 2815 26715 2835
rect 26735 2815 26765 2835
rect 26785 2815 26815 2835
rect 26835 2815 26865 2835
rect 26885 2815 26915 2835
rect 26935 2815 26965 2835
rect 26985 2815 27015 2835
rect 27035 2815 27065 2835
rect 27085 2815 27115 2835
rect 27135 2815 27165 2835
rect 27185 2815 27215 2835
rect 27235 2815 27265 2835
rect 27285 2815 27315 2835
rect 27335 2815 27365 2835
rect 27385 2815 27415 2835
rect 27435 2815 27465 2835
rect 27485 2815 27515 2835
rect 27535 2815 27565 2835
rect 27585 2815 27615 2835
rect 27635 2815 27665 2835
rect 27685 2815 27715 2835
rect 27735 2815 27765 2835
rect 27785 2815 27815 2835
rect 27835 2815 27865 2835
rect 27885 2815 27915 2835
rect 27935 2815 27965 2835
rect 27985 2815 28015 2835
rect 28035 2815 28065 2835
rect 28085 2815 28115 2835
rect 28135 2815 28165 2835
rect 28185 2815 28215 2835
rect 28235 2815 28265 2835
rect 28285 2815 28315 2835
rect 28335 2815 28365 2835
rect 28385 2815 28415 2835
rect 28435 2815 28465 2835
rect 28485 2815 28515 2835
rect 28535 2815 28565 2835
rect 28585 2815 28615 2835
rect 28635 2815 28665 2835
rect 28685 2815 28715 2835
rect 28735 2815 28765 2835
rect 28785 2815 28815 2835
rect 28835 2815 28865 2835
rect 28885 2815 28915 2835
rect 28935 2815 28965 2835
rect 28985 2815 29015 2835
rect 29035 2815 29065 2835
rect 29085 2815 29115 2835
rect 29135 2815 29165 2835
rect 29185 2815 29215 2835
rect 29235 2815 29265 2835
rect 29285 2815 29315 2835
rect 29335 2815 29365 2835
rect 29385 2815 29415 2835
rect 29435 2815 29465 2835
rect 29485 2815 29515 2835
rect 29535 2815 29565 2835
rect 29585 2815 29615 2835
rect 29635 2815 29665 2835
rect 29685 2815 29715 2835
rect 29735 2815 29765 2835
rect 29785 2815 29815 2835
rect 29835 2815 29865 2835
rect 29885 2815 29915 2835
rect 29935 2815 29965 2835
rect 29985 2815 30015 2835
rect 30035 2815 30065 2835
rect 30085 2815 30115 2835
rect 30135 2815 30165 2835
rect 30185 2815 30215 2835
rect 30235 2815 30265 2835
rect 30285 2815 30315 2835
rect 30335 2815 30365 2835
rect 30385 2815 30415 2835
rect 30435 2815 30465 2835
rect 30485 2815 30515 2835
rect 30535 2815 30565 2835
rect 30585 2815 30615 2835
rect 30635 2815 30665 2835
rect 30685 2815 30715 2835
rect 30735 2815 30765 2835
rect 30785 2815 30815 2835
rect 30835 2815 30865 2835
rect 30885 2815 30915 2835
rect 30935 2815 30965 2835
rect 30985 2815 31015 2835
rect 31035 2815 31065 2835
rect 31085 2815 31115 2835
rect 31135 2815 31165 2835
rect 31185 2815 31215 2835
rect 31235 2815 31265 2835
rect 31285 2815 31315 2835
rect 31335 2815 31365 2835
rect 31385 2815 31415 2835
rect 31435 2815 31465 2835
rect 31485 2815 31515 2835
rect 31535 2815 31565 2835
rect 31585 2815 31615 2835
rect 31635 2815 31665 2835
rect 31685 2815 31715 2835
rect 31735 2815 31765 2835
rect 31785 2815 31815 2835
rect 31835 2815 31865 2835
rect 31885 2815 31915 2835
rect 31935 2815 31965 2835
rect 31985 2815 32015 2835
rect 32035 2815 32065 2835
rect 32085 2815 32100 2835
rect -900 2800 32100 2815
rect -900 2035 28800 2050
rect -900 2015 -885 2035
rect -865 2015 -835 2035
rect -815 2015 -785 2035
rect -765 2015 -735 2035
rect -715 2015 -685 2035
rect -665 2015 -635 2035
rect -615 2015 -585 2035
rect -565 2015 -535 2035
rect -515 2015 -485 2035
rect -465 2015 -435 2035
rect -415 2015 -385 2035
rect -365 2015 -335 2035
rect -315 2015 -285 2035
rect -265 2015 -235 2035
rect -215 2015 -185 2035
rect -165 2015 -135 2035
rect -115 2015 -85 2035
rect -65 2015 -35 2035
rect -15 2015 15 2035
rect 35 2015 65 2035
rect 85 2015 115 2035
rect 135 2015 165 2035
rect 185 2015 215 2035
rect 235 2015 265 2035
rect 285 2015 315 2035
rect 335 2015 365 2035
rect 385 2015 415 2035
rect 435 2015 465 2035
rect 485 2015 515 2035
rect 535 2015 565 2035
rect 585 2015 615 2035
rect 635 2015 665 2035
rect 685 2015 715 2035
rect 735 2015 765 2035
rect 785 2015 815 2035
rect 835 2015 865 2035
rect 885 2015 915 2035
rect 935 2015 965 2035
rect 985 2015 1015 2035
rect 1035 2015 1065 2035
rect 1085 2015 1115 2035
rect 1135 2015 1165 2035
rect 1185 2015 1215 2035
rect 1235 2015 1265 2035
rect 1285 2015 1315 2035
rect 1335 2015 1365 2035
rect 1385 2015 1415 2035
rect 1435 2015 1465 2035
rect 1485 2015 1515 2035
rect 1535 2015 1565 2035
rect 1585 2015 1615 2035
rect 1635 2015 1665 2035
rect 1685 2015 1715 2035
rect 1735 2015 1765 2035
rect 1785 2015 1815 2035
rect 1835 2015 1865 2035
rect 1885 2015 1915 2035
rect 1935 2015 1965 2035
rect 1985 2015 2015 2035
rect 2035 2015 2065 2035
rect 2085 2015 2115 2035
rect 2135 2015 2165 2035
rect 2185 2015 2215 2035
rect 2235 2015 2265 2035
rect 2285 2015 2315 2035
rect 2335 2015 2365 2035
rect 2385 2015 2415 2035
rect 2435 2015 2465 2035
rect 2485 2015 2515 2035
rect 2535 2015 2565 2035
rect 2585 2015 2615 2035
rect 2635 2015 2665 2035
rect 2685 2015 2715 2035
rect 2735 2015 2765 2035
rect 2785 2015 2815 2035
rect 2835 2015 2865 2035
rect 2885 2015 2915 2035
rect 2935 2015 2965 2035
rect 2985 2015 3015 2035
rect 3035 2015 3065 2035
rect 3085 2015 3115 2035
rect 3135 2015 3165 2035
rect 3185 2015 3215 2035
rect 3235 2015 3265 2035
rect 3285 2015 3315 2035
rect 3335 2015 3365 2035
rect 3385 2015 3415 2035
rect 3435 2015 3465 2035
rect 3485 2015 3515 2035
rect 3535 2015 3565 2035
rect 3585 2015 3615 2035
rect 3635 2015 3665 2035
rect 3685 2015 3715 2035
rect 3735 2015 3765 2035
rect 3785 2015 3815 2035
rect 3835 2015 3865 2035
rect 3885 2015 3915 2035
rect 3935 2015 3965 2035
rect 3985 2015 4015 2035
rect 4035 2015 4065 2035
rect 4085 2015 4115 2035
rect 4135 2015 4165 2035
rect 4185 2015 4215 2035
rect 4235 2015 4265 2035
rect 4285 2015 4315 2035
rect 4335 2015 4365 2035
rect 4385 2015 4415 2035
rect 4435 2015 4465 2035
rect 4485 2015 4515 2035
rect 4535 2015 4565 2035
rect 4585 2015 4615 2035
rect 4635 2015 4665 2035
rect 4685 2015 4715 2035
rect 4735 2015 4765 2035
rect 4785 2015 4815 2035
rect 4835 2015 4865 2035
rect 4885 2015 4915 2035
rect 4935 2015 4965 2035
rect 4985 2015 5015 2035
rect 5035 2015 5065 2035
rect 5085 2015 5115 2035
rect 5135 2015 5165 2035
rect 5185 2015 5215 2035
rect 5235 2015 5265 2035
rect 5285 2015 5315 2035
rect 5335 2015 5365 2035
rect 5385 2015 5415 2035
rect 5435 2015 5465 2035
rect 5485 2015 5515 2035
rect 5535 2015 5565 2035
rect 5585 2015 5615 2035
rect 5635 2015 5665 2035
rect 5685 2015 5715 2035
rect 5735 2015 5765 2035
rect 5785 2015 5815 2035
rect 5835 2015 5865 2035
rect 5885 2015 5915 2035
rect 5935 2015 5965 2035
rect 5985 2015 6015 2035
rect 6035 2015 6065 2035
rect 6085 2015 6115 2035
rect 6135 2015 6165 2035
rect 6185 2015 6215 2035
rect 6235 2015 6265 2035
rect 6285 2015 6315 2035
rect 6335 2015 6365 2035
rect 6385 2015 6415 2035
rect 6435 2015 6465 2035
rect 6485 2015 6515 2035
rect 6535 2015 6565 2035
rect 6585 2015 6615 2035
rect 6635 2015 6665 2035
rect 6685 2015 6715 2035
rect 6735 2015 6765 2035
rect 6785 2015 6815 2035
rect 6835 2015 6865 2035
rect 6885 2015 6915 2035
rect 6935 2015 6965 2035
rect 6985 2015 7015 2035
rect 7035 2015 7065 2035
rect 7085 2015 7115 2035
rect 7135 2015 7165 2035
rect 7185 2015 7215 2035
rect 7235 2015 7265 2035
rect 7285 2015 7315 2035
rect 7335 2015 7365 2035
rect 7385 2015 7415 2035
rect 7435 2015 7465 2035
rect 7485 2015 7515 2035
rect 7535 2015 7565 2035
rect 7585 2015 7615 2035
rect 7635 2015 7665 2035
rect 7685 2015 7715 2035
rect 7735 2015 7765 2035
rect 7785 2015 7815 2035
rect 7835 2015 7865 2035
rect 7885 2015 7915 2035
rect 7935 2015 7965 2035
rect 7985 2015 8015 2035
rect 8035 2015 8065 2035
rect 8085 2015 8115 2035
rect 8135 2015 8165 2035
rect 8185 2015 8215 2035
rect 8235 2015 8265 2035
rect 8285 2015 8315 2035
rect 8335 2015 8365 2035
rect 8385 2015 8415 2035
rect 8435 2015 8465 2035
rect 8485 2015 8515 2035
rect 8535 2015 8565 2035
rect 8585 2015 8615 2035
rect 8635 2015 8665 2035
rect 8685 2015 8715 2035
rect 8735 2015 8765 2035
rect 8785 2015 8815 2035
rect 8835 2015 8865 2035
rect 8885 2015 8915 2035
rect 8935 2015 8965 2035
rect 8985 2015 9015 2035
rect 9035 2015 9065 2035
rect 9085 2015 9115 2035
rect 9135 2015 9165 2035
rect 9185 2015 9215 2035
rect 9235 2015 9265 2035
rect 9285 2015 9315 2035
rect 9335 2015 9365 2035
rect 9385 2015 9415 2035
rect 9435 2015 9465 2035
rect 9485 2015 9515 2035
rect 9535 2015 9565 2035
rect 9585 2015 9615 2035
rect 9635 2015 9665 2035
rect 9685 2015 9715 2035
rect 9735 2015 9765 2035
rect 9785 2015 9815 2035
rect 9835 2015 9865 2035
rect 9885 2015 9915 2035
rect 9935 2015 9965 2035
rect 9985 2015 10015 2035
rect 10035 2015 10065 2035
rect 10085 2015 10115 2035
rect 10135 2015 10165 2035
rect 10185 2015 10215 2035
rect 10235 2015 10265 2035
rect 10285 2015 10315 2035
rect 10335 2015 10365 2035
rect 10385 2015 10415 2035
rect 10435 2015 10465 2035
rect 10485 2015 10515 2035
rect 10535 2015 10565 2035
rect 10585 2015 10615 2035
rect 10635 2015 10665 2035
rect 10685 2015 10715 2035
rect 10735 2015 10765 2035
rect 10785 2015 10815 2035
rect 10835 2015 10865 2035
rect 10885 2015 10915 2035
rect 10935 2015 10965 2035
rect 10985 2015 11015 2035
rect 11035 2015 11065 2035
rect 11085 2015 11115 2035
rect 11135 2015 11165 2035
rect 11185 2015 11215 2035
rect 11235 2015 11265 2035
rect 11285 2015 11315 2035
rect 11335 2015 11365 2035
rect 11385 2015 11415 2035
rect 11435 2015 11465 2035
rect 11485 2015 11515 2035
rect 11535 2015 11565 2035
rect 11585 2015 11615 2035
rect 11635 2015 11665 2035
rect 11685 2015 11715 2035
rect 11735 2015 11765 2035
rect 11785 2015 11815 2035
rect 11835 2015 11865 2035
rect 11885 2015 11915 2035
rect 11935 2015 11965 2035
rect 11985 2015 12015 2035
rect 12035 2015 12065 2035
rect 12085 2015 12115 2035
rect 12135 2015 12165 2035
rect 12185 2015 12215 2035
rect 12235 2015 12265 2035
rect 12285 2015 12315 2035
rect 12335 2015 12365 2035
rect 12385 2015 12415 2035
rect 12435 2015 12465 2035
rect 12485 2015 12515 2035
rect 12535 2015 12565 2035
rect 12585 2015 12615 2035
rect 12635 2015 12665 2035
rect 12685 2015 12715 2035
rect 12735 2015 12765 2035
rect 12785 2015 12815 2035
rect 12835 2015 12865 2035
rect 12885 2015 12915 2035
rect 12935 2015 12965 2035
rect 12985 2015 13015 2035
rect 13035 2015 13065 2035
rect 13085 2015 13115 2035
rect 13135 2015 13165 2035
rect 13185 2015 13215 2035
rect 13235 2015 13265 2035
rect 13285 2015 13315 2035
rect 13335 2015 13365 2035
rect 13385 2015 13415 2035
rect 13435 2015 13465 2035
rect 13485 2015 13515 2035
rect 13535 2015 13565 2035
rect 13585 2015 13615 2035
rect 13635 2015 13665 2035
rect 13685 2015 13715 2035
rect 13735 2015 13765 2035
rect 13785 2015 13815 2035
rect 13835 2015 13865 2035
rect 13885 2015 13915 2035
rect 13935 2015 13965 2035
rect 13985 2015 14015 2035
rect 14035 2015 14065 2035
rect 14085 2015 14115 2035
rect 14135 2015 14165 2035
rect 14185 2015 14215 2035
rect 14235 2015 14265 2035
rect 14285 2015 14315 2035
rect 14335 2015 14365 2035
rect 14385 2015 14415 2035
rect 14435 2015 14465 2035
rect 14485 2015 14515 2035
rect 14535 2015 14565 2035
rect 14585 2015 14615 2035
rect 14635 2015 14665 2035
rect 14685 2015 14715 2035
rect 14735 2015 14765 2035
rect 14785 2015 14815 2035
rect 14835 2015 14865 2035
rect 14885 2015 14915 2035
rect 14935 2015 14965 2035
rect 14985 2015 15015 2035
rect 15035 2015 15065 2035
rect 15085 2015 15115 2035
rect 15135 2015 15165 2035
rect 15185 2015 15215 2035
rect 15235 2015 15265 2035
rect 15285 2015 15315 2035
rect 15335 2015 15365 2035
rect 15385 2015 15415 2035
rect 15435 2015 15465 2035
rect 15485 2015 15515 2035
rect 15535 2015 15565 2035
rect 15585 2015 15615 2035
rect 15635 2015 15665 2035
rect 15685 2015 15715 2035
rect 15735 2015 15765 2035
rect 15785 2015 15815 2035
rect 15835 2015 15865 2035
rect 15885 2015 15915 2035
rect 15935 2015 15965 2035
rect 15985 2015 16015 2035
rect 16035 2015 16065 2035
rect 16085 2015 16115 2035
rect 16135 2015 16165 2035
rect 16185 2015 16215 2035
rect 16235 2015 16265 2035
rect 16285 2015 16315 2035
rect 16335 2015 16365 2035
rect 16385 2015 16415 2035
rect 16435 2015 16465 2035
rect 16485 2015 16515 2035
rect 16535 2015 16565 2035
rect 16585 2015 16615 2035
rect 16635 2015 16665 2035
rect 16685 2015 16715 2035
rect 16735 2015 16765 2035
rect 16785 2015 16815 2035
rect 16835 2015 16865 2035
rect 16885 2015 16915 2035
rect 16935 2015 16965 2035
rect 16985 2015 17015 2035
rect 17035 2015 17065 2035
rect 17085 2015 17115 2035
rect 17135 2015 17165 2035
rect 17185 2015 17215 2035
rect 17235 2015 17265 2035
rect 17285 2015 17315 2035
rect 17335 2015 17365 2035
rect 17385 2015 17415 2035
rect 17435 2015 17465 2035
rect 17485 2015 17515 2035
rect 17535 2015 17565 2035
rect 17585 2015 17615 2035
rect 17635 2015 17665 2035
rect 17685 2015 17715 2035
rect 17735 2015 17765 2035
rect 17785 2015 17815 2035
rect 17835 2015 17865 2035
rect 17885 2015 17915 2035
rect 17935 2015 17965 2035
rect 17985 2015 18015 2035
rect 18035 2015 18065 2035
rect 18085 2015 18115 2035
rect 18135 2015 18165 2035
rect 18185 2015 18215 2035
rect 18235 2015 18265 2035
rect 18285 2015 18315 2035
rect 18335 2015 18365 2035
rect 18385 2015 18415 2035
rect 18435 2015 18465 2035
rect 18485 2015 18515 2035
rect 18535 2015 18565 2035
rect 18585 2015 18615 2035
rect 18635 2015 18665 2035
rect 18685 2015 18715 2035
rect 18735 2015 18765 2035
rect 18785 2015 18815 2035
rect 18835 2015 18865 2035
rect 18885 2015 18915 2035
rect 18935 2015 18965 2035
rect 18985 2015 19015 2035
rect 19035 2015 19065 2035
rect 19085 2015 19115 2035
rect 19135 2015 19165 2035
rect 19185 2015 19215 2035
rect 19235 2015 19265 2035
rect 19285 2015 19315 2035
rect 19335 2015 19365 2035
rect 19385 2015 19415 2035
rect 19435 2015 19465 2035
rect 19485 2015 19515 2035
rect 19535 2015 19565 2035
rect 19585 2015 19615 2035
rect 19635 2015 19665 2035
rect 19685 2015 19715 2035
rect 19735 2015 19765 2035
rect 19785 2015 19815 2035
rect 19835 2015 19865 2035
rect 19885 2015 19915 2035
rect 19935 2015 19965 2035
rect 19985 2015 20015 2035
rect 20035 2015 20065 2035
rect 20085 2015 20115 2035
rect 20135 2015 20165 2035
rect 20185 2015 20215 2035
rect 20235 2015 20265 2035
rect 20285 2015 20315 2035
rect 20335 2015 20365 2035
rect 20385 2015 20415 2035
rect 20435 2015 20465 2035
rect 20485 2015 20515 2035
rect 20535 2015 20565 2035
rect 20585 2015 20615 2035
rect 20635 2015 20665 2035
rect 20685 2015 20715 2035
rect 20735 2015 20765 2035
rect 20785 2015 20815 2035
rect 20835 2015 20865 2035
rect 20885 2015 20915 2035
rect 20935 2015 20965 2035
rect 20985 2015 21015 2035
rect 21035 2015 21065 2035
rect 21085 2015 21115 2035
rect 21135 2015 21165 2035
rect 21185 2015 21215 2035
rect 21235 2015 21265 2035
rect 21285 2015 21315 2035
rect 21335 2015 21365 2035
rect 21385 2015 21415 2035
rect 21435 2015 21465 2035
rect 21485 2015 21515 2035
rect 21535 2015 21565 2035
rect 21585 2015 21615 2035
rect 21635 2015 21665 2035
rect 21685 2015 21715 2035
rect 21735 2015 21765 2035
rect 21785 2015 21815 2035
rect 21835 2015 21865 2035
rect 21885 2015 21915 2035
rect 21935 2015 21965 2035
rect 21985 2015 22015 2035
rect 22035 2015 22065 2035
rect 22085 2015 22115 2035
rect 22135 2015 22165 2035
rect 22185 2015 22215 2035
rect 22235 2015 22265 2035
rect 22285 2015 22315 2035
rect 22335 2015 22365 2035
rect 22385 2015 22415 2035
rect 22435 2015 22465 2035
rect 22485 2015 22515 2035
rect 22535 2015 22565 2035
rect 22585 2015 22615 2035
rect 22635 2015 22665 2035
rect 22685 2015 22715 2035
rect 22735 2015 22765 2035
rect 22785 2015 22815 2035
rect 22835 2015 22865 2035
rect 22885 2015 22915 2035
rect 22935 2015 22965 2035
rect 22985 2015 23015 2035
rect 23035 2015 23065 2035
rect 23085 2015 23115 2035
rect 23135 2015 23165 2035
rect 23185 2015 23215 2035
rect 23235 2015 23265 2035
rect 23285 2015 23315 2035
rect 23335 2015 23365 2035
rect 23385 2015 23415 2035
rect 23435 2015 23465 2035
rect 23485 2015 23515 2035
rect 23535 2015 23565 2035
rect 23585 2015 23615 2035
rect 23635 2015 23665 2035
rect 23685 2015 23715 2035
rect 23735 2015 23765 2035
rect 23785 2015 23815 2035
rect 23835 2015 23865 2035
rect 23885 2015 23915 2035
rect 23935 2015 23965 2035
rect 23985 2015 24015 2035
rect 24035 2015 24065 2035
rect 24085 2015 24115 2035
rect 24135 2015 24165 2035
rect 24185 2015 24215 2035
rect 24235 2015 24265 2035
rect 24285 2015 24315 2035
rect 24335 2015 24365 2035
rect 24385 2015 24415 2035
rect 24435 2015 24465 2035
rect 24485 2015 24515 2035
rect 24535 2015 24565 2035
rect 24585 2015 24615 2035
rect 24635 2015 24665 2035
rect 24685 2015 24715 2035
rect 24735 2015 24765 2035
rect 24785 2015 24815 2035
rect 24835 2015 24865 2035
rect 24885 2015 24915 2035
rect 24935 2015 24965 2035
rect 24985 2015 25015 2035
rect 25035 2015 25065 2035
rect 25085 2015 25115 2035
rect 25135 2015 25165 2035
rect 25185 2015 25215 2035
rect 25235 2015 25265 2035
rect 25285 2015 25315 2035
rect 25335 2015 25365 2035
rect 25385 2015 25415 2035
rect 25435 2015 25465 2035
rect 25485 2015 25515 2035
rect 25535 2015 25565 2035
rect 25585 2015 25615 2035
rect 25635 2015 25665 2035
rect 25685 2015 25715 2035
rect 25735 2015 25765 2035
rect 25785 2015 25815 2035
rect 25835 2015 25865 2035
rect 25885 2015 25915 2035
rect 25935 2015 25965 2035
rect 25985 2015 26015 2035
rect 26035 2015 26065 2035
rect 26085 2015 26115 2035
rect 26135 2015 26165 2035
rect 26185 2015 26215 2035
rect 26235 2015 26265 2035
rect 26285 2015 26315 2035
rect 26335 2015 26365 2035
rect 26385 2015 26415 2035
rect 26435 2015 26465 2035
rect 26485 2015 26515 2035
rect 26535 2015 26565 2035
rect 26585 2015 26615 2035
rect 26635 2015 26665 2035
rect 26685 2015 26715 2035
rect 26735 2015 26765 2035
rect 26785 2015 26815 2035
rect 26835 2015 26865 2035
rect 26885 2015 26915 2035
rect 26935 2015 26965 2035
rect 26985 2015 27015 2035
rect 27035 2015 27065 2035
rect 27085 2015 27115 2035
rect 27135 2015 27165 2035
rect 27185 2015 27215 2035
rect 27235 2015 27265 2035
rect 27285 2015 27315 2035
rect 27335 2015 27365 2035
rect 27385 2015 27415 2035
rect 27435 2015 27465 2035
rect 27485 2015 27515 2035
rect 27535 2015 27565 2035
rect 27585 2015 27615 2035
rect 27635 2015 27665 2035
rect 27685 2015 27715 2035
rect 27735 2015 27765 2035
rect 27785 2015 27815 2035
rect 27835 2015 27865 2035
rect 27885 2015 27915 2035
rect 27935 2015 27965 2035
rect 27985 2015 28015 2035
rect 28035 2015 28065 2035
rect 28085 2015 28115 2035
rect 28135 2015 28165 2035
rect 28185 2015 28215 2035
rect 28235 2015 28265 2035
rect 28285 2015 28315 2035
rect 28335 2015 28365 2035
rect 28385 2015 28415 2035
rect 28435 2015 28465 2035
rect 28485 2015 28515 2035
rect 28535 2015 28565 2035
rect 28585 2015 28615 2035
rect 28635 2015 28665 2035
rect 28685 2015 28715 2035
rect 28735 2015 28765 2035
rect 28785 2015 28800 2035
rect -900 2000 28800 2015
rect -650 1685 28800 1700
rect -650 1665 -635 1685
rect -615 1665 -585 1685
rect -565 1665 -535 1685
rect -515 1665 -485 1685
rect -465 1665 -435 1685
rect -415 1665 -385 1685
rect -365 1665 -335 1685
rect -315 1665 -285 1685
rect -265 1665 -235 1685
rect -215 1665 -185 1685
rect -165 1665 -135 1685
rect -115 1665 -85 1685
rect -65 1665 -35 1685
rect -15 1665 15 1685
rect 35 1665 65 1685
rect 85 1665 115 1685
rect 135 1665 165 1685
rect 185 1665 215 1685
rect 235 1665 265 1685
rect 285 1665 315 1685
rect 335 1665 365 1685
rect 385 1665 415 1685
rect 435 1665 465 1685
rect 485 1665 515 1685
rect 535 1665 565 1685
rect 585 1665 615 1685
rect 635 1665 665 1685
rect 685 1665 715 1685
rect 735 1665 765 1685
rect 785 1665 815 1685
rect 835 1665 865 1685
rect 885 1665 915 1685
rect 935 1665 965 1685
rect 985 1665 1015 1685
rect 1035 1665 1065 1685
rect 1085 1665 1115 1685
rect 1135 1665 1165 1685
rect 1185 1665 1215 1685
rect 1235 1665 1265 1685
rect 1285 1665 1315 1685
rect 1335 1665 1365 1685
rect 1385 1665 1415 1685
rect 1435 1665 1465 1685
rect 1485 1665 1515 1685
rect 1535 1665 1565 1685
rect 1585 1665 1615 1685
rect 1635 1665 1665 1685
rect 1685 1665 1715 1685
rect 1735 1665 1765 1685
rect 1785 1665 1815 1685
rect 1835 1665 1865 1685
rect 1885 1665 1915 1685
rect 1935 1665 1965 1685
rect 1985 1665 2015 1685
rect 2035 1665 2065 1685
rect 2085 1665 2115 1685
rect 2135 1665 2165 1685
rect 2185 1665 2215 1685
rect 2235 1665 2265 1685
rect 2285 1665 2315 1685
rect 2335 1665 2365 1685
rect 2385 1665 2415 1685
rect 2435 1665 2465 1685
rect 2485 1665 2515 1685
rect 2535 1665 2565 1685
rect 2585 1665 2615 1685
rect 2635 1665 2665 1685
rect 2685 1665 2715 1685
rect 2735 1665 2765 1685
rect 2785 1665 2815 1685
rect 2835 1665 2865 1685
rect 2885 1665 2915 1685
rect 2935 1665 2965 1685
rect 2985 1665 3015 1685
rect 3035 1665 3065 1685
rect 3085 1665 3115 1685
rect 3135 1665 3165 1685
rect 3185 1665 3215 1685
rect 3235 1665 3265 1685
rect 3285 1665 3315 1685
rect 3335 1665 3365 1685
rect 3385 1665 3415 1685
rect 3435 1665 3465 1685
rect 3485 1665 3515 1685
rect 3535 1665 3565 1685
rect 3585 1665 3615 1685
rect 3635 1665 3665 1685
rect 3685 1665 3715 1685
rect 3735 1665 3765 1685
rect 3785 1665 3815 1685
rect 3835 1665 3865 1685
rect 3885 1665 3915 1685
rect 3935 1665 3965 1685
rect 3985 1665 4015 1685
rect 4035 1665 4065 1685
rect 4085 1665 4115 1685
rect 4135 1665 4165 1685
rect 4185 1665 4215 1685
rect 4235 1665 4265 1685
rect 4285 1665 4315 1685
rect 4335 1665 4365 1685
rect 4385 1665 4415 1685
rect 4435 1665 4465 1685
rect 4485 1665 4515 1685
rect 4535 1665 4565 1685
rect 4585 1665 4615 1685
rect 4635 1665 4665 1685
rect 4685 1665 4715 1685
rect 4735 1665 4765 1685
rect 4785 1665 4815 1685
rect 4835 1665 4865 1685
rect 4885 1665 4915 1685
rect 4935 1665 4965 1685
rect 4985 1665 5015 1685
rect 5035 1665 5065 1685
rect 5085 1665 5115 1685
rect 5135 1665 5165 1685
rect 5185 1665 5215 1685
rect 5235 1665 5265 1685
rect 5285 1665 5315 1685
rect 5335 1665 5365 1685
rect 5385 1665 5415 1685
rect 5435 1665 5465 1685
rect 5485 1665 5515 1685
rect 5535 1665 5565 1685
rect 5585 1665 5615 1685
rect 5635 1665 5665 1685
rect 5685 1665 5715 1685
rect 5735 1665 5765 1685
rect 5785 1665 5815 1685
rect 5835 1665 5865 1685
rect 5885 1665 5915 1685
rect 5935 1665 5965 1685
rect 5985 1665 6015 1685
rect 6035 1665 6065 1685
rect 6085 1665 6115 1685
rect 6135 1665 6165 1685
rect 6185 1665 6215 1685
rect 6235 1665 6265 1685
rect 6285 1665 6315 1685
rect 6335 1665 6365 1685
rect 6385 1665 6415 1685
rect 6435 1665 6465 1685
rect 6485 1665 6515 1685
rect 6535 1665 6565 1685
rect 6585 1665 6615 1685
rect 6635 1665 6665 1685
rect 6685 1665 6715 1685
rect 6735 1665 6765 1685
rect 6785 1665 6815 1685
rect 6835 1665 6865 1685
rect 6885 1665 6915 1685
rect 6935 1665 6965 1685
rect 6985 1665 7015 1685
rect 7035 1665 7065 1685
rect 7085 1665 7115 1685
rect 7135 1665 7165 1685
rect 7185 1665 7215 1685
rect 7235 1665 7265 1685
rect 7285 1665 7315 1685
rect 7335 1665 7365 1685
rect 7385 1665 7415 1685
rect 7435 1665 7465 1685
rect 7485 1665 7515 1685
rect 7535 1665 7565 1685
rect 7585 1665 7615 1685
rect 7635 1665 7665 1685
rect 7685 1665 7715 1685
rect 7735 1665 7765 1685
rect 7785 1665 7815 1685
rect 7835 1665 7865 1685
rect 7885 1665 7915 1685
rect 7935 1665 7965 1685
rect 7985 1665 8015 1685
rect 8035 1665 8065 1685
rect 8085 1665 8115 1685
rect 8135 1665 8165 1685
rect 8185 1665 8215 1685
rect 8235 1665 8265 1685
rect 8285 1665 8315 1685
rect 8335 1665 8365 1685
rect 8385 1665 8415 1685
rect 8435 1665 8465 1685
rect 8485 1665 8515 1685
rect 8535 1665 8565 1685
rect 8585 1665 8615 1685
rect 8635 1665 8665 1685
rect 8685 1665 8715 1685
rect 8735 1665 8765 1685
rect 8785 1665 8815 1685
rect 8835 1665 8865 1685
rect 8885 1665 8915 1685
rect 8935 1665 8965 1685
rect 8985 1665 9015 1685
rect 9035 1665 9065 1685
rect 9085 1665 9115 1685
rect 9135 1665 9165 1685
rect 9185 1665 9215 1685
rect 9235 1665 9265 1685
rect 9285 1665 9315 1685
rect 9335 1665 9365 1685
rect 9385 1665 9415 1685
rect 9435 1665 9465 1685
rect 9485 1665 9515 1685
rect 9535 1665 9565 1685
rect 9585 1665 9615 1685
rect 9635 1665 9665 1685
rect 9685 1665 9715 1685
rect 9735 1665 9765 1685
rect 9785 1665 9815 1685
rect 9835 1665 9865 1685
rect 9885 1665 9915 1685
rect 9935 1665 9965 1685
rect 9985 1665 10015 1685
rect 10035 1665 10065 1685
rect 10085 1665 10115 1685
rect 10135 1665 10165 1685
rect 10185 1665 10215 1685
rect 10235 1665 10265 1685
rect 10285 1665 10315 1685
rect 10335 1665 10365 1685
rect 10385 1665 10415 1685
rect 10435 1665 10465 1685
rect 10485 1665 10515 1685
rect 10535 1665 10565 1685
rect 10585 1665 10615 1685
rect 10635 1665 10665 1685
rect 10685 1665 10715 1685
rect 10735 1665 10765 1685
rect 10785 1665 10815 1685
rect 10835 1665 10865 1685
rect 10885 1665 10915 1685
rect 10935 1665 10965 1685
rect 10985 1665 11015 1685
rect 11035 1665 11065 1685
rect 11085 1665 11115 1685
rect 11135 1665 11165 1685
rect 11185 1665 11215 1685
rect 11235 1665 11265 1685
rect 11285 1665 11315 1685
rect 11335 1665 11365 1685
rect 11385 1665 11415 1685
rect 11435 1665 11465 1685
rect 11485 1665 11515 1685
rect 11535 1665 11565 1685
rect 11585 1665 11615 1685
rect 11635 1665 11665 1685
rect 11685 1665 11715 1685
rect 11735 1665 11765 1685
rect 11785 1665 11815 1685
rect 11835 1665 11865 1685
rect 11885 1665 11915 1685
rect 11935 1665 11965 1685
rect 11985 1665 12015 1685
rect 12035 1665 12065 1685
rect 12085 1665 12115 1685
rect 12135 1665 12165 1685
rect 12185 1665 12215 1685
rect 12235 1665 12265 1685
rect 12285 1665 12315 1685
rect 12335 1665 12365 1685
rect 12385 1665 12415 1685
rect 12435 1665 12465 1685
rect 12485 1665 12515 1685
rect 12535 1665 12565 1685
rect 12585 1665 12615 1685
rect 12635 1665 12665 1685
rect 12685 1665 12715 1685
rect 12735 1665 12765 1685
rect 12785 1665 12815 1685
rect 12835 1665 12865 1685
rect 12885 1665 12915 1685
rect 12935 1665 12965 1685
rect 12985 1665 13015 1685
rect 13035 1665 13065 1685
rect 13085 1665 13115 1685
rect 13135 1665 13165 1685
rect 13185 1665 13215 1685
rect 13235 1665 13265 1685
rect 13285 1665 13315 1685
rect 13335 1665 13365 1685
rect 13385 1665 13415 1685
rect 13435 1665 13465 1685
rect 13485 1665 13515 1685
rect 13535 1665 13565 1685
rect 13585 1665 13615 1685
rect 13635 1665 13665 1685
rect 13685 1665 13715 1685
rect 13735 1665 13765 1685
rect 13785 1665 13815 1685
rect 13835 1665 13865 1685
rect 13885 1665 13915 1685
rect 13935 1665 13965 1685
rect 13985 1665 14015 1685
rect 14035 1665 14065 1685
rect 14085 1665 14115 1685
rect 14135 1665 14165 1685
rect 14185 1665 14215 1685
rect 14235 1665 14265 1685
rect 14285 1665 14315 1685
rect 14335 1665 14365 1685
rect 14385 1665 14415 1685
rect 14435 1665 14465 1685
rect 14485 1665 14515 1685
rect 14535 1665 14565 1685
rect 14585 1665 14615 1685
rect 14635 1665 14665 1685
rect 14685 1665 14715 1685
rect 14735 1665 14765 1685
rect 14785 1665 14815 1685
rect 14835 1665 14865 1685
rect 14885 1665 14915 1685
rect 14935 1665 14965 1685
rect 14985 1665 15015 1685
rect 15035 1665 15065 1685
rect 15085 1665 15115 1685
rect 15135 1665 15165 1685
rect 15185 1665 15215 1685
rect 15235 1665 15265 1685
rect 15285 1665 15315 1685
rect 15335 1665 15365 1685
rect 15385 1665 15415 1685
rect 15435 1665 15465 1685
rect 15485 1665 15515 1685
rect 15535 1665 15565 1685
rect 15585 1665 15615 1685
rect 15635 1665 15665 1685
rect 15685 1665 15715 1685
rect 15735 1665 15765 1685
rect 15785 1665 15815 1685
rect 15835 1665 15865 1685
rect 15885 1665 15915 1685
rect 15935 1665 15965 1685
rect 15985 1665 16015 1685
rect 16035 1665 16065 1685
rect 16085 1665 16115 1685
rect 16135 1665 16165 1685
rect 16185 1665 16215 1685
rect 16235 1665 16265 1685
rect 16285 1665 16315 1685
rect 16335 1665 16365 1685
rect 16385 1665 16415 1685
rect 16435 1665 16465 1685
rect 16485 1665 16515 1685
rect 16535 1665 16565 1685
rect 16585 1665 16615 1685
rect 16635 1665 16665 1685
rect 16685 1665 16715 1685
rect 16735 1665 16765 1685
rect 16785 1665 16815 1685
rect 16835 1665 16865 1685
rect 16885 1665 16915 1685
rect 16935 1665 16965 1685
rect 16985 1665 17015 1685
rect 17035 1665 17065 1685
rect 17085 1665 17115 1685
rect 17135 1665 17165 1685
rect 17185 1665 17215 1685
rect 17235 1665 17265 1685
rect 17285 1665 17315 1685
rect 17335 1665 17365 1685
rect 17385 1665 17415 1685
rect 17435 1665 17465 1685
rect 17485 1665 17515 1685
rect 17535 1665 17565 1685
rect 17585 1665 17615 1685
rect 17635 1665 17665 1685
rect 17685 1665 17715 1685
rect 17735 1665 17765 1685
rect 17785 1665 17815 1685
rect 17835 1665 17865 1685
rect 17885 1665 17915 1685
rect 17935 1665 17965 1685
rect 17985 1665 18015 1685
rect 18035 1665 18065 1685
rect 18085 1665 18115 1685
rect 18135 1665 18165 1685
rect 18185 1665 18215 1685
rect 18235 1665 18265 1685
rect 18285 1665 18315 1685
rect 18335 1665 18365 1685
rect 18385 1665 18415 1685
rect 18435 1665 18465 1685
rect 18485 1665 18515 1685
rect 18535 1665 18565 1685
rect 18585 1665 18615 1685
rect 18635 1665 18665 1685
rect 18685 1665 18715 1685
rect 18735 1665 18765 1685
rect 18785 1665 18815 1685
rect 18835 1665 18865 1685
rect 18885 1665 18915 1685
rect 18935 1665 18965 1685
rect 18985 1665 19015 1685
rect 19035 1665 19065 1685
rect 19085 1665 19115 1685
rect 19135 1665 19165 1685
rect 19185 1665 19215 1685
rect 19235 1665 19265 1685
rect 19285 1665 19315 1685
rect 19335 1665 19365 1685
rect 19385 1665 19415 1685
rect 19435 1665 19465 1685
rect 19485 1665 19515 1685
rect 19535 1665 19565 1685
rect 19585 1665 19615 1685
rect 19635 1665 19665 1685
rect 19685 1665 19715 1685
rect 19735 1665 19765 1685
rect 19785 1665 19815 1685
rect 19835 1665 19865 1685
rect 19885 1665 19915 1685
rect 19935 1665 19965 1685
rect 19985 1665 20015 1685
rect 20035 1665 20065 1685
rect 20085 1665 20115 1685
rect 20135 1665 20165 1685
rect 20185 1665 20215 1685
rect 20235 1665 20265 1685
rect 20285 1665 20315 1685
rect 20335 1665 20365 1685
rect 20385 1665 20415 1685
rect 20435 1665 20465 1685
rect 20485 1665 20515 1685
rect 20535 1665 20565 1685
rect 20585 1665 20615 1685
rect 20635 1665 20665 1685
rect 20685 1665 20715 1685
rect 20735 1665 20765 1685
rect 20785 1665 20815 1685
rect 20835 1665 20865 1685
rect 20885 1665 20915 1685
rect 20935 1665 20965 1685
rect 20985 1665 21015 1685
rect 21035 1665 21065 1685
rect 21085 1665 21115 1685
rect 21135 1665 21165 1685
rect 21185 1665 21215 1685
rect 21235 1665 21265 1685
rect 21285 1665 21315 1685
rect 21335 1665 21365 1685
rect 21385 1665 21415 1685
rect 21435 1665 21465 1685
rect 21485 1665 21515 1685
rect 21535 1665 21565 1685
rect 21585 1665 21615 1685
rect 21635 1665 21665 1685
rect 21685 1665 21715 1685
rect 21735 1665 21765 1685
rect 21785 1665 21815 1685
rect 21835 1665 21865 1685
rect 21885 1665 21915 1685
rect 21935 1665 21965 1685
rect 21985 1665 22015 1685
rect 22035 1665 22065 1685
rect 22085 1665 22115 1685
rect 22135 1665 22165 1685
rect 22185 1665 22215 1685
rect 22235 1665 22265 1685
rect 22285 1665 22315 1685
rect 22335 1665 22365 1685
rect 22385 1665 22415 1685
rect 22435 1665 22465 1685
rect 22485 1665 22515 1685
rect 22535 1665 22565 1685
rect 22585 1665 22615 1685
rect 22635 1665 22665 1685
rect 22685 1665 22715 1685
rect 22735 1665 22765 1685
rect 22785 1665 22815 1685
rect 22835 1665 22865 1685
rect 22885 1665 22915 1685
rect 22935 1665 22965 1685
rect 22985 1665 23015 1685
rect 23035 1665 23065 1685
rect 23085 1665 23115 1685
rect 23135 1665 23165 1685
rect 23185 1665 23215 1685
rect 23235 1665 23265 1685
rect 23285 1665 23315 1685
rect 23335 1665 23365 1685
rect 23385 1665 23415 1685
rect 23435 1665 23465 1685
rect 23485 1665 23515 1685
rect 23535 1665 23565 1685
rect 23585 1665 23615 1685
rect 23635 1665 23665 1685
rect 23685 1665 23715 1685
rect 23735 1665 23765 1685
rect 23785 1665 23815 1685
rect 23835 1665 23865 1685
rect 23885 1665 23915 1685
rect 23935 1665 23965 1685
rect 23985 1665 24015 1685
rect 24035 1665 24065 1685
rect 24085 1665 24115 1685
rect 24135 1665 24165 1685
rect 24185 1665 24215 1685
rect 24235 1665 24265 1685
rect 24285 1665 24315 1685
rect 24335 1665 24365 1685
rect 24385 1665 24415 1685
rect 24435 1665 24465 1685
rect 24485 1665 24515 1685
rect 24535 1665 24565 1685
rect 24585 1665 24615 1685
rect 24635 1665 24665 1685
rect 24685 1665 24715 1685
rect 24735 1665 24765 1685
rect 24785 1665 24815 1685
rect 24835 1665 24865 1685
rect 24885 1665 24915 1685
rect 24935 1665 24965 1685
rect 24985 1665 25015 1685
rect 25035 1665 25065 1685
rect 25085 1665 25115 1685
rect 25135 1665 25165 1685
rect 25185 1665 25215 1685
rect 25235 1665 25265 1685
rect 25285 1665 25315 1685
rect 25335 1665 25365 1685
rect 25385 1665 25415 1685
rect 25435 1665 25465 1685
rect 25485 1665 25515 1685
rect 25535 1665 25565 1685
rect 25585 1665 25615 1685
rect 25635 1665 25665 1685
rect 25685 1665 25715 1685
rect 25735 1665 25765 1685
rect 25785 1665 25815 1685
rect 25835 1665 25865 1685
rect 25885 1665 25915 1685
rect 25935 1665 25965 1685
rect 25985 1665 26015 1685
rect 26035 1665 26065 1685
rect 26085 1665 26115 1685
rect 26135 1665 26165 1685
rect 26185 1665 26215 1685
rect 26235 1665 26265 1685
rect 26285 1665 26315 1685
rect 26335 1665 26365 1685
rect 26385 1665 26415 1685
rect 26435 1665 26465 1685
rect 26485 1665 26515 1685
rect 26535 1665 26565 1685
rect 26585 1665 26615 1685
rect 26635 1665 26665 1685
rect 26685 1665 26715 1685
rect 26735 1665 26765 1685
rect 26785 1665 26815 1685
rect 26835 1665 26865 1685
rect 26885 1665 26915 1685
rect 26935 1665 26965 1685
rect 26985 1665 27015 1685
rect 27035 1665 27065 1685
rect 27085 1665 27115 1685
rect 27135 1665 27165 1685
rect 27185 1665 27215 1685
rect 27235 1665 27265 1685
rect 27285 1665 27315 1685
rect 27335 1665 27365 1685
rect 27385 1665 27415 1685
rect 27435 1665 27465 1685
rect 27485 1665 27515 1685
rect 27535 1665 27565 1685
rect 27585 1665 27615 1685
rect 27635 1665 27665 1685
rect 27685 1665 27715 1685
rect 27735 1665 27765 1685
rect 27785 1665 27815 1685
rect 27835 1665 27865 1685
rect 27885 1665 27915 1685
rect 27935 1665 27965 1685
rect 27985 1665 28015 1685
rect 28035 1665 28065 1685
rect 28085 1665 28115 1685
rect 28135 1665 28165 1685
rect 28185 1665 28215 1685
rect 28235 1665 28265 1685
rect 28285 1665 28315 1685
rect 28335 1665 28365 1685
rect 28385 1665 28415 1685
rect 28435 1665 28465 1685
rect 28485 1665 28515 1685
rect 28535 1665 28565 1685
rect 28585 1665 28615 1685
rect 28635 1665 28665 1685
rect 28685 1665 28715 1685
rect 28735 1665 28765 1685
rect 28785 1665 28800 1685
rect -650 1650 28800 1665
rect -650 -15 28800 0
rect -650 -35 -635 -15
rect -615 -35 -585 -15
rect -565 -35 -535 -15
rect -515 -35 -485 -15
rect -465 -35 -435 -15
rect -415 -35 -385 -15
rect -365 -35 -335 -15
rect -315 -35 -285 -15
rect -265 -35 -235 -15
rect -215 -35 -185 -15
rect -165 -35 -135 -15
rect -115 -35 -85 -15
rect -65 -35 -35 -15
rect -15 -35 15 -15
rect 35 -35 65 -15
rect 85 -35 115 -15
rect 135 -35 165 -15
rect 185 -35 215 -15
rect 235 -35 265 -15
rect 285 -35 315 -15
rect 335 -35 365 -15
rect 385 -35 415 -15
rect 435 -35 465 -15
rect 485 -35 515 -15
rect 535 -35 565 -15
rect 585 -35 615 -15
rect 635 -35 665 -15
rect 685 -35 715 -15
rect 735 -35 765 -15
rect 785 -35 815 -15
rect 835 -35 865 -15
rect 885 -35 915 -15
rect 935 -35 965 -15
rect 985 -35 1015 -15
rect 1035 -35 1065 -15
rect 1085 -35 1115 -15
rect 1135 -35 1165 -15
rect 1185 -35 1215 -15
rect 1235 -35 1265 -15
rect 1285 -35 1315 -15
rect 1335 -35 1365 -15
rect 1385 -35 1415 -15
rect 1435 -35 1465 -15
rect 1485 -35 1515 -15
rect 1535 -35 1565 -15
rect 1585 -35 1615 -15
rect 1635 -35 1665 -15
rect 1685 -35 1715 -15
rect 1735 -35 1765 -15
rect 1785 -35 1815 -15
rect 1835 -35 1865 -15
rect 1885 -35 1915 -15
rect 1935 -35 1965 -15
rect 1985 -35 2015 -15
rect 2035 -35 2065 -15
rect 2085 -35 2115 -15
rect 2135 -35 2165 -15
rect 2185 -35 2215 -15
rect 2235 -35 2265 -15
rect 2285 -35 2315 -15
rect 2335 -35 2365 -15
rect 2385 -35 2415 -15
rect 2435 -35 2465 -15
rect 2485 -35 2515 -15
rect 2535 -35 2565 -15
rect 2585 -35 2615 -15
rect 2635 -35 2665 -15
rect 2685 -35 2715 -15
rect 2735 -35 2765 -15
rect 2785 -35 2815 -15
rect 2835 -35 2865 -15
rect 2885 -35 2915 -15
rect 2935 -35 2965 -15
rect 2985 -35 3015 -15
rect 3035 -35 3065 -15
rect 3085 -35 3115 -15
rect 3135 -35 3165 -15
rect 3185 -35 3215 -15
rect 3235 -35 3265 -15
rect 3285 -35 3315 -15
rect 3335 -35 3365 -15
rect 3385 -35 3415 -15
rect 3435 -35 3465 -15
rect 3485 -35 3515 -15
rect 3535 -35 3565 -15
rect 3585 -35 3615 -15
rect 3635 -35 3665 -15
rect 3685 -35 3715 -15
rect 3735 -35 3765 -15
rect 3785 -35 3815 -15
rect 3835 -35 3865 -15
rect 3885 -35 3915 -15
rect 3935 -35 3965 -15
rect 3985 -35 4015 -15
rect 4035 -35 4065 -15
rect 4085 -35 4115 -15
rect 4135 -35 4165 -15
rect 4185 -35 4215 -15
rect 4235 -35 4265 -15
rect 4285 -35 4315 -15
rect 4335 -35 4365 -15
rect 4385 -35 4415 -15
rect 4435 -35 4465 -15
rect 4485 -35 4515 -15
rect 4535 -35 4565 -15
rect 4585 -35 4615 -15
rect 4635 -35 4665 -15
rect 4685 -35 4715 -15
rect 4735 -35 4765 -15
rect 4785 -35 4815 -15
rect 4835 -35 4865 -15
rect 4885 -35 4915 -15
rect 4935 -35 4965 -15
rect 4985 -35 5015 -15
rect 5035 -35 5065 -15
rect 5085 -35 5115 -15
rect 5135 -35 5165 -15
rect 5185 -35 5215 -15
rect 5235 -35 5265 -15
rect 5285 -35 5315 -15
rect 5335 -35 5365 -15
rect 5385 -35 5415 -15
rect 5435 -35 5465 -15
rect 5485 -35 5515 -15
rect 5535 -35 5565 -15
rect 5585 -35 5615 -15
rect 5635 -35 5665 -15
rect 5685 -35 5715 -15
rect 5735 -35 5765 -15
rect 5785 -35 5815 -15
rect 5835 -35 5865 -15
rect 5885 -35 5915 -15
rect 5935 -35 5965 -15
rect 5985 -35 6015 -15
rect 6035 -35 6065 -15
rect 6085 -35 6115 -15
rect 6135 -35 6165 -15
rect 6185 -35 6215 -15
rect 6235 -35 6265 -15
rect 6285 -35 6315 -15
rect 6335 -35 6365 -15
rect 6385 -35 6415 -15
rect 6435 -35 6465 -15
rect 6485 -35 6515 -15
rect 6535 -35 6565 -15
rect 6585 -35 6615 -15
rect 6635 -35 6665 -15
rect 6685 -35 6715 -15
rect 6735 -35 6765 -15
rect 6785 -35 6815 -15
rect 6835 -35 6865 -15
rect 6885 -35 6915 -15
rect 6935 -35 6965 -15
rect 6985 -35 7015 -15
rect 7035 -35 7065 -15
rect 7085 -35 7115 -15
rect 7135 -35 7165 -15
rect 7185 -35 7215 -15
rect 7235 -35 7265 -15
rect 7285 -35 7315 -15
rect 7335 -35 7365 -15
rect 7385 -35 7415 -15
rect 7435 -35 7465 -15
rect 7485 -35 7515 -15
rect 7535 -35 7565 -15
rect 7585 -35 7615 -15
rect 7635 -35 7665 -15
rect 7685 -35 7715 -15
rect 7735 -35 7765 -15
rect 7785 -35 7815 -15
rect 7835 -35 7865 -15
rect 7885 -35 7915 -15
rect 7935 -35 7965 -15
rect 7985 -35 8015 -15
rect 8035 -35 8065 -15
rect 8085 -35 8115 -15
rect 8135 -35 8165 -15
rect 8185 -35 8215 -15
rect 8235 -35 8265 -15
rect 8285 -35 8315 -15
rect 8335 -35 8365 -15
rect 8385 -35 8415 -15
rect 8435 -35 8465 -15
rect 8485 -35 8515 -15
rect 8535 -35 8565 -15
rect 8585 -35 8615 -15
rect 8635 -35 8665 -15
rect 8685 -35 8715 -15
rect 8735 -35 8765 -15
rect 8785 -35 8815 -15
rect 8835 -35 8865 -15
rect 8885 -35 8915 -15
rect 8935 -35 8965 -15
rect 8985 -35 9015 -15
rect 9035 -35 9065 -15
rect 9085 -35 9115 -15
rect 9135 -35 9165 -15
rect 9185 -35 9215 -15
rect 9235 -35 9265 -15
rect 9285 -35 9315 -15
rect 9335 -35 9365 -15
rect 9385 -35 9415 -15
rect 9435 -35 9465 -15
rect 9485 -35 9515 -15
rect 9535 -35 9565 -15
rect 9585 -35 9615 -15
rect 9635 -35 9665 -15
rect 9685 -35 9715 -15
rect 9735 -35 9765 -15
rect 9785 -35 9815 -15
rect 9835 -35 9865 -15
rect 9885 -35 9915 -15
rect 9935 -35 9965 -15
rect 9985 -35 10015 -15
rect 10035 -35 10065 -15
rect 10085 -35 10115 -15
rect 10135 -35 10165 -15
rect 10185 -35 10215 -15
rect 10235 -35 10265 -15
rect 10285 -35 10315 -15
rect 10335 -35 10365 -15
rect 10385 -35 10415 -15
rect 10435 -35 10465 -15
rect 10485 -35 10515 -15
rect 10535 -35 10565 -15
rect 10585 -35 10615 -15
rect 10635 -35 10665 -15
rect 10685 -35 10715 -15
rect 10735 -35 10765 -15
rect 10785 -35 10815 -15
rect 10835 -35 10865 -15
rect 10885 -35 10915 -15
rect 10935 -35 10965 -15
rect 10985 -35 11015 -15
rect 11035 -35 11065 -15
rect 11085 -35 11115 -15
rect 11135 -35 11165 -15
rect 11185 -35 11215 -15
rect 11235 -35 11265 -15
rect 11285 -35 11315 -15
rect 11335 -35 11365 -15
rect 11385 -35 11415 -15
rect 11435 -35 11465 -15
rect 11485 -35 11515 -15
rect 11535 -35 11565 -15
rect 11585 -35 11615 -15
rect 11635 -35 11665 -15
rect 11685 -35 11715 -15
rect 11735 -35 11765 -15
rect 11785 -35 11815 -15
rect 11835 -35 11865 -15
rect 11885 -35 11915 -15
rect 11935 -35 11965 -15
rect 11985 -35 12015 -15
rect 12035 -35 12065 -15
rect 12085 -35 12115 -15
rect 12135 -35 12165 -15
rect 12185 -35 12215 -15
rect 12235 -35 12265 -15
rect 12285 -35 12315 -15
rect 12335 -35 12365 -15
rect 12385 -35 12415 -15
rect 12435 -35 12465 -15
rect 12485 -35 12515 -15
rect 12535 -35 12565 -15
rect 12585 -35 12615 -15
rect 12635 -35 12665 -15
rect 12685 -35 12715 -15
rect 12735 -35 12765 -15
rect 12785 -35 12815 -15
rect 12835 -35 12865 -15
rect 12885 -35 12915 -15
rect 12935 -35 12965 -15
rect 12985 -35 13015 -15
rect 13035 -35 13065 -15
rect 13085 -35 13115 -15
rect 13135 -35 13165 -15
rect 13185 -35 13215 -15
rect 13235 -35 13265 -15
rect 13285 -35 13315 -15
rect 13335 -35 13365 -15
rect 13385 -35 13415 -15
rect 13435 -35 13465 -15
rect 13485 -35 13515 -15
rect 13535 -35 13565 -15
rect 13585 -35 13615 -15
rect 13635 -35 13665 -15
rect 13685 -35 13715 -15
rect 13735 -35 13765 -15
rect 13785 -35 13815 -15
rect 13835 -35 13865 -15
rect 13885 -35 13915 -15
rect 13935 -35 13965 -15
rect 13985 -35 14015 -15
rect 14035 -35 14065 -15
rect 14085 -35 14115 -15
rect 14135 -35 14165 -15
rect 14185 -35 14215 -15
rect 14235 -35 14265 -15
rect 14285 -35 14315 -15
rect 14335 -35 14365 -15
rect 14385 -35 14415 -15
rect 14435 -35 14465 -15
rect 14485 -35 14515 -15
rect 14535 -35 14565 -15
rect 14585 -35 14615 -15
rect 14635 -35 14665 -15
rect 14685 -35 14715 -15
rect 14735 -35 14765 -15
rect 14785 -35 14815 -15
rect 14835 -35 14865 -15
rect 14885 -35 14915 -15
rect 14935 -35 14965 -15
rect 14985 -35 15015 -15
rect 15035 -35 15065 -15
rect 15085 -35 15115 -15
rect 15135 -35 15165 -15
rect 15185 -35 15215 -15
rect 15235 -35 15265 -15
rect 15285 -35 15315 -15
rect 15335 -35 15365 -15
rect 15385 -35 15415 -15
rect 15435 -35 15465 -15
rect 15485 -35 15515 -15
rect 15535 -35 15565 -15
rect 15585 -35 15615 -15
rect 15635 -35 15665 -15
rect 15685 -35 15715 -15
rect 15735 -35 15765 -15
rect 15785 -35 15815 -15
rect 15835 -35 15865 -15
rect 15885 -35 15915 -15
rect 15935 -35 15965 -15
rect 15985 -35 16015 -15
rect 16035 -35 16065 -15
rect 16085 -35 16115 -15
rect 16135 -35 16165 -15
rect 16185 -35 16215 -15
rect 16235 -35 16265 -15
rect 16285 -35 16315 -15
rect 16335 -35 16365 -15
rect 16385 -35 16415 -15
rect 16435 -35 16465 -15
rect 16485 -35 16515 -15
rect 16535 -35 16565 -15
rect 16585 -35 16615 -15
rect 16635 -35 16665 -15
rect 16685 -35 16715 -15
rect 16735 -35 16765 -15
rect 16785 -35 16815 -15
rect 16835 -35 16865 -15
rect 16885 -35 16915 -15
rect 16935 -35 16965 -15
rect 16985 -35 17015 -15
rect 17035 -35 17065 -15
rect 17085 -35 17115 -15
rect 17135 -35 17165 -15
rect 17185 -35 17215 -15
rect 17235 -35 17265 -15
rect 17285 -35 17315 -15
rect 17335 -35 17365 -15
rect 17385 -35 17415 -15
rect 17435 -35 17465 -15
rect 17485 -35 17515 -15
rect 17535 -35 17565 -15
rect 17585 -35 17615 -15
rect 17635 -35 17665 -15
rect 17685 -35 17715 -15
rect 17735 -35 17765 -15
rect 17785 -35 17815 -15
rect 17835 -35 17865 -15
rect 17885 -35 17915 -15
rect 17935 -35 17965 -15
rect 17985 -35 18015 -15
rect 18035 -35 18065 -15
rect 18085 -35 18115 -15
rect 18135 -35 18165 -15
rect 18185 -35 18215 -15
rect 18235 -35 18265 -15
rect 18285 -35 18315 -15
rect 18335 -35 18365 -15
rect 18385 -35 18415 -15
rect 18435 -35 18465 -15
rect 18485 -35 18515 -15
rect 18535 -35 18565 -15
rect 18585 -35 18615 -15
rect 18635 -35 18665 -15
rect 18685 -35 18715 -15
rect 18735 -35 18765 -15
rect 18785 -35 18815 -15
rect 18835 -35 18865 -15
rect 18885 -35 18915 -15
rect 18935 -35 18965 -15
rect 18985 -35 19015 -15
rect 19035 -35 19065 -15
rect 19085 -35 19115 -15
rect 19135 -35 19165 -15
rect 19185 -35 19215 -15
rect 19235 -35 19265 -15
rect 19285 -35 19315 -15
rect 19335 -35 19365 -15
rect 19385 -35 19415 -15
rect 19435 -35 19465 -15
rect 19485 -35 19515 -15
rect 19535 -35 19565 -15
rect 19585 -35 19615 -15
rect 19635 -35 19665 -15
rect 19685 -35 19715 -15
rect 19735 -35 19765 -15
rect 19785 -35 19815 -15
rect 19835 -35 19865 -15
rect 19885 -35 19915 -15
rect 19935 -35 19965 -15
rect 19985 -35 20015 -15
rect 20035 -35 20065 -15
rect 20085 -35 20115 -15
rect 20135 -35 20165 -15
rect 20185 -35 20215 -15
rect 20235 -35 20265 -15
rect 20285 -35 20315 -15
rect 20335 -35 20365 -15
rect 20385 -35 20415 -15
rect 20435 -35 20465 -15
rect 20485 -35 20515 -15
rect 20535 -35 20565 -15
rect 20585 -35 20615 -15
rect 20635 -35 20665 -15
rect 20685 -35 20715 -15
rect 20735 -35 20765 -15
rect 20785 -35 20815 -15
rect 20835 -35 20865 -15
rect 20885 -35 20915 -15
rect 20935 -35 20965 -15
rect 20985 -35 21015 -15
rect 21035 -35 21065 -15
rect 21085 -35 21115 -15
rect 21135 -35 21165 -15
rect 21185 -35 21215 -15
rect 21235 -35 21265 -15
rect 21285 -35 21315 -15
rect 21335 -35 21365 -15
rect 21385 -35 21415 -15
rect 21435 -35 21465 -15
rect 21485 -35 21515 -15
rect 21535 -35 21565 -15
rect 21585 -35 21615 -15
rect 21635 -35 21665 -15
rect 21685 -35 21715 -15
rect 21735 -35 21765 -15
rect 21785 -35 21815 -15
rect 21835 -35 21865 -15
rect 21885 -35 21915 -15
rect 21935 -35 21965 -15
rect 21985 -35 22015 -15
rect 22035 -35 22065 -15
rect 22085 -35 22115 -15
rect 22135 -35 22165 -15
rect 22185 -35 22215 -15
rect 22235 -35 22265 -15
rect 22285 -35 22315 -15
rect 22335 -35 22365 -15
rect 22385 -35 22415 -15
rect 22435 -35 22465 -15
rect 22485 -35 22515 -15
rect 22535 -35 22565 -15
rect 22585 -35 22615 -15
rect 22635 -35 22665 -15
rect 22685 -35 22715 -15
rect 22735 -35 22765 -15
rect 22785 -35 22815 -15
rect 22835 -35 22865 -15
rect 22885 -35 22915 -15
rect 22935 -35 22965 -15
rect 22985 -35 23015 -15
rect 23035 -35 23065 -15
rect 23085 -35 23115 -15
rect 23135 -35 23165 -15
rect 23185 -35 23215 -15
rect 23235 -35 23265 -15
rect 23285 -35 23315 -15
rect 23335 -35 23365 -15
rect 23385 -35 23415 -15
rect 23435 -35 23465 -15
rect 23485 -35 23515 -15
rect 23535 -35 23565 -15
rect 23585 -35 23615 -15
rect 23635 -35 23665 -15
rect 23685 -35 23715 -15
rect 23735 -35 23765 -15
rect 23785 -35 23815 -15
rect 23835 -35 23865 -15
rect 23885 -35 23915 -15
rect 23935 -35 23965 -15
rect 23985 -35 24015 -15
rect 24035 -35 24065 -15
rect 24085 -35 24115 -15
rect 24135 -35 24165 -15
rect 24185 -35 24215 -15
rect 24235 -35 24265 -15
rect 24285 -35 24315 -15
rect 24335 -35 24365 -15
rect 24385 -35 24415 -15
rect 24435 -35 24465 -15
rect 24485 -35 24515 -15
rect 24535 -35 24565 -15
rect 24585 -35 24615 -15
rect 24635 -35 24665 -15
rect 24685 -35 24715 -15
rect 24735 -35 24765 -15
rect 24785 -35 24815 -15
rect 24835 -35 24865 -15
rect 24885 -35 24915 -15
rect 24935 -35 24965 -15
rect 24985 -35 25015 -15
rect 25035 -35 25065 -15
rect 25085 -35 25115 -15
rect 25135 -35 25165 -15
rect 25185 -35 25215 -15
rect 25235 -35 25265 -15
rect 25285 -35 25315 -15
rect 25335 -35 25365 -15
rect 25385 -35 25415 -15
rect 25435 -35 25465 -15
rect 25485 -35 25515 -15
rect 25535 -35 25565 -15
rect 25585 -35 25615 -15
rect 25635 -35 25665 -15
rect 25685 -35 25715 -15
rect 25735 -35 25765 -15
rect 25785 -35 25815 -15
rect 25835 -35 25865 -15
rect 25885 -35 25915 -15
rect 25935 -35 25965 -15
rect 25985 -35 26015 -15
rect 26035 -35 26065 -15
rect 26085 -35 26115 -15
rect 26135 -35 26165 -15
rect 26185 -35 26215 -15
rect 26235 -35 26265 -15
rect 26285 -35 26315 -15
rect 26335 -35 26365 -15
rect 26385 -35 26415 -15
rect 26435 -35 26465 -15
rect 26485 -35 26515 -15
rect 26535 -35 26565 -15
rect 26585 -35 26615 -15
rect 26635 -35 26665 -15
rect 26685 -35 26715 -15
rect 26735 -35 26765 -15
rect 26785 -35 26815 -15
rect 26835 -35 26865 -15
rect 26885 -35 26915 -15
rect 26935 -35 26965 -15
rect 26985 -35 27015 -15
rect 27035 -35 27065 -15
rect 27085 -35 27115 -15
rect 27135 -35 27165 -15
rect 27185 -35 27215 -15
rect 27235 -35 27265 -15
rect 27285 -35 27315 -15
rect 27335 -35 27365 -15
rect 27385 -35 27415 -15
rect 27435 -35 27465 -15
rect 27485 -35 27515 -15
rect 27535 -35 27565 -15
rect 27585 -35 27615 -15
rect 27635 -35 27665 -15
rect 27685 -35 27715 -15
rect 27735 -35 27765 -15
rect 27785 -35 27815 -15
rect 27835 -35 27865 -15
rect 27885 -35 27915 -15
rect 27935 -35 27965 -15
rect 27985 -35 28015 -15
rect 28035 -35 28065 -15
rect 28085 -35 28115 -15
rect 28135 -35 28165 -15
rect 28185 -35 28215 -15
rect 28235 -35 28265 -15
rect 28285 -35 28315 -15
rect 28335 -35 28365 -15
rect 28385 -35 28415 -15
rect 28435 -35 28465 -15
rect 28485 -35 28515 -15
rect 28535 -35 28565 -15
rect 28585 -35 28615 -15
rect 28635 -35 28665 -15
rect 28685 -35 28715 -15
rect 28735 -35 28765 -15
rect 28785 -35 28800 -15
rect -650 -50 28800 -35
rect -650 -1715 28800 -1700
rect -650 -1735 -635 -1715
rect -615 -1735 -585 -1715
rect -565 -1735 -535 -1715
rect -515 -1735 -485 -1715
rect -465 -1735 -435 -1715
rect -415 -1735 -385 -1715
rect -365 -1735 -335 -1715
rect -315 -1735 -285 -1715
rect -265 -1735 -235 -1715
rect -215 -1735 -185 -1715
rect -165 -1735 -135 -1715
rect -115 -1735 -85 -1715
rect -65 -1735 -35 -1715
rect -15 -1735 15 -1715
rect 35 -1735 65 -1715
rect 85 -1735 115 -1715
rect 135 -1735 165 -1715
rect 185 -1735 215 -1715
rect 235 -1735 265 -1715
rect 285 -1735 315 -1715
rect 335 -1735 365 -1715
rect 385 -1735 415 -1715
rect 435 -1735 465 -1715
rect 485 -1735 515 -1715
rect 535 -1735 565 -1715
rect 585 -1735 615 -1715
rect 635 -1735 665 -1715
rect 685 -1735 715 -1715
rect 735 -1735 765 -1715
rect 785 -1735 815 -1715
rect 835 -1735 865 -1715
rect 885 -1735 915 -1715
rect 935 -1735 965 -1715
rect 985 -1735 1015 -1715
rect 1035 -1735 1065 -1715
rect 1085 -1735 1115 -1715
rect 1135 -1735 1165 -1715
rect 1185 -1735 1215 -1715
rect 1235 -1735 1265 -1715
rect 1285 -1735 1315 -1715
rect 1335 -1735 1365 -1715
rect 1385 -1735 1415 -1715
rect 1435 -1735 1465 -1715
rect 1485 -1735 1515 -1715
rect 1535 -1735 1565 -1715
rect 1585 -1735 1615 -1715
rect 1635 -1735 1665 -1715
rect 1685 -1735 1715 -1715
rect 1735 -1735 1765 -1715
rect 1785 -1735 1815 -1715
rect 1835 -1735 1865 -1715
rect 1885 -1735 1915 -1715
rect 1935 -1735 1965 -1715
rect 1985 -1735 2015 -1715
rect 2035 -1735 2065 -1715
rect 2085 -1735 2115 -1715
rect 2135 -1735 2165 -1715
rect 2185 -1735 2215 -1715
rect 2235 -1735 2265 -1715
rect 2285 -1735 2315 -1715
rect 2335 -1735 2365 -1715
rect 2385 -1735 2415 -1715
rect 2435 -1735 2465 -1715
rect 2485 -1735 2515 -1715
rect 2535 -1735 2565 -1715
rect 2585 -1735 2615 -1715
rect 2635 -1735 2665 -1715
rect 2685 -1735 2715 -1715
rect 2735 -1735 2765 -1715
rect 2785 -1735 2815 -1715
rect 2835 -1735 2865 -1715
rect 2885 -1735 2915 -1715
rect 2935 -1735 2965 -1715
rect 2985 -1735 3015 -1715
rect 3035 -1735 3065 -1715
rect 3085 -1735 3115 -1715
rect 3135 -1735 3165 -1715
rect 3185 -1735 3215 -1715
rect 3235 -1735 3265 -1715
rect 3285 -1735 3315 -1715
rect 3335 -1735 3365 -1715
rect 3385 -1735 3415 -1715
rect 3435 -1735 3465 -1715
rect 3485 -1735 3515 -1715
rect 3535 -1735 3565 -1715
rect 3585 -1735 3615 -1715
rect 3635 -1735 3665 -1715
rect 3685 -1735 3715 -1715
rect 3735 -1735 3765 -1715
rect 3785 -1735 3815 -1715
rect 3835 -1735 3865 -1715
rect 3885 -1735 3915 -1715
rect 3935 -1735 3965 -1715
rect 3985 -1735 4015 -1715
rect 4035 -1735 4065 -1715
rect 4085 -1735 4115 -1715
rect 4135 -1735 4165 -1715
rect 4185 -1735 4215 -1715
rect 4235 -1735 4265 -1715
rect 4285 -1735 4315 -1715
rect 4335 -1735 4365 -1715
rect 4385 -1735 4415 -1715
rect 4435 -1735 4465 -1715
rect 4485 -1735 4515 -1715
rect 4535 -1735 4565 -1715
rect 4585 -1735 4615 -1715
rect 4635 -1735 4665 -1715
rect 4685 -1735 4715 -1715
rect 4735 -1735 4765 -1715
rect 4785 -1735 4815 -1715
rect 4835 -1735 4865 -1715
rect 4885 -1735 4915 -1715
rect 4935 -1735 4965 -1715
rect 4985 -1735 5015 -1715
rect 5035 -1735 5065 -1715
rect 5085 -1735 5115 -1715
rect 5135 -1735 5165 -1715
rect 5185 -1735 5215 -1715
rect 5235 -1735 5265 -1715
rect 5285 -1735 5315 -1715
rect 5335 -1735 5365 -1715
rect 5385 -1735 5415 -1715
rect 5435 -1735 5465 -1715
rect 5485 -1735 5515 -1715
rect 5535 -1735 5565 -1715
rect 5585 -1735 5615 -1715
rect 5635 -1735 5665 -1715
rect 5685 -1735 5715 -1715
rect 5735 -1735 5765 -1715
rect 5785 -1735 5815 -1715
rect 5835 -1735 5865 -1715
rect 5885 -1735 5915 -1715
rect 5935 -1735 5965 -1715
rect 5985 -1735 6015 -1715
rect 6035 -1735 6065 -1715
rect 6085 -1735 6115 -1715
rect 6135 -1735 6165 -1715
rect 6185 -1735 6215 -1715
rect 6235 -1735 6265 -1715
rect 6285 -1735 6315 -1715
rect 6335 -1735 6365 -1715
rect 6385 -1735 6415 -1715
rect 6435 -1735 6465 -1715
rect 6485 -1735 6515 -1715
rect 6535 -1735 6565 -1715
rect 6585 -1735 6615 -1715
rect 6635 -1735 6665 -1715
rect 6685 -1735 6715 -1715
rect 6735 -1735 6765 -1715
rect 6785 -1735 6815 -1715
rect 6835 -1735 6865 -1715
rect 6885 -1735 6915 -1715
rect 6935 -1735 6965 -1715
rect 6985 -1735 7015 -1715
rect 7035 -1735 7065 -1715
rect 7085 -1735 7115 -1715
rect 7135 -1735 7165 -1715
rect 7185 -1735 7215 -1715
rect 7235 -1735 7265 -1715
rect 7285 -1735 7315 -1715
rect 7335 -1735 7365 -1715
rect 7385 -1735 7415 -1715
rect 7435 -1735 7465 -1715
rect 7485 -1735 7515 -1715
rect 7535 -1735 7565 -1715
rect 7585 -1735 7615 -1715
rect 7635 -1735 7665 -1715
rect 7685 -1735 7715 -1715
rect 7735 -1735 7765 -1715
rect 7785 -1735 7815 -1715
rect 7835 -1735 7865 -1715
rect 7885 -1735 7915 -1715
rect 7935 -1735 7965 -1715
rect 7985 -1735 8015 -1715
rect 8035 -1735 8065 -1715
rect 8085 -1735 8115 -1715
rect 8135 -1735 8165 -1715
rect 8185 -1735 8215 -1715
rect 8235 -1735 8265 -1715
rect 8285 -1735 8315 -1715
rect 8335 -1735 8365 -1715
rect 8385 -1735 8415 -1715
rect 8435 -1735 8465 -1715
rect 8485 -1735 8515 -1715
rect 8535 -1735 8565 -1715
rect 8585 -1735 8615 -1715
rect 8635 -1735 8665 -1715
rect 8685 -1735 8715 -1715
rect 8735 -1735 8765 -1715
rect 8785 -1735 8815 -1715
rect 8835 -1735 8865 -1715
rect 8885 -1735 8915 -1715
rect 8935 -1735 8965 -1715
rect 8985 -1735 9015 -1715
rect 9035 -1735 9065 -1715
rect 9085 -1735 9115 -1715
rect 9135 -1735 9165 -1715
rect 9185 -1735 9215 -1715
rect 9235 -1735 9265 -1715
rect 9285 -1735 9315 -1715
rect 9335 -1735 9365 -1715
rect 9385 -1735 9415 -1715
rect 9435 -1735 9465 -1715
rect 9485 -1735 9515 -1715
rect 9535 -1735 9565 -1715
rect 9585 -1735 9615 -1715
rect 9635 -1735 9665 -1715
rect 9685 -1735 9715 -1715
rect 9735 -1735 9765 -1715
rect 9785 -1735 9815 -1715
rect 9835 -1735 9865 -1715
rect 9885 -1735 9915 -1715
rect 9935 -1735 9965 -1715
rect 9985 -1735 10015 -1715
rect 10035 -1735 10065 -1715
rect 10085 -1735 10115 -1715
rect 10135 -1735 10165 -1715
rect 10185 -1735 10215 -1715
rect 10235 -1735 10265 -1715
rect 10285 -1735 10315 -1715
rect 10335 -1735 10365 -1715
rect 10385 -1735 10415 -1715
rect 10435 -1735 10465 -1715
rect 10485 -1735 10515 -1715
rect 10535 -1735 10565 -1715
rect 10585 -1735 10615 -1715
rect 10635 -1735 10665 -1715
rect 10685 -1735 10715 -1715
rect 10735 -1735 10765 -1715
rect 10785 -1735 10815 -1715
rect 10835 -1735 10865 -1715
rect 10885 -1735 10915 -1715
rect 10935 -1735 10965 -1715
rect 10985 -1735 11015 -1715
rect 11035 -1735 11065 -1715
rect 11085 -1735 11115 -1715
rect 11135 -1735 11165 -1715
rect 11185 -1735 11215 -1715
rect 11235 -1735 11265 -1715
rect 11285 -1735 11315 -1715
rect 11335 -1735 11365 -1715
rect 11385 -1735 11415 -1715
rect 11435 -1735 11465 -1715
rect 11485 -1735 11515 -1715
rect 11535 -1735 11565 -1715
rect 11585 -1735 11615 -1715
rect 11635 -1735 11665 -1715
rect 11685 -1735 11715 -1715
rect 11735 -1735 11765 -1715
rect 11785 -1735 11815 -1715
rect 11835 -1735 11865 -1715
rect 11885 -1735 11915 -1715
rect 11935 -1735 11965 -1715
rect 11985 -1735 12015 -1715
rect 12035 -1735 12065 -1715
rect 12085 -1735 12115 -1715
rect 12135 -1735 12165 -1715
rect 12185 -1735 12215 -1715
rect 12235 -1735 12265 -1715
rect 12285 -1735 12315 -1715
rect 12335 -1735 12365 -1715
rect 12385 -1735 12415 -1715
rect 12435 -1735 12465 -1715
rect 12485 -1735 12515 -1715
rect 12535 -1735 12565 -1715
rect 12585 -1735 12615 -1715
rect 12635 -1735 12665 -1715
rect 12685 -1735 12715 -1715
rect 12735 -1735 12765 -1715
rect 12785 -1735 12815 -1715
rect 12835 -1735 12865 -1715
rect 12885 -1735 12915 -1715
rect 12935 -1735 12965 -1715
rect 12985 -1735 13015 -1715
rect 13035 -1735 13065 -1715
rect 13085 -1735 13115 -1715
rect 13135 -1735 13165 -1715
rect 13185 -1735 13215 -1715
rect 13235 -1735 13265 -1715
rect 13285 -1735 13315 -1715
rect 13335 -1735 13365 -1715
rect 13385 -1735 13415 -1715
rect 13435 -1735 13465 -1715
rect 13485 -1735 13515 -1715
rect 13535 -1735 13565 -1715
rect 13585 -1735 13615 -1715
rect 13635 -1735 13665 -1715
rect 13685 -1735 13715 -1715
rect 13735 -1735 13765 -1715
rect 13785 -1735 13815 -1715
rect 13835 -1735 13865 -1715
rect 13885 -1735 13915 -1715
rect 13935 -1735 13965 -1715
rect 13985 -1735 14015 -1715
rect 14035 -1735 14065 -1715
rect 14085 -1735 14115 -1715
rect 14135 -1735 14165 -1715
rect 14185 -1735 14215 -1715
rect 14235 -1735 14265 -1715
rect 14285 -1735 14315 -1715
rect 14335 -1735 14365 -1715
rect 14385 -1735 14415 -1715
rect 14435 -1735 14465 -1715
rect 14485 -1735 14515 -1715
rect 14535 -1735 14565 -1715
rect 14585 -1735 14615 -1715
rect 14635 -1735 14665 -1715
rect 14685 -1735 14715 -1715
rect 14735 -1735 14765 -1715
rect 14785 -1735 14815 -1715
rect 14835 -1735 14865 -1715
rect 14885 -1735 14915 -1715
rect 14935 -1735 14965 -1715
rect 14985 -1735 15015 -1715
rect 15035 -1735 15065 -1715
rect 15085 -1735 15115 -1715
rect 15135 -1735 15165 -1715
rect 15185 -1735 15215 -1715
rect 15235 -1735 15265 -1715
rect 15285 -1735 15315 -1715
rect 15335 -1735 15365 -1715
rect 15385 -1735 15415 -1715
rect 15435 -1735 15465 -1715
rect 15485 -1735 15515 -1715
rect 15535 -1735 15565 -1715
rect 15585 -1735 15615 -1715
rect 15635 -1735 15665 -1715
rect 15685 -1735 15715 -1715
rect 15735 -1735 15765 -1715
rect 15785 -1735 15815 -1715
rect 15835 -1735 15865 -1715
rect 15885 -1735 15915 -1715
rect 15935 -1735 15965 -1715
rect 15985 -1735 16015 -1715
rect 16035 -1735 16065 -1715
rect 16085 -1735 16115 -1715
rect 16135 -1735 16165 -1715
rect 16185 -1735 16215 -1715
rect 16235 -1735 16265 -1715
rect 16285 -1735 16315 -1715
rect 16335 -1735 16365 -1715
rect 16385 -1735 16415 -1715
rect 16435 -1735 16465 -1715
rect 16485 -1735 16515 -1715
rect 16535 -1735 16565 -1715
rect 16585 -1735 16615 -1715
rect 16635 -1735 16665 -1715
rect 16685 -1735 16715 -1715
rect 16735 -1735 16765 -1715
rect 16785 -1735 16815 -1715
rect 16835 -1735 16865 -1715
rect 16885 -1735 16915 -1715
rect 16935 -1735 16965 -1715
rect 16985 -1735 17015 -1715
rect 17035 -1735 17065 -1715
rect 17085 -1735 17115 -1715
rect 17135 -1735 17165 -1715
rect 17185 -1735 17215 -1715
rect 17235 -1735 17265 -1715
rect 17285 -1735 17315 -1715
rect 17335 -1735 17365 -1715
rect 17385 -1735 17415 -1715
rect 17435 -1735 17465 -1715
rect 17485 -1735 17515 -1715
rect 17535 -1735 17565 -1715
rect 17585 -1735 17615 -1715
rect 17635 -1735 17665 -1715
rect 17685 -1735 17715 -1715
rect 17735 -1735 17765 -1715
rect 17785 -1735 17815 -1715
rect 17835 -1735 17865 -1715
rect 17885 -1735 17915 -1715
rect 17935 -1735 17965 -1715
rect 17985 -1735 18015 -1715
rect 18035 -1735 18065 -1715
rect 18085 -1735 18115 -1715
rect 18135 -1735 18165 -1715
rect 18185 -1735 18215 -1715
rect 18235 -1735 18265 -1715
rect 18285 -1735 18315 -1715
rect 18335 -1735 18365 -1715
rect 18385 -1735 18415 -1715
rect 18435 -1735 18465 -1715
rect 18485 -1735 18515 -1715
rect 18535 -1735 18565 -1715
rect 18585 -1735 18615 -1715
rect 18635 -1735 18665 -1715
rect 18685 -1735 18715 -1715
rect 18735 -1735 18765 -1715
rect 18785 -1735 18815 -1715
rect 18835 -1735 18865 -1715
rect 18885 -1735 18915 -1715
rect 18935 -1735 18965 -1715
rect 18985 -1735 19015 -1715
rect 19035 -1735 19065 -1715
rect 19085 -1735 19115 -1715
rect 19135 -1735 19165 -1715
rect 19185 -1735 19215 -1715
rect 19235 -1735 19265 -1715
rect 19285 -1735 19315 -1715
rect 19335 -1735 19365 -1715
rect 19385 -1735 19415 -1715
rect 19435 -1735 19465 -1715
rect 19485 -1735 19515 -1715
rect 19535 -1735 19565 -1715
rect 19585 -1735 19615 -1715
rect 19635 -1735 19665 -1715
rect 19685 -1735 19715 -1715
rect 19735 -1735 19765 -1715
rect 19785 -1735 19815 -1715
rect 19835 -1735 19865 -1715
rect 19885 -1735 19915 -1715
rect 19935 -1735 19965 -1715
rect 19985 -1735 20015 -1715
rect 20035 -1735 20065 -1715
rect 20085 -1735 20115 -1715
rect 20135 -1735 20165 -1715
rect 20185 -1735 20215 -1715
rect 20235 -1735 20265 -1715
rect 20285 -1735 20315 -1715
rect 20335 -1735 20365 -1715
rect 20385 -1735 20415 -1715
rect 20435 -1735 20465 -1715
rect 20485 -1735 20515 -1715
rect 20535 -1735 20565 -1715
rect 20585 -1735 20615 -1715
rect 20635 -1735 20665 -1715
rect 20685 -1735 20715 -1715
rect 20735 -1735 20765 -1715
rect 20785 -1735 20815 -1715
rect 20835 -1735 20865 -1715
rect 20885 -1735 20915 -1715
rect 20935 -1735 20965 -1715
rect 20985 -1735 21015 -1715
rect 21035 -1735 21065 -1715
rect 21085 -1735 21115 -1715
rect 21135 -1735 21165 -1715
rect 21185 -1735 21215 -1715
rect 21235 -1735 21265 -1715
rect 21285 -1735 21315 -1715
rect 21335 -1735 21365 -1715
rect 21385 -1735 21415 -1715
rect 21435 -1735 21465 -1715
rect 21485 -1735 21515 -1715
rect 21535 -1735 21565 -1715
rect 21585 -1735 21615 -1715
rect 21635 -1735 21665 -1715
rect 21685 -1735 21715 -1715
rect 21735 -1735 21765 -1715
rect 21785 -1735 21815 -1715
rect 21835 -1735 21865 -1715
rect 21885 -1735 21915 -1715
rect 21935 -1735 21965 -1715
rect 21985 -1735 22015 -1715
rect 22035 -1735 22065 -1715
rect 22085 -1735 22115 -1715
rect 22135 -1735 22165 -1715
rect 22185 -1735 22215 -1715
rect 22235 -1735 22265 -1715
rect 22285 -1735 22315 -1715
rect 22335 -1735 22365 -1715
rect 22385 -1735 22415 -1715
rect 22435 -1735 22465 -1715
rect 22485 -1735 22515 -1715
rect 22535 -1735 22565 -1715
rect 22585 -1735 22615 -1715
rect 22635 -1735 22665 -1715
rect 22685 -1735 22715 -1715
rect 22735 -1735 22765 -1715
rect 22785 -1735 22815 -1715
rect 22835 -1735 22865 -1715
rect 22885 -1735 22915 -1715
rect 22935 -1735 22965 -1715
rect 22985 -1735 23015 -1715
rect 23035 -1735 23065 -1715
rect 23085 -1735 23115 -1715
rect 23135 -1735 23165 -1715
rect 23185 -1735 23215 -1715
rect 23235 -1735 23265 -1715
rect 23285 -1735 23315 -1715
rect 23335 -1735 23365 -1715
rect 23385 -1735 23415 -1715
rect 23435 -1735 23465 -1715
rect 23485 -1735 23515 -1715
rect 23535 -1735 23565 -1715
rect 23585 -1735 23615 -1715
rect 23635 -1735 23665 -1715
rect 23685 -1735 23715 -1715
rect 23735 -1735 23765 -1715
rect 23785 -1735 23815 -1715
rect 23835 -1735 23865 -1715
rect 23885 -1735 23915 -1715
rect 23935 -1735 23965 -1715
rect 23985 -1735 24015 -1715
rect 24035 -1735 24065 -1715
rect 24085 -1735 24115 -1715
rect 24135 -1735 24165 -1715
rect 24185 -1735 24215 -1715
rect 24235 -1735 24265 -1715
rect 24285 -1735 24315 -1715
rect 24335 -1735 24365 -1715
rect 24385 -1735 24415 -1715
rect 24435 -1735 24465 -1715
rect 24485 -1735 24515 -1715
rect 24535 -1735 24565 -1715
rect 24585 -1735 24615 -1715
rect 24635 -1735 24665 -1715
rect 24685 -1735 24715 -1715
rect 24735 -1735 24765 -1715
rect 24785 -1735 24815 -1715
rect 24835 -1735 24865 -1715
rect 24885 -1735 24915 -1715
rect 24935 -1735 24965 -1715
rect 24985 -1735 25015 -1715
rect 25035 -1735 25065 -1715
rect 25085 -1735 25115 -1715
rect 25135 -1735 25165 -1715
rect 25185 -1735 25215 -1715
rect 25235 -1735 25265 -1715
rect 25285 -1735 25315 -1715
rect 25335 -1735 25365 -1715
rect 25385 -1735 25415 -1715
rect 25435 -1735 25465 -1715
rect 25485 -1735 25515 -1715
rect 25535 -1735 25565 -1715
rect 25585 -1735 25615 -1715
rect 25635 -1735 25665 -1715
rect 25685 -1735 25715 -1715
rect 25735 -1735 25765 -1715
rect 25785 -1735 25815 -1715
rect 25835 -1735 25865 -1715
rect 25885 -1735 25915 -1715
rect 25935 -1735 25965 -1715
rect 25985 -1735 26015 -1715
rect 26035 -1735 26065 -1715
rect 26085 -1735 26115 -1715
rect 26135 -1735 26165 -1715
rect 26185 -1735 26215 -1715
rect 26235 -1735 26265 -1715
rect 26285 -1735 26315 -1715
rect 26335 -1735 26365 -1715
rect 26385 -1735 26415 -1715
rect 26435 -1735 26465 -1715
rect 26485 -1735 26515 -1715
rect 26535 -1735 26565 -1715
rect 26585 -1735 26615 -1715
rect 26635 -1735 26665 -1715
rect 26685 -1735 26715 -1715
rect 26735 -1735 26765 -1715
rect 26785 -1735 26815 -1715
rect 26835 -1735 26865 -1715
rect 26885 -1735 26915 -1715
rect 26935 -1735 26965 -1715
rect 26985 -1735 27015 -1715
rect 27035 -1735 27065 -1715
rect 27085 -1735 27115 -1715
rect 27135 -1735 27165 -1715
rect 27185 -1735 27215 -1715
rect 27235 -1735 27265 -1715
rect 27285 -1735 27315 -1715
rect 27335 -1735 27365 -1715
rect 27385 -1735 27415 -1715
rect 27435 -1735 27465 -1715
rect 27485 -1735 27515 -1715
rect 27535 -1735 27565 -1715
rect 27585 -1735 27615 -1715
rect 27635 -1735 27665 -1715
rect 27685 -1735 27715 -1715
rect 27735 -1735 27765 -1715
rect 27785 -1735 27815 -1715
rect 27835 -1735 27865 -1715
rect 27885 -1735 27915 -1715
rect 27935 -1735 27965 -1715
rect 27985 -1735 28015 -1715
rect 28035 -1735 28065 -1715
rect 28085 -1735 28115 -1715
rect 28135 -1735 28165 -1715
rect 28185 -1735 28215 -1715
rect 28235 -1735 28265 -1715
rect 28285 -1735 28315 -1715
rect 28335 -1735 28365 -1715
rect 28385 -1735 28415 -1715
rect 28435 -1735 28465 -1715
rect 28485 -1735 28515 -1715
rect 28535 -1735 28565 -1715
rect 28585 -1735 28615 -1715
rect 28635 -1735 28665 -1715
rect 28685 -1735 28715 -1715
rect 28735 -1735 28765 -1715
rect 28785 -1735 28800 -1715
rect -650 -1750 28800 -1735
<< mvnsubdiff >>
rect -650 5585 32100 5600
rect -650 5565 -635 5585
rect -615 5565 -585 5585
rect -565 5565 -535 5585
rect -515 5565 -485 5585
rect -465 5565 -435 5585
rect -415 5565 -385 5585
rect -365 5565 -335 5585
rect -315 5565 -285 5585
rect -265 5565 -235 5585
rect -215 5565 -185 5585
rect -165 5565 -135 5585
rect -115 5565 -85 5585
rect -65 5565 -35 5585
rect -15 5565 15 5585
rect 35 5565 65 5585
rect 85 5565 115 5585
rect 135 5565 165 5585
rect 185 5565 215 5585
rect 235 5565 265 5585
rect 285 5565 315 5585
rect 335 5565 365 5585
rect 385 5565 415 5585
rect 435 5565 465 5585
rect 485 5565 515 5585
rect 535 5565 565 5585
rect 585 5565 615 5585
rect 635 5565 665 5585
rect 685 5565 715 5585
rect 735 5565 765 5585
rect 785 5565 815 5585
rect 835 5565 865 5585
rect 885 5565 915 5585
rect 935 5565 965 5585
rect 985 5565 1015 5585
rect 1035 5565 1065 5585
rect 1085 5565 1115 5585
rect 1135 5565 1165 5585
rect 1185 5565 1215 5585
rect 1235 5565 1265 5585
rect 1285 5565 1315 5585
rect 1335 5565 1365 5585
rect 1385 5565 1415 5585
rect 1435 5565 1465 5585
rect 1485 5565 1515 5585
rect 1535 5565 1565 5585
rect 1585 5565 1615 5585
rect 1635 5565 1665 5585
rect 1685 5565 1715 5585
rect 1735 5565 1765 5585
rect 1785 5565 1815 5585
rect 1835 5565 1865 5585
rect 1885 5565 1915 5585
rect 1935 5565 1965 5585
rect 1985 5565 2015 5585
rect 2035 5565 2065 5585
rect 2085 5565 2115 5585
rect 2135 5565 2165 5585
rect 2185 5565 2215 5585
rect 2235 5565 2265 5585
rect 2285 5565 2315 5585
rect 2335 5565 2365 5585
rect 2385 5565 2415 5585
rect 2435 5565 2465 5585
rect 2485 5565 2515 5585
rect 2535 5565 2565 5585
rect 2585 5565 2615 5585
rect 2635 5565 2665 5585
rect 2685 5565 2715 5585
rect 2735 5565 2765 5585
rect 2785 5565 2815 5585
rect 2835 5565 2865 5585
rect 2885 5565 2915 5585
rect 2935 5565 2965 5585
rect 2985 5565 3015 5585
rect 3035 5565 3065 5585
rect 3085 5565 3115 5585
rect 3135 5565 3165 5585
rect 3185 5565 3215 5585
rect 3235 5565 3265 5585
rect 3285 5565 3315 5585
rect 3335 5565 3365 5585
rect 3385 5565 3415 5585
rect 3435 5565 3465 5585
rect 3485 5565 3515 5585
rect 3535 5565 3565 5585
rect 3585 5565 3615 5585
rect 3635 5565 3665 5585
rect 3685 5565 3715 5585
rect 3735 5565 3765 5585
rect 3785 5565 3815 5585
rect 3835 5565 3865 5585
rect 3885 5565 3915 5585
rect 3935 5565 3965 5585
rect 3985 5565 4015 5585
rect 4035 5565 4065 5585
rect 4085 5565 4115 5585
rect 4135 5565 4165 5585
rect 4185 5565 4215 5585
rect 4235 5565 4265 5585
rect 4285 5565 4315 5585
rect 4335 5565 4365 5585
rect 4385 5565 4415 5585
rect 4435 5565 4465 5585
rect 4485 5565 4515 5585
rect 4535 5565 4565 5585
rect 4585 5565 4615 5585
rect 4635 5565 4665 5585
rect 4685 5565 4715 5585
rect 4735 5565 4765 5585
rect 4785 5565 4815 5585
rect 4835 5565 4865 5585
rect 4885 5565 4915 5585
rect 4935 5565 4965 5585
rect 4985 5565 5015 5585
rect 5035 5565 5065 5585
rect 5085 5565 5115 5585
rect 5135 5565 5165 5585
rect 5185 5565 5215 5585
rect 5235 5565 5265 5585
rect 5285 5565 5315 5585
rect 5335 5565 5365 5585
rect 5385 5565 5415 5585
rect 5435 5565 5465 5585
rect 5485 5565 5515 5585
rect 5535 5565 5565 5585
rect 5585 5565 5615 5585
rect 5635 5565 5665 5585
rect 5685 5565 5715 5585
rect 5735 5565 5765 5585
rect 5785 5565 5815 5585
rect 5835 5565 5865 5585
rect 5885 5565 5915 5585
rect 5935 5565 5965 5585
rect 5985 5565 6015 5585
rect 6035 5565 6065 5585
rect 6085 5565 6115 5585
rect 6135 5565 6165 5585
rect 6185 5565 6215 5585
rect 6235 5565 6265 5585
rect 6285 5565 6315 5585
rect 6335 5565 6365 5585
rect 6385 5565 6415 5585
rect 6435 5565 6465 5585
rect 6485 5565 6515 5585
rect 6535 5565 6565 5585
rect 6585 5565 6615 5585
rect 6635 5565 6665 5585
rect 6685 5565 6715 5585
rect 6735 5565 6765 5585
rect 6785 5565 6815 5585
rect 6835 5565 6865 5585
rect 6885 5565 6915 5585
rect 6935 5565 6965 5585
rect 6985 5565 7015 5585
rect 7035 5565 7065 5585
rect 7085 5565 7115 5585
rect 7135 5565 7165 5585
rect 7185 5565 7215 5585
rect 7235 5565 7265 5585
rect 7285 5565 7315 5585
rect 7335 5565 7365 5585
rect 7385 5565 7415 5585
rect 7435 5565 7465 5585
rect 7485 5565 7515 5585
rect 7535 5565 7565 5585
rect 7585 5565 7615 5585
rect 7635 5565 7665 5585
rect 7685 5565 7715 5585
rect 7735 5565 7765 5585
rect 7785 5565 7815 5585
rect 7835 5565 7865 5585
rect 7885 5565 7915 5585
rect 7935 5565 7965 5585
rect 7985 5565 8015 5585
rect 8035 5565 8065 5585
rect 8085 5565 8115 5585
rect 8135 5565 8165 5585
rect 8185 5565 8215 5585
rect 8235 5565 8265 5585
rect 8285 5565 8315 5585
rect 8335 5565 8365 5585
rect 8385 5565 8415 5585
rect 8435 5565 8465 5585
rect 8485 5565 8515 5585
rect 8535 5565 8565 5585
rect 8585 5565 8615 5585
rect 8635 5565 8665 5585
rect 8685 5565 8715 5585
rect 8735 5565 8765 5585
rect 8785 5565 8815 5585
rect 8835 5565 8865 5585
rect 8885 5565 8915 5585
rect 8935 5565 8965 5585
rect 8985 5565 9015 5585
rect 9035 5565 9065 5585
rect 9085 5565 9115 5585
rect 9135 5565 9165 5585
rect 9185 5565 9215 5585
rect 9235 5565 9265 5585
rect 9285 5565 9315 5585
rect 9335 5565 9365 5585
rect 9385 5565 9415 5585
rect 9435 5565 9465 5585
rect 9485 5565 9515 5585
rect 9535 5565 9565 5585
rect 9585 5565 9615 5585
rect 9635 5565 9665 5585
rect 9685 5565 9715 5585
rect 9735 5565 9765 5585
rect 9785 5565 9815 5585
rect 9835 5565 9865 5585
rect 9885 5565 9915 5585
rect 9935 5565 9965 5585
rect 9985 5565 10015 5585
rect 10035 5565 10065 5585
rect 10085 5565 10115 5585
rect 10135 5565 10165 5585
rect 10185 5565 10215 5585
rect 10235 5565 10265 5585
rect 10285 5565 10315 5585
rect 10335 5565 10365 5585
rect 10385 5565 10415 5585
rect 10435 5565 10465 5585
rect 10485 5565 10515 5585
rect 10535 5565 10565 5585
rect 10585 5565 10615 5585
rect 10635 5565 10665 5585
rect 10685 5565 10715 5585
rect 10735 5565 10765 5585
rect 10785 5565 10815 5585
rect 10835 5565 10865 5585
rect 10885 5565 10915 5585
rect 10935 5565 10965 5585
rect 10985 5565 11015 5585
rect 11035 5565 11065 5585
rect 11085 5565 11115 5585
rect 11135 5565 11165 5585
rect 11185 5565 11215 5585
rect 11235 5565 11265 5585
rect 11285 5565 11315 5585
rect 11335 5565 11365 5585
rect 11385 5565 11415 5585
rect 11435 5565 11465 5585
rect 11485 5565 11515 5585
rect 11535 5565 11565 5585
rect 11585 5565 11615 5585
rect 11635 5565 11665 5585
rect 11685 5565 11715 5585
rect 11735 5565 11765 5585
rect 11785 5565 11815 5585
rect 11835 5565 11865 5585
rect 11885 5565 11915 5585
rect 11935 5565 11965 5585
rect 11985 5565 12015 5585
rect 12035 5565 12065 5585
rect 12085 5565 12115 5585
rect 12135 5565 12165 5585
rect 12185 5565 12215 5585
rect 12235 5565 12265 5585
rect 12285 5565 12315 5585
rect 12335 5565 12365 5585
rect 12385 5565 12415 5585
rect 12435 5565 12465 5585
rect 12485 5565 12515 5585
rect 12535 5565 12565 5585
rect 12585 5565 12615 5585
rect 12635 5565 12665 5585
rect 12685 5565 12715 5585
rect 12735 5565 12765 5585
rect 12785 5565 12815 5585
rect 12835 5565 12865 5585
rect 12885 5565 12915 5585
rect 12935 5565 12965 5585
rect 12985 5565 13015 5585
rect 13035 5565 13065 5585
rect 13085 5565 13115 5585
rect 13135 5565 13165 5585
rect 13185 5565 13215 5585
rect 13235 5565 13265 5585
rect 13285 5565 13315 5585
rect 13335 5565 13365 5585
rect 13385 5565 13415 5585
rect 13435 5565 13465 5585
rect 13485 5565 13515 5585
rect 13535 5565 13565 5585
rect 13585 5565 13615 5585
rect 13635 5565 13665 5585
rect 13685 5565 13715 5585
rect 13735 5565 13765 5585
rect 13785 5565 13815 5585
rect 13835 5565 13865 5585
rect 13885 5565 13915 5585
rect 13935 5565 13965 5585
rect 13985 5565 14015 5585
rect 14035 5565 14065 5585
rect 14085 5565 14115 5585
rect 14135 5565 14165 5585
rect 14185 5565 14215 5585
rect 14235 5565 14265 5585
rect 14285 5565 14315 5585
rect 14335 5565 14365 5585
rect 14385 5565 14415 5585
rect 14435 5565 14465 5585
rect 14485 5565 14515 5585
rect 14535 5565 14565 5585
rect 14585 5565 14615 5585
rect 14635 5565 14665 5585
rect 14685 5565 14715 5585
rect 14735 5565 14765 5585
rect 14785 5565 14815 5585
rect 14835 5565 14865 5585
rect 14885 5565 14915 5585
rect 14935 5565 14965 5585
rect 14985 5565 15015 5585
rect 15035 5565 15065 5585
rect 15085 5565 15115 5585
rect 15135 5565 15165 5585
rect 15185 5565 15215 5585
rect 15235 5565 15265 5585
rect 15285 5565 15315 5585
rect 15335 5565 15365 5585
rect 15385 5565 15415 5585
rect 15435 5565 15465 5585
rect 15485 5565 15515 5585
rect 15535 5565 15565 5585
rect 15585 5565 15615 5585
rect 15635 5565 15665 5585
rect 15685 5565 15715 5585
rect 15735 5565 15765 5585
rect 15785 5565 15815 5585
rect 15835 5565 15865 5585
rect 15885 5565 15915 5585
rect 15935 5565 15965 5585
rect 15985 5565 16015 5585
rect 16035 5565 16065 5585
rect 16085 5565 16115 5585
rect 16135 5565 16165 5585
rect 16185 5565 16215 5585
rect 16235 5565 16265 5585
rect 16285 5565 16315 5585
rect 16335 5565 16365 5585
rect 16385 5565 16415 5585
rect 16435 5565 16465 5585
rect 16485 5565 16515 5585
rect 16535 5565 16565 5585
rect 16585 5565 16615 5585
rect 16635 5565 16665 5585
rect 16685 5565 16715 5585
rect 16735 5565 16765 5585
rect 16785 5565 16815 5585
rect 16835 5565 16865 5585
rect 16885 5565 16915 5585
rect 16935 5565 16965 5585
rect 16985 5565 17015 5585
rect 17035 5565 17065 5585
rect 17085 5565 17115 5585
rect 17135 5565 17165 5585
rect 17185 5565 17215 5585
rect 17235 5565 17265 5585
rect 17285 5565 17315 5585
rect 17335 5565 17365 5585
rect 17385 5565 17415 5585
rect 17435 5565 17465 5585
rect 17485 5565 17515 5585
rect 17535 5565 17565 5585
rect 17585 5565 17615 5585
rect 17635 5565 17665 5585
rect 17685 5565 17715 5585
rect 17735 5565 17765 5585
rect 17785 5565 17815 5585
rect 17835 5565 17865 5585
rect 17885 5565 17915 5585
rect 17935 5565 17965 5585
rect 17985 5565 18015 5585
rect 18035 5565 18065 5585
rect 18085 5565 18115 5585
rect 18135 5565 18165 5585
rect 18185 5565 18215 5585
rect 18235 5565 18265 5585
rect 18285 5565 18315 5585
rect 18335 5565 18365 5585
rect 18385 5565 18415 5585
rect 18435 5565 18465 5585
rect 18485 5565 18515 5585
rect 18535 5565 18565 5585
rect 18585 5565 18615 5585
rect 18635 5565 18665 5585
rect 18685 5565 18715 5585
rect 18735 5565 18765 5585
rect 18785 5565 18815 5585
rect 18835 5565 18865 5585
rect 18885 5565 18915 5585
rect 18935 5565 18965 5585
rect 18985 5565 19015 5585
rect 19035 5565 19065 5585
rect 19085 5565 19115 5585
rect 19135 5565 19165 5585
rect 19185 5565 19215 5585
rect 19235 5565 19265 5585
rect 19285 5565 19315 5585
rect 19335 5565 19365 5585
rect 19385 5565 19415 5585
rect 19435 5565 19465 5585
rect 19485 5565 19515 5585
rect 19535 5565 19565 5585
rect 19585 5565 19615 5585
rect 19635 5565 19665 5585
rect 19685 5565 19715 5585
rect 19735 5565 19765 5585
rect 19785 5565 19815 5585
rect 19835 5565 19865 5585
rect 19885 5565 19915 5585
rect 19935 5565 19965 5585
rect 19985 5565 20015 5585
rect 20035 5565 20065 5585
rect 20085 5565 20115 5585
rect 20135 5565 20165 5585
rect 20185 5565 20215 5585
rect 20235 5565 20265 5585
rect 20285 5565 20315 5585
rect 20335 5565 20365 5585
rect 20385 5565 20415 5585
rect 20435 5565 20465 5585
rect 20485 5565 20515 5585
rect 20535 5565 20565 5585
rect 20585 5565 20615 5585
rect 20635 5565 20665 5585
rect 20685 5565 20715 5585
rect 20735 5565 20765 5585
rect 20785 5565 20815 5585
rect 20835 5565 20865 5585
rect 20885 5565 20915 5585
rect 20935 5565 20965 5585
rect 20985 5565 21015 5585
rect 21035 5565 21065 5585
rect 21085 5565 21115 5585
rect 21135 5565 21165 5585
rect 21185 5565 21215 5585
rect 21235 5565 21265 5585
rect 21285 5565 21315 5585
rect 21335 5565 21365 5585
rect 21385 5565 21415 5585
rect 21435 5565 21465 5585
rect 21485 5565 21515 5585
rect 21535 5565 21565 5585
rect 21585 5565 21615 5585
rect 21635 5565 21665 5585
rect 21685 5565 21715 5585
rect 21735 5565 21765 5585
rect 21785 5565 21815 5585
rect 21835 5565 21865 5585
rect 21885 5565 21915 5585
rect 21935 5565 21965 5585
rect 21985 5565 22015 5585
rect 22035 5565 22065 5585
rect 22085 5565 22115 5585
rect 22135 5565 22165 5585
rect 22185 5565 22215 5585
rect 22235 5565 22265 5585
rect 22285 5565 22315 5585
rect 22335 5565 22365 5585
rect 22385 5565 22415 5585
rect 22435 5565 22465 5585
rect 22485 5565 22515 5585
rect 22535 5565 22565 5585
rect 22585 5565 22615 5585
rect 22635 5565 22665 5585
rect 22685 5565 22715 5585
rect 22735 5565 22765 5585
rect 22785 5565 22815 5585
rect 22835 5565 22865 5585
rect 22885 5565 22915 5585
rect 22935 5565 22965 5585
rect 22985 5565 23015 5585
rect 23035 5565 23065 5585
rect 23085 5565 23115 5585
rect 23135 5565 23165 5585
rect 23185 5565 23215 5585
rect 23235 5565 23265 5585
rect 23285 5565 23315 5585
rect 23335 5565 23365 5585
rect 23385 5565 23415 5585
rect 23435 5565 23465 5585
rect 23485 5565 23515 5585
rect 23535 5565 23565 5585
rect 23585 5565 23615 5585
rect 23635 5565 23665 5585
rect 23685 5565 23715 5585
rect 23735 5565 23765 5585
rect 23785 5565 23815 5585
rect 23835 5565 23865 5585
rect 23885 5565 23915 5585
rect 23935 5565 23965 5585
rect 23985 5565 24015 5585
rect 24035 5565 24065 5585
rect 24085 5565 24115 5585
rect 24135 5565 24165 5585
rect 24185 5565 24215 5585
rect 24235 5565 24265 5585
rect 24285 5565 24315 5585
rect 24335 5565 24365 5585
rect 24385 5565 24415 5585
rect 24435 5565 24465 5585
rect 24485 5565 24515 5585
rect 24535 5565 24565 5585
rect 24585 5565 24615 5585
rect 24635 5565 24665 5585
rect 24685 5565 24715 5585
rect 24735 5565 24765 5585
rect 24785 5565 24815 5585
rect 24835 5565 24865 5585
rect 24885 5565 24915 5585
rect 24935 5565 24965 5585
rect 24985 5565 25015 5585
rect 25035 5565 25065 5585
rect 25085 5565 25115 5585
rect 25135 5565 25165 5585
rect 25185 5565 25215 5585
rect 25235 5565 25265 5585
rect 25285 5565 25315 5585
rect 25335 5565 25365 5585
rect 25385 5565 25415 5585
rect 25435 5565 25465 5585
rect 25485 5565 25515 5585
rect 25535 5565 25565 5585
rect 25585 5565 25615 5585
rect 25635 5565 25665 5585
rect 25685 5565 25715 5585
rect 25735 5565 25765 5585
rect 25785 5565 25815 5585
rect 25835 5565 25865 5585
rect 25885 5565 25915 5585
rect 25935 5565 25965 5585
rect 25985 5565 26015 5585
rect 26035 5565 26065 5585
rect 26085 5565 26115 5585
rect 26135 5565 26165 5585
rect 26185 5565 26215 5585
rect 26235 5565 26265 5585
rect 26285 5565 26315 5585
rect 26335 5565 26365 5585
rect 26385 5565 26415 5585
rect 26435 5565 26465 5585
rect 26485 5565 26515 5585
rect 26535 5565 26565 5585
rect 26585 5565 26615 5585
rect 26635 5565 26665 5585
rect 26685 5565 26715 5585
rect 26735 5565 26765 5585
rect 26785 5565 26815 5585
rect 26835 5565 26865 5585
rect 26885 5565 26915 5585
rect 26935 5565 26965 5585
rect 26985 5565 27015 5585
rect 27035 5565 27065 5585
rect 27085 5565 27115 5585
rect 27135 5565 27165 5585
rect 27185 5565 27215 5585
rect 27235 5565 27265 5585
rect 27285 5565 27315 5585
rect 27335 5565 27365 5585
rect 27385 5565 27415 5585
rect 27435 5565 27465 5585
rect 27485 5565 27515 5585
rect 27535 5565 27565 5585
rect 27585 5565 27615 5585
rect 27635 5565 27665 5585
rect 27685 5565 27715 5585
rect 27735 5565 27765 5585
rect 27785 5565 27815 5585
rect 27835 5565 27865 5585
rect 27885 5565 27915 5585
rect 27935 5565 27965 5585
rect 27985 5565 28015 5585
rect 28035 5565 28065 5585
rect 28085 5565 28115 5585
rect 28135 5565 28165 5585
rect 28185 5565 28215 5585
rect 28235 5565 28265 5585
rect 28285 5565 28315 5585
rect 28335 5565 28365 5585
rect 28385 5565 28415 5585
rect 28435 5565 28465 5585
rect 28485 5565 28515 5585
rect 28535 5565 28565 5585
rect 28585 5565 28615 5585
rect 28635 5565 28665 5585
rect 28685 5565 28715 5585
rect 28735 5565 28765 5585
rect 28785 5565 28815 5585
rect 28835 5565 28865 5585
rect 28885 5565 28915 5585
rect 28935 5565 28965 5585
rect 28985 5565 29015 5585
rect 29035 5565 29065 5585
rect 29085 5565 29115 5585
rect 29135 5565 29165 5585
rect 29185 5565 29215 5585
rect 29235 5565 29265 5585
rect 29285 5565 29315 5585
rect 29335 5565 29365 5585
rect 29385 5565 29415 5585
rect 29435 5565 29465 5585
rect 29485 5565 29515 5585
rect 29535 5565 29565 5585
rect 29585 5565 29615 5585
rect 29635 5565 29665 5585
rect 29685 5565 29715 5585
rect 29735 5565 29765 5585
rect 29785 5565 29815 5585
rect 29835 5565 29865 5585
rect 29885 5565 29915 5585
rect 29935 5565 29965 5585
rect 29985 5565 30015 5585
rect 30035 5565 30065 5585
rect 30085 5565 30115 5585
rect 30135 5565 30165 5585
rect 30185 5565 30215 5585
rect 30235 5565 30265 5585
rect 30285 5565 30315 5585
rect 30335 5565 30365 5585
rect 30385 5565 30415 5585
rect 30435 5565 30465 5585
rect 30485 5565 30515 5585
rect 30535 5565 30565 5585
rect 30585 5565 30615 5585
rect 30635 5565 30665 5585
rect 30685 5565 30715 5585
rect 30735 5565 30765 5585
rect 30785 5565 30815 5585
rect 30835 5565 30865 5585
rect 30885 5565 30915 5585
rect 30935 5565 30965 5585
rect 30985 5565 31015 5585
rect 31035 5565 31065 5585
rect 31085 5565 31115 5585
rect 31135 5565 31165 5585
rect 31185 5565 31215 5585
rect 31235 5565 31265 5585
rect 31285 5565 31315 5585
rect 31335 5565 31365 5585
rect 31385 5565 31415 5585
rect 31435 5565 31465 5585
rect 31485 5565 31515 5585
rect 31535 5565 31565 5585
rect 31585 5565 31615 5585
rect 31635 5565 31665 5585
rect 31685 5565 31715 5585
rect 31735 5565 31765 5585
rect 31785 5565 31815 5585
rect 31835 5565 31865 5585
rect 31885 5565 31915 5585
rect 31935 5565 31965 5585
rect 31985 5565 32015 5585
rect 32035 5565 32065 5585
rect 32085 5565 32100 5585
rect -650 5550 32100 5565
rect -650 4285 32100 4300
rect -650 4265 -635 4285
rect -615 4265 -585 4285
rect -565 4265 -535 4285
rect -515 4265 -485 4285
rect -465 4265 -435 4285
rect -415 4265 -385 4285
rect -365 4265 -335 4285
rect -315 4265 -285 4285
rect -265 4265 -235 4285
rect -215 4265 -185 4285
rect -165 4265 -135 4285
rect -115 4265 -85 4285
rect -65 4265 -35 4285
rect -15 4265 15 4285
rect 35 4265 65 4285
rect 85 4265 115 4285
rect 135 4265 165 4285
rect 185 4265 215 4285
rect 235 4265 265 4285
rect 285 4265 315 4285
rect 335 4265 365 4285
rect 385 4265 415 4285
rect 435 4265 465 4285
rect 485 4265 515 4285
rect 535 4265 565 4285
rect 585 4265 615 4285
rect 635 4265 665 4285
rect 685 4265 715 4285
rect 735 4265 765 4285
rect 785 4265 815 4285
rect 835 4265 865 4285
rect 885 4265 915 4285
rect 935 4265 965 4285
rect 985 4265 1015 4285
rect 1035 4265 1065 4285
rect 1085 4265 1115 4285
rect 1135 4265 1165 4285
rect 1185 4265 1215 4285
rect 1235 4265 1265 4285
rect 1285 4265 1315 4285
rect 1335 4265 1365 4285
rect 1385 4265 1415 4285
rect 1435 4265 1465 4285
rect 1485 4265 1515 4285
rect 1535 4265 1565 4285
rect 1585 4265 1615 4285
rect 1635 4265 1665 4285
rect 1685 4265 1715 4285
rect 1735 4265 1765 4285
rect 1785 4265 1815 4285
rect 1835 4265 1865 4285
rect 1885 4265 1915 4285
rect 1935 4265 1965 4285
rect 1985 4265 2015 4285
rect 2035 4265 2065 4285
rect 2085 4265 2115 4285
rect 2135 4265 2165 4285
rect 2185 4265 2215 4285
rect 2235 4265 2265 4285
rect 2285 4265 2315 4285
rect 2335 4265 2365 4285
rect 2385 4265 2415 4285
rect 2435 4265 2465 4285
rect 2485 4265 2515 4285
rect 2535 4265 2565 4285
rect 2585 4265 2615 4285
rect 2635 4265 2665 4285
rect 2685 4265 2715 4285
rect 2735 4265 2765 4285
rect 2785 4265 2815 4285
rect 2835 4265 2865 4285
rect 2885 4265 2915 4285
rect 2935 4265 2965 4285
rect 2985 4265 3015 4285
rect 3035 4265 3065 4285
rect 3085 4265 3115 4285
rect 3135 4265 3165 4285
rect 3185 4265 3215 4285
rect 3235 4265 3265 4285
rect 3285 4265 3315 4285
rect 3335 4265 3365 4285
rect 3385 4265 3415 4285
rect 3435 4265 3465 4285
rect 3485 4265 3515 4285
rect 3535 4265 3565 4285
rect 3585 4265 3615 4285
rect 3635 4265 3665 4285
rect 3685 4265 3715 4285
rect 3735 4265 3765 4285
rect 3785 4265 3815 4285
rect 3835 4265 3865 4285
rect 3885 4265 3915 4285
rect 3935 4265 3965 4285
rect 3985 4265 4015 4285
rect 4035 4265 4065 4285
rect 4085 4265 4115 4285
rect 4135 4265 4165 4285
rect 4185 4265 4215 4285
rect 4235 4265 4265 4285
rect 4285 4265 4315 4285
rect 4335 4265 4365 4285
rect 4385 4265 4415 4285
rect 4435 4265 4465 4285
rect 4485 4265 4515 4285
rect 4535 4265 4565 4285
rect 4585 4265 4615 4285
rect 4635 4265 4665 4285
rect 4685 4265 4715 4285
rect 4735 4265 4765 4285
rect 4785 4265 4815 4285
rect 4835 4265 4865 4285
rect 4885 4265 4915 4285
rect 4935 4265 4965 4285
rect 4985 4265 5015 4285
rect 5035 4265 5065 4285
rect 5085 4265 5115 4285
rect 5135 4265 5165 4285
rect 5185 4265 5215 4285
rect 5235 4265 5265 4285
rect 5285 4265 5315 4285
rect 5335 4265 5365 4285
rect 5385 4265 5415 4285
rect 5435 4265 5465 4285
rect 5485 4265 5515 4285
rect 5535 4265 5565 4285
rect 5585 4265 5615 4285
rect 5635 4265 5665 4285
rect 5685 4265 5715 4285
rect 5735 4265 5765 4285
rect 5785 4265 5815 4285
rect 5835 4265 5865 4285
rect 5885 4265 5915 4285
rect 5935 4265 5965 4285
rect 5985 4265 6015 4285
rect 6035 4265 6065 4285
rect 6085 4265 6115 4285
rect 6135 4265 6165 4285
rect 6185 4265 6215 4285
rect 6235 4265 6265 4285
rect 6285 4265 6315 4285
rect 6335 4265 6365 4285
rect 6385 4265 6415 4285
rect 6435 4265 6465 4285
rect 6485 4265 6515 4285
rect 6535 4265 6565 4285
rect 6585 4265 6615 4285
rect 6635 4265 6665 4285
rect 6685 4265 6715 4285
rect 6735 4265 6765 4285
rect 6785 4265 6815 4285
rect 6835 4265 6865 4285
rect 6885 4265 6915 4285
rect 6935 4265 6965 4285
rect 6985 4265 7015 4285
rect 7035 4265 7065 4285
rect 7085 4265 7115 4285
rect 7135 4265 7165 4285
rect 7185 4265 7215 4285
rect 7235 4265 7265 4285
rect 7285 4265 7315 4285
rect 7335 4265 7365 4285
rect 7385 4265 7415 4285
rect 7435 4265 7465 4285
rect 7485 4265 7515 4285
rect 7535 4265 7565 4285
rect 7585 4265 7615 4285
rect 7635 4265 7665 4285
rect 7685 4265 7715 4285
rect 7735 4265 7765 4285
rect 7785 4265 7815 4285
rect 7835 4265 7865 4285
rect 7885 4265 7915 4285
rect 7935 4265 7965 4285
rect 7985 4265 8015 4285
rect 8035 4265 8065 4285
rect 8085 4265 8115 4285
rect 8135 4265 8165 4285
rect 8185 4265 8215 4285
rect 8235 4265 8265 4285
rect 8285 4265 8315 4285
rect 8335 4265 8365 4285
rect 8385 4265 8415 4285
rect 8435 4265 8465 4285
rect 8485 4265 8515 4285
rect 8535 4265 8565 4285
rect 8585 4265 8615 4285
rect 8635 4265 8665 4285
rect 8685 4265 8715 4285
rect 8735 4265 8765 4285
rect 8785 4265 8815 4285
rect 8835 4265 8865 4285
rect 8885 4265 8915 4285
rect 8935 4265 8965 4285
rect 8985 4265 9015 4285
rect 9035 4265 9065 4285
rect 9085 4265 9115 4285
rect 9135 4265 9165 4285
rect 9185 4265 9215 4285
rect 9235 4265 9265 4285
rect 9285 4265 9315 4285
rect 9335 4265 9365 4285
rect 9385 4265 9415 4285
rect 9435 4265 9465 4285
rect 9485 4265 9515 4285
rect 9535 4265 9565 4285
rect 9585 4265 9615 4285
rect 9635 4265 9665 4285
rect 9685 4265 9715 4285
rect 9735 4265 9765 4285
rect 9785 4265 9815 4285
rect 9835 4265 9865 4285
rect 9885 4265 9915 4285
rect 9935 4265 9965 4285
rect 9985 4265 10015 4285
rect 10035 4265 10065 4285
rect 10085 4265 10115 4285
rect 10135 4265 10165 4285
rect 10185 4265 10215 4285
rect 10235 4265 10265 4285
rect 10285 4265 10315 4285
rect 10335 4265 10365 4285
rect 10385 4265 10415 4285
rect 10435 4265 10465 4285
rect 10485 4265 10515 4285
rect 10535 4265 10565 4285
rect 10585 4265 10615 4285
rect 10635 4265 10665 4285
rect 10685 4265 10715 4285
rect 10735 4265 10765 4285
rect 10785 4265 10815 4285
rect 10835 4265 10865 4285
rect 10885 4265 10915 4285
rect 10935 4265 10965 4285
rect 10985 4265 11015 4285
rect 11035 4265 11065 4285
rect 11085 4265 11115 4285
rect 11135 4265 11165 4285
rect 11185 4265 11215 4285
rect 11235 4265 11265 4285
rect 11285 4265 11315 4285
rect 11335 4265 11365 4285
rect 11385 4265 11415 4285
rect 11435 4265 11465 4285
rect 11485 4265 11515 4285
rect 11535 4265 11565 4285
rect 11585 4265 11615 4285
rect 11635 4265 11665 4285
rect 11685 4265 11715 4285
rect 11735 4265 11765 4285
rect 11785 4265 11815 4285
rect 11835 4265 11865 4285
rect 11885 4265 11915 4285
rect 11935 4265 11965 4285
rect 11985 4265 12015 4285
rect 12035 4265 12065 4285
rect 12085 4265 12115 4285
rect 12135 4265 12165 4285
rect 12185 4265 12215 4285
rect 12235 4265 12265 4285
rect 12285 4265 12315 4285
rect 12335 4265 12365 4285
rect 12385 4265 12415 4285
rect 12435 4265 12465 4285
rect 12485 4265 12515 4285
rect 12535 4265 12565 4285
rect 12585 4265 12615 4285
rect 12635 4265 12665 4285
rect 12685 4265 12715 4285
rect 12735 4265 12765 4285
rect 12785 4265 12815 4285
rect 12835 4265 12865 4285
rect 12885 4265 12915 4285
rect 12935 4265 12965 4285
rect 12985 4265 13015 4285
rect 13035 4265 13065 4285
rect 13085 4265 13115 4285
rect 13135 4265 13165 4285
rect 13185 4265 13215 4285
rect 13235 4265 13265 4285
rect 13285 4265 13315 4285
rect 13335 4265 13365 4285
rect 13385 4265 13415 4285
rect 13435 4265 13465 4285
rect 13485 4265 13515 4285
rect 13535 4265 13565 4285
rect 13585 4265 13615 4285
rect 13635 4265 13665 4285
rect 13685 4265 13715 4285
rect 13735 4265 13765 4285
rect 13785 4265 13815 4285
rect 13835 4265 13865 4285
rect 13885 4265 13915 4285
rect 13935 4265 13965 4285
rect 13985 4265 14015 4285
rect 14035 4265 14065 4285
rect 14085 4265 14115 4285
rect 14135 4265 14165 4285
rect 14185 4265 14215 4285
rect 14235 4265 14265 4285
rect 14285 4265 14315 4285
rect 14335 4265 14365 4285
rect 14385 4265 14415 4285
rect 14435 4265 14465 4285
rect 14485 4265 14515 4285
rect 14535 4265 14565 4285
rect 14585 4265 14615 4285
rect 14635 4265 14665 4285
rect 14685 4265 14715 4285
rect 14735 4265 14765 4285
rect 14785 4265 14815 4285
rect 14835 4265 14865 4285
rect 14885 4265 14915 4285
rect 14935 4265 14965 4285
rect 14985 4265 15015 4285
rect 15035 4265 15065 4285
rect 15085 4265 15115 4285
rect 15135 4265 15165 4285
rect 15185 4265 15215 4285
rect 15235 4265 15265 4285
rect 15285 4265 15315 4285
rect 15335 4265 15365 4285
rect 15385 4265 15415 4285
rect 15435 4265 15465 4285
rect 15485 4265 15515 4285
rect 15535 4265 15565 4285
rect 15585 4265 15615 4285
rect 15635 4265 15665 4285
rect 15685 4265 15715 4285
rect 15735 4265 15765 4285
rect 15785 4265 15815 4285
rect 15835 4265 15865 4285
rect 15885 4265 15915 4285
rect 15935 4265 15965 4285
rect 15985 4265 16015 4285
rect 16035 4265 16065 4285
rect 16085 4265 16115 4285
rect 16135 4265 16165 4285
rect 16185 4265 16215 4285
rect 16235 4265 16265 4285
rect 16285 4265 16315 4285
rect 16335 4265 16365 4285
rect 16385 4265 16415 4285
rect 16435 4265 16465 4285
rect 16485 4265 16515 4285
rect 16535 4265 16565 4285
rect 16585 4265 16615 4285
rect 16635 4265 16665 4285
rect 16685 4265 16715 4285
rect 16735 4265 16765 4285
rect 16785 4265 16815 4285
rect 16835 4265 16865 4285
rect 16885 4265 16915 4285
rect 16935 4265 16965 4285
rect 16985 4265 17015 4285
rect 17035 4265 17065 4285
rect 17085 4265 17115 4285
rect 17135 4265 17165 4285
rect 17185 4265 17215 4285
rect 17235 4265 17265 4285
rect 17285 4265 17315 4285
rect 17335 4265 17365 4285
rect 17385 4265 17415 4285
rect 17435 4265 17465 4285
rect 17485 4265 17515 4285
rect 17535 4265 17565 4285
rect 17585 4265 17615 4285
rect 17635 4265 17665 4285
rect 17685 4265 17715 4285
rect 17735 4265 17765 4285
rect 17785 4265 17815 4285
rect 17835 4265 17865 4285
rect 17885 4265 17915 4285
rect 17935 4265 17965 4285
rect 17985 4265 18015 4285
rect 18035 4265 18065 4285
rect 18085 4265 18115 4285
rect 18135 4265 18165 4285
rect 18185 4265 18215 4285
rect 18235 4265 18265 4285
rect 18285 4265 18315 4285
rect 18335 4265 18365 4285
rect 18385 4265 18415 4285
rect 18435 4265 18465 4285
rect 18485 4265 18515 4285
rect 18535 4265 18565 4285
rect 18585 4265 18615 4285
rect 18635 4265 18665 4285
rect 18685 4265 18715 4285
rect 18735 4265 18765 4285
rect 18785 4265 18815 4285
rect 18835 4265 18865 4285
rect 18885 4265 18915 4285
rect 18935 4265 18965 4285
rect 18985 4265 19015 4285
rect 19035 4265 19065 4285
rect 19085 4265 19115 4285
rect 19135 4265 19165 4285
rect 19185 4265 19215 4285
rect 19235 4265 19265 4285
rect 19285 4265 19315 4285
rect 19335 4265 19365 4285
rect 19385 4265 19415 4285
rect 19435 4265 19465 4285
rect 19485 4265 19515 4285
rect 19535 4265 19565 4285
rect 19585 4265 19615 4285
rect 19635 4265 19665 4285
rect 19685 4265 19715 4285
rect 19735 4265 19765 4285
rect 19785 4265 19815 4285
rect 19835 4265 19865 4285
rect 19885 4265 19915 4285
rect 19935 4265 19965 4285
rect 19985 4265 20015 4285
rect 20035 4265 20065 4285
rect 20085 4265 20115 4285
rect 20135 4265 20165 4285
rect 20185 4265 20215 4285
rect 20235 4265 20265 4285
rect 20285 4265 20315 4285
rect 20335 4265 20365 4285
rect 20385 4265 20415 4285
rect 20435 4265 20465 4285
rect 20485 4265 20515 4285
rect 20535 4265 20565 4285
rect 20585 4265 20615 4285
rect 20635 4265 20665 4285
rect 20685 4265 20715 4285
rect 20735 4265 20765 4285
rect 20785 4265 20815 4285
rect 20835 4265 20865 4285
rect 20885 4265 20915 4285
rect 20935 4265 20965 4285
rect 20985 4265 21015 4285
rect 21035 4265 21065 4285
rect 21085 4265 21115 4285
rect 21135 4265 21165 4285
rect 21185 4265 21215 4285
rect 21235 4265 21265 4285
rect 21285 4265 21315 4285
rect 21335 4265 21365 4285
rect 21385 4265 21415 4285
rect 21435 4265 21465 4285
rect 21485 4265 21515 4285
rect 21535 4265 21565 4285
rect 21585 4265 21615 4285
rect 21635 4265 21665 4285
rect 21685 4265 21715 4285
rect 21735 4265 21765 4285
rect 21785 4265 21815 4285
rect 21835 4265 21865 4285
rect 21885 4265 21915 4285
rect 21935 4265 21965 4285
rect 21985 4265 22015 4285
rect 22035 4265 22065 4285
rect 22085 4265 22115 4285
rect 22135 4265 22165 4285
rect 22185 4265 22215 4285
rect 22235 4265 22265 4285
rect 22285 4265 22315 4285
rect 22335 4265 22365 4285
rect 22385 4265 22415 4285
rect 22435 4265 22465 4285
rect 22485 4265 22515 4285
rect 22535 4265 22565 4285
rect 22585 4265 22615 4285
rect 22635 4265 22665 4285
rect 22685 4265 22715 4285
rect 22735 4265 22765 4285
rect 22785 4265 22815 4285
rect 22835 4265 22865 4285
rect 22885 4265 22915 4285
rect 22935 4265 22965 4285
rect 22985 4265 23015 4285
rect 23035 4265 23065 4285
rect 23085 4265 23115 4285
rect 23135 4265 23165 4285
rect 23185 4265 23215 4285
rect 23235 4265 23265 4285
rect 23285 4265 23315 4285
rect 23335 4265 23365 4285
rect 23385 4265 23415 4285
rect 23435 4265 23465 4285
rect 23485 4265 23515 4285
rect 23535 4265 23565 4285
rect 23585 4265 23615 4285
rect 23635 4265 23665 4285
rect 23685 4265 23715 4285
rect 23735 4265 23765 4285
rect 23785 4265 23815 4285
rect 23835 4265 23865 4285
rect 23885 4265 23915 4285
rect 23935 4265 23965 4285
rect 23985 4265 24015 4285
rect 24035 4265 24065 4285
rect 24085 4265 24115 4285
rect 24135 4265 24165 4285
rect 24185 4265 24215 4285
rect 24235 4265 24265 4285
rect 24285 4265 24315 4285
rect 24335 4265 24365 4285
rect 24385 4265 24415 4285
rect 24435 4265 24465 4285
rect 24485 4265 24515 4285
rect 24535 4265 24565 4285
rect 24585 4265 24615 4285
rect 24635 4265 24665 4285
rect 24685 4265 24715 4285
rect 24735 4265 24765 4285
rect 24785 4265 24815 4285
rect 24835 4265 24865 4285
rect 24885 4265 24915 4285
rect 24935 4265 24965 4285
rect 24985 4265 25015 4285
rect 25035 4265 25065 4285
rect 25085 4265 25115 4285
rect 25135 4265 25165 4285
rect 25185 4265 25215 4285
rect 25235 4265 25265 4285
rect 25285 4265 25315 4285
rect 25335 4265 25365 4285
rect 25385 4265 25415 4285
rect 25435 4265 25465 4285
rect 25485 4265 25515 4285
rect 25535 4265 25565 4285
rect 25585 4265 25615 4285
rect 25635 4265 25665 4285
rect 25685 4265 25715 4285
rect 25735 4265 25765 4285
rect 25785 4265 25815 4285
rect 25835 4265 25865 4285
rect 25885 4265 25915 4285
rect 25935 4265 25965 4285
rect 25985 4265 26015 4285
rect 26035 4265 26065 4285
rect 26085 4265 26115 4285
rect 26135 4265 26165 4285
rect 26185 4265 26215 4285
rect 26235 4265 26265 4285
rect 26285 4265 26315 4285
rect 26335 4265 26365 4285
rect 26385 4265 26415 4285
rect 26435 4265 26465 4285
rect 26485 4265 26515 4285
rect 26535 4265 26565 4285
rect 26585 4265 26615 4285
rect 26635 4265 26665 4285
rect 26685 4265 26715 4285
rect 26735 4265 26765 4285
rect 26785 4265 26815 4285
rect 26835 4265 26865 4285
rect 26885 4265 26915 4285
rect 26935 4265 26965 4285
rect 26985 4265 27015 4285
rect 27035 4265 27065 4285
rect 27085 4265 27115 4285
rect 27135 4265 27165 4285
rect 27185 4265 27215 4285
rect 27235 4265 27265 4285
rect 27285 4265 27315 4285
rect 27335 4265 27365 4285
rect 27385 4265 27415 4285
rect 27435 4265 27465 4285
rect 27485 4265 27515 4285
rect 27535 4265 27565 4285
rect 27585 4265 27615 4285
rect 27635 4265 27665 4285
rect 27685 4265 27715 4285
rect 27735 4265 27765 4285
rect 27785 4265 27815 4285
rect 27835 4265 27865 4285
rect 27885 4265 27915 4285
rect 27935 4265 27965 4285
rect 27985 4265 28015 4285
rect 28035 4265 28065 4285
rect 28085 4265 28115 4285
rect 28135 4265 28165 4285
rect 28185 4265 28215 4285
rect 28235 4265 28265 4285
rect 28285 4265 28315 4285
rect 28335 4265 28365 4285
rect 28385 4265 28415 4285
rect 28435 4265 28465 4285
rect 28485 4265 28515 4285
rect 28535 4265 28565 4285
rect 28585 4265 28615 4285
rect 28635 4265 28665 4285
rect 28685 4265 28715 4285
rect 28735 4265 28765 4285
rect 28785 4265 28815 4285
rect 28835 4265 28865 4285
rect 28885 4265 28915 4285
rect 28935 4265 28965 4285
rect 28985 4265 29015 4285
rect 29035 4265 29065 4285
rect 29085 4265 29115 4285
rect 29135 4265 29165 4285
rect 29185 4265 29215 4285
rect 29235 4265 29265 4285
rect 29285 4265 29315 4285
rect 29335 4265 29365 4285
rect 29385 4265 29415 4285
rect 29435 4265 29465 4285
rect 29485 4265 29515 4285
rect 29535 4265 29565 4285
rect 29585 4265 29615 4285
rect 29635 4265 29665 4285
rect 29685 4265 29715 4285
rect 29735 4265 29765 4285
rect 29785 4265 29815 4285
rect 29835 4265 29865 4285
rect 29885 4265 29915 4285
rect 29935 4265 29965 4285
rect 29985 4265 30015 4285
rect 30035 4265 30065 4285
rect 30085 4265 30115 4285
rect 30135 4265 30165 4285
rect 30185 4265 30215 4285
rect 30235 4265 30265 4285
rect 30285 4265 30315 4285
rect 30335 4265 30365 4285
rect 30385 4265 30415 4285
rect 30435 4265 30465 4285
rect 30485 4265 30515 4285
rect 30535 4265 30565 4285
rect 30585 4265 30615 4285
rect 30635 4265 30665 4285
rect 30685 4265 30715 4285
rect 30735 4265 30765 4285
rect 30785 4265 30815 4285
rect 30835 4265 30865 4285
rect 30885 4265 30915 4285
rect 30935 4265 30965 4285
rect 30985 4265 31015 4285
rect 31035 4265 31065 4285
rect 31085 4265 31115 4285
rect 31135 4265 31165 4285
rect 31185 4265 31215 4285
rect 31235 4265 31265 4285
rect 31285 4265 31315 4285
rect 31335 4265 31365 4285
rect 31385 4265 31415 4285
rect 31435 4265 31465 4285
rect 31485 4265 31515 4285
rect 31535 4265 31565 4285
rect 31585 4265 31615 4285
rect 31635 4265 31665 4285
rect 31685 4265 31715 4285
rect 31735 4265 31765 4285
rect 31785 4265 31815 4285
rect 31835 4265 31865 4285
rect 31885 4265 31915 4285
rect 31935 4265 31965 4285
rect 31985 4265 32015 4285
rect 32035 4265 32065 4285
rect 32085 4265 32100 4285
rect -650 4250 32100 4265
rect -650 2985 32100 3000
rect -650 2965 -635 2985
rect -615 2965 -585 2985
rect -565 2965 -535 2985
rect -515 2965 -485 2985
rect -465 2965 -435 2985
rect -415 2965 -385 2985
rect -365 2965 -335 2985
rect -315 2965 -285 2985
rect -265 2965 -235 2985
rect -215 2965 -185 2985
rect -165 2965 -135 2985
rect -115 2965 -85 2985
rect -65 2965 -35 2985
rect -15 2965 15 2985
rect 35 2965 65 2985
rect 85 2965 115 2985
rect 135 2965 165 2985
rect 185 2965 215 2985
rect 235 2965 265 2985
rect 285 2965 315 2985
rect 335 2965 365 2985
rect 385 2965 415 2985
rect 435 2965 465 2985
rect 485 2965 515 2985
rect 535 2965 565 2985
rect 585 2965 615 2985
rect 635 2965 665 2985
rect 685 2965 715 2985
rect 735 2965 765 2985
rect 785 2965 815 2985
rect 835 2965 865 2985
rect 885 2965 915 2985
rect 935 2965 965 2985
rect 985 2965 1015 2985
rect 1035 2965 1065 2985
rect 1085 2965 1115 2985
rect 1135 2965 1165 2985
rect 1185 2965 1215 2985
rect 1235 2965 1265 2985
rect 1285 2965 1315 2985
rect 1335 2965 1365 2985
rect 1385 2965 1415 2985
rect 1435 2965 1465 2985
rect 1485 2965 1515 2985
rect 1535 2965 1565 2985
rect 1585 2965 1615 2985
rect 1635 2965 1665 2985
rect 1685 2965 1715 2985
rect 1735 2965 1765 2985
rect 1785 2965 1815 2985
rect 1835 2965 1865 2985
rect 1885 2965 1915 2985
rect 1935 2965 1965 2985
rect 1985 2965 2015 2985
rect 2035 2965 2065 2985
rect 2085 2965 2115 2985
rect 2135 2965 2165 2985
rect 2185 2965 2215 2985
rect 2235 2965 2265 2985
rect 2285 2965 2315 2985
rect 2335 2965 2365 2985
rect 2385 2965 2415 2985
rect 2435 2965 2465 2985
rect 2485 2965 2515 2985
rect 2535 2965 2565 2985
rect 2585 2965 2615 2985
rect 2635 2965 2665 2985
rect 2685 2965 2715 2985
rect 2735 2965 2765 2985
rect 2785 2965 2815 2985
rect 2835 2965 2865 2985
rect 2885 2965 2915 2985
rect 2935 2965 2965 2985
rect 2985 2965 3015 2985
rect 3035 2965 3065 2985
rect 3085 2965 3115 2985
rect 3135 2965 3165 2985
rect 3185 2965 3215 2985
rect 3235 2965 3265 2985
rect 3285 2965 3315 2985
rect 3335 2965 3365 2985
rect 3385 2965 3415 2985
rect 3435 2965 3465 2985
rect 3485 2965 3515 2985
rect 3535 2965 3565 2985
rect 3585 2965 3615 2985
rect 3635 2965 3665 2985
rect 3685 2965 3715 2985
rect 3735 2965 3765 2985
rect 3785 2965 3815 2985
rect 3835 2965 3865 2985
rect 3885 2965 3915 2985
rect 3935 2965 3965 2985
rect 3985 2965 4015 2985
rect 4035 2965 4065 2985
rect 4085 2965 4115 2985
rect 4135 2965 4165 2985
rect 4185 2965 4215 2985
rect 4235 2965 4265 2985
rect 4285 2965 4315 2985
rect 4335 2965 4365 2985
rect 4385 2965 4415 2985
rect 4435 2965 4465 2985
rect 4485 2965 4515 2985
rect 4535 2965 4565 2985
rect 4585 2965 4615 2985
rect 4635 2965 4665 2985
rect 4685 2965 4715 2985
rect 4735 2965 4765 2985
rect 4785 2965 4815 2985
rect 4835 2965 4865 2985
rect 4885 2965 4915 2985
rect 4935 2965 4965 2985
rect 4985 2965 5015 2985
rect 5035 2965 5065 2985
rect 5085 2965 5115 2985
rect 5135 2965 5165 2985
rect 5185 2965 5215 2985
rect 5235 2965 5265 2985
rect 5285 2965 5315 2985
rect 5335 2965 5365 2985
rect 5385 2965 5415 2985
rect 5435 2965 5465 2985
rect 5485 2965 5515 2985
rect 5535 2965 5565 2985
rect 5585 2965 5615 2985
rect 5635 2965 5665 2985
rect 5685 2965 5715 2985
rect 5735 2965 5765 2985
rect 5785 2965 5815 2985
rect 5835 2965 5865 2985
rect 5885 2965 5915 2985
rect 5935 2965 5965 2985
rect 5985 2965 6015 2985
rect 6035 2965 6065 2985
rect 6085 2965 6115 2985
rect 6135 2965 6165 2985
rect 6185 2965 6215 2985
rect 6235 2965 6265 2985
rect 6285 2965 6315 2985
rect 6335 2965 6365 2985
rect 6385 2965 6415 2985
rect 6435 2965 6465 2985
rect 6485 2965 6515 2985
rect 6535 2965 6565 2985
rect 6585 2965 6615 2985
rect 6635 2965 6665 2985
rect 6685 2965 6715 2985
rect 6735 2965 6765 2985
rect 6785 2965 6815 2985
rect 6835 2965 6865 2985
rect 6885 2965 6915 2985
rect 6935 2965 6965 2985
rect 6985 2965 7015 2985
rect 7035 2965 7065 2985
rect 7085 2965 7115 2985
rect 7135 2965 7165 2985
rect 7185 2965 7215 2985
rect 7235 2965 7265 2985
rect 7285 2965 7315 2985
rect 7335 2965 7365 2985
rect 7385 2965 7415 2985
rect 7435 2965 7465 2985
rect 7485 2965 7515 2985
rect 7535 2965 7565 2985
rect 7585 2965 7615 2985
rect 7635 2965 7665 2985
rect 7685 2965 7715 2985
rect 7735 2965 7765 2985
rect 7785 2965 7815 2985
rect 7835 2965 7865 2985
rect 7885 2965 7915 2985
rect 7935 2965 7965 2985
rect 7985 2965 8015 2985
rect 8035 2965 8065 2985
rect 8085 2965 8115 2985
rect 8135 2965 8165 2985
rect 8185 2965 8215 2985
rect 8235 2965 8265 2985
rect 8285 2965 8315 2985
rect 8335 2965 8365 2985
rect 8385 2965 8415 2985
rect 8435 2965 8465 2985
rect 8485 2965 8515 2985
rect 8535 2965 8565 2985
rect 8585 2965 8615 2985
rect 8635 2965 8665 2985
rect 8685 2965 8715 2985
rect 8735 2965 8765 2985
rect 8785 2965 8815 2985
rect 8835 2965 8865 2985
rect 8885 2965 8915 2985
rect 8935 2965 8965 2985
rect 8985 2965 9015 2985
rect 9035 2965 9065 2985
rect 9085 2965 9115 2985
rect 9135 2965 9165 2985
rect 9185 2965 9215 2985
rect 9235 2965 9265 2985
rect 9285 2965 9315 2985
rect 9335 2965 9365 2985
rect 9385 2965 9415 2985
rect 9435 2965 9465 2985
rect 9485 2965 9515 2985
rect 9535 2965 9565 2985
rect 9585 2965 9615 2985
rect 9635 2965 9665 2985
rect 9685 2965 9715 2985
rect 9735 2965 9765 2985
rect 9785 2965 9815 2985
rect 9835 2965 9865 2985
rect 9885 2965 9915 2985
rect 9935 2965 9965 2985
rect 9985 2965 10015 2985
rect 10035 2965 10065 2985
rect 10085 2965 10115 2985
rect 10135 2965 10165 2985
rect 10185 2965 10215 2985
rect 10235 2965 10265 2985
rect 10285 2965 10315 2985
rect 10335 2965 10365 2985
rect 10385 2965 10415 2985
rect 10435 2965 10465 2985
rect 10485 2965 10515 2985
rect 10535 2965 10565 2985
rect 10585 2965 10615 2985
rect 10635 2965 10665 2985
rect 10685 2965 10715 2985
rect 10735 2965 10765 2985
rect 10785 2965 10815 2985
rect 10835 2965 10865 2985
rect 10885 2965 10915 2985
rect 10935 2965 10965 2985
rect 10985 2965 11015 2985
rect 11035 2965 11065 2985
rect 11085 2965 11115 2985
rect 11135 2965 11165 2985
rect 11185 2965 11215 2985
rect 11235 2965 11265 2985
rect 11285 2965 11315 2985
rect 11335 2965 11365 2985
rect 11385 2965 11415 2985
rect 11435 2965 11465 2985
rect 11485 2965 11515 2985
rect 11535 2965 11565 2985
rect 11585 2965 11615 2985
rect 11635 2965 11665 2985
rect 11685 2965 11715 2985
rect 11735 2965 11765 2985
rect 11785 2965 11815 2985
rect 11835 2965 11865 2985
rect 11885 2965 11915 2985
rect 11935 2965 11965 2985
rect 11985 2965 12015 2985
rect 12035 2965 12065 2985
rect 12085 2965 12115 2985
rect 12135 2965 12165 2985
rect 12185 2965 12215 2985
rect 12235 2965 12265 2985
rect 12285 2965 12315 2985
rect 12335 2965 12365 2985
rect 12385 2965 12415 2985
rect 12435 2965 12465 2985
rect 12485 2965 12515 2985
rect 12535 2965 12565 2985
rect 12585 2965 12615 2985
rect 12635 2965 12665 2985
rect 12685 2965 12715 2985
rect 12735 2965 12765 2985
rect 12785 2965 12815 2985
rect 12835 2965 12865 2985
rect 12885 2965 12915 2985
rect 12935 2965 12965 2985
rect 12985 2965 13015 2985
rect 13035 2965 13065 2985
rect 13085 2965 13115 2985
rect 13135 2965 13165 2985
rect 13185 2965 13215 2985
rect 13235 2965 13265 2985
rect 13285 2965 13315 2985
rect 13335 2965 13365 2985
rect 13385 2965 13415 2985
rect 13435 2965 13465 2985
rect 13485 2965 13515 2985
rect 13535 2965 13565 2985
rect 13585 2965 13615 2985
rect 13635 2965 13665 2985
rect 13685 2965 13715 2985
rect 13735 2965 13765 2985
rect 13785 2965 13815 2985
rect 13835 2965 13865 2985
rect 13885 2965 13915 2985
rect 13935 2965 13965 2985
rect 13985 2965 14015 2985
rect 14035 2965 14065 2985
rect 14085 2965 14115 2985
rect 14135 2965 14165 2985
rect 14185 2965 14215 2985
rect 14235 2965 14265 2985
rect 14285 2965 14315 2985
rect 14335 2965 14365 2985
rect 14385 2965 14415 2985
rect 14435 2965 14465 2985
rect 14485 2965 14515 2985
rect 14535 2965 14565 2985
rect 14585 2965 14615 2985
rect 14635 2965 14665 2985
rect 14685 2965 14715 2985
rect 14735 2965 14765 2985
rect 14785 2965 14815 2985
rect 14835 2965 14865 2985
rect 14885 2965 14915 2985
rect 14935 2965 14965 2985
rect 14985 2965 15015 2985
rect 15035 2965 15065 2985
rect 15085 2965 15115 2985
rect 15135 2965 15165 2985
rect 15185 2965 15215 2985
rect 15235 2965 15265 2985
rect 15285 2965 15315 2985
rect 15335 2965 15365 2985
rect 15385 2965 15415 2985
rect 15435 2965 15465 2985
rect 15485 2965 15515 2985
rect 15535 2965 15565 2985
rect 15585 2965 15615 2985
rect 15635 2965 15665 2985
rect 15685 2965 15715 2985
rect 15735 2965 15765 2985
rect 15785 2965 15815 2985
rect 15835 2965 15865 2985
rect 15885 2965 15915 2985
rect 15935 2965 15965 2985
rect 15985 2965 16015 2985
rect 16035 2965 16065 2985
rect 16085 2965 16115 2985
rect 16135 2965 16165 2985
rect 16185 2965 16215 2985
rect 16235 2965 16265 2985
rect 16285 2965 16315 2985
rect 16335 2965 16365 2985
rect 16385 2965 16415 2985
rect 16435 2965 16465 2985
rect 16485 2965 16515 2985
rect 16535 2965 16565 2985
rect 16585 2965 16615 2985
rect 16635 2965 16665 2985
rect 16685 2965 16715 2985
rect 16735 2965 16765 2985
rect 16785 2965 16815 2985
rect 16835 2965 16865 2985
rect 16885 2965 16915 2985
rect 16935 2965 16965 2985
rect 16985 2965 17015 2985
rect 17035 2965 17065 2985
rect 17085 2965 17115 2985
rect 17135 2965 17165 2985
rect 17185 2965 17215 2985
rect 17235 2965 17265 2985
rect 17285 2965 17315 2985
rect 17335 2965 17365 2985
rect 17385 2965 17415 2985
rect 17435 2965 17465 2985
rect 17485 2965 17515 2985
rect 17535 2965 17565 2985
rect 17585 2965 17615 2985
rect 17635 2965 17665 2985
rect 17685 2965 17715 2985
rect 17735 2965 17765 2985
rect 17785 2965 17815 2985
rect 17835 2965 17865 2985
rect 17885 2965 17915 2985
rect 17935 2965 17965 2985
rect 17985 2965 18015 2985
rect 18035 2965 18065 2985
rect 18085 2965 18115 2985
rect 18135 2965 18165 2985
rect 18185 2965 18215 2985
rect 18235 2965 18265 2985
rect 18285 2965 18315 2985
rect 18335 2965 18365 2985
rect 18385 2965 18415 2985
rect 18435 2965 18465 2985
rect 18485 2965 18515 2985
rect 18535 2965 18565 2985
rect 18585 2965 18615 2985
rect 18635 2965 18665 2985
rect 18685 2965 18715 2985
rect 18735 2965 18765 2985
rect 18785 2965 18815 2985
rect 18835 2965 18865 2985
rect 18885 2965 18915 2985
rect 18935 2965 18965 2985
rect 18985 2965 19015 2985
rect 19035 2965 19065 2985
rect 19085 2965 19115 2985
rect 19135 2965 19165 2985
rect 19185 2965 19215 2985
rect 19235 2965 19265 2985
rect 19285 2965 19315 2985
rect 19335 2965 19365 2985
rect 19385 2965 19415 2985
rect 19435 2965 19465 2985
rect 19485 2965 19515 2985
rect 19535 2965 19565 2985
rect 19585 2965 19615 2985
rect 19635 2965 19665 2985
rect 19685 2965 19715 2985
rect 19735 2965 19765 2985
rect 19785 2965 19815 2985
rect 19835 2965 19865 2985
rect 19885 2965 19915 2985
rect 19935 2965 19965 2985
rect 19985 2965 20015 2985
rect 20035 2965 20065 2985
rect 20085 2965 20115 2985
rect 20135 2965 20165 2985
rect 20185 2965 20215 2985
rect 20235 2965 20265 2985
rect 20285 2965 20315 2985
rect 20335 2965 20365 2985
rect 20385 2965 20415 2985
rect 20435 2965 20465 2985
rect 20485 2965 20515 2985
rect 20535 2965 20565 2985
rect 20585 2965 20615 2985
rect 20635 2965 20665 2985
rect 20685 2965 20715 2985
rect 20735 2965 20765 2985
rect 20785 2965 20815 2985
rect 20835 2965 20865 2985
rect 20885 2965 20915 2985
rect 20935 2965 20965 2985
rect 20985 2965 21015 2985
rect 21035 2965 21065 2985
rect 21085 2965 21115 2985
rect 21135 2965 21165 2985
rect 21185 2965 21215 2985
rect 21235 2965 21265 2985
rect 21285 2965 21315 2985
rect 21335 2965 21365 2985
rect 21385 2965 21415 2985
rect 21435 2965 21465 2985
rect 21485 2965 21515 2985
rect 21535 2965 21565 2985
rect 21585 2965 21615 2985
rect 21635 2965 21665 2985
rect 21685 2965 21715 2985
rect 21735 2965 21765 2985
rect 21785 2965 21815 2985
rect 21835 2965 21865 2985
rect 21885 2965 21915 2985
rect 21935 2965 21965 2985
rect 21985 2965 22015 2985
rect 22035 2965 22065 2985
rect 22085 2965 22115 2985
rect 22135 2965 22165 2985
rect 22185 2965 22215 2985
rect 22235 2965 22265 2985
rect 22285 2965 22315 2985
rect 22335 2965 22365 2985
rect 22385 2965 22415 2985
rect 22435 2965 22465 2985
rect 22485 2965 22515 2985
rect 22535 2965 22565 2985
rect 22585 2965 22615 2985
rect 22635 2965 22665 2985
rect 22685 2965 22715 2985
rect 22735 2965 22765 2985
rect 22785 2965 22815 2985
rect 22835 2965 22865 2985
rect 22885 2965 22915 2985
rect 22935 2965 22965 2985
rect 22985 2965 23015 2985
rect 23035 2965 23065 2985
rect 23085 2965 23115 2985
rect 23135 2965 23165 2985
rect 23185 2965 23215 2985
rect 23235 2965 23265 2985
rect 23285 2965 23315 2985
rect 23335 2965 23365 2985
rect 23385 2965 23415 2985
rect 23435 2965 23465 2985
rect 23485 2965 23515 2985
rect 23535 2965 23565 2985
rect 23585 2965 23615 2985
rect 23635 2965 23665 2985
rect 23685 2965 23715 2985
rect 23735 2965 23765 2985
rect 23785 2965 23815 2985
rect 23835 2965 23865 2985
rect 23885 2965 23915 2985
rect 23935 2965 23965 2985
rect 23985 2965 24015 2985
rect 24035 2965 24065 2985
rect 24085 2965 24115 2985
rect 24135 2965 24165 2985
rect 24185 2965 24215 2985
rect 24235 2965 24265 2985
rect 24285 2965 24315 2985
rect 24335 2965 24365 2985
rect 24385 2965 24415 2985
rect 24435 2965 24465 2985
rect 24485 2965 24515 2985
rect 24535 2965 24565 2985
rect 24585 2965 24615 2985
rect 24635 2965 24665 2985
rect 24685 2965 24715 2985
rect 24735 2965 24765 2985
rect 24785 2965 24815 2985
rect 24835 2965 24865 2985
rect 24885 2965 24915 2985
rect 24935 2965 24965 2985
rect 24985 2965 25015 2985
rect 25035 2965 25065 2985
rect 25085 2965 25115 2985
rect 25135 2965 25165 2985
rect 25185 2965 25215 2985
rect 25235 2965 25265 2985
rect 25285 2965 25315 2985
rect 25335 2965 25365 2985
rect 25385 2965 25415 2985
rect 25435 2965 25465 2985
rect 25485 2965 25515 2985
rect 25535 2965 25565 2985
rect 25585 2965 25615 2985
rect 25635 2965 25665 2985
rect 25685 2965 25715 2985
rect 25735 2965 25765 2985
rect 25785 2965 25815 2985
rect 25835 2965 25865 2985
rect 25885 2965 25915 2985
rect 25935 2965 25965 2985
rect 25985 2965 26015 2985
rect 26035 2965 26065 2985
rect 26085 2965 26115 2985
rect 26135 2965 26165 2985
rect 26185 2965 26215 2985
rect 26235 2965 26265 2985
rect 26285 2965 26315 2985
rect 26335 2965 26365 2985
rect 26385 2965 26415 2985
rect 26435 2965 26465 2985
rect 26485 2965 26515 2985
rect 26535 2965 26565 2985
rect 26585 2965 26615 2985
rect 26635 2965 26665 2985
rect 26685 2965 26715 2985
rect 26735 2965 26765 2985
rect 26785 2965 26815 2985
rect 26835 2965 26865 2985
rect 26885 2965 26915 2985
rect 26935 2965 26965 2985
rect 26985 2965 27015 2985
rect 27035 2965 27065 2985
rect 27085 2965 27115 2985
rect 27135 2965 27165 2985
rect 27185 2965 27215 2985
rect 27235 2965 27265 2985
rect 27285 2965 27315 2985
rect 27335 2965 27365 2985
rect 27385 2965 27415 2985
rect 27435 2965 27465 2985
rect 27485 2965 27515 2985
rect 27535 2965 27565 2985
rect 27585 2965 27615 2985
rect 27635 2965 27665 2985
rect 27685 2965 27715 2985
rect 27735 2965 27765 2985
rect 27785 2965 27815 2985
rect 27835 2965 27865 2985
rect 27885 2965 27915 2985
rect 27935 2965 27965 2985
rect 27985 2965 28015 2985
rect 28035 2965 28065 2985
rect 28085 2965 28115 2985
rect 28135 2965 28165 2985
rect 28185 2965 28215 2985
rect 28235 2965 28265 2985
rect 28285 2965 28315 2985
rect 28335 2965 28365 2985
rect 28385 2965 28415 2985
rect 28435 2965 28465 2985
rect 28485 2965 28515 2985
rect 28535 2965 28565 2985
rect 28585 2965 28615 2985
rect 28635 2965 28665 2985
rect 28685 2965 28715 2985
rect 28735 2965 28765 2985
rect 28785 2965 28815 2985
rect 28835 2965 28865 2985
rect 28885 2965 28915 2985
rect 28935 2965 28965 2985
rect 28985 2965 29015 2985
rect 29035 2965 29065 2985
rect 29085 2965 29115 2985
rect 29135 2965 29165 2985
rect 29185 2965 29215 2985
rect 29235 2965 29265 2985
rect 29285 2965 29315 2985
rect 29335 2965 29365 2985
rect 29385 2965 29415 2985
rect 29435 2965 29465 2985
rect 29485 2965 29515 2985
rect 29535 2965 29565 2985
rect 29585 2965 29615 2985
rect 29635 2965 29665 2985
rect 29685 2965 29715 2985
rect 29735 2965 29765 2985
rect 29785 2965 29815 2985
rect 29835 2965 29865 2985
rect 29885 2965 29915 2985
rect 29935 2965 29965 2985
rect 29985 2965 30015 2985
rect 30035 2965 30065 2985
rect 30085 2965 30115 2985
rect 30135 2965 30165 2985
rect 30185 2965 30215 2985
rect 30235 2965 30265 2985
rect 30285 2965 30315 2985
rect 30335 2965 30365 2985
rect 30385 2965 30415 2985
rect 30435 2965 30465 2985
rect 30485 2965 30515 2985
rect 30535 2965 30565 2985
rect 30585 2965 30615 2985
rect 30635 2965 30665 2985
rect 30685 2965 30715 2985
rect 30735 2965 30765 2985
rect 30785 2965 30815 2985
rect 30835 2965 30865 2985
rect 30885 2965 30915 2985
rect 30935 2965 30965 2985
rect 30985 2965 31015 2985
rect 31035 2965 31065 2985
rect 31085 2965 31115 2985
rect 31135 2965 31165 2985
rect 31185 2965 31215 2985
rect 31235 2965 31265 2985
rect 31285 2965 31315 2985
rect 31335 2965 31365 2985
rect 31385 2965 31415 2985
rect 31435 2965 31465 2985
rect 31485 2965 31515 2985
rect 31535 2965 31565 2985
rect 31585 2965 31615 2985
rect 31635 2965 31665 2985
rect 31685 2965 31715 2985
rect 31735 2965 31765 2985
rect 31785 2965 31815 2985
rect 31835 2965 31865 2985
rect 31885 2965 31915 2985
rect 31935 2965 31965 2985
rect 31985 2965 32015 2985
rect 32035 2965 32065 2985
rect 32085 2965 32100 2985
rect -650 2950 32100 2965
rect -650 1835 28800 1850
rect -650 1815 -635 1835
rect -615 1815 -585 1835
rect -565 1815 -535 1835
rect -515 1815 -485 1835
rect -465 1815 -435 1835
rect -415 1815 -385 1835
rect -365 1815 -335 1835
rect -315 1815 -285 1835
rect -265 1815 -235 1835
rect -215 1815 -185 1835
rect -165 1815 -135 1835
rect -115 1815 -85 1835
rect -65 1815 -35 1835
rect -15 1815 15 1835
rect 35 1815 65 1835
rect 85 1815 115 1835
rect 135 1815 165 1835
rect 185 1815 215 1835
rect 235 1815 265 1835
rect 285 1815 315 1835
rect 335 1815 365 1835
rect 385 1815 415 1835
rect 435 1815 465 1835
rect 485 1815 515 1835
rect 535 1815 565 1835
rect 585 1815 615 1835
rect 635 1815 665 1835
rect 685 1815 715 1835
rect 735 1815 765 1835
rect 785 1815 815 1835
rect 835 1815 865 1835
rect 885 1815 915 1835
rect 935 1815 965 1835
rect 985 1815 1015 1835
rect 1035 1815 1065 1835
rect 1085 1815 1115 1835
rect 1135 1815 1165 1835
rect 1185 1815 1215 1835
rect 1235 1815 1265 1835
rect 1285 1815 1315 1835
rect 1335 1815 1365 1835
rect 1385 1815 1415 1835
rect 1435 1815 1465 1835
rect 1485 1815 1515 1835
rect 1535 1815 1565 1835
rect 1585 1815 1615 1835
rect 1635 1815 1665 1835
rect 1685 1815 1715 1835
rect 1735 1815 1765 1835
rect 1785 1815 1815 1835
rect 1835 1815 1865 1835
rect 1885 1815 1915 1835
rect 1935 1815 1965 1835
rect 1985 1815 2015 1835
rect 2035 1815 2065 1835
rect 2085 1815 2115 1835
rect 2135 1815 2165 1835
rect 2185 1815 2215 1835
rect 2235 1815 2265 1835
rect 2285 1815 2315 1835
rect 2335 1815 2365 1835
rect 2385 1815 2415 1835
rect 2435 1815 2465 1835
rect 2485 1815 2515 1835
rect 2535 1815 2565 1835
rect 2585 1815 2615 1835
rect 2635 1815 2665 1835
rect 2685 1815 2715 1835
rect 2735 1815 2765 1835
rect 2785 1815 2815 1835
rect 2835 1815 2865 1835
rect 2885 1815 2915 1835
rect 2935 1815 2965 1835
rect 2985 1815 3015 1835
rect 3035 1815 3065 1835
rect 3085 1815 3115 1835
rect 3135 1815 3165 1835
rect 3185 1815 3215 1835
rect 3235 1815 3265 1835
rect 3285 1815 3315 1835
rect 3335 1815 3365 1835
rect 3385 1815 3415 1835
rect 3435 1815 3465 1835
rect 3485 1815 3515 1835
rect 3535 1815 3565 1835
rect 3585 1815 3615 1835
rect 3635 1815 3665 1835
rect 3685 1815 3715 1835
rect 3735 1815 3765 1835
rect 3785 1815 3815 1835
rect 3835 1815 3865 1835
rect 3885 1815 3915 1835
rect 3935 1815 3965 1835
rect 3985 1815 4015 1835
rect 4035 1815 4065 1835
rect 4085 1815 4115 1835
rect 4135 1815 4165 1835
rect 4185 1815 4215 1835
rect 4235 1815 4265 1835
rect 4285 1815 4315 1835
rect 4335 1815 4365 1835
rect 4385 1815 4415 1835
rect 4435 1815 4465 1835
rect 4485 1815 4515 1835
rect 4535 1815 4565 1835
rect 4585 1815 4615 1835
rect 4635 1815 4665 1835
rect 4685 1815 4715 1835
rect 4735 1815 4765 1835
rect 4785 1815 4815 1835
rect 4835 1815 4865 1835
rect 4885 1815 4915 1835
rect 4935 1815 4965 1835
rect 4985 1815 5015 1835
rect 5035 1815 5065 1835
rect 5085 1815 5115 1835
rect 5135 1815 5165 1835
rect 5185 1815 5215 1835
rect 5235 1815 5265 1835
rect 5285 1815 5315 1835
rect 5335 1815 5365 1835
rect 5385 1815 5415 1835
rect 5435 1815 5465 1835
rect 5485 1815 5515 1835
rect 5535 1815 5565 1835
rect 5585 1815 5615 1835
rect 5635 1815 5665 1835
rect 5685 1815 5715 1835
rect 5735 1815 5765 1835
rect 5785 1815 5815 1835
rect 5835 1815 5865 1835
rect 5885 1815 5915 1835
rect 5935 1815 5965 1835
rect 5985 1815 6015 1835
rect 6035 1815 6065 1835
rect 6085 1815 6115 1835
rect 6135 1815 6165 1835
rect 6185 1815 6215 1835
rect 6235 1815 6265 1835
rect 6285 1815 6315 1835
rect 6335 1815 6365 1835
rect 6385 1815 6415 1835
rect 6435 1815 6465 1835
rect 6485 1815 6515 1835
rect 6535 1815 6565 1835
rect 6585 1815 6615 1835
rect 6635 1815 6665 1835
rect 6685 1815 6715 1835
rect 6735 1815 6765 1835
rect 6785 1815 6815 1835
rect 6835 1815 6865 1835
rect 6885 1815 6915 1835
rect 6935 1815 6965 1835
rect 6985 1815 7015 1835
rect 7035 1815 7065 1835
rect 7085 1815 7115 1835
rect 7135 1815 7165 1835
rect 7185 1815 7215 1835
rect 7235 1815 7265 1835
rect 7285 1815 7315 1835
rect 7335 1815 7365 1835
rect 7385 1815 7415 1835
rect 7435 1815 7465 1835
rect 7485 1815 7515 1835
rect 7535 1815 7565 1835
rect 7585 1815 7615 1835
rect 7635 1815 7665 1835
rect 7685 1815 7715 1835
rect 7735 1815 7765 1835
rect 7785 1815 7815 1835
rect 7835 1815 7865 1835
rect 7885 1815 7915 1835
rect 7935 1815 7965 1835
rect 7985 1815 8015 1835
rect 8035 1815 8065 1835
rect 8085 1815 8115 1835
rect 8135 1815 8165 1835
rect 8185 1815 8215 1835
rect 8235 1815 8265 1835
rect 8285 1815 8315 1835
rect 8335 1815 8365 1835
rect 8385 1815 8415 1835
rect 8435 1815 8465 1835
rect 8485 1815 8515 1835
rect 8535 1815 8565 1835
rect 8585 1815 8615 1835
rect 8635 1815 8665 1835
rect 8685 1815 8715 1835
rect 8735 1815 8765 1835
rect 8785 1815 8815 1835
rect 8835 1815 8865 1835
rect 8885 1815 8915 1835
rect 8935 1815 8965 1835
rect 8985 1815 9015 1835
rect 9035 1815 9065 1835
rect 9085 1815 9115 1835
rect 9135 1815 9165 1835
rect 9185 1815 9215 1835
rect 9235 1815 9265 1835
rect 9285 1815 9315 1835
rect 9335 1815 9365 1835
rect 9385 1815 9415 1835
rect 9435 1815 9465 1835
rect 9485 1815 9515 1835
rect 9535 1815 9565 1835
rect 9585 1815 9615 1835
rect 9635 1815 9665 1835
rect 9685 1815 9715 1835
rect 9735 1815 9765 1835
rect 9785 1815 9815 1835
rect 9835 1815 9865 1835
rect 9885 1815 9915 1835
rect 9935 1815 9965 1835
rect 9985 1815 10015 1835
rect 10035 1815 10065 1835
rect 10085 1815 10115 1835
rect 10135 1815 10165 1835
rect 10185 1815 10215 1835
rect 10235 1815 10265 1835
rect 10285 1815 10315 1835
rect 10335 1815 10365 1835
rect 10385 1815 10415 1835
rect 10435 1815 10465 1835
rect 10485 1815 10515 1835
rect 10535 1815 10565 1835
rect 10585 1815 10615 1835
rect 10635 1815 10665 1835
rect 10685 1815 10715 1835
rect 10735 1815 10765 1835
rect 10785 1815 10815 1835
rect 10835 1815 10865 1835
rect 10885 1815 10915 1835
rect 10935 1815 10965 1835
rect 10985 1815 11015 1835
rect 11035 1815 11065 1835
rect 11085 1815 11115 1835
rect 11135 1815 11165 1835
rect 11185 1815 11215 1835
rect 11235 1815 11265 1835
rect 11285 1815 11315 1835
rect 11335 1815 11365 1835
rect 11385 1815 11415 1835
rect 11435 1815 11465 1835
rect 11485 1815 11515 1835
rect 11535 1815 11565 1835
rect 11585 1815 11615 1835
rect 11635 1815 11665 1835
rect 11685 1815 11715 1835
rect 11735 1815 11765 1835
rect 11785 1815 11815 1835
rect 11835 1815 11865 1835
rect 11885 1815 11915 1835
rect 11935 1815 11965 1835
rect 11985 1815 12015 1835
rect 12035 1815 12065 1835
rect 12085 1815 12115 1835
rect 12135 1815 12165 1835
rect 12185 1815 12215 1835
rect 12235 1815 12265 1835
rect 12285 1815 12315 1835
rect 12335 1815 12365 1835
rect 12385 1815 12415 1835
rect 12435 1815 12465 1835
rect 12485 1815 12515 1835
rect 12535 1815 12565 1835
rect 12585 1815 12615 1835
rect 12635 1815 12665 1835
rect 12685 1815 12715 1835
rect 12735 1815 12765 1835
rect 12785 1815 12815 1835
rect 12835 1815 12865 1835
rect 12885 1815 12915 1835
rect 12935 1815 12965 1835
rect 12985 1815 13015 1835
rect 13035 1815 13065 1835
rect 13085 1815 13115 1835
rect 13135 1815 13165 1835
rect 13185 1815 13215 1835
rect 13235 1815 13265 1835
rect 13285 1815 13315 1835
rect 13335 1815 13365 1835
rect 13385 1815 13415 1835
rect 13435 1815 13465 1835
rect 13485 1815 13515 1835
rect 13535 1815 13565 1835
rect 13585 1815 13615 1835
rect 13635 1815 13665 1835
rect 13685 1815 13715 1835
rect 13735 1815 13765 1835
rect 13785 1815 13815 1835
rect 13835 1815 13865 1835
rect 13885 1815 13915 1835
rect 13935 1815 13965 1835
rect 13985 1815 14015 1835
rect 14035 1815 14065 1835
rect 14085 1815 14115 1835
rect 14135 1815 14165 1835
rect 14185 1815 14215 1835
rect 14235 1815 14265 1835
rect 14285 1815 14315 1835
rect 14335 1815 14365 1835
rect 14385 1815 14415 1835
rect 14435 1815 14465 1835
rect 14485 1815 14515 1835
rect 14535 1815 14565 1835
rect 14585 1815 14615 1835
rect 14635 1815 14665 1835
rect 14685 1815 14715 1835
rect 14735 1815 14765 1835
rect 14785 1815 14815 1835
rect 14835 1815 14865 1835
rect 14885 1815 14915 1835
rect 14935 1815 14965 1835
rect 14985 1815 15015 1835
rect 15035 1815 15065 1835
rect 15085 1815 15115 1835
rect 15135 1815 15165 1835
rect 15185 1815 15215 1835
rect 15235 1815 15265 1835
rect 15285 1815 15315 1835
rect 15335 1815 15365 1835
rect 15385 1815 15415 1835
rect 15435 1815 15465 1835
rect 15485 1815 15515 1835
rect 15535 1815 15565 1835
rect 15585 1815 15615 1835
rect 15635 1815 15665 1835
rect 15685 1815 15715 1835
rect 15735 1815 15765 1835
rect 15785 1815 15815 1835
rect 15835 1815 15865 1835
rect 15885 1815 15915 1835
rect 15935 1815 15965 1835
rect 15985 1815 16015 1835
rect 16035 1815 16065 1835
rect 16085 1815 16115 1835
rect 16135 1815 16165 1835
rect 16185 1815 16215 1835
rect 16235 1815 16265 1835
rect 16285 1815 16315 1835
rect 16335 1815 16365 1835
rect 16385 1815 16415 1835
rect 16435 1815 16465 1835
rect 16485 1815 16515 1835
rect 16535 1815 16565 1835
rect 16585 1815 16615 1835
rect 16635 1815 16665 1835
rect 16685 1815 16715 1835
rect 16735 1815 16765 1835
rect 16785 1815 16815 1835
rect 16835 1815 16865 1835
rect 16885 1815 16915 1835
rect 16935 1815 16965 1835
rect 16985 1815 17015 1835
rect 17035 1815 17065 1835
rect 17085 1815 17115 1835
rect 17135 1815 17165 1835
rect 17185 1815 17215 1835
rect 17235 1815 17265 1835
rect 17285 1815 17315 1835
rect 17335 1815 17365 1835
rect 17385 1815 17415 1835
rect 17435 1815 17465 1835
rect 17485 1815 17515 1835
rect 17535 1815 17565 1835
rect 17585 1815 17615 1835
rect 17635 1815 17665 1835
rect 17685 1815 17715 1835
rect 17735 1815 17765 1835
rect 17785 1815 17815 1835
rect 17835 1815 17865 1835
rect 17885 1815 17915 1835
rect 17935 1815 17965 1835
rect 17985 1815 18015 1835
rect 18035 1815 18065 1835
rect 18085 1815 18115 1835
rect 18135 1815 18165 1835
rect 18185 1815 18215 1835
rect 18235 1815 18265 1835
rect 18285 1815 18315 1835
rect 18335 1815 18365 1835
rect 18385 1815 18415 1835
rect 18435 1815 18465 1835
rect 18485 1815 18515 1835
rect 18535 1815 18565 1835
rect 18585 1815 18615 1835
rect 18635 1815 18665 1835
rect 18685 1815 18715 1835
rect 18735 1815 18765 1835
rect 18785 1815 18815 1835
rect 18835 1815 18865 1835
rect 18885 1815 18915 1835
rect 18935 1815 18965 1835
rect 18985 1815 19015 1835
rect 19035 1815 19065 1835
rect 19085 1815 19115 1835
rect 19135 1815 19165 1835
rect 19185 1815 19215 1835
rect 19235 1815 19265 1835
rect 19285 1815 19315 1835
rect 19335 1815 19365 1835
rect 19385 1815 19415 1835
rect 19435 1815 19465 1835
rect 19485 1815 19515 1835
rect 19535 1815 19565 1835
rect 19585 1815 19615 1835
rect 19635 1815 19665 1835
rect 19685 1815 19715 1835
rect 19735 1815 19765 1835
rect 19785 1815 19815 1835
rect 19835 1815 19865 1835
rect 19885 1815 19915 1835
rect 19935 1815 19965 1835
rect 19985 1815 20015 1835
rect 20035 1815 20065 1835
rect 20085 1815 20115 1835
rect 20135 1815 20165 1835
rect 20185 1815 20215 1835
rect 20235 1815 20265 1835
rect 20285 1815 20315 1835
rect 20335 1815 20365 1835
rect 20385 1815 20415 1835
rect 20435 1815 20465 1835
rect 20485 1815 20515 1835
rect 20535 1815 20565 1835
rect 20585 1815 20615 1835
rect 20635 1815 20665 1835
rect 20685 1815 20715 1835
rect 20735 1815 20765 1835
rect 20785 1815 20815 1835
rect 20835 1815 20865 1835
rect 20885 1815 20915 1835
rect 20935 1815 20965 1835
rect 20985 1815 21015 1835
rect 21035 1815 21065 1835
rect 21085 1815 21115 1835
rect 21135 1815 21165 1835
rect 21185 1815 21215 1835
rect 21235 1815 21265 1835
rect 21285 1815 21315 1835
rect 21335 1815 21365 1835
rect 21385 1815 21415 1835
rect 21435 1815 21465 1835
rect 21485 1815 21515 1835
rect 21535 1815 21565 1835
rect 21585 1815 21615 1835
rect 21635 1815 21665 1835
rect 21685 1815 21715 1835
rect 21735 1815 21765 1835
rect 21785 1815 21815 1835
rect 21835 1815 21865 1835
rect 21885 1815 21915 1835
rect 21935 1815 21965 1835
rect 21985 1815 22015 1835
rect 22035 1815 22065 1835
rect 22085 1815 22115 1835
rect 22135 1815 22165 1835
rect 22185 1815 22215 1835
rect 22235 1815 22265 1835
rect 22285 1815 22315 1835
rect 22335 1815 22365 1835
rect 22385 1815 22415 1835
rect 22435 1815 22465 1835
rect 22485 1815 22515 1835
rect 22535 1815 22565 1835
rect 22585 1815 22615 1835
rect 22635 1815 22665 1835
rect 22685 1815 22715 1835
rect 22735 1815 22765 1835
rect 22785 1815 22815 1835
rect 22835 1815 22865 1835
rect 22885 1815 22915 1835
rect 22935 1815 22965 1835
rect 22985 1815 23015 1835
rect 23035 1815 23065 1835
rect 23085 1815 23115 1835
rect 23135 1815 23165 1835
rect 23185 1815 23215 1835
rect 23235 1815 23265 1835
rect 23285 1815 23315 1835
rect 23335 1815 23365 1835
rect 23385 1815 23415 1835
rect 23435 1815 23465 1835
rect 23485 1815 23515 1835
rect 23535 1815 23565 1835
rect 23585 1815 23615 1835
rect 23635 1815 23665 1835
rect 23685 1815 23715 1835
rect 23735 1815 23765 1835
rect 23785 1815 23815 1835
rect 23835 1815 23865 1835
rect 23885 1815 23915 1835
rect 23935 1815 23965 1835
rect 23985 1815 24015 1835
rect 24035 1815 24065 1835
rect 24085 1815 24115 1835
rect 24135 1815 24165 1835
rect 24185 1815 24215 1835
rect 24235 1815 24265 1835
rect 24285 1815 24315 1835
rect 24335 1815 24365 1835
rect 24385 1815 24415 1835
rect 24435 1815 24465 1835
rect 24485 1815 24515 1835
rect 24535 1815 24565 1835
rect 24585 1815 24615 1835
rect 24635 1815 24665 1835
rect 24685 1815 24715 1835
rect 24735 1815 24765 1835
rect 24785 1815 24815 1835
rect 24835 1815 24865 1835
rect 24885 1815 24915 1835
rect 24935 1815 24965 1835
rect 24985 1815 25015 1835
rect 25035 1815 25065 1835
rect 25085 1815 25115 1835
rect 25135 1815 25165 1835
rect 25185 1815 25215 1835
rect 25235 1815 25265 1835
rect 25285 1815 25315 1835
rect 25335 1815 25365 1835
rect 25385 1815 25415 1835
rect 25435 1815 25465 1835
rect 25485 1815 25515 1835
rect 25535 1815 25565 1835
rect 25585 1815 25615 1835
rect 25635 1815 25665 1835
rect 25685 1815 25715 1835
rect 25735 1815 25765 1835
rect 25785 1815 25815 1835
rect 25835 1815 25865 1835
rect 25885 1815 25915 1835
rect 25935 1815 25965 1835
rect 25985 1815 26015 1835
rect 26035 1815 26065 1835
rect 26085 1815 26115 1835
rect 26135 1815 26165 1835
rect 26185 1815 26215 1835
rect 26235 1815 26265 1835
rect 26285 1815 26315 1835
rect 26335 1815 26365 1835
rect 26385 1815 26415 1835
rect 26435 1815 26465 1835
rect 26485 1815 26515 1835
rect 26535 1815 26565 1835
rect 26585 1815 26615 1835
rect 26635 1815 26665 1835
rect 26685 1815 26715 1835
rect 26735 1815 26765 1835
rect 26785 1815 26815 1835
rect 26835 1815 26865 1835
rect 26885 1815 26915 1835
rect 26935 1815 26965 1835
rect 26985 1815 27015 1835
rect 27035 1815 27065 1835
rect 27085 1815 27115 1835
rect 27135 1815 27165 1835
rect 27185 1815 27215 1835
rect 27235 1815 27265 1835
rect 27285 1815 27315 1835
rect 27335 1815 27365 1835
rect 27385 1815 27415 1835
rect 27435 1815 27465 1835
rect 27485 1815 27515 1835
rect 27535 1815 27565 1835
rect 27585 1815 27615 1835
rect 27635 1815 27665 1835
rect 27685 1815 27715 1835
rect 27735 1815 27765 1835
rect 27785 1815 27815 1835
rect 27835 1815 27865 1835
rect 27885 1815 27915 1835
rect 27935 1815 27965 1835
rect 27985 1815 28015 1835
rect 28035 1815 28065 1835
rect 28085 1815 28115 1835
rect 28135 1815 28165 1835
rect 28185 1815 28215 1835
rect 28235 1815 28265 1835
rect 28285 1815 28315 1835
rect 28335 1815 28365 1835
rect 28385 1815 28415 1835
rect 28435 1815 28465 1835
rect 28485 1815 28515 1835
rect 28535 1815 28565 1835
rect 28585 1815 28615 1835
rect 28635 1815 28665 1835
rect 28685 1815 28715 1835
rect 28735 1815 28765 1835
rect 28785 1815 28800 1835
rect -650 1800 28800 1815
rect -650 -1865 28800 -1850
rect -650 -1885 -635 -1865
rect -615 -1885 -585 -1865
rect -565 -1885 -535 -1865
rect -515 -1885 -485 -1865
rect -465 -1885 -435 -1865
rect -415 -1885 -385 -1865
rect -365 -1885 -335 -1865
rect -315 -1885 -285 -1865
rect -265 -1885 -235 -1865
rect -215 -1885 -185 -1865
rect -165 -1885 -135 -1865
rect -115 -1885 -85 -1865
rect -65 -1885 -35 -1865
rect -15 -1885 15 -1865
rect 35 -1885 65 -1865
rect 85 -1885 115 -1865
rect 135 -1885 165 -1865
rect 185 -1885 215 -1865
rect 235 -1885 265 -1865
rect 285 -1885 315 -1865
rect 335 -1885 365 -1865
rect 385 -1885 415 -1865
rect 435 -1885 465 -1865
rect 485 -1885 515 -1865
rect 535 -1885 565 -1865
rect 585 -1885 615 -1865
rect 635 -1885 665 -1865
rect 685 -1885 715 -1865
rect 735 -1885 765 -1865
rect 785 -1885 815 -1865
rect 835 -1885 865 -1865
rect 885 -1885 915 -1865
rect 935 -1885 965 -1865
rect 985 -1885 1015 -1865
rect 1035 -1885 1065 -1865
rect 1085 -1885 1115 -1865
rect 1135 -1885 1165 -1865
rect 1185 -1885 1215 -1865
rect 1235 -1885 1265 -1865
rect 1285 -1885 1315 -1865
rect 1335 -1885 1365 -1865
rect 1385 -1885 1415 -1865
rect 1435 -1885 1465 -1865
rect 1485 -1885 1515 -1865
rect 1535 -1885 1565 -1865
rect 1585 -1885 1615 -1865
rect 1635 -1885 1665 -1865
rect 1685 -1885 1715 -1865
rect 1735 -1885 1765 -1865
rect 1785 -1885 1815 -1865
rect 1835 -1885 1865 -1865
rect 1885 -1885 1915 -1865
rect 1935 -1885 1965 -1865
rect 1985 -1885 2015 -1865
rect 2035 -1885 2065 -1865
rect 2085 -1885 2115 -1865
rect 2135 -1885 2165 -1865
rect 2185 -1885 2215 -1865
rect 2235 -1885 2265 -1865
rect 2285 -1885 2315 -1865
rect 2335 -1885 2365 -1865
rect 2385 -1885 2415 -1865
rect 2435 -1885 2465 -1865
rect 2485 -1885 2515 -1865
rect 2535 -1885 2565 -1865
rect 2585 -1885 2615 -1865
rect 2635 -1885 2665 -1865
rect 2685 -1885 2715 -1865
rect 2735 -1885 2765 -1865
rect 2785 -1885 2815 -1865
rect 2835 -1885 2865 -1865
rect 2885 -1885 2915 -1865
rect 2935 -1885 2965 -1865
rect 2985 -1885 3015 -1865
rect 3035 -1885 3065 -1865
rect 3085 -1885 3115 -1865
rect 3135 -1885 3165 -1865
rect 3185 -1885 3215 -1865
rect 3235 -1885 3265 -1865
rect 3285 -1885 3315 -1865
rect 3335 -1885 3365 -1865
rect 3385 -1885 3415 -1865
rect 3435 -1885 3465 -1865
rect 3485 -1885 3515 -1865
rect 3535 -1885 3565 -1865
rect 3585 -1885 3615 -1865
rect 3635 -1885 3665 -1865
rect 3685 -1885 3715 -1865
rect 3735 -1885 3765 -1865
rect 3785 -1885 3815 -1865
rect 3835 -1885 3865 -1865
rect 3885 -1885 3915 -1865
rect 3935 -1885 3965 -1865
rect 3985 -1885 4015 -1865
rect 4035 -1885 4065 -1865
rect 4085 -1885 4115 -1865
rect 4135 -1885 4165 -1865
rect 4185 -1885 4215 -1865
rect 4235 -1885 4265 -1865
rect 4285 -1885 4315 -1865
rect 4335 -1885 4365 -1865
rect 4385 -1885 4415 -1865
rect 4435 -1885 4465 -1865
rect 4485 -1885 4515 -1865
rect 4535 -1885 4565 -1865
rect 4585 -1885 4615 -1865
rect 4635 -1885 4665 -1865
rect 4685 -1885 4715 -1865
rect 4735 -1885 4765 -1865
rect 4785 -1885 4815 -1865
rect 4835 -1885 4865 -1865
rect 4885 -1885 4915 -1865
rect 4935 -1885 4965 -1865
rect 4985 -1885 5015 -1865
rect 5035 -1885 5065 -1865
rect 5085 -1885 5115 -1865
rect 5135 -1885 5165 -1865
rect 5185 -1885 5215 -1865
rect 5235 -1885 5265 -1865
rect 5285 -1885 5315 -1865
rect 5335 -1885 5365 -1865
rect 5385 -1885 5415 -1865
rect 5435 -1885 5465 -1865
rect 5485 -1885 5515 -1865
rect 5535 -1885 5565 -1865
rect 5585 -1885 5615 -1865
rect 5635 -1885 5665 -1865
rect 5685 -1885 5715 -1865
rect 5735 -1885 5765 -1865
rect 5785 -1885 5815 -1865
rect 5835 -1885 5865 -1865
rect 5885 -1885 5915 -1865
rect 5935 -1885 5965 -1865
rect 5985 -1885 6015 -1865
rect 6035 -1885 6065 -1865
rect 6085 -1885 6115 -1865
rect 6135 -1885 6165 -1865
rect 6185 -1885 6215 -1865
rect 6235 -1885 6265 -1865
rect 6285 -1885 6315 -1865
rect 6335 -1885 6365 -1865
rect 6385 -1885 6415 -1865
rect 6435 -1885 6465 -1865
rect 6485 -1885 6515 -1865
rect 6535 -1885 6565 -1865
rect 6585 -1885 6615 -1865
rect 6635 -1885 6665 -1865
rect 6685 -1885 6715 -1865
rect 6735 -1885 6765 -1865
rect 6785 -1885 6815 -1865
rect 6835 -1885 6865 -1865
rect 6885 -1885 6915 -1865
rect 6935 -1885 6965 -1865
rect 6985 -1885 7015 -1865
rect 7035 -1885 7065 -1865
rect 7085 -1885 7115 -1865
rect 7135 -1885 7165 -1865
rect 7185 -1885 7215 -1865
rect 7235 -1885 7265 -1865
rect 7285 -1885 7315 -1865
rect 7335 -1885 7365 -1865
rect 7385 -1885 7415 -1865
rect 7435 -1885 7465 -1865
rect 7485 -1885 7515 -1865
rect 7535 -1885 7565 -1865
rect 7585 -1885 7615 -1865
rect 7635 -1885 7665 -1865
rect 7685 -1885 7715 -1865
rect 7735 -1885 7765 -1865
rect 7785 -1885 7815 -1865
rect 7835 -1885 7865 -1865
rect 7885 -1885 7915 -1865
rect 7935 -1885 7965 -1865
rect 7985 -1885 8015 -1865
rect 8035 -1885 8065 -1865
rect 8085 -1885 8115 -1865
rect 8135 -1885 8165 -1865
rect 8185 -1885 8215 -1865
rect 8235 -1885 8265 -1865
rect 8285 -1885 8315 -1865
rect 8335 -1885 8365 -1865
rect 8385 -1885 8415 -1865
rect 8435 -1885 8465 -1865
rect 8485 -1885 8515 -1865
rect 8535 -1885 8565 -1865
rect 8585 -1885 8615 -1865
rect 8635 -1885 8665 -1865
rect 8685 -1885 8715 -1865
rect 8735 -1885 8765 -1865
rect 8785 -1885 8815 -1865
rect 8835 -1885 8865 -1865
rect 8885 -1885 8915 -1865
rect 8935 -1885 8965 -1865
rect 8985 -1885 9015 -1865
rect 9035 -1885 9065 -1865
rect 9085 -1885 9115 -1865
rect 9135 -1885 9165 -1865
rect 9185 -1885 9215 -1865
rect 9235 -1885 9265 -1865
rect 9285 -1885 9315 -1865
rect 9335 -1885 9365 -1865
rect 9385 -1885 9415 -1865
rect 9435 -1885 9465 -1865
rect 9485 -1885 9515 -1865
rect 9535 -1885 9565 -1865
rect 9585 -1885 9615 -1865
rect 9635 -1885 9665 -1865
rect 9685 -1885 9715 -1865
rect 9735 -1885 9765 -1865
rect 9785 -1885 9815 -1865
rect 9835 -1885 9865 -1865
rect 9885 -1885 9915 -1865
rect 9935 -1885 9965 -1865
rect 9985 -1885 10015 -1865
rect 10035 -1885 10065 -1865
rect 10085 -1885 10115 -1865
rect 10135 -1885 10165 -1865
rect 10185 -1885 10215 -1865
rect 10235 -1885 10265 -1865
rect 10285 -1885 10315 -1865
rect 10335 -1885 10365 -1865
rect 10385 -1885 10415 -1865
rect 10435 -1885 10465 -1865
rect 10485 -1885 10515 -1865
rect 10535 -1885 10565 -1865
rect 10585 -1885 10615 -1865
rect 10635 -1885 10665 -1865
rect 10685 -1885 10715 -1865
rect 10735 -1885 10765 -1865
rect 10785 -1885 10815 -1865
rect 10835 -1885 10865 -1865
rect 10885 -1885 10915 -1865
rect 10935 -1885 10965 -1865
rect 10985 -1885 11015 -1865
rect 11035 -1885 11065 -1865
rect 11085 -1885 11115 -1865
rect 11135 -1885 11165 -1865
rect 11185 -1885 11215 -1865
rect 11235 -1885 11265 -1865
rect 11285 -1885 11315 -1865
rect 11335 -1885 11365 -1865
rect 11385 -1885 11415 -1865
rect 11435 -1885 11465 -1865
rect 11485 -1885 11515 -1865
rect 11535 -1885 11565 -1865
rect 11585 -1885 11615 -1865
rect 11635 -1885 11665 -1865
rect 11685 -1885 11715 -1865
rect 11735 -1885 11765 -1865
rect 11785 -1885 11815 -1865
rect 11835 -1885 11865 -1865
rect 11885 -1885 11915 -1865
rect 11935 -1885 11965 -1865
rect 11985 -1885 12015 -1865
rect 12035 -1885 12065 -1865
rect 12085 -1885 12115 -1865
rect 12135 -1885 12165 -1865
rect 12185 -1885 12215 -1865
rect 12235 -1885 12265 -1865
rect 12285 -1885 12315 -1865
rect 12335 -1885 12365 -1865
rect 12385 -1885 12415 -1865
rect 12435 -1885 12465 -1865
rect 12485 -1885 12515 -1865
rect 12535 -1885 12565 -1865
rect 12585 -1885 12615 -1865
rect 12635 -1885 12665 -1865
rect 12685 -1885 12715 -1865
rect 12735 -1885 12765 -1865
rect 12785 -1885 12815 -1865
rect 12835 -1885 12865 -1865
rect 12885 -1885 12915 -1865
rect 12935 -1885 12965 -1865
rect 12985 -1885 13015 -1865
rect 13035 -1885 13065 -1865
rect 13085 -1885 13115 -1865
rect 13135 -1885 13165 -1865
rect 13185 -1885 13215 -1865
rect 13235 -1885 13265 -1865
rect 13285 -1885 13315 -1865
rect 13335 -1885 13365 -1865
rect 13385 -1885 13415 -1865
rect 13435 -1885 13465 -1865
rect 13485 -1885 13515 -1865
rect 13535 -1885 13565 -1865
rect 13585 -1885 13615 -1865
rect 13635 -1885 13665 -1865
rect 13685 -1885 13715 -1865
rect 13735 -1885 13765 -1865
rect 13785 -1885 13815 -1865
rect 13835 -1885 13865 -1865
rect 13885 -1885 13915 -1865
rect 13935 -1885 13965 -1865
rect 13985 -1885 14015 -1865
rect 14035 -1885 14065 -1865
rect 14085 -1885 14115 -1865
rect 14135 -1885 14165 -1865
rect 14185 -1885 14215 -1865
rect 14235 -1885 14265 -1865
rect 14285 -1885 14315 -1865
rect 14335 -1885 14365 -1865
rect 14385 -1885 14415 -1865
rect 14435 -1885 14465 -1865
rect 14485 -1885 14515 -1865
rect 14535 -1885 14565 -1865
rect 14585 -1885 14615 -1865
rect 14635 -1885 14665 -1865
rect 14685 -1885 14715 -1865
rect 14735 -1885 14765 -1865
rect 14785 -1885 14815 -1865
rect 14835 -1885 14865 -1865
rect 14885 -1885 14915 -1865
rect 14935 -1885 14965 -1865
rect 14985 -1885 15015 -1865
rect 15035 -1885 15065 -1865
rect 15085 -1885 15115 -1865
rect 15135 -1885 15165 -1865
rect 15185 -1885 15215 -1865
rect 15235 -1885 15265 -1865
rect 15285 -1885 15315 -1865
rect 15335 -1885 15365 -1865
rect 15385 -1885 15415 -1865
rect 15435 -1885 15465 -1865
rect 15485 -1885 15515 -1865
rect 15535 -1885 15565 -1865
rect 15585 -1885 15615 -1865
rect 15635 -1885 15665 -1865
rect 15685 -1885 15715 -1865
rect 15735 -1885 15765 -1865
rect 15785 -1885 15815 -1865
rect 15835 -1885 15865 -1865
rect 15885 -1885 15915 -1865
rect 15935 -1885 15965 -1865
rect 15985 -1885 16015 -1865
rect 16035 -1885 16065 -1865
rect 16085 -1885 16115 -1865
rect 16135 -1885 16165 -1865
rect 16185 -1885 16215 -1865
rect 16235 -1885 16265 -1865
rect 16285 -1885 16315 -1865
rect 16335 -1885 16365 -1865
rect 16385 -1885 16415 -1865
rect 16435 -1885 16465 -1865
rect 16485 -1885 16515 -1865
rect 16535 -1885 16565 -1865
rect 16585 -1885 16615 -1865
rect 16635 -1885 16665 -1865
rect 16685 -1885 16715 -1865
rect 16735 -1885 16765 -1865
rect 16785 -1885 16815 -1865
rect 16835 -1885 16865 -1865
rect 16885 -1885 16915 -1865
rect 16935 -1885 16965 -1865
rect 16985 -1885 17015 -1865
rect 17035 -1885 17065 -1865
rect 17085 -1885 17115 -1865
rect 17135 -1885 17165 -1865
rect 17185 -1885 17215 -1865
rect 17235 -1885 17265 -1865
rect 17285 -1885 17315 -1865
rect 17335 -1885 17365 -1865
rect 17385 -1885 17415 -1865
rect 17435 -1885 17465 -1865
rect 17485 -1885 17515 -1865
rect 17535 -1885 17565 -1865
rect 17585 -1885 17615 -1865
rect 17635 -1885 17665 -1865
rect 17685 -1885 17715 -1865
rect 17735 -1885 17765 -1865
rect 17785 -1885 17815 -1865
rect 17835 -1885 17865 -1865
rect 17885 -1885 17915 -1865
rect 17935 -1885 17965 -1865
rect 17985 -1885 18015 -1865
rect 18035 -1885 18065 -1865
rect 18085 -1885 18115 -1865
rect 18135 -1885 18165 -1865
rect 18185 -1885 18215 -1865
rect 18235 -1885 18265 -1865
rect 18285 -1885 18315 -1865
rect 18335 -1885 18365 -1865
rect 18385 -1885 18415 -1865
rect 18435 -1885 18465 -1865
rect 18485 -1885 18515 -1865
rect 18535 -1885 18565 -1865
rect 18585 -1885 18615 -1865
rect 18635 -1885 18665 -1865
rect 18685 -1885 18715 -1865
rect 18735 -1885 18765 -1865
rect 18785 -1885 18815 -1865
rect 18835 -1885 18865 -1865
rect 18885 -1885 18915 -1865
rect 18935 -1885 18965 -1865
rect 18985 -1885 19015 -1865
rect 19035 -1885 19065 -1865
rect 19085 -1885 19115 -1865
rect 19135 -1885 19165 -1865
rect 19185 -1885 19215 -1865
rect 19235 -1885 19265 -1865
rect 19285 -1885 19315 -1865
rect 19335 -1885 19365 -1865
rect 19385 -1885 19415 -1865
rect 19435 -1885 19465 -1865
rect 19485 -1885 19515 -1865
rect 19535 -1885 19565 -1865
rect 19585 -1885 19615 -1865
rect 19635 -1885 19665 -1865
rect 19685 -1885 19715 -1865
rect 19735 -1885 19765 -1865
rect 19785 -1885 19815 -1865
rect 19835 -1885 19865 -1865
rect 19885 -1885 19915 -1865
rect 19935 -1885 19965 -1865
rect 19985 -1885 20015 -1865
rect 20035 -1885 20065 -1865
rect 20085 -1885 20115 -1865
rect 20135 -1885 20165 -1865
rect 20185 -1885 20215 -1865
rect 20235 -1885 20265 -1865
rect 20285 -1885 20315 -1865
rect 20335 -1885 20365 -1865
rect 20385 -1885 20415 -1865
rect 20435 -1885 20465 -1865
rect 20485 -1885 20515 -1865
rect 20535 -1885 20565 -1865
rect 20585 -1885 20615 -1865
rect 20635 -1885 20665 -1865
rect 20685 -1885 20715 -1865
rect 20735 -1885 20765 -1865
rect 20785 -1885 20815 -1865
rect 20835 -1885 20865 -1865
rect 20885 -1885 20915 -1865
rect 20935 -1885 20965 -1865
rect 20985 -1885 21015 -1865
rect 21035 -1885 21065 -1865
rect 21085 -1885 21115 -1865
rect 21135 -1885 21165 -1865
rect 21185 -1885 21215 -1865
rect 21235 -1885 21265 -1865
rect 21285 -1885 21315 -1865
rect 21335 -1885 21365 -1865
rect 21385 -1885 21415 -1865
rect 21435 -1885 21465 -1865
rect 21485 -1885 21515 -1865
rect 21535 -1885 21565 -1865
rect 21585 -1885 21615 -1865
rect 21635 -1885 21665 -1865
rect 21685 -1885 21715 -1865
rect 21735 -1885 21765 -1865
rect 21785 -1885 21815 -1865
rect 21835 -1885 21865 -1865
rect 21885 -1885 21915 -1865
rect 21935 -1885 21965 -1865
rect 21985 -1885 22015 -1865
rect 22035 -1885 22065 -1865
rect 22085 -1885 22115 -1865
rect 22135 -1885 22165 -1865
rect 22185 -1885 22215 -1865
rect 22235 -1885 22265 -1865
rect 22285 -1885 22315 -1865
rect 22335 -1885 22365 -1865
rect 22385 -1885 22415 -1865
rect 22435 -1885 22465 -1865
rect 22485 -1885 22515 -1865
rect 22535 -1885 22565 -1865
rect 22585 -1885 22615 -1865
rect 22635 -1885 22665 -1865
rect 22685 -1885 22715 -1865
rect 22735 -1885 22765 -1865
rect 22785 -1885 22815 -1865
rect 22835 -1885 22865 -1865
rect 22885 -1885 22915 -1865
rect 22935 -1885 22965 -1865
rect 22985 -1885 23015 -1865
rect 23035 -1885 23065 -1865
rect 23085 -1885 23115 -1865
rect 23135 -1885 23165 -1865
rect 23185 -1885 23215 -1865
rect 23235 -1885 23265 -1865
rect 23285 -1885 23315 -1865
rect 23335 -1885 23365 -1865
rect 23385 -1885 23415 -1865
rect 23435 -1885 23465 -1865
rect 23485 -1885 23515 -1865
rect 23535 -1885 23565 -1865
rect 23585 -1885 23615 -1865
rect 23635 -1885 23665 -1865
rect 23685 -1885 23715 -1865
rect 23735 -1885 23765 -1865
rect 23785 -1885 23815 -1865
rect 23835 -1885 23865 -1865
rect 23885 -1885 23915 -1865
rect 23935 -1885 23965 -1865
rect 23985 -1885 24015 -1865
rect 24035 -1885 24065 -1865
rect 24085 -1885 24115 -1865
rect 24135 -1885 24165 -1865
rect 24185 -1885 24215 -1865
rect 24235 -1885 24265 -1865
rect 24285 -1885 24315 -1865
rect 24335 -1885 24365 -1865
rect 24385 -1885 24415 -1865
rect 24435 -1885 24465 -1865
rect 24485 -1885 24515 -1865
rect 24535 -1885 24565 -1865
rect 24585 -1885 24615 -1865
rect 24635 -1885 24665 -1865
rect 24685 -1885 24715 -1865
rect 24735 -1885 24765 -1865
rect 24785 -1885 24815 -1865
rect 24835 -1885 24865 -1865
rect 24885 -1885 24915 -1865
rect 24935 -1885 24965 -1865
rect 24985 -1885 25015 -1865
rect 25035 -1885 25065 -1865
rect 25085 -1885 25115 -1865
rect 25135 -1885 25165 -1865
rect 25185 -1885 25215 -1865
rect 25235 -1885 25265 -1865
rect 25285 -1885 25315 -1865
rect 25335 -1885 25365 -1865
rect 25385 -1885 25415 -1865
rect 25435 -1885 25465 -1865
rect 25485 -1885 25515 -1865
rect 25535 -1885 25565 -1865
rect 25585 -1885 25615 -1865
rect 25635 -1885 25665 -1865
rect 25685 -1885 25715 -1865
rect 25735 -1885 25765 -1865
rect 25785 -1885 25815 -1865
rect 25835 -1885 25865 -1865
rect 25885 -1885 25915 -1865
rect 25935 -1885 25965 -1865
rect 25985 -1885 26015 -1865
rect 26035 -1885 26065 -1865
rect 26085 -1885 26115 -1865
rect 26135 -1885 26165 -1865
rect 26185 -1885 26215 -1865
rect 26235 -1885 26265 -1865
rect 26285 -1885 26315 -1865
rect 26335 -1885 26365 -1865
rect 26385 -1885 26415 -1865
rect 26435 -1885 26465 -1865
rect 26485 -1885 26515 -1865
rect 26535 -1885 26565 -1865
rect 26585 -1885 26615 -1865
rect 26635 -1885 26665 -1865
rect 26685 -1885 26715 -1865
rect 26735 -1885 26765 -1865
rect 26785 -1885 26815 -1865
rect 26835 -1885 26865 -1865
rect 26885 -1885 26915 -1865
rect 26935 -1885 26965 -1865
rect 26985 -1885 27015 -1865
rect 27035 -1885 27065 -1865
rect 27085 -1885 27115 -1865
rect 27135 -1885 27165 -1865
rect 27185 -1885 27215 -1865
rect 27235 -1885 27265 -1865
rect 27285 -1885 27315 -1865
rect 27335 -1885 27365 -1865
rect 27385 -1885 27415 -1865
rect 27435 -1885 27465 -1865
rect 27485 -1885 27515 -1865
rect 27535 -1885 27565 -1865
rect 27585 -1885 27615 -1865
rect 27635 -1885 27665 -1865
rect 27685 -1885 27715 -1865
rect 27735 -1885 27765 -1865
rect 27785 -1885 27815 -1865
rect 27835 -1885 27865 -1865
rect 27885 -1885 27915 -1865
rect 27935 -1885 27965 -1865
rect 27985 -1885 28015 -1865
rect 28035 -1885 28065 -1865
rect 28085 -1885 28115 -1865
rect 28135 -1885 28165 -1865
rect 28185 -1885 28215 -1865
rect 28235 -1885 28265 -1865
rect 28285 -1885 28315 -1865
rect 28335 -1885 28365 -1865
rect 28385 -1885 28415 -1865
rect 28435 -1885 28465 -1865
rect 28485 -1885 28515 -1865
rect 28535 -1885 28565 -1865
rect 28585 -1885 28615 -1865
rect 28635 -1885 28665 -1865
rect 28685 -1885 28715 -1865
rect 28735 -1885 28765 -1865
rect 28785 -1885 28800 -1865
rect -650 -1900 28800 -1885
<< mvpsubdiffcont >>
rect -885 2815 -865 2835
rect -835 2815 -815 2835
rect -785 2815 -765 2835
rect -735 2815 -715 2835
rect -685 2815 -665 2835
rect -635 2815 -615 2835
rect -585 2815 -565 2835
rect -535 2815 -515 2835
rect -485 2815 -465 2835
rect -435 2815 -415 2835
rect -385 2815 -365 2835
rect -335 2815 -315 2835
rect -285 2815 -265 2835
rect -235 2815 -215 2835
rect -185 2815 -165 2835
rect -135 2815 -115 2835
rect -85 2815 -65 2835
rect -35 2815 -15 2835
rect 15 2815 35 2835
rect 65 2815 85 2835
rect 115 2815 135 2835
rect 165 2815 185 2835
rect 215 2815 235 2835
rect 265 2815 285 2835
rect 315 2815 335 2835
rect 365 2815 385 2835
rect 415 2815 435 2835
rect 465 2815 485 2835
rect 515 2815 535 2835
rect 565 2815 585 2835
rect 615 2815 635 2835
rect 665 2815 685 2835
rect 715 2815 735 2835
rect 765 2815 785 2835
rect 815 2815 835 2835
rect 865 2815 885 2835
rect 915 2815 935 2835
rect 965 2815 985 2835
rect 1015 2815 1035 2835
rect 1065 2815 1085 2835
rect 1115 2815 1135 2835
rect 1165 2815 1185 2835
rect 1215 2815 1235 2835
rect 1265 2815 1285 2835
rect 1315 2815 1335 2835
rect 1365 2815 1385 2835
rect 1415 2815 1435 2835
rect 1465 2815 1485 2835
rect 1515 2815 1535 2835
rect 1565 2815 1585 2835
rect 1615 2815 1635 2835
rect 1665 2815 1685 2835
rect 1715 2815 1735 2835
rect 1765 2815 1785 2835
rect 1815 2815 1835 2835
rect 1865 2815 1885 2835
rect 1915 2815 1935 2835
rect 1965 2815 1985 2835
rect 2015 2815 2035 2835
rect 2065 2815 2085 2835
rect 2115 2815 2135 2835
rect 2165 2815 2185 2835
rect 2215 2815 2235 2835
rect 2265 2815 2285 2835
rect 2315 2815 2335 2835
rect 2365 2815 2385 2835
rect 2415 2815 2435 2835
rect 2465 2815 2485 2835
rect 2515 2815 2535 2835
rect 2565 2815 2585 2835
rect 2615 2815 2635 2835
rect 2665 2815 2685 2835
rect 2715 2815 2735 2835
rect 2765 2815 2785 2835
rect 2815 2815 2835 2835
rect 2865 2815 2885 2835
rect 2915 2815 2935 2835
rect 2965 2815 2985 2835
rect 3015 2815 3035 2835
rect 3065 2815 3085 2835
rect 3115 2815 3135 2835
rect 3165 2815 3185 2835
rect 3215 2815 3235 2835
rect 3265 2815 3285 2835
rect 3315 2815 3335 2835
rect 3365 2815 3385 2835
rect 3415 2815 3435 2835
rect 3465 2815 3485 2835
rect 3515 2815 3535 2835
rect 3565 2815 3585 2835
rect 3615 2815 3635 2835
rect 3665 2815 3685 2835
rect 3715 2815 3735 2835
rect 3765 2815 3785 2835
rect 3815 2815 3835 2835
rect 3865 2815 3885 2835
rect 3915 2815 3935 2835
rect 3965 2815 3985 2835
rect 4015 2815 4035 2835
rect 4065 2815 4085 2835
rect 4115 2815 4135 2835
rect 4165 2815 4185 2835
rect 4215 2815 4235 2835
rect 4265 2815 4285 2835
rect 4315 2815 4335 2835
rect 4365 2815 4385 2835
rect 4415 2815 4435 2835
rect 4465 2815 4485 2835
rect 4515 2815 4535 2835
rect 4565 2815 4585 2835
rect 4615 2815 4635 2835
rect 4665 2815 4685 2835
rect 4715 2815 4735 2835
rect 4765 2815 4785 2835
rect 4815 2815 4835 2835
rect 4865 2815 4885 2835
rect 4915 2815 4935 2835
rect 4965 2815 4985 2835
rect 5015 2815 5035 2835
rect 5065 2815 5085 2835
rect 5115 2815 5135 2835
rect 5165 2815 5185 2835
rect 5215 2815 5235 2835
rect 5265 2815 5285 2835
rect 5315 2815 5335 2835
rect 5365 2815 5385 2835
rect 5415 2815 5435 2835
rect 5465 2815 5485 2835
rect 5515 2815 5535 2835
rect 5565 2815 5585 2835
rect 5615 2815 5635 2835
rect 5665 2815 5685 2835
rect 5715 2815 5735 2835
rect 5765 2815 5785 2835
rect 5815 2815 5835 2835
rect 5865 2815 5885 2835
rect 5915 2815 5935 2835
rect 5965 2815 5985 2835
rect 6015 2815 6035 2835
rect 6065 2815 6085 2835
rect 6115 2815 6135 2835
rect 6165 2815 6185 2835
rect 6215 2815 6235 2835
rect 6265 2815 6285 2835
rect 6315 2815 6335 2835
rect 6365 2815 6385 2835
rect 6415 2815 6435 2835
rect 6465 2815 6485 2835
rect 6515 2815 6535 2835
rect 6565 2815 6585 2835
rect 6615 2815 6635 2835
rect 6665 2815 6685 2835
rect 6715 2815 6735 2835
rect 6765 2815 6785 2835
rect 6815 2815 6835 2835
rect 6865 2815 6885 2835
rect 6915 2815 6935 2835
rect 6965 2815 6985 2835
rect 7015 2815 7035 2835
rect 7065 2815 7085 2835
rect 7115 2815 7135 2835
rect 7165 2815 7185 2835
rect 7215 2815 7235 2835
rect 7265 2815 7285 2835
rect 7315 2815 7335 2835
rect 7365 2815 7385 2835
rect 7415 2815 7435 2835
rect 7465 2815 7485 2835
rect 7515 2815 7535 2835
rect 7565 2815 7585 2835
rect 7615 2815 7635 2835
rect 7665 2815 7685 2835
rect 7715 2815 7735 2835
rect 7765 2815 7785 2835
rect 7815 2815 7835 2835
rect 7865 2815 7885 2835
rect 7915 2815 7935 2835
rect 7965 2815 7985 2835
rect 8015 2815 8035 2835
rect 8065 2815 8085 2835
rect 8115 2815 8135 2835
rect 8165 2815 8185 2835
rect 8215 2815 8235 2835
rect 8265 2815 8285 2835
rect 8315 2815 8335 2835
rect 8365 2815 8385 2835
rect 8415 2815 8435 2835
rect 8465 2815 8485 2835
rect 8515 2815 8535 2835
rect 8565 2815 8585 2835
rect 8615 2815 8635 2835
rect 8665 2815 8685 2835
rect 8715 2815 8735 2835
rect 8765 2815 8785 2835
rect 8815 2815 8835 2835
rect 8865 2815 8885 2835
rect 8915 2815 8935 2835
rect 8965 2815 8985 2835
rect 9015 2815 9035 2835
rect 9065 2815 9085 2835
rect 9115 2815 9135 2835
rect 9165 2815 9185 2835
rect 9215 2815 9235 2835
rect 9265 2815 9285 2835
rect 9315 2815 9335 2835
rect 9365 2815 9385 2835
rect 9415 2815 9435 2835
rect 9465 2815 9485 2835
rect 9515 2815 9535 2835
rect 9565 2815 9585 2835
rect 9615 2815 9635 2835
rect 9665 2815 9685 2835
rect 9715 2815 9735 2835
rect 9765 2815 9785 2835
rect 9815 2815 9835 2835
rect 9865 2815 9885 2835
rect 9915 2815 9935 2835
rect 9965 2815 9985 2835
rect 10015 2815 10035 2835
rect 10065 2815 10085 2835
rect 10115 2815 10135 2835
rect 10165 2815 10185 2835
rect 10215 2815 10235 2835
rect 10265 2815 10285 2835
rect 10315 2815 10335 2835
rect 10365 2815 10385 2835
rect 10415 2815 10435 2835
rect 10465 2815 10485 2835
rect 10515 2815 10535 2835
rect 10565 2815 10585 2835
rect 10615 2815 10635 2835
rect 10665 2815 10685 2835
rect 10715 2815 10735 2835
rect 10765 2815 10785 2835
rect 10815 2815 10835 2835
rect 10865 2815 10885 2835
rect 10915 2815 10935 2835
rect 10965 2815 10985 2835
rect 11015 2815 11035 2835
rect 11065 2815 11085 2835
rect 11115 2815 11135 2835
rect 11165 2815 11185 2835
rect 11215 2815 11235 2835
rect 11265 2815 11285 2835
rect 11315 2815 11335 2835
rect 11365 2815 11385 2835
rect 11415 2815 11435 2835
rect 11465 2815 11485 2835
rect 11515 2815 11535 2835
rect 11565 2815 11585 2835
rect 11615 2815 11635 2835
rect 11665 2815 11685 2835
rect 11715 2815 11735 2835
rect 11765 2815 11785 2835
rect 11815 2815 11835 2835
rect 11865 2815 11885 2835
rect 11915 2815 11935 2835
rect 11965 2815 11985 2835
rect 12015 2815 12035 2835
rect 12065 2815 12085 2835
rect 12115 2815 12135 2835
rect 12165 2815 12185 2835
rect 12215 2815 12235 2835
rect 12265 2815 12285 2835
rect 12315 2815 12335 2835
rect 12365 2815 12385 2835
rect 12415 2815 12435 2835
rect 12465 2815 12485 2835
rect 12515 2815 12535 2835
rect 12565 2815 12585 2835
rect 12615 2815 12635 2835
rect 12665 2815 12685 2835
rect 12715 2815 12735 2835
rect 12765 2815 12785 2835
rect 12815 2815 12835 2835
rect 12865 2815 12885 2835
rect 12915 2815 12935 2835
rect 12965 2815 12985 2835
rect 13015 2815 13035 2835
rect 13065 2815 13085 2835
rect 13115 2815 13135 2835
rect 13165 2815 13185 2835
rect 13215 2815 13235 2835
rect 13265 2815 13285 2835
rect 13315 2815 13335 2835
rect 13365 2815 13385 2835
rect 13415 2815 13435 2835
rect 13465 2815 13485 2835
rect 13515 2815 13535 2835
rect 13565 2815 13585 2835
rect 13615 2815 13635 2835
rect 13665 2815 13685 2835
rect 13715 2815 13735 2835
rect 13765 2815 13785 2835
rect 13815 2815 13835 2835
rect 13865 2815 13885 2835
rect 13915 2815 13935 2835
rect 13965 2815 13985 2835
rect 14015 2815 14035 2835
rect 14065 2815 14085 2835
rect 14115 2815 14135 2835
rect 14165 2815 14185 2835
rect 14215 2815 14235 2835
rect 14265 2815 14285 2835
rect 14315 2815 14335 2835
rect 14365 2815 14385 2835
rect 14415 2815 14435 2835
rect 14465 2815 14485 2835
rect 14515 2815 14535 2835
rect 14565 2815 14585 2835
rect 14615 2815 14635 2835
rect 14665 2815 14685 2835
rect 14715 2815 14735 2835
rect 14765 2815 14785 2835
rect 14815 2815 14835 2835
rect 14865 2815 14885 2835
rect 14915 2815 14935 2835
rect 14965 2815 14985 2835
rect 15015 2815 15035 2835
rect 15065 2815 15085 2835
rect 15115 2815 15135 2835
rect 15165 2815 15185 2835
rect 15215 2815 15235 2835
rect 15265 2815 15285 2835
rect 15315 2815 15335 2835
rect 15365 2815 15385 2835
rect 15415 2815 15435 2835
rect 15465 2815 15485 2835
rect 15515 2815 15535 2835
rect 15565 2815 15585 2835
rect 15615 2815 15635 2835
rect 15665 2815 15685 2835
rect 15715 2815 15735 2835
rect 15765 2815 15785 2835
rect 15815 2815 15835 2835
rect 15865 2815 15885 2835
rect 15915 2815 15935 2835
rect 15965 2815 15985 2835
rect 16015 2815 16035 2835
rect 16065 2815 16085 2835
rect 16115 2815 16135 2835
rect 16165 2815 16185 2835
rect 16215 2815 16235 2835
rect 16265 2815 16285 2835
rect 16315 2815 16335 2835
rect 16365 2815 16385 2835
rect 16415 2815 16435 2835
rect 16465 2815 16485 2835
rect 16515 2815 16535 2835
rect 16565 2815 16585 2835
rect 16615 2815 16635 2835
rect 16665 2815 16685 2835
rect 16715 2815 16735 2835
rect 16765 2815 16785 2835
rect 16815 2815 16835 2835
rect 16865 2815 16885 2835
rect 16915 2815 16935 2835
rect 16965 2815 16985 2835
rect 17015 2815 17035 2835
rect 17065 2815 17085 2835
rect 17115 2815 17135 2835
rect 17165 2815 17185 2835
rect 17215 2815 17235 2835
rect 17265 2815 17285 2835
rect 17315 2815 17335 2835
rect 17365 2815 17385 2835
rect 17415 2815 17435 2835
rect 17465 2815 17485 2835
rect 17515 2815 17535 2835
rect 17565 2815 17585 2835
rect 17615 2815 17635 2835
rect 17665 2815 17685 2835
rect 17715 2815 17735 2835
rect 17765 2815 17785 2835
rect 17815 2815 17835 2835
rect 17865 2815 17885 2835
rect 17915 2815 17935 2835
rect 17965 2815 17985 2835
rect 18015 2815 18035 2835
rect 18065 2815 18085 2835
rect 18115 2815 18135 2835
rect 18165 2815 18185 2835
rect 18215 2815 18235 2835
rect 18265 2815 18285 2835
rect 18315 2815 18335 2835
rect 18365 2815 18385 2835
rect 18415 2815 18435 2835
rect 18465 2815 18485 2835
rect 18515 2815 18535 2835
rect 18565 2815 18585 2835
rect 18615 2815 18635 2835
rect 18665 2815 18685 2835
rect 18715 2815 18735 2835
rect 18765 2815 18785 2835
rect 18815 2815 18835 2835
rect 18865 2815 18885 2835
rect 18915 2815 18935 2835
rect 18965 2815 18985 2835
rect 19015 2815 19035 2835
rect 19065 2815 19085 2835
rect 19115 2815 19135 2835
rect 19165 2815 19185 2835
rect 19215 2815 19235 2835
rect 19265 2815 19285 2835
rect 19315 2815 19335 2835
rect 19365 2815 19385 2835
rect 19415 2815 19435 2835
rect 19465 2815 19485 2835
rect 19515 2815 19535 2835
rect 19565 2815 19585 2835
rect 19615 2815 19635 2835
rect 19665 2815 19685 2835
rect 19715 2815 19735 2835
rect 19765 2815 19785 2835
rect 19815 2815 19835 2835
rect 19865 2815 19885 2835
rect 19915 2815 19935 2835
rect 19965 2815 19985 2835
rect 20015 2815 20035 2835
rect 20065 2815 20085 2835
rect 20115 2815 20135 2835
rect 20165 2815 20185 2835
rect 20215 2815 20235 2835
rect 20265 2815 20285 2835
rect 20315 2815 20335 2835
rect 20365 2815 20385 2835
rect 20415 2815 20435 2835
rect 20465 2815 20485 2835
rect 20515 2815 20535 2835
rect 20565 2815 20585 2835
rect 20615 2815 20635 2835
rect 20665 2815 20685 2835
rect 20715 2815 20735 2835
rect 20765 2815 20785 2835
rect 20815 2815 20835 2835
rect 20865 2815 20885 2835
rect 20915 2815 20935 2835
rect 20965 2815 20985 2835
rect 21015 2815 21035 2835
rect 21065 2815 21085 2835
rect 21115 2815 21135 2835
rect 21165 2815 21185 2835
rect 21215 2815 21235 2835
rect 21265 2815 21285 2835
rect 21315 2815 21335 2835
rect 21365 2815 21385 2835
rect 21415 2815 21435 2835
rect 21465 2815 21485 2835
rect 21515 2815 21535 2835
rect 21565 2815 21585 2835
rect 21615 2815 21635 2835
rect 21665 2815 21685 2835
rect 21715 2815 21735 2835
rect 21765 2815 21785 2835
rect 21815 2815 21835 2835
rect 21865 2815 21885 2835
rect 21915 2815 21935 2835
rect 21965 2815 21985 2835
rect 22015 2815 22035 2835
rect 22065 2815 22085 2835
rect 22115 2815 22135 2835
rect 22165 2815 22185 2835
rect 22215 2815 22235 2835
rect 22265 2815 22285 2835
rect 22315 2815 22335 2835
rect 22365 2815 22385 2835
rect 22415 2815 22435 2835
rect 22465 2815 22485 2835
rect 22515 2815 22535 2835
rect 22565 2815 22585 2835
rect 22615 2815 22635 2835
rect 22665 2815 22685 2835
rect 22715 2815 22735 2835
rect 22765 2815 22785 2835
rect 22815 2815 22835 2835
rect 22865 2815 22885 2835
rect 22915 2815 22935 2835
rect 22965 2815 22985 2835
rect 23015 2815 23035 2835
rect 23065 2815 23085 2835
rect 23115 2815 23135 2835
rect 23165 2815 23185 2835
rect 23215 2815 23235 2835
rect 23265 2815 23285 2835
rect 23315 2815 23335 2835
rect 23365 2815 23385 2835
rect 23415 2815 23435 2835
rect 23465 2815 23485 2835
rect 23515 2815 23535 2835
rect 23565 2815 23585 2835
rect 23615 2815 23635 2835
rect 23665 2815 23685 2835
rect 23715 2815 23735 2835
rect 23765 2815 23785 2835
rect 23815 2815 23835 2835
rect 23865 2815 23885 2835
rect 23915 2815 23935 2835
rect 23965 2815 23985 2835
rect 24015 2815 24035 2835
rect 24065 2815 24085 2835
rect 24115 2815 24135 2835
rect 24165 2815 24185 2835
rect 24215 2815 24235 2835
rect 24265 2815 24285 2835
rect 24315 2815 24335 2835
rect 24365 2815 24385 2835
rect 24415 2815 24435 2835
rect 24465 2815 24485 2835
rect 24515 2815 24535 2835
rect 24565 2815 24585 2835
rect 24615 2815 24635 2835
rect 24665 2815 24685 2835
rect 24715 2815 24735 2835
rect 24765 2815 24785 2835
rect 24815 2815 24835 2835
rect 24865 2815 24885 2835
rect 24915 2815 24935 2835
rect 24965 2815 24985 2835
rect 25015 2815 25035 2835
rect 25065 2815 25085 2835
rect 25115 2815 25135 2835
rect 25165 2815 25185 2835
rect 25215 2815 25235 2835
rect 25265 2815 25285 2835
rect 25315 2815 25335 2835
rect 25365 2815 25385 2835
rect 25415 2815 25435 2835
rect 25465 2815 25485 2835
rect 25515 2815 25535 2835
rect 25565 2815 25585 2835
rect 25615 2815 25635 2835
rect 25665 2815 25685 2835
rect 25715 2815 25735 2835
rect 25765 2815 25785 2835
rect 25815 2815 25835 2835
rect 25865 2815 25885 2835
rect 25915 2815 25935 2835
rect 25965 2815 25985 2835
rect 26015 2815 26035 2835
rect 26065 2815 26085 2835
rect 26115 2815 26135 2835
rect 26165 2815 26185 2835
rect 26215 2815 26235 2835
rect 26265 2815 26285 2835
rect 26315 2815 26335 2835
rect 26365 2815 26385 2835
rect 26415 2815 26435 2835
rect 26465 2815 26485 2835
rect 26515 2815 26535 2835
rect 26565 2815 26585 2835
rect 26615 2815 26635 2835
rect 26665 2815 26685 2835
rect 26715 2815 26735 2835
rect 26765 2815 26785 2835
rect 26815 2815 26835 2835
rect 26865 2815 26885 2835
rect 26915 2815 26935 2835
rect 26965 2815 26985 2835
rect 27015 2815 27035 2835
rect 27065 2815 27085 2835
rect 27115 2815 27135 2835
rect 27165 2815 27185 2835
rect 27215 2815 27235 2835
rect 27265 2815 27285 2835
rect 27315 2815 27335 2835
rect 27365 2815 27385 2835
rect 27415 2815 27435 2835
rect 27465 2815 27485 2835
rect 27515 2815 27535 2835
rect 27565 2815 27585 2835
rect 27615 2815 27635 2835
rect 27665 2815 27685 2835
rect 27715 2815 27735 2835
rect 27765 2815 27785 2835
rect 27815 2815 27835 2835
rect 27865 2815 27885 2835
rect 27915 2815 27935 2835
rect 27965 2815 27985 2835
rect 28015 2815 28035 2835
rect 28065 2815 28085 2835
rect 28115 2815 28135 2835
rect 28165 2815 28185 2835
rect 28215 2815 28235 2835
rect 28265 2815 28285 2835
rect 28315 2815 28335 2835
rect 28365 2815 28385 2835
rect 28415 2815 28435 2835
rect 28465 2815 28485 2835
rect 28515 2815 28535 2835
rect 28565 2815 28585 2835
rect 28615 2815 28635 2835
rect 28665 2815 28685 2835
rect 28715 2815 28735 2835
rect 28765 2815 28785 2835
rect 28815 2815 28835 2835
rect 28865 2815 28885 2835
rect 28915 2815 28935 2835
rect 28965 2815 28985 2835
rect 29015 2815 29035 2835
rect 29065 2815 29085 2835
rect 29115 2815 29135 2835
rect 29165 2815 29185 2835
rect 29215 2815 29235 2835
rect 29265 2815 29285 2835
rect 29315 2815 29335 2835
rect 29365 2815 29385 2835
rect 29415 2815 29435 2835
rect 29465 2815 29485 2835
rect 29515 2815 29535 2835
rect 29565 2815 29585 2835
rect 29615 2815 29635 2835
rect 29665 2815 29685 2835
rect 29715 2815 29735 2835
rect 29765 2815 29785 2835
rect 29815 2815 29835 2835
rect 29865 2815 29885 2835
rect 29915 2815 29935 2835
rect 29965 2815 29985 2835
rect 30015 2815 30035 2835
rect 30065 2815 30085 2835
rect 30115 2815 30135 2835
rect 30165 2815 30185 2835
rect 30215 2815 30235 2835
rect 30265 2815 30285 2835
rect 30315 2815 30335 2835
rect 30365 2815 30385 2835
rect 30415 2815 30435 2835
rect 30465 2815 30485 2835
rect 30515 2815 30535 2835
rect 30565 2815 30585 2835
rect 30615 2815 30635 2835
rect 30665 2815 30685 2835
rect 30715 2815 30735 2835
rect 30765 2815 30785 2835
rect 30815 2815 30835 2835
rect 30865 2815 30885 2835
rect 30915 2815 30935 2835
rect 30965 2815 30985 2835
rect 31015 2815 31035 2835
rect 31065 2815 31085 2835
rect 31115 2815 31135 2835
rect 31165 2815 31185 2835
rect 31215 2815 31235 2835
rect 31265 2815 31285 2835
rect 31315 2815 31335 2835
rect 31365 2815 31385 2835
rect 31415 2815 31435 2835
rect 31465 2815 31485 2835
rect 31515 2815 31535 2835
rect 31565 2815 31585 2835
rect 31615 2815 31635 2835
rect 31665 2815 31685 2835
rect 31715 2815 31735 2835
rect 31765 2815 31785 2835
rect 31815 2815 31835 2835
rect 31865 2815 31885 2835
rect 31915 2815 31935 2835
rect 31965 2815 31985 2835
rect 32015 2815 32035 2835
rect 32065 2815 32085 2835
rect -885 2015 -865 2035
rect -835 2015 -815 2035
rect -785 2015 -765 2035
rect -735 2015 -715 2035
rect -685 2015 -665 2035
rect -635 2015 -615 2035
rect -585 2015 -565 2035
rect -535 2015 -515 2035
rect -485 2015 -465 2035
rect -435 2015 -415 2035
rect -385 2015 -365 2035
rect -335 2015 -315 2035
rect -285 2015 -265 2035
rect -235 2015 -215 2035
rect -185 2015 -165 2035
rect -135 2015 -115 2035
rect -85 2015 -65 2035
rect -35 2015 -15 2035
rect 15 2015 35 2035
rect 65 2015 85 2035
rect 115 2015 135 2035
rect 165 2015 185 2035
rect 215 2015 235 2035
rect 265 2015 285 2035
rect 315 2015 335 2035
rect 365 2015 385 2035
rect 415 2015 435 2035
rect 465 2015 485 2035
rect 515 2015 535 2035
rect 565 2015 585 2035
rect 615 2015 635 2035
rect 665 2015 685 2035
rect 715 2015 735 2035
rect 765 2015 785 2035
rect 815 2015 835 2035
rect 865 2015 885 2035
rect 915 2015 935 2035
rect 965 2015 985 2035
rect 1015 2015 1035 2035
rect 1065 2015 1085 2035
rect 1115 2015 1135 2035
rect 1165 2015 1185 2035
rect 1215 2015 1235 2035
rect 1265 2015 1285 2035
rect 1315 2015 1335 2035
rect 1365 2015 1385 2035
rect 1415 2015 1435 2035
rect 1465 2015 1485 2035
rect 1515 2015 1535 2035
rect 1565 2015 1585 2035
rect 1615 2015 1635 2035
rect 1665 2015 1685 2035
rect 1715 2015 1735 2035
rect 1765 2015 1785 2035
rect 1815 2015 1835 2035
rect 1865 2015 1885 2035
rect 1915 2015 1935 2035
rect 1965 2015 1985 2035
rect 2015 2015 2035 2035
rect 2065 2015 2085 2035
rect 2115 2015 2135 2035
rect 2165 2015 2185 2035
rect 2215 2015 2235 2035
rect 2265 2015 2285 2035
rect 2315 2015 2335 2035
rect 2365 2015 2385 2035
rect 2415 2015 2435 2035
rect 2465 2015 2485 2035
rect 2515 2015 2535 2035
rect 2565 2015 2585 2035
rect 2615 2015 2635 2035
rect 2665 2015 2685 2035
rect 2715 2015 2735 2035
rect 2765 2015 2785 2035
rect 2815 2015 2835 2035
rect 2865 2015 2885 2035
rect 2915 2015 2935 2035
rect 2965 2015 2985 2035
rect 3015 2015 3035 2035
rect 3065 2015 3085 2035
rect 3115 2015 3135 2035
rect 3165 2015 3185 2035
rect 3215 2015 3235 2035
rect 3265 2015 3285 2035
rect 3315 2015 3335 2035
rect 3365 2015 3385 2035
rect 3415 2015 3435 2035
rect 3465 2015 3485 2035
rect 3515 2015 3535 2035
rect 3565 2015 3585 2035
rect 3615 2015 3635 2035
rect 3665 2015 3685 2035
rect 3715 2015 3735 2035
rect 3765 2015 3785 2035
rect 3815 2015 3835 2035
rect 3865 2015 3885 2035
rect 3915 2015 3935 2035
rect 3965 2015 3985 2035
rect 4015 2015 4035 2035
rect 4065 2015 4085 2035
rect 4115 2015 4135 2035
rect 4165 2015 4185 2035
rect 4215 2015 4235 2035
rect 4265 2015 4285 2035
rect 4315 2015 4335 2035
rect 4365 2015 4385 2035
rect 4415 2015 4435 2035
rect 4465 2015 4485 2035
rect 4515 2015 4535 2035
rect 4565 2015 4585 2035
rect 4615 2015 4635 2035
rect 4665 2015 4685 2035
rect 4715 2015 4735 2035
rect 4765 2015 4785 2035
rect 4815 2015 4835 2035
rect 4865 2015 4885 2035
rect 4915 2015 4935 2035
rect 4965 2015 4985 2035
rect 5015 2015 5035 2035
rect 5065 2015 5085 2035
rect 5115 2015 5135 2035
rect 5165 2015 5185 2035
rect 5215 2015 5235 2035
rect 5265 2015 5285 2035
rect 5315 2015 5335 2035
rect 5365 2015 5385 2035
rect 5415 2015 5435 2035
rect 5465 2015 5485 2035
rect 5515 2015 5535 2035
rect 5565 2015 5585 2035
rect 5615 2015 5635 2035
rect 5665 2015 5685 2035
rect 5715 2015 5735 2035
rect 5765 2015 5785 2035
rect 5815 2015 5835 2035
rect 5865 2015 5885 2035
rect 5915 2015 5935 2035
rect 5965 2015 5985 2035
rect 6015 2015 6035 2035
rect 6065 2015 6085 2035
rect 6115 2015 6135 2035
rect 6165 2015 6185 2035
rect 6215 2015 6235 2035
rect 6265 2015 6285 2035
rect 6315 2015 6335 2035
rect 6365 2015 6385 2035
rect 6415 2015 6435 2035
rect 6465 2015 6485 2035
rect 6515 2015 6535 2035
rect 6565 2015 6585 2035
rect 6615 2015 6635 2035
rect 6665 2015 6685 2035
rect 6715 2015 6735 2035
rect 6765 2015 6785 2035
rect 6815 2015 6835 2035
rect 6865 2015 6885 2035
rect 6915 2015 6935 2035
rect 6965 2015 6985 2035
rect 7015 2015 7035 2035
rect 7065 2015 7085 2035
rect 7115 2015 7135 2035
rect 7165 2015 7185 2035
rect 7215 2015 7235 2035
rect 7265 2015 7285 2035
rect 7315 2015 7335 2035
rect 7365 2015 7385 2035
rect 7415 2015 7435 2035
rect 7465 2015 7485 2035
rect 7515 2015 7535 2035
rect 7565 2015 7585 2035
rect 7615 2015 7635 2035
rect 7665 2015 7685 2035
rect 7715 2015 7735 2035
rect 7765 2015 7785 2035
rect 7815 2015 7835 2035
rect 7865 2015 7885 2035
rect 7915 2015 7935 2035
rect 7965 2015 7985 2035
rect 8015 2015 8035 2035
rect 8065 2015 8085 2035
rect 8115 2015 8135 2035
rect 8165 2015 8185 2035
rect 8215 2015 8235 2035
rect 8265 2015 8285 2035
rect 8315 2015 8335 2035
rect 8365 2015 8385 2035
rect 8415 2015 8435 2035
rect 8465 2015 8485 2035
rect 8515 2015 8535 2035
rect 8565 2015 8585 2035
rect 8615 2015 8635 2035
rect 8665 2015 8685 2035
rect 8715 2015 8735 2035
rect 8765 2015 8785 2035
rect 8815 2015 8835 2035
rect 8865 2015 8885 2035
rect 8915 2015 8935 2035
rect 8965 2015 8985 2035
rect 9015 2015 9035 2035
rect 9065 2015 9085 2035
rect 9115 2015 9135 2035
rect 9165 2015 9185 2035
rect 9215 2015 9235 2035
rect 9265 2015 9285 2035
rect 9315 2015 9335 2035
rect 9365 2015 9385 2035
rect 9415 2015 9435 2035
rect 9465 2015 9485 2035
rect 9515 2015 9535 2035
rect 9565 2015 9585 2035
rect 9615 2015 9635 2035
rect 9665 2015 9685 2035
rect 9715 2015 9735 2035
rect 9765 2015 9785 2035
rect 9815 2015 9835 2035
rect 9865 2015 9885 2035
rect 9915 2015 9935 2035
rect 9965 2015 9985 2035
rect 10015 2015 10035 2035
rect 10065 2015 10085 2035
rect 10115 2015 10135 2035
rect 10165 2015 10185 2035
rect 10215 2015 10235 2035
rect 10265 2015 10285 2035
rect 10315 2015 10335 2035
rect 10365 2015 10385 2035
rect 10415 2015 10435 2035
rect 10465 2015 10485 2035
rect 10515 2015 10535 2035
rect 10565 2015 10585 2035
rect 10615 2015 10635 2035
rect 10665 2015 10685 2035
rect 10715 2015 10735 2035
rect 10765 2015 10785 2035
rect 10815 2015 10835 2035
rect 10865 2015 10885 2035
rect 10915 2015 10935 2035
rect 10965 2015 10985 2035
rect 11015 2015 11035 2035
rect 11065 2015 11085 2035
rect 11115 2015 11135 2035
rect 11165 2015 11185 2035
rect 11215 2015 11235 2035
rect 11265 2015 11285 2035
rect 11315 2015 11335 2035
rect 11365 2015 11385 2035
rect 11415 2015 11435 2035
rect 11465 2015 11485 2035
rect 11515 2015 11535 2035
rect 11565 2015 11585 2035
rect 11615 2015 11635 2035
rect 11665 2015 11685 2035
rect 11715 2015 11735 2035
rect 11765 2015 11785 2035
rect 11815 2015 11835 2035
rect 11865 2015 11885 2035
rect 11915 2015 11935 2035
rect 11965 2015 11985 2035
rect 12015 2015 12035 2035
rect 12065 2015 12085 2035
rect 12115 2015 12135 2035
rect 12165 2015 12185 2035
rect 12215 2015 12235 2035
rect 12265 2015 12285 2035
rect 12315 2015 12335 2035
rect 12365 2015 12385 2035
rect 12415 2015 12435 2035
rect 12465 2015 12485 2035
rect 12515 2015 12535 2035
rect 12565 2015 12585 2035
rect 12615 2015 12635 2035
rect 12665 2015 12685 2035
rect 12715 2015 12735 2035
rect 12765 2015 12785 2035
rect 12815 2015 12835 2035
rect 12865 2015 12885 2035
rect 12915 2015 12935 2035
rect 12965 2015 12985 2035
rect 13015 2015 13035 2035
rect 13065 2015 13085 2035
rect 13115 2015 13135 2035
rect 13165 2015 13185 2035
rect 13215 2015 13235 2035
rect 13265 2015 13285 2035
rect 13315 2015 13335 2035
rect 13365 2015 13385 2035
rect 13415 2015 13435 2035
rect 13465 2015 13485 2035
rect 13515 2015 13535 2035
rect 13565 2015 13585 2035
rect 13615 2015 13635 2035
rect 13665 2015 13685 2035
rect 13715 2015 13735 2035
rect 13765 2015 13785 2035
rect 13815 2015 13835 2035
rect 13865 2015 13885 2035
rect 13915 2015 13935 2035
rect 13965 2015 13985 2035
rect 14015 2015 14035 2035
rect 14065 2015 14085 2035
rect 14115 2015 14135 2035
rect 14165 2015 14185 2035
rect 14215 2015 14235 2035
rect 14265 2015 14285 2035
rect 14315 2015 14335 2035
rect 14365 2015 14385 2035
rect 14415 2015 14435 2035
rect 14465 2015 14485 2035
rect 14515 2015 14535 2035
rect 14565 2015 14585 2035
rect 14615 2015 14635 2035
rect 14665 2015 14685 2035
rect 14715 2015 14735 2035
rect 14765 2015 14785 2035
rect 14815 2015 14835 2035
rect 14865 2015 14885 2035
rect 14915 2015 14935 2035
rect 14965 2015 14985 2035
rect 15015 2015 15035 2035
rect 15065 2015 15085 2035
rect 15115 2015 15135 2035
rect 15165 2015 15185 2035
rect 15215 2015 15235 2035
rect 15265 2015 15285 2035
rect 15315 2015 15335 2035
rect 15365 2015 15385 2035
rect 15415 2015 15435 2035
rect 15465 2015 15485 2035
rect 15515 2015 15535 2035
rect 15565 2015 15585 2035
rect 15615 2015 15635 2035
rect 15665 2015 15685 2035
rect 15715 2015 15735 2035
rect 15765 2015 15785 2035
rect 15815 2015 15835 2035
rect 15865 2015 15885 2035
rect 15915 2015 15935 2035
rect 15965 2015 15985 2035
rect 16015 2015 16035 2035
rect 16065 2015 16085 2035
rect 16115 2015 16135 2035
rect 16165 2015 16185 2035
rect 16215 2015 16235 2035
rect 16265 2015 16285 2035
rect 16315 2015 16335 2035
rect 16365 2015 16385 2035
rect 16415 2015 16435 2035
rect 16465 2015 16485 2035
rect 16515 2015 16535 2035
rect 16565 2015 16585 2035
rect 16615 2015 16635 2035
rect 16665 2015 16685 2035
rect 16715 2015 16735 2035
rect 16765 2015 16785 2035
rect 16815 2015 16835 2035
rect 16865 2015 16885 2035
rect 16915 2015 16935 2035
rect 16965 2015 16985 2035
rect 17015 2015 17035 2035
rect 17065 2015 17085 2035
rect 17115 2015 17135 2035
rect 17165 2015 17185 2035
rect 17215 2015 17235 2035
rect 17265 2015 17285 2035
rect 17315 2015 17335 2035
rect 17365 2015 17385 2035
rect 17415 2015 17435 2035
rect 17465 2015 17485 2035
rect 17515 2015 17535 2035
rect 17565 2015 17585 2035
rect 17615 2015 17635 2035
rect 17665 2015 17685 2035
rect 17715 2015 17735 2035
rect 17765 2015 17785 2035
rect 17815 2015 17835 2035
rect 17865 2015 17885 2035
rect 17915 2015 17935 2035
rect 17965 2015 17985 2035
rect 18015 2015 18035 2035
rect 18065 2015 18085 2035
rect 18115 2015 18135 2035
rect 18165 2015 18185 2035
rect 18215 2015 18235 2035
rect 18265 2015 18285 2035
rect 18315 2015 18335 2035
rect 18365 2015 18385 2035
rect 18415 2015 18435 2035
rect 18465 2015 18485 2035
rect 18515 2015 18535 2035
rect 18565 2015 18585 2035
rect 18615 2015 18635 2035
rect 18665 2015 18685 2035
rect 18715 2015 18735 2035
rect 18765 2015 18785 2035
rect 18815 2015 18835 2035
rect 18865 2015 18885 2035
rect 18915 2015 18935 2035
rect 18965 2015 18985 2035
rect 19015 2015 19035 2035
rect 19065 2015 19085 2035
rect 19115 2015 19135 2035
rect 19165 2015 19185 2035
rect 19215 2015 19235 2035
rect 19265 2015 19285 2035
rect 19315 2015 19335 2035
rect 19365 2015 19385 2035
rect 19415 2015 19435 2035
rect 19465 2015 19485 2035
rect 19515 2015 19535 2035
rect 19565 2015 19585 2035
rect 19615 2015 19635 2035
rect 19665 2015 19685 2035
rect 19715 2015 19735 2035
rect 19765 2015 19785 2035
rect 19815 2015 19835 2035
rect 19865 2015 19885 2035
rect 19915 2015 19935 2035
rect 19965 2015 19985 2035
rect 20015 2015 20035 2035
rect 20065 2015 20085 2035
rect 20115 2015 20135 2035
rect 20165 2015 20185 2035
rect 20215 2015 20235 2035
rect 20265 2015 20285 2035
rect 20315 2015 20335 2035
rect 20365 2015 20385 2035
rect 20415 2015 20435 2035
rect 20465 2015 20485 2035
rect 20515 2015 20535 2035
rect 20565 2015 20585 2035
rect 20615 2015 20635 2035
rect 20665 2015 20685 2035
rect 20715 2015 20735 2035
rect 20765 2015 20785 2035
rect 20815 2015 20835 2035
rect 20865 2015 20885 2035
rect 20915 2015 20935 2035
rect 20965 2015 20985 2035
rect 21015 2015 21035 2035
rect 21065 2015 21085 2035
rect 21115 2015 21135 2035
rect 21165 2015 21185 2035
rect 21215 2015 21235 2035
rect 21265 2015 21285 2035
rect 21315 2015 21335 2035
rect 21365 2015 21385 2035
rect 21415 2015 21435 2035
rect 21465 2015 21485 2035
rect 21515 2015 21535 2035
rect 21565 2015 21585 2035
rect 21615 2015 21635 2035
rect 21665 2015 21685 2035
rect 21715 2015 21735 2035
rect 21765 2015 21785 2035
rect 21815 2015 21835 2035
rect 21865 2015 21885 2035
rect 21915 2015 21935 2035
rect 21965 2015 21985 2035
rect 22015 2015 22035 2035
rect 22065 2015 22085 2035
rect 22115 2015 22135 2035
rect 22165 2015 22185 2035
rect 22215 2015 22235 2035
rect 22265 2015 22285 2035
rect 22315 2015 22335 2035
rect 22365 2015 22385 2035
rect 22415 2015 22435 2035
rect 22465 2015 22485 2035
rect 22515 2015 22535 2035
rect 22565 2015 22585 2035
rect 22615 2015 22635 2035
rect 22665 2015 22685 2035
rect 22715 2015 22735 2035
rect 22765 2015 22785 2035
rect 22815 2015 22835 2035
rect 22865 2015 22885 2035
rect 22915 2015 22935 2035
rect 22965 2015 22985 2035
rect 23015 2015 23035 2035
rect 23065 2015 23085 2035
rect 23115 2015 23135 2035
rect 23165 2015 23185 2035
rect 23215 2015 23235 2035
rect 23265 2015 23285 2035
rect 23315 2015 23335 2035
rect 23365 2015 23385 2035
rect 23415 2015 23435 2035
rect 23465 2015 23485 2035
rect 23515 2015 23535 2035
rect 23565 2015 23585 2035
rect 23615 2015 23635 2035
rect 23665 2015 23685 2035
rect 23715 2015 23735 2035
rect 23765 2015 23785 2035
rect 23815 2015 23835 2035
rect 23865 2015 23885 2035
rect 23915 2015 23935 2035
rect 23965 2015 23985 2035
rect 24015 2015 24035 2035
rect 24065 2015 24085 2035
rect 24115 2015 24135 2035
rect 24165 2015 24185 2035
rect 24215 2015 24235 2035
rect 24265 2015 24285 2035
rect 24315 2015 24335 2035
rect 24365 2015 24385 2035
rect 24415 2015 24435 2035
rect 24465 2015 24485 2035
rect 24515 2015 24535 2035
rect 24565 2015 24585 2035
rect 24615 2015 24635 2035
rect 24665 2015 24685 2035
rect 24715 2015 24735 2035
rect 24765 2015 24785 2035
rect 24815 2015 24835 2035
rect 24865 2015 24885 2035
rect 24915 2015 24935 2035
rect 24965 2015 24985 2035
rect 25015 2015 25035 2035
rect 25065 2015 25085 2035
rect 25115 2015 25135 2035
rect 25165 2015 25185 2035
rect 25215 2015 25235 2035
rect 25265 2015 25285 2035
rect 25315 2015 25335 2035
rect 25365 2015 25385 2035
rect 25415 2015 25435 2035
rect 25465 2015 25485 2035
rect 25515 2015 25535 2035
rect 25565 2015 25585 2035
rect 25615 2015 25635 2035
rect 25665 2015 25685 2035
rect 25715 2015 25735 2035
rect 25765 2015 25785 2035
rect 25815 2015 25835 2035
rect 25865 2015 25885 2035
rect 25915 2015 25935 2035
rect 25965 2015 25985 2035
rect 26015 2015 26035 2035
rect 26065 2015 26085 2035
rect 26115 2015 26135 2035
rect 26165 2015 26185 2035
rect 26215 2015 26235 2035
rect 26265 2015 26285 2035
rect 26315 2015 26335 2035
rect 26365 2015 26385 2035
rect 26415 2015 26435 2035
rect 26465 2015 26485 2035
rect 26515 2015 26535 2035
rect 26565 2015 26585 2035
rect 26615 2015 26635 2035
rect 26665 2015 26685 2035
rect 26715 2015 26735 2035
rect 26765 2015 26785 2035
rect 26815 2015 26835 2035
rect 26865 2015 26885 2035
rect 26915 2015 26935 2035
rect 26965 2015 26985 2035
rect 27015 2015 27035 2035
rect 27065 2015 27085 2035
rect 27115 2015 27135 2035
rect 27165 2015 27185 2035
rect 27215 2015 27235 2035
rect 27265 2015 27285 2035
rect 27315 2015 27335 2035
rect 27365 2015 27385 2035
rect 27415 2015 27435 2035
rect 27465 2015 27485 2035
rect 27515 2015 27535 2035
rect 27565 2015 27585 2035
rect 27615 2015 27635 2035
rect 27665 2015 27685 2035
rect 27715 2015 27735 2035
rect 27765 2015 27785 2035
rect 27815 2015 27835 2035
rect 27865 2015 27885 2035
rect 27915 2015 27935 2035
rect 27965 2015 27985 2035
rect 28015 2015 28035 2035
rect 28065 2015 28085 2035
rect 28115 2015 28135 2035
rect 28165 2015 28185 2035
rect 28215 2015 28235 2035
rect 28265 2015 28285 2035
rect 28315 2015 28335 2035
rect 28365 2015 28385 2035
rect 28415 2015 28435 2035
rect 28465 2015 28485 2035
rect 28515 2015 28535 2035
rect 28565 2015 28585 2035
rect 28615 2015 28635 2035
rect 28665 2015 28685 2035
rect 28715 2015 28735 2035
rect 28765 2015 28785 2035
rect -635 1665 -615 1685
rect -585 1665 -565 1685
rect -535 1665 -515 1685
rect -485 1665 -465 1685
rect -435 1665 -415 1685
rect -385 1665 -365 1685
rect -335 1665 -315 1685
rect -285 1665 -265 1685
rect -235 1665 -215 1685
rect -185 1665 -165 1685
rect -135 1665 -115 1685
rect -85 1665 -65 1685
rect -35 1665 -15 1685
rect 15 1665 35 1685
rect 65 1665 85 1685
rect 115 1665 135 1685
rect 165 1665 185 1685
rect 215 1665 235 1685
rect 265 1665 285 1685
rect 315 1665 335 1685
rect 365 1665 385 1685
rect 415 1665 435 1685
rect 465 1665 485 1685
rect 515 1665 535 1685
rect 565 1665 585 1685
rect 615 1665 635 1685
rect 665 1665 685 1685
rect 715 1665 735 1685
rect 765 1665 785 1685
rect 815 1665 835 1685
rect 865 1665 885 1685
rect 915 1665 935 1685
rect 965 1665 985 1685
rect 1015 1665 1035 1685
rect 1065 1665 1085 1685
rect 1115 1665 1135 1685
rect 1165 1665 1185 1685
rect 1215 1665 1235 1685
rect 1265 1665 1285 1685
rect 1315 1665 1335 1685
rect 1365 1665 1385 1685
rect 1415 1665 1435 1685
rect 1465 1665 1485 1685
rect 1515 1665 1535 1685
rect 1565 1665 1585 1685
rect 1615 1665 1635 1685
rect 1665 1665 1685 1685
rect 1715 1665 1735 1685
rect 1765 1665 1785 1685
rect 1815 1665 1835 1685
rect 1865 1665 1885 1685
rect 1915 1665 1935 1685
rect 1965 1665 1985 1685
rect 2015 1665 2035 1685
rect 2065 1665 2085 1685
rect 2115 1665 2135 1685
rect 2165 1665 2185 1685
rect 2215 1665 2235 1685
rect 2265 1665 2285 1685
rect 2315 1665 2335 1685
rect 2365 1665 2385 1685
rect 2415 1665 2435 1685
rect 2465 1665 2485 1685
rect 2515 1665 2535 1685
rect 2565 1665 2585 1685
rect 2615 1665 2635 1685
rect 2665 1665 2685 1685
rect 2715 1665 2735 1685
rect 2765 1665 2785 1685
rect 2815 1665 2835 1685
rect 2865 1665 2885 1685
rect 2915 1665 2935 1685
rect 2965 1665 2985 1685
rect 3015 1665 3035 1685
rect 3065 1665 3085 1685
rect 3115 1665 3135 1685
rect 3165 1665 3185 1685
rect 3215 1665 3235 1685
rect 3265 1665 3285 1685
rect 3315 1665 3335 1685
rect 3365 1665 3385 1685
rect 3415 1665 3435 1685
rect 3465 1665 3485 1685
rect 3515 1665 3535 1685
rect 3565 1665 3585 1685
rect 3615 1665 3635 1685
rect 3665 1665 3685 1685
rect 3715 1665 3735 1685
rect 3765 1665 3785 1685
rect 3815 1665 3835 1685
rect 3865 1665 3885 1685
rect 3915 1665 3935 1685
rect 3965 1665 3985 1685
rect 4015 1665 4035 1685
rect 4065 1665 4085 1685
rect 4115 1665 4135 1685
rect 4165 1665 4185 1685
rect 4215 1665 4235 1685
rect 4265 1665 4285 1685
rect 4315 1665 4335 1685
rect 4365 1665 4385 1685
rect 4415 1665 4435 1685
rect 4465 1665 4485 1685
rect 4515 1665 4535 1685
rect 4565 1665 4585 1685
rect 4615 1665 4635 1685
rect 4665 1665 4685 1685
rect 4715 1665 4735 1685
rect 4765 1665 4785 1685
rect 4815 1665 4835 1685
rect 4865 1665 4885 1685
rect 4915 1665 4935 1685
rect 4965 1665 4985 1685
rect 5015 1665 5035 1685
rect 5065 1665 5085 1685
rect 5115 1665 5135 1685
rect 5165 1665 5185 1685
rect 5215 1665 5235 1685
rect 5265 1665 5285 1685
rect 5315 1665 5335 1685
rect 5365 1665 5385 1685
rect 5415 1665 5435 1685
rect 5465 1665 5485 1685
rect 5515 1665 5535 1685
rect 5565 1665 5585 1685
rect 5615 1665 5635 1685
rect 5665 1665 5685 1685
rect 5715 1665 5735 1685
rect 5765 1665 5785 1685
rect 5815 1665 5835 1685
rect 5865 1665 5885 1685
rect 5915 1665 5935 1685
rect 5965 1665 5985 1685
rect 6015 1665 6035 1685
rect 6065 1665 6085 1685
rect 6115 1665 6135 1685
rect 6165 1665 6185 1685
rect 6215 1665 6235 1685
rect 6265 1665 6285 1685
rect 6315 1665 6335 1685
rect 6365 1665 6385 1685
rect 6415 1665 6435 1685
rect 6465 1665 6485 1685
rect 6515 1665 6535 1685
rect 6565 1665 6585 1685
rect 6615 1665 6635 1685
rect 6665 1665 6685 1685
rect 6715 1665 6735 1685
rect 6765 1665 6785 1685
rect 6815 1665 6835 1685
rect 6865 1665 6885 1685
rect 6915 1665 6935 1685
rect 6965 1665 6985 1685
rect 7015 1665 7035 1685
rect 7065 1665 7085 1685
rect 7115 1665 7135 1685
rect 7165 1665 7185 1685
rect 7215 1665 7235 1685
rect 7265 1665 7285 1685
rect 7315 1665 7335 1685
rect 7365 1665 7385 1685
rect 7415 1665 7435 1685
rect 7465 1665 7485 1685
rect 7515 1665 7535 1685
rect 7565 1665 7585 1685
rect 7615 1665 7635 1685
rect 7665 1665 7685 1685
rect 7715 1665 7735 1685
rect 7765 1665 7785 1685
rect 7815 1665 7835 1685
rect 7865 1665 7885 1685
rect 7915 1665 7935 1685
rect 7965 1665 7985 1685
rect 8015 1665 8035 1685
rect 8065 1665 8085 1685
rect 8115 1665 8135 1685
rect 8165 1665 8185 1685
rect 8215 1665 8235 1685
rect 8265 1665 8285 1685
rect 8315 1665 8335 1685
rect 8365 1665 8385 1685
rect 8415 1665 8435 1685
rect 8465 1665 8485 1685
rect 8515 1665 8535 1685
rect 8565 1665 8585 1685
rect 8615 1665 8635 1685
rect 8665 1665 8685 1685
rect 8715 1665 8735 1685
rect 8765 1665 8785 1685
rect 8815 1665 8835 1685
rect 8865 1665 8885 1685
rect 8915 1665 8935 1685
rect 8965 1665 8985 1685
rect 9015 1665 9035 1685
rect 9065 1665 9085 1685
rect 9115 1665 9135 1685
rect 9165 1665 9185 1685
rect 9215 1665 9235 1685
rect 9265 1665 9285 1685
rect 9315 1665 9335 1685
rect 9365 1665 9385 1685
rect 9415 1665 9435 1685
rect 9465 1665 9485 1685
rect 9515 1665 9535 1685
rect 9565 1665 9585 1685
rect 9615 1665 9635 1685
rect 9665 1665 9685 1685
rect 9715 1665 9735 1685
rect 9765 1665 9785 1685
rect 9815 1665 9835 1685
rect 9865 1665 9885 1685
rect 9915 1665 9935 1685
rect 9965 1665 9985 1685
rect 10015 1665 10035 1685
rect 10065 1665 10085 1685
rect 10115 1665 10135 1685
rect 10165 1665 10185 1685
rect 10215 1665 10235 1685
rect 10265 1665 10285 1685
rect 10315 1665 10335 1685
rect 10365 1665 10385 1685
rect 10415 1665 10435 1685
rect 10465 1665 10485 1685
rect 10515 1665 10535 1685
rect 10565 1665 10585 1685
rect 10615 1665 10635 1685
rect 10665 1665 10685 1685
rect 10715 1665 10735 1685
rect 10765 1665 10785 1685
rect 10815 1665 10835 1685
rect 10865 1665 10885 1685
rect 10915 1665 10935 1685
rect 10965 1665 10985 1685
rect 11015 1665 11035 1685
rect 11065 1665 11085 1685
rect 11115 1665 11135 1685
rect 11165 1665 11185 1685
rect 11215 1665 11235 1685
rect 11265 1665 11285 1685
rect 11315 1665 11335 1685
rect 11365 1665 11385 1685
rect 11415 1665 11435 1685
rect 11465 1665 11485 1685
rect 11515 1665 11535 1685
rect 11565 1665 11585 1685
rect 11615 1665 11635 1685
rect 11665 1665 11685 1685
rect 11715 1665 11735 1685
rect 11765 1665 11785 1685
rect 11815 1665 11835 1685
rect 11865 1665 11885 1685
rect 11915 1665 11935 1685
rect 11965 1665 11985 1685
rect 12015 1665 12035 1685
rect 12065 1665 12085 1685
rect 12115 1665 12135 1685
rect 12165 1665 12185 1685
rect 12215 1665 12235 1685
rect 12265 1665 12285 1685
rect 12315 1665 12335 1685
rect 12365 1665 12385 1685
rect 12415 1665 12435 1685
rect 12465 1665 12485 1685
rect 12515 1665 12535 1685
rect 12565 1665 12585 1685
rect 12615 1665 12635 1685
rect 12665 1665 12685 1685
rect 12715 1665 12735 1685
rect 12765 1665 12785 1685
rect 12815 1665 12835 1685
rect 12865 1665 12885 1685
rect 12915 1665 12935 1685
rect 12965 1665 12985 1685
rect 13015 1665 13035 1685
rect 13065 1665 13085 1685
rect 13115 1665 13135 1685
rect 13165 1665 13185 1685
rect 13215 1665 13235 1685
rect 13265 1665 13285 1685
rect 13315 1665 13335 1685
rect 13365 1665 13385 1685
rect 13415 1665 13435 1685
rect 13465 1665 13485 1685
rect 13515 1665 13535 1685
rect 13565 1665 13585 1685
rect 13615 1665 13635 1685
rect 13665 1665 13685 1685
rect 13715 1665 13735 1685
rect 13765 1665 13785 1685
rect 13815 1665 13835 1685
rect 13865 1665 13885 1685
rect 13915 1665 13935 1685
rect 13965 1665 13985 1685
rect 14015 1665 14035 1685
rect 14065 1665 14085 1685
rect 14115 1665 14135 1685
rect 14165 1665 14185 1685
rect 14215 1665 14235 1685
rect 14265 1665 14285 1685
rect 14315 1665 14335 1685
rect 14365 1665 14385 1685
rect 14415 1665 14435 1685
rect 14465 1665 14485 1685
rect 14515 1665 14535 1685
rect 14565 1665 14585 1685
rect 14615 1665 14635 1685
rect 14665 1665 14685 1685
rect 14715 1665 14735 1685
rect 14765 1665 14785 1685
rect 14815 1665 14835 1685
rect 14865 1665 14885 1685
rect 14915 1665 14935 1685
rect 14965 1665 14985 1685
rect 15015 1665 15035 1685
rect 15065 1665 15085 1685
rect 15115 1665 15135 1685
rect 15165 1665 15185 1685
rect 15215 1665 15235 1685
rect 15265 1665 15285 1685
rect 15315 1665 15335 1685
rect 15365 1665 15385 1685
rect 15415 1665 15435 1685
rect 15465 1665 15485 1685
rect 15515 1665 15535 1685
rect 15565 1665 15585 1685
rect 15615 1665 15635 1685
rect 15665 1665 15685 1685
rect 15715 1665 15735 1685
rect 15765 1665 15785 1685
rect 15815 1665 15835 1685
rect 15865 1665 15885 1685
rect 15915 1665 15935 1685
rect 15965 1665 15985 1685
rect 16015 1665 16035 1685
rect 16065 1665 16085 1685
rect 16115 1665 16135 1685
rect 16165 1665 16185 1685
rect 16215 1665 16235 1685
rect 16265 1665 16285 1685
rect 16315 1665 16335 1685
rect 16365 1665 16385 1685
rect 16415 1665 16435 1685
rect 16465 1665 16485 1685
rect 16515 1665 16535 1685
rect 16565 1665 16585 1685
rect 16615 1665 16635 1685
rect 16665 1665 16685 1685
rect 16715 1665 16735 1685
rect 16765 1665 16785 1685
rect 16815 1665 16835 1685
rect 16865 1665 16885 1685
rect 16915 1665 16935 1685
rect 16965 1665 16985 1685
rect 17015 1665 17035 1685
rect 17065 1665 17085 1685
rect 17115 1665 17135 1685
rect 17165 1665 17185 1685
rect 17215 1665 17235 1685
rect 17265 1665 17285 1685
rect 17315 1665 17335 1685
rect 17365 1665 17385 1685
rect 17415 1665 17435 1685
rect 17465 1665 17485 1685
rect 17515 1665 17535 1685
rect 17565 1665 17585 1685
rect 17615 1665 17635 1685
rect 17665 1665 17685 1685
rect 17715 1665 17735 1685
rect 17765 1665 17785 1685
rect 17815 1665 17835 1685
rect 17865 1665 17885 1685
rect 17915 1665 17935 1685
rect 17965 1665 17985 1685
rect 18015 1665 18035 1685
rect 18065 1665 18085 1685
rect 18115 1665 18135 1685
rect 18165 1665 18185 1685
rect 18215 1665 18235 1685
rect 18265 1665 18285 1685
rect 18315 1665 18335 1685
rect 18365 1665 18385 1685
rect 18415 1665 18435 1685
rect 18465 1665 18485 1685
rect 18515 1665 18535 1685
rect 18565 1665 18585 1685
rect 18615 1665 18635 1685
rect 18665 1665 18685 1685
rect 18715 1665 18735 1685
rect 18765 1665 18785 1685
rect 18815 1665 18835 1685
rect 18865 1665 18885 1685
rect 18915 1665 18935 1685
rect 18965 1665 18985 1685
rect 19015 1665 19035 1685
rect 19065 1665 19085 1685
rect 19115 1665 19135 1685
rect 19165 1665 19185 1685
rect 19215 1665 19235 1685
rect 19265 1665 19285 1685
rect 19315 1665 19335 1685
rect 19365 1665 19385 1685
rect 19415 1665 19435 1685
rect 19465 1665 19485 1685
rect 19515 1665 19535 1685
rect 19565 1665 19585 1685
rect 19615 1665 19635 1685
rect 19665 1665 19685 1685
rect 19715 1665 19735 1685
rect 19765 1665 19785 1685
rect 19815 1665 19835 1685
rect 19865 1665 19885 1685
rect 19915 1665 19935 1685
rect 19965 1665 19985 1685
rect 20015 1665 20035 1685
rect 20065 1665 20085 1685
rect 20115 1665 20135 1685
rect 20165 1665 20185 1685
rect 20215 1665 20235 1685
rect 20265 1665 20285 1685
rect 20315 1665 20335 1685
rect 20365 1665 20385 1685
rect 20415 1665 20435 1685
rect 20465 1665 20485 1685
rect 20515 1665 20535 1685
rect 20565 1665 20585 1685
rect 20615 1665 20635 1685
rect 20665 1665 20685 1685
rect 20715 1665 20735 1685
rect 20765 1665 20785 1685
rect 20815 1665 20835 1685
rect 20865 1665 20885 1685
rect 20915 1665 20935 1685
rect 20965 1665 20985 1685
rect 21015 1665 21035 1685
rect 21065 1665 21085 1685
rect 21115 1665 21135 1685
rect 21165 1665 21185 1685
rect 21215 1665 21235 1685
rect 21265 1665 21285 1685
rect 21315 1665 21335 1685
rect 21365 1665 21385 1685
rect 21415 1665 21435 1685
rect 21465 1665 21485 1685
rect 21515 1665 21535 1685
rect 21565 1665 21585 1685
rect 21615 1665 21635 1685
rect 21665 1665 21685 1685
rect 21715 1665 21735 1685
rect 21765 1665 21785 1685
rect 21815 1665 21835 1685
rect 21865 1665 21885 1685
rect 21915 1665 21935 1685
rect 21965 1665 21985 1685
rect 22015 1665 22035 1685
rect 22065 1665 22085 1685
rect 22115 1665 22135 1685
rect 22165 1665 22185 1685
rect 22215 1665 22235 1685
rect 22265 1665 22285 1685
rect 22315 1665 22335 1685
rect 22365 1665 22385 1685
rect 22415 1665 22435 1685
rect 22465 1665 22485 1685
rect 22515 1665 22535 1685
rect 22565 1665 22585 1685
rect 22615 1665 22635 1685
rect 22665 1665 22685 1685
rect 22715 1665 22735 1685
rect 22765 1665 22785 1685
rect 22815 1665 22835 1685
rect 22865 1665 22885 1685
rect 22915 1665 22935 1685
rect 22965 1665 22985 1685
rect 23015 1665 23035 1685
rect 23065 1665 23085 1685
rect 23115 1665 23135 1685
rect 23165 1665 23185 1685
rect 23215 1665 23235 1685
rect 23265 1665 23285 1685
rect 23315 1665 23335 1685
rect 23365 1665 23385 1685
rect 23415 1665 23435 1685
rect 23465 1665 23485 1685
rect 23515 1665 23535 1685
rect 23565 1665 23585 1685
rect 23615 1665 23635 1685
rect 23665 1665 23685 1685
rect 23715 1665 23735 1685
rect 23765 1665 23785 1685
rect 23815 1665 23835 1685
rect 23865 1665 23885 1685
rect 23915 1665 23935 1685
rect 23965 1665 23985 1685
rect 24015 1665 24035 1685
rect 24065 1665 24085 1685
rect 24115 1665 24135 1685
rect 24165 1665 24185 1685
rect 24215 1665 24235 1685
rect 24265 1665 24285 1685
rect 24315 1665 24335 1685
rect 24365 1665 24385 1685
rect 24415 1665 24435 1685
rect 24465 1665 24485 1685
rect 24515 1665 24535 1685
rect 24565 1665 24585 1685
rect 24615 1665 24635 1685
rect 24665 1665 24685 1685
rect 24715 1665 24735 1685
rect 24765 1665 24785 1685
rect 24815 1665 24835 1685
rect 24865 1665 24885 1685
rect 24915 1665 24935 1685
rect 24965 1665 24985 1685
rect 25015 1665 25035 1685
rect 25065 1665 25085 1685
rect 25115 1665 25135 1685
rect 25165 1665 25185 1685
rect 25215 1665 25235 1685
rect 25265 1665 25285 1685
rect 25315 1665 25335 1685
rect 25365 1665 25385 1685
rect 25415 1665 25435 1685
rect 25465 1665 25485 1685
rect 25515 1665 25535 1685
rect 25565 1665 25585 1685
rect 25615 1665 25635 1685
rect 25665 1665 25685 1685
rect 25715 1665 25735 1685
rect 25765 1665 25785 1685
rect 25815 1665 25835 1685
rect 25865 1665 25885 1685
rect 25915 1665 25935 1685
rect 25965 1665 25985 1685
rect 26015 1665 26035 1685
rect 26065 1665 26085 1685
rect 26115 1665 26135 1685
rect 26165 1665 26185 1685
rect 26215 1665 26235 1685
rect 26265 1665 26285 1685
rect 26315 1665 26335 1685
rect 26365 1665 26385 1685
rect 26415 1665 26435 1685
rect 26465 1665 26485 1685
rect 26515 1665 26535 1685
rect 26565 1665 26585 1685
rect 26615 1665 26635 1685
rect 26665 1665 26685 1685
rect 26715 1665 26735 1685
rect 26765 1665 26785 1685
rect 26815 1665 26835 1685
rect 26865 1665 26885 1685
rect 26915 1665 26935 1685
rect 26965 1665 26985 1685
rect 27015 1665 27035 1685
rect 27065 1665 27085 1685
rect 27115 1665 27135 1685
rect 27165 1665 27185 1685
rect 27215 1665 27235 1685
rect 27265 1665 27285 1685
rect 27315 1665 27335 1685
rect 27365 1665 27385 1685
rect 27415 1665 27435 1685
rect 27465 1665 27485 1685
rect 27515 1665 27535 1685
rect 27565 1665 27585 1685
rect 27615 1665 27635 1685
rect 27665 1665 27685 1685
rect 27715 1665 27735 1685
rect 27765 1665 27785 1685
rect 27815 1665 27835 1685
rect 27865 1665 27885 1685
rect 27915 1665 27935 1685
rect 27965 1665 27985 1685
rect 28015 1665 28035 1685
rect 28065 1665 28085 1685
rect 28115 1665 28135 1685
rect 28165 1665 28185 1685
rect 28215 1665 28235 1685
rect 28265 1665 28285 1685
rect 28315 1665 28335 1685
rect 28365 1665 28385 1685
rect 28415 1665 28435 1685
rect 28465 1665 28485 1685
rect 28515 1665 28535 1685
rect 28565 1665 28585 1685
rect 28615 1665 28635 1685
rect 28665 1665 28685 1685
rect 28715 1665 28735 1685
rect 28765 1665 28785 1685
rect -635 -35 -615 -15
rect -585 -35 -565 -15
rect -535 -35 -515 -15
rect -485 -35 -465 -15
rect -435 -35 -415 -15
rect -385 -35 -365 -15
rect -335 -35 -315 -15
rect -285 -35 -265 -15
rect -235 -35 -215 -15
rect -185 -35 -165 -15
rect -135 -35 -115 -15
rect -85 -35 -65 -15
rect -35 -35 -15 -15
rect 15 -35 35 -15
rect 65 -35 85 -15
rect 115 -35 135 -15
rect 165 -35 185 -15
rect 215 -35 235 -15
rect 265 -35 285 -15
rect 315 -35 335 -15
rect 365 -35 385 -15
rect 415 -35 435 -15
rect 465 -35 485 -15
rect 515 -35 535 -15
rect 565 -35 585 -15
rect 615 -35 635 -15
rect 665 -35 685 -15
rect 715 -35 735 -15
rect 765 -35 785 -15
rect 815 -35 835 -15
rect 865 -35 885 -15
rect 915 -35 935 -15
rect 965 -35 985 -15
rect 1015 -35 1035 -15
rect 1065 -35 1085 -15
rect 1115 -35 1135 -15
rect 1165 -35 1185 -15
rect 1215 -35 1235 -15
rect 1265 -35 1285 -15
rect 1315 -35 1335 -15
rect 1365 -35 1385 -15
rect 1415 -35 1435 -15
rect 1465 -35 1485 -15
rect 1515 -35 1535 -15
rect 1565 -35 1585 -15
rect 1615 -35 1635 -15
rect 1665 -35 1685 -15
rect 1715 -35 1735 -15
rect 1765 -35 1785 -15
rect 1815 -35 1835 -15
rect 1865 -35 1885 -15
rect 1915 -35 1935 -15
rect 1965 -35 1985 -15
rect 2015 -35 2035 -15
rect 2065 -35 2085 -15
rect 2115 -35 2135 -15
rect 2165 -35 2185 -15
rect 2215 -35 2235 -15
rect 2265 -35 2285 -15
rect 2315 -35 2335 -15
rect 2365 -35 2385 -15
rect 2415 -35 2435 -15
rect 2465 -35 2485 -15
rect 2515 -35 2535 -15
rect 2565 -35 2585 -15
rect 2615 -35 2635 -15
rect 2665 -35 2685 -15
rect 2715 -35 2735 -15
rect 2765 -35 2785 -15
rect 2815 -35 2835 -15
rect 2865 -35 2885 -15
rect 2915 -35 2935 -15
rect 2965 -35 2985 -15
rect 3015 -35 3035 -15
rect 3065 -35 3085 -15
rect 3115 -35 3135 -15
rect 3165 -35 3185 -15
rect 3215 -35 3235 -15
rect 3265 -35 3285 -15
rect 3315 -35 3335 -15
rect 3365 -35 3385 -15
rect 3415 -35 3435 -15
rect 3465 -35 3485 -15
rect 3515 -35 3535 -15
rect 3565 -35 3585 -15
rect 3615 -35 3635 -15
rect 3665 -35 3685 -15
rect 3715 -35 3735 -15
rect 3765 -35 3785 -15
rect 3815 -35 3835 -15
rect 3865 -35 3885 -15
rect 3915 -35 3935 -15
rect 3965 -35 3985 -15
rect 4015 -35 4035 -15
rect 4065 -35 4085 -15
rect 4115 -35 4135 -15
rect 4165 -35 4185 -15
rect 4215 -35 4235 -15
rect 4265 -35 4285 -15
rect 4315 -35 4335 -15
rect 4365 -35 4385 -15
rect 4415 -35 4435 -15
rect 4465 -35 4485 -15
rect 4515 -35 4535 -15
rect 4565 -35 4585 -15
rect 4615 -35 4635 -15
rect 4665 -35 4685 -15
rect 4715 -35 4735 -15
rect 4765 -35 4785 -15
rect 4815 -35 4835 -15
rect 4865 -35 4885 -15
rect 4915 -35 4935 -15
rect 4965 -35 4985 -15
rect 5015 -35 5035 -15
rect 5065 -35 5085 -15
rect 5115 -35 5135 -15
rect 5165 -35 5185 -15
rect 5215 -35 5235 -15
rect 5265 -35 5285 -15
rect 5315 -35 5335 -15
rect 5365 -35 5385 -15
rect 5415 -35 5435 -15
rect 5465 -35 5485 -15
rect 5515 -35 5535 -15
rect 5565 -35 5585 -15
rect 5615 -35 5635 -15
rect 5665 -35 5685 -15
rect 5715 -35 5735 -15
rect 5765 -35 5785 -15
rect 5815 -35 5835 -15
rect 5865 -35 5885 -15
rect 5915 -35 5935 -15
rect 5965 -35 5985 -15
rect 6015 -35 6035 -15
rect 6065 -35 6085 -15
rect 6115 -35 6135 -15
rect 6165 -35 6185 -15
rect 6215 -35 6235 -15
rect 6265 -35 6285 -15
rect 6315 -35 6335 -15
rect 6365 -35 6385 -15
rect 6415 -35 6435 -15
rect 6465 -35 6485 -15
rect 6515 -35 6535 -15
rect 6565 -35 6585 -15
rect 6615 -35 6635 -15
rect 6665 -35 6685 -15
rect 6715 -35 6735 -15
rect 6765 -35 6785 -15
rect 6815 -35 6835 -15
rect 6865 -35 6885 -15
rect 6915 -35 6935 -15
rect 6965 -35 6985 -15
rect 7015 -35 7035 -15
rect 7065 -35 7085 -15
rect 7115 -35 7135 -15
rect 7165 -35 7185 -15
rect 7215 -35 7235 -15
rect 7265 -35 7285 -15
rect 7315 -35 7335 -15
rect 7365 -35 7385 -15
rect 7415 -35 7435 -15
rect 7465 -35 7485 -15
rect 7515 -35 7535 -15
rect 7565 -35 7585 -15
rect 7615 -35 7635 -15
rect 7665 -35 7685 -15
rect 7715 -35 7735 -15
rect 7765 -35 7785 -15
rect 7815 -35 7835 -15
rect 7865 -35 7885 -15
rect 7915 -35 7935 -15
rect 7965 -35 7985 -15
rect 8015 -35 8035 -15
rect 8065 -35 8085 -15
rect 8115 -35 8135 -15
rect 8165 -35 8185 -15
rect 8215 -35 8235 -15
rect 8265 -35 8285 -15
rect 8315 -35 8335 -15
rect 8365 -35 8385 -15
rect 8415 -35 8435 -15
rect 8465 -35 8485 -15
rect 8515 -35 8535 -15
rect 8565 -35 8585 -15
rect 8615 -35 8635 -15
rect 8665 -35 8685 -15
rect 8715 -35 8735 -15
rect 8765 -35 8785 -15
rect 8815 -35 8835 -15
rect 8865 -35 8885 -15
rect 8915 -35 8935 -15
rect 8965 -35 8985 -15
rect 9015 -35 9035 -15
rect 9065 -35 9085 -15
rect 9115 -35 9135 -15
rect 9165 -35 9185 -15
rect 9215 -35 9235 -15
rect 9265 -35 9285 -15
rect 9315 -35 9335 -15
rect 9365 -35 9385 -15
rect 9415 -35 9435 -15
rect 9465 -35 9485 -15
rect 9515 -35 9535 -15
rect 9565 -35 9585 -15
rect 9615 -35 9635 -15
rect 9665 -35 9685 -15
rect 9715 -35 9735 -15
rect 9765 -35 9785 -15
rect 9815 -35 9835 -15
rect 9865 -35 9885 -15
rect 9915 -35 9935 -15
rect 9965 -35 9985 -15
rect 10015 -35 10035 -15
rect 10065 -35 10085 -15
rect 10115 -35 10135 -15
rect 10165 -35 10185 -15
rect 10215 -35 10235 -15
rect 10265 -35 10285 -15
rect 10315 -35 10335 -15
rect 10365 -35 10385 -15
rect 10415 -35 10435 -15
rect 10465 -35 10485 -15
rect 10515 -35 10535 -15
rect 10565 -35 10585 -15
rect 10615 -35 10635 -15
rect 10665 -35 10685 -15
rect 10715 -35 10735 -15
rect 10765 -35 10785 -15
rect 10815 -35 10835 -15
rect 10865 -35 10885 -15
rect 10915 -35 10935 -15
rect 10965 -35 10985 -15
rect 11015 -35 11035 -15
rect 11065 -35 11085 -15
rect 11115 -35 11135 -15
rect 11165 -35 11185 -15
rect 11215 -35 11235 -15
rect 11265 -35 11285 -15
rect 11315 -35 11335 -15
rect 11365 -35 11385 -15
rect 11415 -35 11435 -15
rect 11465 -35 11485 -15
rect 11515 -35 11535 -15
rect 11565 -35 11585 -15
rect 11615 -35 11635 -15
rect 11665 -35 11685 -15
rect 11715 -35 11735 -15
rect 11765 -35 11785 -15
rect 11815 -35 11835 -15
rect 11865 -35 11885 -15
rect 11915 -35 11935 -15
rect 11965 -35 11985 -15
rect 12015 -35 12035 -15
rect 12065 -35 12085 -15
rect 12115 -35 12135 -15
rect 12165 -35 12185 -15
rect 12215 -35 12235 -15
rect 12265 -35 12285 -15
rect 12315 -35 12335 -15
rect 12365 -35 12385 -15
rect 12415 -35 12435 -15
rect 12465 -35 12485 -15
rect 12515 -35 12535 -15
rect 12565 -35 12585 -15
rect 12615 -35 12635 -15
rect 12665 -35 12685 -15
rect 12715 -35 12735 -15
rect 12765 -35 12785 -15
rect 12815 -35 12835 -15
rect 12865 -35 12885 -15
rect 12915 -35 12935 -15
rect 12965 -35 12985 -15
rect 13015 -35 13035 -15
rect 13065 -35 13085 -15
rect 13115 -35 13135 -15
rect 13165 -35 13185 -15
rect 13215 -35 13235 -15
rect 13265 -35 13285 -15
rect 13315 -35 13335 -15
rect 13365 -35 13385 -15
rect 13415 -35 13435 -15
rect 13465 -35 13485 -15
rect 13515 -35 13535 -15
rect 13565 -35 13585 -15
rect 13615 -35 13635 -15
rect 13665 -35 13685 -15
rect 13715 -35 13735 -15
rect 13765 -35 13785 -15
rect 13815 -35 13835 -15
rect 13865 -35 13885 -15
rect 13915 -35 13935 -15
rect 13965 -35 13985 -15
rect 14015 -35 14035 -15
rect 14065 -35 14085 -15
rect 14115 -35 14135 -15
rect 14165 -35 14185 -15
rect 14215 -35 14235 -15
rect 14265 -35 14285 -15
rect 14315 -35 14335 -15
rect 14365 -35 14385 -15
rect 14415 -35 14435 -15
rect 14465 -35 14485 -15
rect 14515 -35 14535 -15
rect 14565 -35 14585 -15
rect 14615 -35 14635 -15
rect 14665 -35 14685 -15
rect 14715 -35 14735 -15
rect 14765 -35 14785 -15
rect 14815 -35 14835 -15
rect 14865 -35 14885 -15
rect 14915 -35 14935 -15
rect 14965 -35 14985 -15
rect 15015 -35 15035 -15
rect 15065 -35 15085 -15
rect 15115 -35 15135 -15
rect 15165 -35 15185 -15
rect 15215 -35 15235 -15
rect 15265 -35 15285 -15
rect 15315 -35 15335 -15
rect 15365 -35 15385 -15
rect 15415 -35 15435 -15
rect 15465 -35 15485 -15
rect 15515 -35 15535 -15
rect 15565 -35 15585 -15
rect 15615 -35 15635 -15
rect 15665 -35 15685 -15
rect 15715 -35 15735 -15
rect 15765 -35 15785 -15
rect 15815 -35 15835 -15
rect 15865 -35 15885 -15
rect 15915 -35 15935 -15
rect 15965 -35 15985 -15
rect 16015 -35 16035 -15
rect 16065 -35 16085 -15
rect 16115 -35 16135 -15
rect 16165 -35 16185 -15
rect 16215 -35 16235 -15
rect 16265 -35 16285 -15
rect 16315 -35 16335 -15
rect 16365 -35 16385 -15
rect 16415 -35 16435 -15
rect 16465 -35 16485 -15
rect 16515 -35 16535 -15
rect 16565 -35 16585 -15
rect 16615 -35 16635 -15
rect 16665 -35 16685 -15
rect 16715 -35 16735 -15
rect 16765 -35 16785 -15
rect 16815 -35 16835 -15
rect 16865 -35 16885 -15
rect 16915 -35 16935 -15
rect 16965 -35 16985 -15
rect 17015 -35 17035 -15
rect 17065 -35 17085 -15
rect 17115 -35 17135 -15
rect 17165 -35 17185 -15
rect 17215 -35 17235 -15
rect 17265 -35 17285 -15
rect 17315 -35 17335 -15
rect 17365 -35 17385 -15
rect 17415 -35 17435 -15
rect 17465 -35 17485 -15
rect 17515 -35 17535 -15
rect 17565 -35 17585 -15
rect 17615 -35 17635 -15
rect 17665 -35 17685 -15
rect 17715 -35 17735 -15
rect 17765 -35 17785 -15
rect 17815 -35 17835 -15
rect 17865 -35 17885 -15
rect 17915 -35 17935 -15
rect 17965 -35 17985 -15
rect 18015 -35 18035 -15
rect 18065 -35 18085 -15
rect 18115 -35 18135 -15
rect 18165 -35 18185 -15
rect 18215 -35 18235 -15
rect 18265 -35 18285 -15
rect 18315 -35 18335 -15
rect 18365 -35 18385 -15
rect 18415 -35 18435 -15
rect 18465 -35 18485 -15
rect 18515 -35 18535 -15
rect 18565 -35 18585 -15
rect 18615 -35 18635 -15
rect 18665 -35 18685 -15
rect 18715 -35 18735 -15
rect 18765 -35 18785 -15
rect 18815 -35 18835 -15
rect 18865 -35 18885 -15
rect 18915 -35 18935 -15
rect 18965 -35 18985 -15
rect 19015 -35 19035 -15
rect 19065 -35 19085 -15
rect 19115 -35 19135 -15
rect 19165 -35 19185 -15
rect 19215 -35 19235 -15
rect 19265 -35 19285 -15
rect 19315 -35 19335 -15
rect 19365 -35 19385 -15
rect 19415 -35 19435 -15
rect 19465 -35 19485 -15
rect 19515 -35 19535 -15
rect 19565 -35 19585 -15
rect 19615 -35 19635 -15
rect 19665 -35 19685 -15
rect 19715 -35 19735 -15
rect 19765 -35 19785 -15
rect 19815 -35 19835 -15
rect 19865 -35 19885 -15
rect 19915 -35 19935 -15
rect 19965 -35 19985 -15
rect 20015 -35 20035 -15
rect 20065 -35 20085 -15
rect 20115 -35 20135 -15
rect 20165 -35 20185 -15
rect 20215 -35 20235 -15
rect 20265 -35 20285 -15
rect 20315 -35 20335 -15
rect 20365 -35 20385 -15
rect 20415 -35 20435 -15
rect 20465 -35 20485 -15
rect 20515 -35 20535 -15
rect 20565 -35 20585 -15
rect 20615 -35 20635 -15
rect 20665 -35 20685 -15
rect 20715 -35 20735 -15
rect 20765 -35 20785 -15
rect 20815 -35 20835 -15
rect 20865 -35 20885 -15
rect 20915 -35 20935 -15
rect 20965 -35 20985 -15
rect 21015 -35 21035 -15
rect 21065 -35 21085 -15
rect 21115 -35 21135 -15
rect 21165 -35 21185 -15
rect 21215 -35 21235 -15
rect 21265 -35 21285 -15
rect 21315 -35 21335 -15
rect 21365 -35 21385 -15
rect 21415 -35 21435 -15
rect 21465 -35 21485 -15
rect 21515 -35 21535 -15
rect 21565 -35 21585 -15
rect 21615 -35 21635 -15
rect 21665 -35 21685 -15
rect 21715 -35 21735 -15
rect 21765 -35 21785 -15
rect 21815 -35 21835 -15
rect 21865 -35 21885 -15
rect 21915 -35 21935 -15
rect 21965 -35 21985 -15
rect 22015 -35 22035 -15
rect 22065 -35 22085 -15
rect 22115 -35 22135 -15
rect 22165 -35 22185 -15
rect 22215 -35 22235 -15
rect 22265 -35 22285 -15
rect 22315 -35 22335 -15
rect 22365 -35 22385 -15
rect 22415 -35 22435 -15
rect 22465 -35 22485 -15
rect 22515 -35 22535 -15
rect 22565 -35 22585 -15
rect 22615 -35 22635 -15
rect 22665 -35 22685 -15
rect 22715 -35 22735 -15
rect 22765 -35 22785 -15
rect 22815 -35 22835 -15
rect 22865 -35 22885 -15
rect 22915 -35 22935 -15
rect 22965 -35 22985 -15
rect 23015 -35 23035 -15
rect 23065 -35 23085 -15
rect 23115 -35 23135 -15
rect 23165 -35 23185 -15
rect 23215 -35 23235 -15
rect 23265 -35 23285 -15
rect 23315 -35 23335 -15
rect 23365 -35 23385 -15
rect 23415 -35 23435 -15
rect 23465 -35 23485 -15
rect 23515 -35 23535 -15
rect 23565 -35 23585 -15
rect 23615 -35 23635 -15
rect 23665 -35 23685 -15
rect 23715 -35 23735 -15
rect 23765 -35 23785 -15
rect 23815 -35 23835 -15
rect 23865 -35 23885 -15
rect 23915 -35 23935 -15
rect 23965 -35 23985 -15
rect 24015 -35 24035 -15
rect 24065 -35 24085 -15
rect 24115 -35 24135 -15
rect 24165 -35 24185 -15
rect 24215 -35 24235 -15
rect 24265 -35 24285 -15
rect 24315 -35 24335 -15
rect 24365 -35 24385 -15
rect 24415 -35 24435 -15
rect 24465 -35 24485 -15
rect 24515 -35 24535 -15
rect 24565 -35 24585 -15
rect 24615 -35 24635 -15
rect 24665 -35 24685 -15
rect 24715 -35 24735 -15
rect 24765 -35 24785 -15
rect 24815 -35 24835 -15
rect 24865 -35 24885 -15
rect 24915 -35 24935 -15
rect 24965 -35 24985 -15
rect 25015 -35 25035 -15
rect 25065 -35 25085 -15
rect 25115 -35 25135 -15
rect 25165 -35 25185 -15
rect 25215 -35 25235 -15
rect 25265 -35 25285 -15
rect 25315 -35 25335 -15
rect 25365 -35 25385 -15
rect 25415 -35 25435 -15
rect 25465 -35 25485 -15
rect 25515 -35 25535 -15
rect 25565 -35 25585 -15
rect 25615 -35 25635 -15
rect 25665 -35 25685 -15
rect 25715 -35 25735 -15
rect 25765 -35 25785 -15
rect 25815 -35 25835 -15
rect 25865 -35 25885 -15
rect 25915 -35 25935 -15
rect 25965 -35 25985 -15
rect 26015 -35 26035 -15
rect 26065 -35 26085 -15
rect 26115 -35 26135 -15
rect 26165 -35 26185 -15
rect 26215 -35 26235 -15
rect 26265 -35 26285 -15
rect 26315 -35 26335 -15
rect 26365 -35 26385 -15
rect 26415 -35 26435 -15
rect 26465 -35 26485 -15
rect 26515 -35 26535 -15
rect 26565 -35 26585 -15
rect 26615 -35 26635 -15
rect 26665 -35 26685 -15
rect 26715 -35 26735 -15
rect 26765 -35 26785 -15
rect 26815 -35 26835 -15
rect 26865 -35 26885 -15
rect 26915 -35 26935 -15
rect 26965 -35 26985 -15
rect 27015 -35 27035 -15
rect 27065 -35 27085 -15
rect 27115 -35 27135 -15
rect 27165 -35 27185 -15
rect 27215 -35 27235 -15
rect 27265 -35 27285 -15
rect 27315 -35 27335 -15
rect 27365 -35 27385 -15
rect 27415 -35 27435 -15
rect 27465 -35 27485 -15
rect 27515 -35 27535 -15
rect 27565 -35 27585 -15
rect 27615 -35 27635 -15
rect 27665 -35 27685 -15
rect 27715 -35 27735 -15
rect 27765 -35 27785 -15
rect 27815 -35 27835 -15
rect 27865 -35 27885 -15
rect 27915 -35 27935 -15
rect 27965 -35 27985 -15
rect 28015 -35 28035 -15
rect 28065 -35 28085 -15
rect 28115 -35 28135 -15
rect 28165 -35 28185 -15
rect 28215 -35 28235 -15
rect 28265 -35 28285 -15
rect 28315 -35 28335 -15
rect 28365 -35 28385 -15
rect 28415 -35 28435 -15
rect 28465 -35 28485 -15
rect 28515 -35 28535 -15
rect 28565 -35 28585 -15
rect 28615 -35 28635 -15
rect 28665 -35 28685 -15
rect 28715 -35 28735 -15
rect 28765 -35 28785 -15
rect -635 -1735 -615 -1715
rect -585 -1735 -565 -1715
rect -535 -1735 -515 -1715
rect -485 -1735 -465 -1715
rect -435 -1735 -415 -1715
rect -385 -1735 -365 -1715
rect -335 -1735 -315 -1715
rect -285 -1735 -265 -1715
rect -235 -1735 -215 -1715
rect -185 -1735 -165 -1715
rect -135 -1735 -115 -1715
rect -85 -1735 -65 -1715
rect -35 -1735 -15 -1715
rect 15 -1735 35 -1715
rect 65 -1735 85 -1715
rect 115 -1735 135 -1715
rect 165 -1735 185 -1715
rect 215 -1735 235 -1715
rect 265 -1735 285 -1715
rect 315 -1735 335 -1715
rect 365 -1735 385 -1715
rect 415 -1735 435 -1715
rect 465 -1735 485 -1715
rect 515 -1735 535 -1715
rect 565 -1735 585 -1715
rect 615 -1735 635 -1715
rect 665 -1735 685 -1715
rect 715 -1735 735 -1715
rect 765 -1735 785 -1715
rect 815 -1735 835 -1715
rect 865 -1735 885 -1715
rect 915 -1735 935 -1715
rect 965 -1735 985 -1715
rect 1015 -1735 1035 -1715
rect 1065 -1735 1085 -1715
rect 1115 -1735 1135 -1715
rect 1165 -1735 1185 -1715
rect 1215 -1735 1235 -1715
rect 1265 -1735 1285 -1715
rect 1315 -1735 1335 -1715
rect 1365 -1735 1385 -1715
rect 1415 -1735 1435 -1715
rect 1465 -1735 1485 -1715
rect 1515 -1735 1535 -1715
rect 1565 -1735 1585 -1715
rect 1615 -1735 1635 -1715
rect 1665 -1735 1685 -1715
rect 1715 -1735 1735 -1715
rect 1765 -1735 1785 -1715
rect 1815 -1735 1835 -1715
rect 1865 -1735 1885 -1715
rect 1915 -1735 1935 -1715
rect 1965 -1735 1985 -1715
rect 2015 -1735 2035 -1715
rect 2065 -1735 2085 -1715
rect 2115 -1735 2135 -1715
rect 2165 -1735 2185 -1715
rect 2215 -1735 2235 -1715
rect 2265 -1735 2285 -1715
rect 2315 -1735 2335 -1715
rect 2365 -1735 2385 -1715
rect 2415 -1735 2435 -1715
rect 2465 -1735 2485 -1715
rect 2515 -1735 2535 -1715
rect 2565 -1735 2585 -1715
rect 2615 -1735 2635 -1715
rect 2665 -1735 2685 -1715
rect 2715 -1735 2735 -1715
rect 2765 -1735 2785 -1715
rect 2815 -1735 2835 -1715
rect 2865 -1735 2885 -1715
rect 2915 -1735 2935 -1715
rect 2965 -1735 2985 -1715
rect 3015 -1735 3035 -1715
rect 3065 -1735 3085 -1715
rect 3115 -1735 3135 -1715
rect 3165 -1735 3185 -1715
rect 3215 -1735 3235 -1715
rect 3265 -1735 3285 -1715
rect 3315 -1735 3335 -1715
rect 3365 -1735 3385 -1715
rect 3415 -1735 3435 -1715
rect 3465 -1735 3485 -1715
rect 3515 -1735 3535 -1715
rect 3565 -1735 3585 -1715
rect 3615 -1735 3635 -1715
rect 3665 -1735 3685 -1715
rect 3715 -1735 3735 -1715
rect 3765 -1735 3785 -1715
rect 3815 -1735 3835 -1715
rect 3865 -1735 3885 -1715
rect 3915 -1735 3935 -1715
rect 3965 -1735 3985 -1715
rect 4015 -1735 4035 -1715
rect 4065 -1735 4085 -1715
rect 4115 -1735 4135 -1715
rect 4165 -1735 4185 -1715
rect 4215 -1735 4235 -1715
rect 4265 -1735 4285 -1715
rect 4315 -1735 4335 -1715
rect 4365 -1735 4385 -1715
rect 4415 -1735 4435 -1715
rect 4465 -1735 4485 -1715
rect 4515 -1735 4535 -1715
rect 4565 -1735 4585 -1715
rect 4615 -1735 4635 -1715
rect 4665 -1735 4685 -1715
rect 4715 -1735 4735 -1715
rect 4765 -1735 4785 -1715
rect 4815 -1735 4835 -1715
rect 4865 -1735 4885 -1715
rect 4915 -1735 4935 -1715
rect 4965 -1735 4985 -1715
rect 5015 -1735 5035 -1715
rect 5065 -1735 5085 -1715
rect 5115 -1735 5135 -1715
rect 5165 -1735 5185 -1715
rect 5215 -1735 5235 -1715
rect 5265 -1735 5285 -1715
rect 5315 -1735 5335 -1715
rect 5365 -1735 5385 -1715
rect 5415 -1735 5435 -1715
rect 5465 -1735 5485 -1715
rect 5515 -1735 5535 -1715
rect 5565 -1735 5585 -1715
rect 5615 -1735 5635 -1715
rect 5665 -1735 5685 -1715
rect 5715 -1735 5735 -1715
rect 5765 -1735 5785 -1715
rect 5815 -1735 5835 -1715
rect 5865 -1735 5885 -1715
rect 5915 -1735 5935 -1715
rect 5965 -1735 5985 -1715
rect 6015 -1735 6035 -1715
rect 6065 -1735 6085 -1715
rect 6115 -1735 6135 -1715
rect 6165 -1735 6185 -1715
rect 6215 -1735 6235 -1715
rect 6265 -1735 6285 -1715
rect 6315 -1735 6335 -1715
rect 6365 -1735 6385 -1715
rect 6415 -1735 6435 -1715
rect 6465 -1735 6485 -1715
rect 6515 -1735 6535 -1715
rect 6565 -1735 6585 -1715
rect 6615 -1735 6635 -1715
rect 6665 -1735 6685 -1715
rect 6715 -1735 6735 -1715
rect 6765 -1735 6785 -1715
rect 6815 -1735 6835 -1715
rect 6865 -1735 6885 -1715
rect 6915 -1735 6935 -1715
rect 6965 -1735 6985 -1715
rect 7015 -1735 7035 -1715
rect 7065 -1735 7085 -1715
rect 7115 -1735 7135 -1715
rect 7165 -1735 7185 -1715
rect 7215 -1735 7235 -1715
rect 7265 -1735 7285 -1715
rect 7315 -1735 7335 -1715
rect 7365 -1735 7385 -1715
rect 7415 -1735 7435 -1715
rect 7465 -1735 7485 -1715
rect 7515 -1735 7535 -1715
rect 7565 -1735 7585 -1715
rect 7615 -1735 7635 -1715
rect 7665 -1735 7685 -1715
rect 7715 -1735 7735 -1715
rect 7765 -1735 7785 -1715
rect 7815 -1735 7835 -1715
rect 7865 -1735 7885 -1715
rect 7915 -1735 7935 -1715
rect 7965 -1735 7985 -1715
rect 8015 -1735 8035 -1715
rect 8065 -1735 8085 -1715
rect 8115 -1735 8135 -1715
rect 8165 -1735 8185 -1715
rect 8215 -1735 8235 -1715
rect 8265 -1735 8285 -1715
rect 8315 -1735 8335 -1715
rect 8365 -1735 8385 -1715
rect 8415 -1735 8435 -1715
rect 8465 -1735 8485 -1715
rect 8515 -1735 8535 -1715
rect 8565 -1735 8585 -1715
rect 8615 -1735 8635 -1715
rect 8665 -1735 8685 -1715
rect 8715 -1735 8735 -1715
rect 8765 -1735 8785 -1715
rect 8815 -1735 8835 -1715
rect 8865 -1735 8885 -1715
rect 8915 -1735 8935 -1715
rect 8965 -1735 8985 -1715
rect 9015 -1735 9035 -1715
rect 9065 -1735 9085 -1715
rect 9115 -1735 9135 -1715
rect 9165 -1735 9185 -1715
rect 9215 -1735 9235 -1715
rect 9265 -1735 9285 -1715
rect 9315 -1735 9335 -1715
rect 9365 -1735 9385 -1715
rect 9415 -1735 9435 -1715
rect 9465 -1735 9485 -1715
rect 9515 -1735 9535 -1715
rect 9565 -1735 9585 -1715
rect 9615 -1735 9635 -1715
rect 9665 -1735 9685 -1715
rect 9715 -1735 9735 -1715
rect 9765 -1735 9785 -1715
rect 9815 -1735 9835 -1715
rect 9865 -1735 9885 -1715
rect 9915 -1735 9935 -1715
rect 9965 -1735 9985 -1715
rect 10015 -1735 10035 -1715
rect 10065 -1735 10085 -1715
rect 10115 -1735 10135 -1715
rect 10165 -1735 10185 -1715
rect 10215 -1735 10235 -1715
rect 10265 -1735 10285 -1715
rect 10315 -1735 10335 -1715
rect 10365 -1735 10385 -1715
rect 10415 -1735 10435 -1715
rect 10465 -1735 10485 -1715
rect 10515 -1735 10535 -1715
rect 10565 -1735 10585 -1715
rect 10615 -1735 10635 -1715
rect 10665 -1735 10685 -1715
rect 10715 -1735 10735 -1715
rect 10765 -1735 10785 -1715
rect 10815 -1735 10835 -1715
rect 10865 -1735 10885 -1715
rect 10915 -1735 10935 -1715
rect 10965 -1735 10985 -1715
rect 11015 -1735 11035 -1715
rect 11065 -1735 11085 -1715
rect 11115 -1735 11135 -1715
rect 11165 -1735 11185 -1715
rect 11215 -1735 11235 -1715
rect 11265 -1735 11285 -1715
rect 11315 -1735 11335 -1715
rect 11365 -1735 11385 -1715
rect 11415 -1735 11435 -1715
rect 11465 -1735 11485 -1715
rect 11515 -1735 11535 -1715
rect 11565 -1735 11585 -1715
rect 11615 -1735 11635 -1715
rect 11665 -1735 11685 -1715
rect 11715 -1735 11735 -1715
rect 11765 -1735 11785 -1715
rect 11815 -1735 11835 -1715
rect 11865 -1735 11885 -1715
rect 11915 -1735 11935 -1715
rect 11965 -1735 11985 -1715
rect 12015 -1735 12035 -1715
rect 12065 -1735 12085 -1715
rect 12115 -1735 12135 -1715
rect 12165 -1735 12185 -1715
rect 12215 -1735 12235 -1715
rect 12265 -1735 12285 -1715
rect 12315 -1735 12335 -1715
rect 12365 -1735 12385 -1715
rect 12415 -1735 12435 -1715
rect 12465 -1735 12485 -1715
rect 12515 -1735 12535 -1715
rect 12565 -1735 12585 -1715
rect 12615 -1735 12635 -1715
rect 12665 -1735 12685 -1715
rect 12715 -1735 12735 -1715
rect 12765 -1735 12785 -1715
rect 12815 -1735 12835 -1715
rect 12865 -1735 12885 -1715
rect 12915 -1735 12935 -1715
rect 12965 -1735 12985 -1715
rect 13015 -1735 13035 -1715
rect 13065 -1735 13085 -1715
rect 13115 -1735 13135 -1715
rect 13165 -1735 13185 -1715
rect 13215 -1735 13235 -1715
rect 13265 -1735 13285 -1715
rect 13315 -1735 13335 -1715
rect 13365 -1735 13385 -1715
rect 13415 -1735 13435 -1715
rect 13465 -1735 13485 -1715
rect 13515 -1735 13535 -1715
rect 13565 -1735 13585 -1715
rect 13615 -1735 13635 -1715
rect 13665 -1735 13685 -1715
rect 13715 -1735 13735 -1715
rect 13765 -1735 13785 -1715
rect 13815 -1735 13835 -1715
rect 13865 -1735 13885 -1715
rect 13915 -1735 13935 -1715
rect 13965 -1735 13985 -1715
rect 14015 -1735 14035 -1715
rect 14065 -1735 14085 -1715
rect 14115 -1735 14135 -1715
rect 14165 -1735 14185 -1715
rect 14215 -1735 14235 -1715
rect 14265 -1735 14285 -1715
rect 14315 -1735 14335 -1715
rect 14365 -1735 14385 -1715
rect 14415 -1735 14435 -1715
rect 14465 -1735 14485 -1715
rect 14515 -1735 14535 -1715
rect 14565 -1735 14585 -1715
rect 14615 -1735 14635 -1715
rect 14665 -1735 14685 -1715
rect 14715 -1735 14735 -1715
rect 14765 -1735 14785 -1715
rect 14815 -1735 14835 -1715
rect 14865 -1735 14885 -1715
rect 14915 -1735 14935 -1715
rect 14965 -1735 14985 -1715
rect 15015 -1735 15035 -1715
rect 15065 -1735 15085 -1715
rect 15115 -1735 15135 -1715
rect 15165 -1735 15185 -1715
rect 15215 -1735 15235 -1715
rect 15265 -1735 15285 -1715
rect 15315 -1735 15335 -1715
rect 15365 -1735 15385 -1715
rect 15415 -1735 15435 -1715
rect 15465 -1735 15485 -1715
rect 15515 -1735 15535 -1715
rect 15565 -1735 15585 -1715
rect 15615 -1735 15635 -1715
rect 15665 -1735 15685 -1715
rect 15715 -1735 15735 -1715
rect 15765 -1735 15785 -1715
rect 15815 -1735 15835 -1715
rect 15865 -1735 15885 -1715
rect 15915 -1735 15935 -1715
rect 15965 -1735 15985 -1715
rect 16015 -1735 16035 -1715
rect 16065 -1735 16085 -1715
rect 16115 -1735 16135 -1715
rect 16165 -1735 16185 -1715
rect 16215 -1735 16235 -1715
rect 16265 -1735 16285 -1715
rect 16315 -1735 16335 -1715
rect 16365 -1735 16385 -1715
rect 16415 -1735 16435 -1715
rect 16465 -1735 16485 -1715
rect 16515 -1735 16535 -1715
rect 16565 -1735 16585 -1715
rect 16615 -1735 16635 -1715
rect 16665 -1735 16685 -1715
rect 16715 -1735 16735 -1715
rect 16765 -1735 16785 -1715
rect 16815 -1735 16835 -1715
rect 16865 -1735 16885 -1715
rect 16915 -1735 16935 -1715
rect 16965 -1735 16985 -1715
rect 17015 -1735 17035 -1715
rect 17065 -1735 17085 -1715
rect 17115 -1735 17135 -1715
rect 17165 -1735 17185 -1715
rect 17215 -1735 17235 -1715
rect 17265 -1735 17285 -1715
rect 17315 -1735 17335 -1715
rect 17365 -1735 17385 -1715
rect 17415 -1735 17435 -1715
rect 17465 -1735 17485 -1715
rect 17515 -1735 17535 -1715
rect 17565 -1735 17585 -1715
rect 17615 -1735 17635 -1715
rect 17665 -1735 17685 -1715
rect 17715 -1735 17735 -1715
rect 17765 -1735 17785 -1715
rect 17815 -1735 17835 -1715
rect 17865 -1735 17885 -1715
rect 17915 -1735 17935 -1715
rect 17965 -1735 17985 -1715
rect 18015 -1735 18035 -1715
rect 18065 -1735 18085 -1715
rect 18115 -1735 18135 -1715
rect 18165 -1735 18185 -1715
rect 18215 -1735 18235 -1715
rect 18265 -1735 18285 -1715
rect 18315 -1735 18335 -1715
rect 18365 -1735 18385 -1715
rect 18415 -1735 18435 -1715
rect 18465 -1735 18485 -1715
rect 18515 -1735 18535 -1715
rect 18565 -1735 18585 -1715
rect 18615 -1735 18635 -1715
rect 18665 -1735 18685 -1715
rect 18715 -1735 18735 -1715
rect 18765 -1735 18785 -1715
rect 18815 -1735 18835 -1715
rect 18865 -1735 18885 -1715
rect 18915 -1735 18935 -1715
rect 18965 -1735 18985 -1715
rect 19015 -1735 19035 -1715
rect 19065 -1735 19085 -1715
rect 19115 -1735 19135 -1715
rect 19165 -1735 19185 -1715
rect 19215 -1735 19235 -1715
rect 19265 -1735 19285 -1715
rect 19315 -1735 19335 -1715
rect 19365 -1735 19385 -1715
rect 19415 -1735 19435 -1715
rect 19465 -1735 19485 -1715
rect 19515 -1735 19535 -1715
rect 19565 -1735 19585 -1715
rect 19615 -1735 19635 -1715
rect 19665 -1735 19685 -1715
rect 19715 -1735 19735 -1715
rect 19765 -1735 19785 -1715
rect 19815 -1735 19835 -1715
rect 19865 -1735 19885 -1715
rect 19915 -1735 19935 -1715
rect 19965 -1735 19985 -1715
rect 20015 -1735 20035 -1715
rect 20065 -1735 20085 -1715
rect 20115 -1735 20135 -1715
rect 20165 -1735 20185 -1715
rect 20215 -1735 20235 -1715
rect 20265 -1735 20285 -1715
rect 20315 -1735 20335 -1715
rect 20365 -1735 20385 -1715
rect 20415 -1735 20435 -1715
rect 20465 -1735 20485 -1715
rect 20515 -1735 20535 -1715
rect 20565 -1735 20585 -1715
rect 20615 -1735 20635 -1715
rect 20665 -1735 20685 -1715
rect 20715 -1735 20735 -1715
rect 20765 -1735 20785 -1715
rect 20815 -1735 20835 -1715
rect 20865 -1735 20885 -1715
rect 20915 -1735 20935 -1715
rect 20965 -1735 20985 -1715
rect 21015 -1735 21035 -1715
rect 21065 -1735 21085 -1715
rect 21115 -1735 21135 -1715
rect 21165 -1735 21185 -1715
rect 21215 -1735 21235 -1715
rect 21265 -1735 21285 -1715
rect 21315 -1735 21335 -1715
rect 21365 -1735 21385 -1715
rect 21415 -1735 21435 -1715
rect 21465 -1735 21485 -1715
rect 21515 -1735 21535 -1715
rect 21565 -1735 21585 -1715
rect 21615 -1735 21635 -1715
rect 21665 -1735 21685 -1715
rect 21715 -1735 21735 -1715
rect 21765 -1735 21785 -1715
rect 21815 -1735 21835 -1715
rect 21865 -1735 21885 -1715
rect 21915 -1735 21935 -1715
rect 21965 -1735 21985 -1715
rect 22015 -1735 22035 -1715
rect 22065 -1735 22085 -1715
rect 22115 -1735 22135 -1715
rect 22165 -1735 22185 -1715
rect 22215 -1735 22235 -1715
rect 22265 -1735 22285 -1715
rect 22315 -1735 22335 -1715
rect 22365 -1735 22385 -1715
rect 22415 -1735 22435 -1715
rect 22465 -1735 22485 -1715
rect 22515 -1735 22535 -1715
rect 22565 -1735 22585 -1715
rect 22615 -1735 22635 -1715
rect 22665 -1735 22685 -1715
rect 22715 -1735 22735 -1715
rect 22765 -1735 22785 -1715
rect 22815 -1735 22835 -1715
rect 22865 -1735 22885 -1715
rect 22915 -1735 22935 -1715
rect 22965 -1735 22985 -1715
rect 23015 -1735 23035 -1715
rect 23065 -1735 23085 -1715
rect 23115 -1735 23135 -1715
rect 23165 -1735 23185 -1715
rect 23215 -1735 23235 -1715
rect 23265 -1735 23285 -1715
rect 23315 -1735 23335 -1715
rect 23365 -1735 23385 -1715
rect 23415 -1735 23435 -1715
rect 23465 -1735 23485 -1715
rect 23515 -1735 23535 -1715
rect 23565 -1735 23585 -1715
rect 23615 -1735 23635 -1715
rect 23665 -1735 23685 -1715
rect 23715 -1735 23735 -1715
rect 23765 -1735 23785 -1715
rect 23815 -1735 23835 -1715
rect 23865 -1735 23885 -1715
rect 23915 -1735 23935 -1715
rect 23965 -1735 23985 -1715
rect 24015 -1735 24035 -1715
rect 24065 -1735 24085 -1715
rect 24115 -1735 24135 -1715
rect 24165 -1735 24185 -1715
rect 24215 -1735 24235 -1715
rect 24265 -1735 24285 -1715
rect 24315 -1735 24335 -1715
rect 24365 -1735 24385 -1715
rect 24415 -1735 24435 -1715
rect 24465 -1735 24485 -1715
rect 24515 -1735 24535 -1715
rect 24565 -1735 24585 -1715
rect 24615 -1735 24635 -1715
rect 24665 -1735 24685 -1715
rect 24715 -1735 24735 -1715
rect 24765 -1735 24785 -1715
rect 24815 -1735 24835 -1715
rect 24865 -1735 24885 -1715
rect 24915 -1735 24935 -1715
rect 24965 -1735 24985 -1715
rect 25015 -1735 25035 -1715
rect 25065 -1735 25085 -1715
rect 25115 -1735 25135 -1715
rect 25165 -1735 25185 -1715
rect 25215 -1735 25235 -1715
rect 25265 -1735 25285 -1715
rect 25315 -1735 25335 -1715
rect 25365 -1735 25385 -1715
rect 25415 -1735 25435 -1715
rect 25465 -1735 25485 -1715
rect 25515 -1735 25535 -1715
rect 25565 -1735 25585 -1715
rect 25615 -1735 25635 -1715
rect 25665 -1735 25685 -1715
rect 25715 -1735 25735 -1715
rect 25765 -1735 25785 -1715
rect 25815 -1735 25835 -1715
rect 25865 -1735 25885 -1715
rect 25915 -1735 25935 -1715
rect 25965 -1735 25985 -1715
rect 26015 -1735 26035 -1715
rect 26065 -1735 26085 -1715
rect 26115 -1735 26135 -1715
rect 26165 -1735 26185 -1715
rect 26215 -1735 26235 -1715
rect 26265 -1735 26285 -1715
rect 26315 -1735 26335 -1715
rect 26365 -1735 26385 -1715
rect 26415 -1735 26435 -1715
rect 26465 -1735 26485 -1715
rect 26515 -1735 26535 -1715
rect 26565 -1735 26585 -1715
rect 26615 -1735 26635 -1715
rect 26665 -1735 26685 -1715
rect 26715 -1735 26735 -1715
rect 26765 -1735 26785 -1715
rect 26815 -1735 26835 -1715
rect 26865 -1735 26885 -1715
rect 26915 -1735 26935 -1715
rect 26965 -1735 26985 -1715
rect 27015 -1735 27035 -1715
rect 27065 -1735 27085 -1715
rect 27115 -1735 27135 -1715
rect 27165 -1735 27185 -1715
rect 27215 -1735 27235 -1715
rect 27265 -1735 27285 -1715
rect 27315 -1735 27335 -1715
rect 27365 -1735 27385 -1715
rect 27415 -1735 27435 -1715
rect 27465 -1735 27485 -1715
rect 27515 -1735 27535 -1715
rect 27565 -1735 27585 -1715
rect 27615 -1735 27635 -1715
rect 27665 -1735 27685 -1715
rect 27715 -1735 27735 -1715
rect 27765 -1735 27785 -1715
rect 27815 -1735 27835 -1715
rect 27865 -1735 27885 -1715
rect 27915 -1735 27935 -1715
rect 27965 -1735 27985 -1715
rect 28015 -1735 28035 -1715
rect 28065 -1735 28085 -1715
rect 28115 -1735 28135 -1715
rect 28165 -1735 28185 -1715
rect 28215 -1735 28235 -1715
rect 28265 -1735 28285 -1715
rect 28315 -1735 28335 -1715
rect 28365 -1735 28385 -1715
rect 28415 -1735 28435 -1715
rect 28465 -1735 28485 -1715
rect 28515 -1735 28535 -1715
rect 28565 -1735 28585 -1715
rect 28615 -1735 28635 -1715
rect 28665 -1735 28685 -1715
rect 28715 -1735 28735 -1715
rect 28765 -1735 28785 -1715
<< mvnsubdiffcont >>
rect -635 5565 -615 5585
rect -585 5565 -565 5585
rect -535 5565 -515 5585
rect -485 5565 -465 5585
rect -435 5565 -415 5585
rect -385 5565 -365 5585
rect -335 5565 -315 5585
rect -285 5565 -265 5585
rect -235 5565 -215 5585
rect -185 5565 -165 5585
rect -135 5565 -115 5585
rect -85 5565 -65 5585
rect -35 5565 -15 5585
rect 15 5565 35 5585
rect 65 5565 85 5585
rect 115 5565 135 5585
rect 165 5565 185 5585
rect 215 5565 235 5585
rect 265 5565 285 5585
rect 315 5565 335 5585
rect 365 5565 385 5585
rect 415 5565 435 5585
rect 465 5565 485 5585
rect 515 5565 535 5585
rect 565 5565 585 5585
rect 615 5565 635 5585
rect 665 5565 685 5585
rect 715 5565 735 5585
rect 765 5565 785 5585
rect 815 5565 835 5585
rect 865 5565 885 5585
rect 915 5565 935 5585
rect 965 5565 985 5585
rect 1015 5565 1035 5585
rect 1065 5565 1085 5585
rect 1115 5565 1135 5585
rect 1165 5565 1185 5585
rect 1215 5565 1235 5585
rect 1265 5565 1285 5585
rect 1315 5565 1335 5585
rect 1365 5565 1385 5585
rect 1415 5565 1435 5585
rect 1465 5565 1485 5585
rect 1515 5565 1535 5585
rect 1565 5565 1585 5585
rect 1615 5565 1635 5585
rect 1665 5565 1685 5585
rect 1715 5565 1735 5585
rect 1765 5565 1785 5585
rect 1815 5565 1835 5585
rect 1865 5565 1885 5585
rect 1915 5565 1935 5585
rect 1965 5565 1985 5585
rect 2015 5565 2035 5585
rect 2065 5565 2085 5585
rect 2115 5565 2135 5585
rect 2165 5565 2185 5585
rect 2215 5565 2235 5585
rect 2265 5565 2285 5585
rect 2315 5565 2335 5585
rect 2365 5565 2385 5585
rect 2415 5565 2435 5585
rect 2465 5565 2485 5585
rect 2515 5565 2535 5585
rect 2565 5565 2585 5585
rect 2615 5565 2635 5585
rect 2665 5565 2685 5585
rect 2715 5565 2735 5585
rect 2765 5565 2785 5585
rect 2815 5565 2835 5585
rect 2865 5565 2885 5585
rect 2915 5565 2935 5585
rect 2965 5565 2985 5585
rect 3015 5565 3035 5585
rect 3065 5565 3085 5585
rect 3115 5565 3135 5585
rect 3165 5565 3185 5585
rect 3215 5565 3235 5585
rect 3265 5565 3285 5585
rect 3315 5565 3335 5585
rect 3365 5565 3385 5585
rect 3415 5565 3435 5585
rect 3465 5565 3485 5585
rect 3515 5565 3535 5585
rect 3565 5565 3585 5585
rect 3615 5565 3635 5585
rect 3665 5565 3685 5585
rect 3715 5565 3735 5585
rect 3765 5565 3785 5585
rect 3815 5565 3835 5585
rect 3865 5565 3885 5585
rect 3915 5565 3935 5585
rect 3965 5565 3985 5585
rect 4015 5565 4035 5585
rect 4065 5565 4085 5585
rect 4115 5565 4135 5585
rect 4165 5565 4185 5585
rect 4215 5565 4235 5585
rect 4265 5565 4285 5585
rect 4315 5565 4335 5585
rect 4365 5565 4385 5585
rect 4415 5565 4435 5585
rect 4465 5565 4485 5585
rect 4515 5565 4535 5585
rect 4565 5565 4585 5585
rect 4615 5565 4635 5585
rect 4665 5565 4685 5585
rect 4715 5565 4735 5585
rect 4765 5565 4785 5585
rect 4815 5565 4835 5585
rect 4865 5565 4885 5585
rect 4915 5565 4935 5585
rect 4965 5565 4985 5585
rect 5015 5565 5035 5585
rect 5065 5565 5085 5585
rect 5115 5565 5135 5585
rect 5165 5565 5185 5585
rect 5215 5565 5235 5585
rect 5265 5565 5285 5585
rect 5315 5565 5335 5585
rect 5365 5565 5385 5585
rect 5415 5565 5435 5585
rect 5465 5565 5485 5585
rect 5515 5565 5535 5585
rect 5565 5565 5585 5585
rect 5615 5565 5635 5585
rect 5665 5565 5685 5585
rect 5715 5565 5735 5585
rect 5765 5565 5785 5585
rect 5815 5565 5835 5585
rect 5865 5565 5885 5585
rect 5915 5565 5935 5585
rect 5965 5565 5985 5585
rect 6015 5565 6035 5585
rect 6065 5565 6085 5585
rect 6115 5565 6135 5585
rect 6165 5565 6185 5585
rect 6215 5565 6235 5585
rect 6265 5565 6285 5585
rect 6315 5565 6335 5585
rect 6365 5565 6385 5585
rect 6415 5565 6435 5585
rect 6465 5565 6485 5585
rect 6515 5565 6535 5585
rect 6565 5565 6585 5585
rect 6615 5565 6635 5585
rect 6665 5565 6685 5585
rect 6715 5565 6735 5585
rect 6765 5565 6785 5585
rect 6815 5565 6835 5585
rect 6865 5565 6885 5585
rect 6915 5565 6935 5585
rect 6965 5565 6985 5585
rect 7015 5565 7035 5585
rect 7065 5565 7085 5585
rect 7115 5565 7135 5585
rect 7165 5565 7185 5585
rect 7215 5565 7235 5585
rect 7265 5565 7285 5585
rect 7315 5565 7335 5585
rect 7365 5565 7385 5585
rect 7415 5565 7435 5585
rect 7465 5565 7485 5585
rect 7515 5565 7535 5585
rect 7565 5565 7585 5585
rect 7615 5565 7635 5585
rect 7665 5565 7685 5585
rect 7715 5565 7735 5585
rect 7765 5565 7785 5585
rect 7815 5565 7835 5585
rect 7865 5565 7885 5585
rect 7915 5565 7935 5585
rect 7965 5565 7985 5585
rect 8015 5565 8035 5585
rect 8065 5565 8085 5585
rect 8115 5565 8135 5585
rect 8165 5565 8185 5585
rect 8215 5565 8235 5585
rect 8265 5565 8285 5585
rect 8315 5565 8335 5585
rect 8365 5565 8385 5585
rect 8415 5565 8435 5585
rect 8465 5565 8485 5585
rect 8515 5565 8535 5585
rect 8565 5565 8585 5585
rect 8615 5565 8635 5585
rect 8665 5565 8685 5585
rect 8715 5565 8735 5585
rect 8765 5565 8785 5585
rect 8815 5565 8835 5585
rect 8865 5565 8885 5585
rect 8915 5565 8935 5585
rect 8965 5565 8985 5585
rect 9015 5565 9035 5585
rect 9065 5565 9085 5585
rect 9115 5565 9135 5585
rect 9165 5565 9185 5585
rect 9215 5565 9235 5585
rect 9265 5565 9285 5585
rect 9315 5565 9335 5585
rect 9365 5565 9385 5585
rect 9415 5565 9435 5585
rect 9465 5565 9485 5585
rect 9515 5565 9535 5585
rect 9565 5565 9585 5585
rect 9615 5565 9635 5585
rect 9665 5565 9685 5585
rect 9715 5565 9735 5585
rect 9765 5565 9785 5585
rect 9815 5565 9835 5585
rect 9865 5565 9885 5585
rect 9915 5565 9935 5585
rect 9965 5565 9985 5585
rect 10015 5565 10035 5585
rect 10065 5565 10085 5585
rect 10115 5565 10135 5585
rect 10165 5565 10185 5585
rect 10215 5565 10235 5585
rect 10265 5565 10285 5585
rect 10315 5565 10335 5585
rect 10365 5565 10385 5585
rect 10415 5565 10435 5585
rect 10465 5565 10485 5585
rect 10515 5565 10535 5585
rect 10565 5565 10585 5585
rect 10615 5565 10635 5585
rect 10665 5565 10685 5585
rect 10715 5565 10735 5585
rect 10765 5565 10785 5585
rect 10815 5565 10835 5585
rect 10865 5565 10885 5585
rect 10915 5565 10935 5585
rect 10965 5565 10985 5585
rect 11015 5565 11035 5585
rect 11065 5565 11085 5585
rect 11115 5565 11135 5585
rect 11165 5565 11185 5585
rect 11215 5565 11235 5585
rect 11265 5565 11285 5585
rect 11315 5565 11335 5585
rect 11365 5565 11385 5585
rect 11415 5565 11435 5585
rect 11465 5565 11485 5585
rect 11515 5565 11535 5585
rect 11565 5565 11585 5585
rect 11615 5565 11635 5585
rect 11665 5565 11685 5585
rect 11715 5565 11735 5585
rect 11765 5565 11785 5585
rect 11815 5565 11835 5585
rect 11865 5565 11885 5585
rect 11915 5565 11935 5585
rect 11965 5565 11985 5585
rect 12015 5565 12035 5585
rect 12065 5565 12085 5585
rect 12115 5565 12135 5585
rect 12165 5565 12185 5585
rect 12215 5565 12235 5585
rect 12265 5565 12285 5585
rect 12315 5565 12335 5585
rect 12365 5565 12385 5585
rect 12415 5565 12435 5585
rect 12465 5565 12485 5585
rect 12515 5565 12535 5585
rect 12565 5565 12585 5585
rect 12615 5565 12635 5585
rect 12665 5565 12685 5585
rect 12715 5565 12735 5585
rect 12765 5565 12785 5585
rect 12815 5565 12835 5585
rect 12865 5565 12885 5585
rect 12915 5565 12935 5585
rect 12965 5565 12985 5585
rect 13015 5565 13035 5585
rect 13065 5565 13085 5585
rect 13115 5565 13135 5585
rect 13165 5565 13185 5585
rect 13215 5565 13235 5585
rect 13265 5565 13285 5585
rect 13315 5565 13335 5585
rect 13365 5565 13385 5585
rect 13415 5565 13435 5585
rect 13465 5565 13485 5585
rect 13515 5565 13535 5585
rect 13565 5565 13585 5585
rect 13615 5565 13635 5585
rect 13665 5565 13685 5585
rect 13715 5565 13735 5585
rect 13765 5565 13785 5585
rect 13815 5565 13835 5585
rect 13865 5565 13885 5585
rect 13915 5565 13935 5585
rect 13965 5565 13985 5585
rect 14015 5565 14035 5585
rect 14065 5565 14085 5585
rect 14115 5565 14135 5585
rect 14165 5565 14185 5585
rect 14215 5565 14235 5585
rect 14265 5565 14285 5585
rect 14315 5565 14335 5585
rect 14365 5565 14385 5585
rect 14415 5565 14435 5585
rect 14465 5565 14485 5585
rect 14515 5565 14535 5585
rect 14565 5565 14585 5585
rect 14615 5565 14635 5585
rect 14665 5565 14685 5585
rect 14715 5565 14735 5585
rect 14765 5565 14785 5585
rect 14815 5565 14835 5585
rect 14865 5565 14885 5585
rect 14915 5565 14935 5585
rect 14965 5565 14985 5585
rect 15015 5565 15035 5585
rect 15065 5565 15085 5585
rect 15115 5565 15135 5585
rect 15165 5565 15185 5585
rect 15215 5565 15235 5585
rect 15265 5565 15285 5585
rect 15315 5565 15335 5585
rect 15365 5565 15385 5585
rect 15415 5565 15435 5585
rect 15465 5565 15485 5585
rect 15515 5565 15535 5585
rect 15565 5565 15585 5585
rect 15615 5565 15635 5585
rect 15665 5565 15685 5585
rect 15715 5565 15735 5585
rect 15765 5565 15785 5585
rect 15815 5565 15835 5585
rect 15865 5565 15885 5585
rect 15915 5565 15935 5585
rect 15965 5565 15985 5585
rect 16015 5565 16035 5585
rect 16065 5565 16085 5585
rect 16115 5565 16135 5585
rect 16165 5565 16185 5585
rect 16215 5565 16235 5585
rect 16265 5565 16285 5585
rect 16315 5565 16335 5585
rect 16365 5565 16385 5585
rect 16415 5565 16435 5585
rect 16465 5565 16485 5585
rect 16515 5565 16535 5585
rect 16565 5565 16585 5585
rect 16615 5565 16635 5585
rect 16665 5565 16685 5585
rect 16715 5565 16735 5585
rect 16765 5565 16785 5585
rect 16815 5565 16835 5585
rect 16865 5565 16885 5585
rect 16915 5565 16935 5585
rect 16965 5565 16985 5585
rect 17015 5565 17035 5585
rect 17065 5565 17085 5585
rect 17115 5565 17135 5585
rect 17165 5565 17185 5585
rect 17215 5565 17235 5585
rect 17265 5565 17285 5585
rect 17315 5565 17335 5585
rect 17365 5565 17385 5585
rect 17415 5565 17435 5585
rect 17465 5565 17485 5585
rect 17515 5565 17535 5585
rect 17565 5565 17585 5585
rect 17615 5565 17635 5585
rect 17665 5565 17685 5585
rect 17715 5565 17735 5585
rect 17765 5565 17785 5585
rect 17815 5565 17835 5585
rect 17865 5565 17885 5585
rect 17915 5565 17935 5585
rect 17965 5565 17985 5585
rect 18015 5565 18035 5585
rect 18065 5565 18085 5585
rect 18115 5565 18135 5585
rect 18165 5565 18185 5585
rect 18215 5565 18235 5585
rect 18265 5565 18285 5585
rect 18315 5565 18335 5585
rect 18365 5565 18385 5585
rect 18415 5565 18435 5585
rect 18465 5565 18485 5585
rect 18515 5565 18535 5585
rect 18565 5565 18585 5585
rect 18615 5565 18635 5585
rect 18665 5565 18685 5585
rect 18715 5565 18735 5585
rect 18765 5565 18785 5585
rect 18815 5565 18835 5585
rect 18865 5565 18885 5585
rect 18915 5565 18935 5585
rect 18965 5565 18985 5585
rect 19015 5565 19035 5585
rect 19065 5565 19085 5585
rect 19115 5565 19135 5585
rect 19165 5565 19185 5585
rect 19215 5565 19235 5585
rect 19265 5565 19285 5585
rect 19315 5565 19335 5585
rect 19365 5565 19385 5585
rect 19415 5565 19435 5585
rect 19465 5565 19485 5585
rect 19515 5565 19535 5585
rect 19565 5565 19585 5585
rect 19615 5565 19635 5585
rect 19665 5565 19685 5585
rect 19715 5565 19735 5585
rect 19765 5565 19785 5585
rect 19815 5565 19835 5585
rect 19865 5565 19885 5585
rect 19915 5565 19935 5585
rect 19965 5565 19985 5585
rect 20015 5565 20035 5585
rect 20065 5565 20085 5585
rect 20115 5565 20135 5585
rect 20165 5565 20185 5585
rect 20215 5565 20235 5585
rect 20265 5565 20285 5585
rect 20315 5565 20335 5585
rect 20365 5565 20385 5585
rect 20415 5565 20435 5585
rect 20465 5565 20485 5585
rect 20515 5565 20535 5585
rect 20565 5565 20585 5585
rect 20615 5565 20635 5585
rect 20665 5565 20685 5585
rect 20715 5565 20735 5585
rect 20765 5565 20785 5585
rect 20815 5565 20835 5585
rect 20865 5565 20885 5585
rect 20915 5565 20935 5585
rect 20965 5565 20985 5585
rect 21015 5565 21035 5585
rect 21065 5565 21085 5585
rect 21115 5565 21135 5585
rect 21165 5565 21185 5585
rect 21215 5565 21235 5585
rect 21265 5565 21285 5585
rect 21315 5565 21335 5585
rect 21365 5565 21385 5585
rect 21415 5565 21435 5585
rect 21465 5565 21485 5585
rect 21515 5565 21535 5585
rect 21565 5565 21585 5585
rect 21615 5565 21635 5585
rect 21665 5565 21685 5585
rect 21715 5565 21735 5585
rect 21765 5565 21785 5585
rect 21815 5565 21835 5585
rect 21865 5565 21885 5585
rect 21915 5565 21935 5585
rect 21965 5565 21985 5585
rect 22015 5565 22035 5585
rect 22065 5565 22085 5585
rect 22115 5565 22135 5585
rect 22165 5565 22185 5585
rect 22215 5565 22235 5585
rect 22265 5565 22285 5585
rect 22315 5565 22335 5585
rect 22365 5565 22385 5585
rect 22415 5565 22435 5585
rect 22465 5565 22485 5585
rect 22515 5565 22535 5585
rect 22565 5565 22585 5585
rect 22615 5565 22635 5585
rect 22665 5565 22685 5585
rect 22715 5565 22735 5585
rect 22765 5565 22785 5585
rect 22815 5565 22835 5585
rect 22865 5565 22885 5585
rect 22915 5565 22935 5585
rect 22965 5565 22985 5585
rect 23015 5565 23035 5585
rect 23065 5565 23085 5585
rect 23115 5565 23135 5585
rect 23165 5565 23185 5585
rect 23215 5565 23235 5585
rect 23265 5565 23285 5585
rect 23315 5565 23335 5585
rect 23365 5565 23385 5585
rect 23415 5565 23435 5585
rect 23465 5565 23485 5585
rect 23515 5565 23535 5585
rect 23565 5565 23585 5585
rect 23615 5565 23635 5585
rect 23665 5565 23685 5585
rect 23715 5565 23735 5585
rect 23765 5565 23785 5585
rect 23815 5565 23835 5585
rect 23865 5565 23885 5585
rect 23915 5565 23935 5585
rect 23965 5565 23985 5585
rect 24015 5565 24035 5585
rect 24065 5565 24085 5585
rect 24115 5565 24135 5585
rect 24165 5565 24185 5585
rect 24215 5565 24235 5585
rect 24265 5565 24285 5585
rect 24315 5565 24335 5585
rect 24365 5565 24385 5585
rect 24415 5565 24435 5585
rect 24465 5565 24485 5585
rect 24515 5565 24535 5585
rect 24565 5565 24585 5585
rect 24615 5565 24635 5585
rect 24665 5565 24685 5585
rect 24715 5565 24735 5585
rect 24765 5565 24785 5585
rect 24815 5565 24835 5585
rect 24865 5565 24885 5585
rect 24915 5565 24935 5585
rect 24965 5565 24985 5585
rect 25015 5565 25035 5585
rect 25065 5565 25085 5585
rect 25115 5565 25135 5585
rect 25165 5565 25185 5585
rect 25215 5565 25235 5585
rect 25265 5565 25285 5585
rect 25315 5565 25335 5585
rect 25365 5565 25385 5585
rect 25415 5565 25435 5585
rect 25465 5565 25485 5585
rect 25515 5565 25535 5585
rect 25565 5565 25585 5585
rect 25615 5565 25635 5585
rect 25665 5565 25685 5585
rect 25715 5565 25735 5585
rect 25765 5565 25785 5585
rect 25815 5565 25835 5585
rect 25865 5565 25885 5585
rect 25915 5565 25935 5585
rect 25965 5565 25985 5585
rect 26015 5565 26035 5585
rect 26065 5565 26085 5585
rect 26115 5565 26135 5585
rect 26165 5565 26185 5585
rect 26215 5565 26235 5585
rect 26265 5565 26285 5585
rect 26315 5565 26335 5585
rect 26365 5565 26385 5585
rect 26415 5565 26435 5585
rect 26465 5565 26485 5585
rect 26515 5565 26535 5585
rect 26565 5565 26585 5585
rect 26615 5565 26635 5585
rect 26665 5565 26685 5585
rect 26715 5565 26735 5585
rect 26765 5565 26785 5585
rect 26815 5565 26835 5585
rect 26865 5565 26885 5585
rect 26915 5565 26935 5585
rect 26965 5565 26985 5585
rect 27015 5565 27035 5585
rect 27065 5565 27085 5585
rect 27115 5565 27135 5585
rect 27165 5565 27185 5585
rect 27215 5565 27235 5585
rect 27265 5565 27285 5585
rect 27315 5565 27335 5585
rect 27365 5565 27385 5585
rect 27415 5565 27435 5585
rect 27465 5565 27485 5585
rect 27515 5565 27535 5585
rect 27565 5565 27585 5585
rect 27615 5565 27635 5585
rect 27665 5565 27685 5585
rect 27715 5565 27735 5585
rect 27765 5565 27785 5585
rect 27815 5565 27835 5585
rect 27865 5565 27885 5585
rect 27915 5565 27935 5585
rect 27965 5565 27985 5585
rect 28015 5565 28035 5585
rect 28065 5565 28085 5585
rect 28115 5565 28135 5585
rect 28165 5565 28185 5585
rect 28215 5565 28235 5585
rect 28265 5565 28285 5585
rect 28315 5565 28335 5585
rect 28365 5565 28385 5585
rect 28415 5565 28435 5585
rect 28465 5565 28485 5585
rect 28515 5565 28535 5585
rect 28565 5565 28585 5585
rect 28615 5565 28635 5585
rect 28665 5565 28685 5585
rect 28715 5565 28735 5585
rect 28765 5565 28785 5585
rect 28815 5565 28835 5585
rect 28865 5565 28885 5585
rect 28915 5565 28935 5585
rect 28965 5565 28985 5585
rect 29015 5565 29035 5585
rect 29065 5565 29085 5585
rect 29115 5565 29135 5585
rect 29165 5565 29185 5585
rect 29215 5565 29235 5585
rect 29265 5565 29285 5585
rect 29315 5565 29335 5585
rect 29365 5565 29385 5585
rect 29415 5565 29435 5585
rect 29465 5565 29485 5585
rect 29515 5565 29535 5585
rect 29565 5565 29585 5585
rect 29615 5565 29635 5585
rect 29665 5565 29685 5585
rect 29715 5565 29735 5585
rect 29765 5565 29785 5585
rect 29815 5565 29835 5585
rect 29865 5565 29885 5585
rect 29915 5565 29935 5585
rect 29965 5565 29985 5585
rect 30015 5565 30035 5585
rect 30065 5565 30085 5585
rect 30115 5565 30135 5585
rect 30165 5565 30185 5585
rect 30215 5565 30235 5585
rect 30265 5565 30285 5585
rect 30315 5565 30335 5585
rect 30365 5565 30385 5585
rect 30415 5565 30435 5585
rect 30465 5565 30485 5585
rect 30515 5565 30535 5585
rect 30565 5565 30585 5585
rect 30615 5565 30635 5585
rect 30665 5565 30685 5585
rect 30715 5565 30735 5585
rect 30765 5565 30785 5585
rect 30815 5565 30835 5585
rect 30865 5565 30885 5585
rect 30915 5565 30935 5585
rect 30965 5565 30985 5585
rect 31015 5565 31035 5585
rect 31065 5565 31085 5585
rect 31115 5565 31135 5585
rect 31165 5565 31185 5585
rect 31215 5565 31235 5585
rect 31265 5565 31285 5585
rect 31315 5565 31335 5585
rect 31365 5565 31385 5585
rect 31415 5565 31435 5585
rect 31465 5565 31485 5585
rect 31515 5565 31535 5585
rect 31565 5565 31585 5585
rect 31615 5565 31635 5585
rect 31665 5565 31685 5585
rect 31715 5565 31735 5585
rect 31765 5565 31785 5585
rect 31815 5565 31835 5585
rect 31865 5565 31885 5585
rect 31915 5565 31935 5585
rect 31965 5565 31985 5585
rect 32015 5565 32035 5585
rect 32065 5565 32085 5585
rect -635 4265 -615 4285
rect -585 4265 -565 4285
rect -535 4265 -515 4285
rect -485 4265 -465 4285
rect -435 4265 -415 4285
rect -385 4265 -365 4285
rect -335 4265 -315 4285
rect -285 4265 -265 4285
rect -235 4265 -215 4285
rect -185 4265 -165 4285
rect -135 4265 -115 4285
rect -85 4265 -65 4285
rect -35 4265 -15 4285
rect 15 4265 35 4285
rect 65 4265 85 4285
rect 115 4265 135 4285
rect 165 4265 185 4285
rect 215 4265 235 4285
rect 265 4265 285 4285
rect 315 4265 335 4285
rect 365 4265 385 4285
rect 415 4265 435 4285
rect 465 4265 485 4285
rect 515 4265 535 4285
rect 565 4265 585 4285
rect 615 4265 635 4285
rect 665 4265 685 4285
rect 715 4265 735 4285
rect 765 4265 785 4285
rect 815 4265 835 4285
rect 865 4265 885 4285
rect 915 4265 935 4285
rect 965 4265 985 4285
rect 1015 4265 1035 4285
rect 1065 4265 1085 4285
rect 1115 4265 1135 4285
rect 1165 4265 1185 4285
rect 1215 4265 1235 4285
rect 1265 4265 1285 4285
rect 1315 4265 1335 4285
rect 1365 4265 1385 4285
rect 1415 4265 1435 4285
rect 1465 4265 1485 4285
rect 1515 4265 1535 4285
rect 1565 4265 1585 4285
rect 1615 4265 1635 4285
rect 1665 4265 1685 4285
rect 1715 4265 1735 4285
rect 1765 4265 1785 4285
rect 1815 4265 1835 4285
rect 1865 4265 1885 4285
rect 1915 4265 1935 4285
rect 1965 4265 1985 4285
rect 2015 4265 2035 4285
rect 2065 4265 2085 4285
rect 2115 4265 2135 4285
rect 2165 4265 2185 4285
rect 2215 4265 2235 4285
rect 2265 4265 2285 4285
rect 2315 4265 2335 4285
rect 2365 4265 2385 4285
rect 2415 4265 2435 4285
rect 2465 4265 2485 4285
rect 2515 4265 2535 4285
rect 2565 4265 2585 4285
rect 2615 4265 2635 4285
rect 2665 4265 2685 4285
rect 2715 4265 2735 4285
rect 2765 4265 2785 4285
rect 2815 4265 2835 4285
rect 2865 4265 2885 4285
rect 2915 4265 2935 4285
rect 2965 4265 2985 4285
rect 3015 4265 3035 4285
rect 3065 4265 3085 4285
rect 3115 4265 3135 4285
rect 3165 4265 3185 4285
rect 3215 4265 3235 4285
rect 3265 4265 3285 4285
rect 3315 4265 3335 4285
rect 3365 4265 3385 4285
rect 3415 4265 3435 4285
rect 3465 4265 3485 4285
rect 3515 4265 3535 4285
rect 3565 4265 3585 4285
rect 3615 4265 3635 4285
rect 3665 4265 3685 4285
rect 3715 4265 3735 4285
rect 3765 4265 3785 4285
rect 3815 4265 3835 4285
rect 3865 4265 3885 4285
rect 3915 4265 3935 4285
rect 3965 4265 3985 4285
rect 4015 4265 4035 4285
rect 4065 4265 4085 4285
rect 4115 4265 4135 4285
rect 4165 4265 4185 4285
rect 4215 4265 4235 4285
rect 4265 4265 4285 4285
rect 4315 4265 4335 4285
rect 4365 4265 4385 4285
rect 4415 4265 4435 4285
rect 4465 4265 4485 4285
rect 4515 4265 4535 4285
rect 4565 4265 4585 4285
rect 4615 4265 4635 4285
rect 4665 4265 4685 4285
rect 4715 4265 4735 4285
rect 4765 4265 4785 4285
rect 4815 4265 4835 4285
rect 4865 4265 4885 4285
rect 4915 4265 4935 4285
rect 4965 4265 4985 4285
rect 5015 4265 5035 4285
rect 5065 4265 5085 4285
rect 5115 4265 5135 4285
rect 5165 4265 5185 4285
rect 5215 4265 5235 4285
rect 5265 4265 5285 4285
rect 5315 4265 5335 4285
rect 5365 4265 5385 4285
rect 5415 4265 5435 4285
rect 5465 4265 5485 4285
rect 5515 4265 5535 4285
rect 5565 4265 5585 4285
rect 5615 4265 5635 4285
rect 5665 4265 5685 4285
rect 5715 4265 5735 4285
rect 5765 4265 5785 4285
rect 5815 4265 5835 4285
rect 5865 4265 5885 4285
rect 5915 4265 5935 4285
rect 5965 4265 5985 4285
rect 6015 4265 6035 4285
rect 6065 4265 6085 4285
rect 6115 4265 6135 4285
rect 6165 4265 6185 4285
rect 6215 4265 6235 4285
rect 6265 4265 6285 4285
rect 6315 4265 6335 4285
rect 6365 4265 6385 4285
rect 6415 4265 6435 4285
rect 6465 4265 6485 4285
rect 6515 4265 6535 4285
rect 6565 4265 6585 4285
rect 6615 4265 6635 4285
rect 6665 4265 6685 4285
rect 6715 4265 6735 4285
rect 6765 4265 6785 4285
rect 6815 4265 6835 4285
rect 6865 4265 6885 4285
rect 6915 4265 6935 4285
rect 6965 4265 6985 4285
rect 7015 4265 7035 4285
rect 7065 4265 7085 4285
rect 7115 4265 7135 4285
rect 7165 4265 7185 4285
rect 7215 4265 7235 4285
rect 7265 4265 7285 4285
rect 7315 4265 7335 4285
rect 7365 4265 7385 4285
rect 7415 4265 7435 4285
rect 7465 4265 7485 4285
rect 7515 4265 7535 4285
rect 7565 4265 7585 4285
rect 7615 4265 7635 4285
rect 7665 4265 7685 4285
rect 7715 4265 7735 4285
rect 7765 4265 7785 4285
rect 7815 4265 7835 4285
rect 7865 4265 7885 4285
rect 7915 4265 7935 4285
rect 7965 4265 7985 4285
rect 8015 4265 8035 4285
rect 8065 4265 8085 4285
rect 8115 4265 8135 4285
rect 8165 4265 8185 4285
rect 8215 4265 8235 4285
rect 8265 4265 8285 4285
rect 8315 4265 8335 4285
rect 8365 4265 8385 4285
rect 8415 4265 8435 4285
rect 8465 4265 8485 4285
rect 8515 4265 8535 4285
rect 8565 4265 8585 4285
rect 8615 4265 8635 4285
rect 8665 4265 8685 4285
rect 8715 4265 8735 4285
rect 8765 4265 8785 4285
rect 8815 4265 8835 4285
rect 8865 4265 8885 4285
rect 8915 4265 8935 4285
rect 8965 4265 8985 4285
rect 9015 4265 9035 4285
rect 9065 4265 9085 4285
rect 9115 4265 9135 4285
rect 9165 4265 9185 4285
rect 9215 4265 9235 4285
rect 9265 4265 9285 4285
rect 9315 4265 9335 4285
rect 9365 4265 9385 4285
rect 9415 4265 9435 4285
rect 9465 4265 9485 4285
rect 9515 4265 9535 4285
rect 9565 4265 9585 4285
rect 9615 4265 9635 4285
rect 9665 4265 9685 4285
rect 9715 4265 9735 4285
rect 9765 4265 9785 4285
rect 9815 4265 9835 4285
rect 9865 4265 9885 4285
rect 9915 4265 9935 4285
rect 9965 4265 9985 4285
rect 10015 4265 10035 4285
rect 10065 4265 10085 4285
rect 10115 4265 10135 4285
rect 10165 4265 10185 4285
rect 10215 4265 10235 4285
rect 10265 4265 10285 4285
rect 10315 4265 10335 4285
rect 10365 4265 10385 4285
rect 10415 4265 10435 4285
rect 10465 4265 10485 4285
rect 10515 4265 10535 4285
rect 10565 4265 10585 4285
rect 10615 4265 10635 4285
rect 10665 4265 10685 4285
rect 10715 4265 10735 4285
rect 10765 4265 10785 4285
rect 10815 4265 10835 4285
rect 10865 4265 10885 4285
rect 10915 4265 10935 4285
rect 10965 4265 10985 4285
rect 11015 4265 11035 4285
rect 11065 4265 11085 4285
rect 11115 4265 11135 4285
rect 11165 4265 11185 4285
rect 11215 4265 11235 4285
rect 11265 4265 11285 4285
rect 11315 4265 11335 4285
rect 11365 4265 11385 4285
rect 11415 4265 11435 4285
rect 11465 4265 11485 4285
rect 11515 4265 11535 4285
rect 11565 4265 11585 4285
rect 11615 4265 11635 4285
rect 11665 4265 11685 4285
rect 11715 4265 11735 4285
rect 11765 4265 11785 4285
rect 11815 4265 11835 4285
rect 11865 4265 11885 4285
rect 11915 4265 11935 4285
rect 11965 4265 11985 4285
rect 12015 4265 12035 4285
rect 12065 4265 12085 4285
rect 12115 4265 12135 4285
rect 12165 4265 12185 4285
rect 12215 4265 12235 4285
rect 12265 4265 12285 4285
rect 12315 4265 12335 4285
rect 12365 4265 12385 4285
rect 12415 4265 12435 4285
rect 12465 4265 12485 4285
rect 12515 4265 12535 4285
rect 12565 4265 12585 4285
rect 12615 4265 12635 4285
rect 12665 4265 12685 4285
rect 12715 4265 12735 4285
rect 12765 4265 12785 4285
rect 12815 4265 12835 4285
rect 12865 4265 12885 4285
rect 12915 4265 12935 4285
rect 12965 4265 12985 4285
rect 13015 4265 13035 4285
rect 13065 4265 13085 4285
rect 13115 4265 13135 4285
rect 13165 4265 13185 4285
rect 13215 4265 13235 4285
rect 13265 4265 13285 4285
rect 13315 4265 13335 4285
rect 13365 4265 13385 4285
rect 13415 4265 13435 4285
rect 13465 4265 13485 4285
rect 13515 4265 13535 4285
rect 13565 4265 13585 4285
rect 13615 4265 13635 4285
rect 13665 4265 13685 4285
rect 13715 4265 13735 4285
rect 13765 4265 13785 4285
rect 13815 4265 13835 4285
rect 13865 4265 13885 4285
rect 13915 4265 13935 4285
rect 13965 4265 13985 4285
rect 14015 4265 14035 4285
rect 14065 4265 14085 4285
rect 14115 4265 14135 4285
rect 14165 4265 14185 4285
rect 14215 4265 14235 4285
rect 14265 4265 14285 4285
rect 14315 4265 14335 4285
rect 14365 4265 14385 4285
rect 14415 4265 14435 4285
rect 14465 4265 14485 4285
rect 14515 4265 14535 4285
rect 14565 4265 14585 4285
rect 14615 4265 14635 4285
rect 14665 4265 14685 4285
rect 14715 4265 14735 4285
rect 14765 4265 14785 4285
rect 14815 4265 14835 4285
rect 14865 4265 14885 4285
rect 14915 4265 14935 4285
rect 14965 4265 14985 4285
rect 15015 4265 15035 4285
rect 15065 4265 15085 4285
rect 15115 4265 15135 4285
rect 15165 4265 15185 4285
rect 15215 4265 15235 4285
rect 15265 4265 15285 4285
rect 15315 4265 15335 4285
rect 15365 4265 15385 4285
rect 15415 4265 15435 4285
rect 15465 4265 15485 4285
rect 15515 4265 15535 4285
rect 15565 4265 15585 4285
rect 15615 4265 15635 4285
rect 15665 4265 15685 4285
rect 15715 4265 15735 4285
rect 15765 4265 15785 4285
rect 15815 4265 15835 4285
rect 15865 4265 15885 4285
rect 15915 4265 15935 4285
rect 15965 4265 15985 4285
rect 16015 4265 16035 4285
rect 16065 4265 16085 4285
rect 16115 4265 16135 4285
rect 16165 4265 16185 4285
rect 16215 4265 16235 4285
rect 16265 4265 16285 4285
rect 16315 4265 16335 4285
rect 16365 4265 16385 4285
rect 16415 4265 16435 4285
rect 16465 4265 16485 4285
rect 16515 4265 16535 4285
rect 16565 4265 16585 4285
rect 16615 4265 16635 4285
rect 16665 4265 16685 4285
rect 16715 4265 16735 4285
rect 16765 4265 16785 4285
rect 16815 4265 16835 4285
rect 16865 4265 16885 4285
rect 16915 4265 16935 4285
rect 16965 4265 16985 4285
rect 17015 4265 17035 4285
rect 17065 4265 17085 4285
rect 17115 4265 17135 4285
rect 17165 4265 17185 4285
rect 17215 4265 17235 4285
rect 17265 4265 17285 4285
rect 17315 4265 17335 4285
rect 17365 4265 17385 4285
rect 17415 4265 17435 4285
rect 17465 4265 17485 4285
rect 17515 4265 17535 4285
rect 17565 4265 17585 4285
rect 17615 4265 17635 4285
rect 17665 4265 17685 4285
rect 17715 4265 17735 4285
rect 17765 4265 17785 4285
rect 17815 4265 17835 4285
rect 17865 4265 17885 4285
rect 17915 4265 17935 4285
rect 17965 4265 17985 4285
rect 18015 4265 18035 4285
rect 18065 4265 18085 4285
rect 18115 4265 18135 4285
rect 18165 4265 18185 4285
rect 18215 4265 18235 4285
rect 18265 4265 18285 4285
rect 18315 4265 18335 4285
rect 18365 4265 18385 4285
rect 18415 4265 18435 4285
rect 18465 4265 18485 4285
rect 18515 4265 18535 4285
rect 18565 4265 18585 4285
rect 18615 4265 18635 4285
rect 18665 4265 18685 4285
rect 18715 4265 18735 4285
rect 18765 4265 18785 4285
rect 18815 4265 18835 4285
rect 18865 4265 18885 4285
rect 18915 4265 18935 4285
rect 18965 4265 18985 4285
rect 19015 4265 19035 4285
rect 19065 4265 19085 4285
rect 19115 4265 19135 4285
rect 19165 4265 19185 4285
rect 19215 4265 19235 4285
rect 19265 4265 19285 4285
rect 19315 4265 19335 4285
rect 19365 4265 19385 4285
rect 19415 4265 19435 4285
rect 19465 4265 19485 4285
rect 19515 4265 19535 4285
rect 19565 4265 19585 4285
rect 19615 4265 19635 4285
rect 19665 4265 19685 4285
rect 19715 4265 19735 4285
rect 19765 4265 19785 4285
rect 19815 4265 19835 4285
rect 19865 4265 19885 4285
rect 19915 4265 19935 4285
rect 19965 4265 19985 4285
rect 20015 4265 20035 4285
rect 20065 4265 20085 4285
rect 20115 4265 20135 4285
rect 20165 4265 20185 4285
rect 20215 4265 20235 4285
rect 20265 4265 20285 4285
rect 20315 4265 20335 4285
rect 20365 4265 20385 4285
rect 20415 4265 20435 4285
rect 20465 4265 20485 4285
rect 20515 4265 20535 4285
rect 20565 4265 20585 4285
rect 20615 4265 20635 4285
rect 20665 4265 20685 4285
rect 20715 4265 20735 4285
rect 20765 4265 20785 4285
rect 20815 4265 20835 4285
rect 20865 4265 20885 4285
rect 20915 4265 20935 4285
rect 20965 4265 20985 4285
rect 21015 4265 21035 4285
rect 21065 4265 21085 4285
rect 21115 4265 21135 4285
rect 21165 4265 21185 4285
rect 21215 4265 21235 4285
rect 21265 4265 21285 4285
rect 21315 4265 21335 4285
rect 21365 4265 21385 4285
rect 21415 4265 21435 4285
rect 21465 4265 21485 4285
rect 21515 4265 21535 4285
rect 21565 4265 21585 4285
rect 21615 4265 21635 4285
rect 21665 4265 21685 4285
rect 21715 4265 21735 4285
rect 21765 4265 21785 4285
rect 21815 4265 21835 4285
rect 21865 4265 21885 4285
rect 21915 4265 21935 4285
rect 21965 4265 21985 4285
rect 22015 4265 22035 4285
rect 22065 4265 22085 4285
rect 22115 4265 22135 4285
rect 22165 4265 22185 4285
rect 22215 4265 22235 4285
rect 22265 4265 22285 4285
rect 22315 4265 22335 4285
rect 22365 4265 22385 4285
rect 22415 4265 22435 4285
rect 22465 4265 22485 4285
rect 22515 4265 22535 4285
rect 22565 4265 22585 4285
rect 22615 4265 22635 4285
rect 22665 4265 22685 4285
rect 22715 4265 22735 4285
rect 22765 4265 22785 4285
rect 22815 4265 22835 4285
rect 22865 4265 22885 4285
rect 22915 4265 22935 4285
rect 22965 4265 22985 4285
rect 23015 4265 23035 4285
rect 23065 4265 23085 4285
rect 23115 4265 23135 4285
rect 23165 4265 23185 4285
rect 23215 4265 23235 4285
rect 23265 4265 23285 4285
rect 23315 4265 23335 4285
rect 23365 4265 23385 4285
rect 23415 4265 23435 4285
rect 23465 4265 23485 4285
rect 23515 4265 23535 4285
rect 23565 4265 23585 4285
rect 23615 4265 23635 4285
rect 23665 4265 23685 4285
rect 23715 4265 23735 4285
rect 23765 4265 23785 4285
rect 23815 4265 23835 4285
rect 23865 4265 23885 4285
rect 23915 4265 23935 4285
rect 23965 4265 23985 4285
rect 24015 4265 24035 4285
rect 24065 4265 24085 4285
rect 24115 4265 24135 4285
rect 24165 4265 24185 4285
rect 24215 4265 24235 4285
rect 24265 4265 24285 4285
rect 24315 4265 24335 4285
rect 24365 4265 24385 4285
rect 24415 4265 24435 4285
rect 24465 4265 24485 4285
rect 24515 4265 24535 4285
rect 24565 4265 24585 4285
rect 24615 4265 24635 4285
rect 24665 4265 24685 4285
rect 24715 4265 24735 4285
rect 24765 4265 24785 4285
rect 24815 4265 24835 4285
rect 24865 4265 24885 4285
rect 24915 4265 24935 4285
rect 24965 4265 24985 4285
rect 25015 4265 25035 4285
rect 25065 4265 25085 4285
rect 25115 4265 25135 4285
rect 25165 4265 25185 4285
rect 25215 4265 25235 4285
rect 25265 4265 25285 4285
rect 25315 4265 25335 4285
rect 25365 4265 25385 4285
rect 25415 4265 25435 4285
rect 25465 4265 25485 4285
rect 25515 4265 25535 4285
rect 25565 4265 25585 4285
rect 25615 4265 25635 4285
rect 25665 4265 25685 4285
rect 25715 4265 25735 4285
rect 25765 4265 25785 4285
rect 25815 4265 25835 4285
rect 25865 4265 25885 4285
rect 25915 4265 25935 4285
rect 25965 4265 25985 4285
rect 26015 4265 26035 4285
rect 26065 4265 26085 4285
rect 26115 4265 26135 4285
rect 26165 4265 26185 4285
rect 26215 4265 26235 4285
rect 26265 4265 26285 4285
rect 26315 4265 26335 4285
rect 26365 4265 26385 4285
rect 26415 4265 26435 4285
rect 26465 4265 26485 4285
rect 26515 4265 26535 4285
rect 26565 4265 26585 4285
rect 26615 4265 26635 4285
rect 26665 4265 26685 4285
rect 26715 4265 26735 4285
rect 26765 4265 26785 4285
rect 26815 4265 26835 4285
rect 26865 4265 26885 4285
rect 26915 4265 26935 4285
rect 26965 4265 26985 4285
rect 27015 4265 27035 4285
rect 27065 4265 27085 4285
rect 27115 4265 27135 4285
rect 27165 4265 27185 4285
rect 27215 4265 27235 4285
rect 27265 4265 27285 4285
rect 27315 4265 27335 4285
rect 27365 4265 27385 4285
rect 27415 4265 27435 4285
rect 27465 4265 27485 4285
rect 27515 4265 27535 4285
rect 27565 4265 27585 4285
rect 27615 4265 27635 4285
rect 27665 4265 27685 4285
rect 27715 4265 27735 4285
rect 27765 4265 27785 4285
rect 27815 4265 27835 4285
rect 27865 4265 27885 4285
rect 27915 4265 27935 4285
rect 27965 4265 27985 4285
rect 28015 4265 28035 4285
rect 28065 4265 28085 4285
rect 28115 4265 28135 4285
rect 28165 4265 28185 4285
rect 28215 4265 28235 4285
rect 28265 4265 28285 4285
rect 28315 4265 28335 4285
rect 28365 4265 28385 4285
rect 28415 4265 28435 4285
rect 28465 4265 28485 4285
rect 28515 4265 28535 4285
rect 28565 4265 28585 4285
rect 28615 4265 28635 4285
rect 28665 4265 28685 4285
rect 28715 4265 28735 4285
rect 28765 4265 28785 4285
rect 28815 4265 28835 4285
rect 28865 4265 28885 4285
rect 28915 4265 28935 4285
rect 28965 4265 28985 4285
rect 29015 4265 29035 4285
rect 29065 4265 29085 4285
rect 29115 4265 29135 4285
rect 29165 4265 29185 4285
rect 29215 4265 29235 4285
rect 29265 4265 29285 4285
rect 29315 4265 29335 4285
rect 29365 4265 29385 4285
rect 29415 4265 29435 4285
rect 29465 4265 29485 4285
rect 29515 4265 29535 4285
rect 29565 4265 29585 4285
rect 29615 4265 29635 4285
rect 29665 4265 29685 4285
rect 29715 4265 29735 4285
rect 29765 4265 29785 4285
rect 29815 4265 29835 4285
rect 29865 4265 29885 4285
rect 29915 4265 29935 4285
rect 29965 4265 29985 4285
rect 30015 4265 30035 4285
rect 30065 4265 30085 4285
rect 30115 4265 30135 4285
rect 30165 4265 30185 4285
rect 30215 4265 30235 4285
rect 30265 4265 30285 4285
rect 30315 4265 30335 4285
rect 30365 4265 30385 4285
rect 30415 4265 30435 4285
rect 30465 4265 30485 4285
rect 30515 4265 30535 4285
rect 30565 4265 30585 4285
rect 30615 4265 30635 4285
rect 30665 4265 30685 4285
rect 30715 4265 30735 4285
rect 30765 4265 30785 4285
rect 30815 4265 30835 4285
rect 30865 4265 30885 4285
rect 30915 4265 30935 4285
rect 30965 4265 30985 4285
rect 31015 4265 31035 4285
rect 31065 4265 31085 4285
rect 31115 4265 31135 4285
rect 31165 4265 31185 4285
rect 31215 4265 31235 4285
rect 31265 4265 31285 4285
rect 31315 4265 31335 4285
rect 31365 4265 31385 4285
rect 31415 4265 31435 4285
rect 31465 4265 31485 4285
rect 31515 4265 31535 4285
rect 31565 4265 31585 4285
rect 31615 4265 31635 4285
rect 31665 4265 31685 4285
rect 31715 4265 31735 4285
rect 31765 4265 31785 4285
rect 31815 4265 31835 4285
rect 31865 4265 31885 4285
rect 31915 4265 31935 4285
rect 31965 4265 31985 4285
rect 32015 4265 32035 4285
rect 32065 4265 32085 4285
rect -635 2965 -615 2985
rect -585 2965 -565 2985
rect -535 2965 -515 2985
rect -485 2965 -465 2985
rect -435 2965 -415 2985
rect -385 2965 -365 2985
rect -335 2965 -315 2985
rect -285 2965 -265 2985
rect -235 2965 -215 2985
rect -185 2965 -165 2985
rect -135 2965 -115 2985
rect -85 2965 -65 2985
rect -35 2965 -15 2985
rect 15 2965 35 2985
rect 65 2965 85 2985
rect 115 2965 135 2985
rect 165 2965 185 2985
rect 215 2965 235 2985
rect 265 2965 285 2985
rect 315 2965 335 2985
rect 365 2965 385 2985
rect 415 2965 435 2985
rect 465 2965 485 2985
rect 515 2965 535 2985
rect 565 2965 585 2985
rect 615 2965 635 2985
rect 665 2965 685 2985
rect 715 2965 735 2985
rect 765 2965 785 2985
rect 815 2965 835 2985
rect 865 2965 885 2985
rect 915 2965 935 2985
rect 965 2965 985 2985
rect 1015 2965 1035 2985
rect 1065 2965 1085 2985
rect 1115 2965 1135 2985
rect 1165 2965 1185 2985
rect 1215 2965 1235 2985
rect 1265 2965 1285 2985
rect 1315 2965 1335 2985
rect 1365 2965 1385 2985
rect 1415 2965 1435 2985
rect 1465 2965 1485 2985
rect 1515 2965 1535 2985
rect 1565 2965 1585 2985
rect 1615 2965 1635 2985
rect 1665 2965 1685 2985
rect 1715 2965 1735 2985
rect 1765 2965 1785 2985
rect 1815 2965 1835 2985
rect 1865 2965 1885 2985
rect 1915 2965 1935 2985
rect 1965 2965 1985 2985
rect 2015 2965 2035 2985
rect 2065 2965 2085 2985
rect 2115 2965 2135 2985
rect 2165 2965 2185 2985
rect 2215 2965 2235 2985
rect 2265 2965 2285 2985
rect 2315 2965 2335 2985
rect 2365 2965 2385 2985
rect 2415 2965 2435 2985
rect 2465 2965 2485 2985
rect 2515 2965 2535 2985
rect 2565 2965 2585 2985
rect 2615 2965 2635 2985
rect 2665 2965 2685 2985
rect 2715 2965 2735 2985
rect 2765 2965 2785 2985
rect 2815 2965 2835 2985
rect 2865 2965 2885 2985
rect 2915 2965 2935 2985
rect 2965 2965 2985 2985
rect 3015 2965 3035 2985
rect 3065 2965 3085 2985
rect 3115 2965 3135 2985
rect 3165 2965 3185 2985
rect 3215 2965 3235 2985
rect 3265 2965 3285 2985
rect 3315 2965 3335 2985
rect 3365 2965 3385 2985
rect 3415 2965 3435 2985
rect 3465 2965 3485 2985
rect 3515 2965 3535 2985
rect 3565 2965 3585 2985
rect 3615 2965 3635 2985
rect 3665 2965 3685 2985
rect 3715 2965 3735 2985
rect 3765 2965 3785 2985
rect 3815 2965 3835 2985
rect 3865 2965 3885 2985
rect 3915 2965 3935 2985
rect 3965 2965 3985 2985
rect 4015 2965 4035 2985
rect 4065 2965 4085 2985
rect 4115 2965 4135 2985
rect 4165 2965 4185 2985
rect 4215 2965 4235 2985
rect 4265 2965 4285 2985
rect 4315 2965 4335 2985
rect 4365 2965 4385 2985
rect 4415 2965 4435 2985
rect 4465 2965 4485 2985
rect 4515 2965 4535 2985
rect 4565 2965 4585 2985
rect 4615 2965 4635 2985
rect 4665 2965 4685 2985
rect 4715 2965 4735 2985
rect 4765 2965 4785 2985
rect 4815 2965 4835 2985
rect 4865 2965 4885 2985
rect 4915 2965 4935 2985
rect 4965 2965 4985 2985
rect 5015 2965 5035 2985
rect 5065 2965 5085 2985
rect 5115 2965 5135 2985
rect 5165 2965 5185 2985
rect 5215 2965 5235 2985
rect 5265 2965 5285 2985
rect 5315 2965 5335 2985
rect 5365 2965 5385 2985
rect 5415 2965 5435 2985
rect 5465 2965 5485 2985
rect 5515 2965 5535 2985
rect 5565 2965 5585 2985
rect 5615 2965 5635 2985
rect 5665 2965 5685 2985
rect 5715 2965 5735 2985
rect 5765 2965 5785 2985
rect 5815 2965 5835 2985
rect 5865 2965 5885 2985
rect 5915 2965 5935 2985
rect 5965 2965 5985 2985
rect 6015 2965 6035 2985
rect 6065 2965 6085 2985
rect 6115 2965 6135 2985
rect 6165 2965 6185 2985
rect 6215 2965 6235 2985
rect 6265 2965 6285 2985
rect 6315 2965 6335 2985
rect 6365 2965 6385 2985
rect 6415 2965 6435 2985
rect 6465 2965 6485 2985
rect 6515 2965 6535 2985
rect 6565 2965 6585 2985
rect 6615 2965 6635 2985
rect 6665 2965 6685 2985
rect 6715 2965 6735 2985
rect 6765 2965 6785 2985
rect 6815 2965 6835 2985
rect 6865 2965 6885 2985
rect 6915 2965 6935 2985
rect 6965 2965 6985 2985
rect 7015 2965 7035 2985
rect 7065 2965 7085 2985
rect 7115 2965 7135 2985
rect 7165 2965 7185 2985
rect 7215 2965 7235 2985
rect 7265 2965 7285 2985
rect 7315 2965 7335 2985
rect 7365 2965 7385 2985
rect 7415 2965 7435 2985
rect 7465 2965 7485 2985
rect 7515 2965 7535 2985
rect 7565 2965 7585 2985
rect 7615 2965 7635 2985
rect 7665 2965 7685 2985
rect 7715 2965 7735 2985
rect 7765 2965 7785 2985
rect 7815 2965 7835 2985
rect 7865 2965 7885 2985
rect 7915 2965 7935 2985
rect 7965 2965 7985 2985
rect 8015 2965 8035 2985
rect 8065 2965 8085 2985
rect 8115 2965 8135 2985
rect 8165 2965 8185 2985
rect 8215 2965 8235 2985
rect 8265 2965 8285 2985
rect 8315 2965 8335 2985
rect 8365 2965 8385 2985
rect 8415 2965 8435 2985
rect 8465 2965 8485 2985
rect 8515 2965 8535 2985
rect 8565 2965 8585 2985
rect 8615 2965 8635 2985
rect 8665 2965 8685 2985
rect 8715 2965 8735 2985
rect 8765 2965 8785 2985
rect 8815 2965 8835 2985
rect 8865 2965 8885 2985
rect 8915 2965 8935 2985
rect 8965 2965 8985 2985
rect 9015 2965 9035 2985
rect 9065 2965 9085 2985
rect 9115 2965 9135 2985
rect 9165 2965 9185 2985
rect 9215 2965 9235 2985
rect 9265 2965 9285 2985
rect 9315 2965 9335 2985
rect 9365 2965 9385 2985
rect 9415 2965 9435 2985
rect 9465 2965 9485 2985
rect 9515 2965 9535 2985
rect 9565 2965 9585 2985
rect 9615 2965 9635 2985
rect 9665 2965 9685 2985
rect 9715 2965 9735 2985
rect 9765 2965 9785 2985
rect 9815 2965 9835 2985
rect 9865 2965 9885 2985
rect 9915 2965 9935 2985
rect 9965 2965 9985 2985
rect 10015 2965 10035 2985
rect 10065 2965 10085 2985
rect 10115 2965 10135 2985
rect 10165 2965 10185 2985
rect 10215 2965 10235 2985
rect 10265 2965 10285 2985
rect 10315 2965 10335 2985
rect 10365 2965 10385 2985
rect 10415 2965 10435 2985
rect 10465 2965 10485 2985
rect 10515 2965 10535 2985
rect 10565 2965 10585 2985
rect 10615 2965 10635 2985
rect 10665 2965 10685 2985
rect 10715 2965 10735 2985
rect 10765 2965 10785 2985
rect 10815 2965 10835 2985
rect 10865 2965 10885 2985
rect 10915 2965 10935 2985
rect 10965 2965 10985 2985
rect 11015 2965 11035 2985
rect 11065 2965 11085 2985
rect 11115 2965 11135 2985
rect 11165 2965 11185 2985
rect 11215 2965 11235 2985
rect 11265 2965 11285 2985
rect 11315 2965 11335 2985
rect 11365 2965 11385 2985
rect 11415 2965 11435 2985
rect 11465 2965 11485 2985
rect 11515 2965 11535 2985
rect 11565 2965 11585 2985
rect 11615 2965 11635 2985
rect 11665 2965 11685 2985
rect 11715 2965 11735 2985
rect 11765 2965 11785 2985
rect 11815 2965 11835 2985
rect 11865 2965 11885 2985
rect 11915 2965 11935 2985
rect 11965 2965 11985 2985
rect 12015 2965 12035 2985
rect 12065 2965 12085 2985
rect 12115 2965 12135 2985
rect 12165 2965 12185 2985
rect 12215 2965 12235 2985
rect 12265 2965 12285 2985
rect 12315 2965 12335 2985
rect 12365 2965 12385 2985
rect 12415 2965 12435 2985
rect 12465 2965 12485 2985
rect 12515 2965 12535 2985
rect 12565 2965 12585 2985
rect 12615 2965 12635 2985
rect 12665 2965 12685 2985
rect 12715 2965 12735 2985
rect 12765 2965 12785 2985
rect 12815 2965 12835 2985
rect 12865 2965 12885 2985
rect 12915 2965 12935 2985
rect 12965 2965 12985 2985
rect 13015 2965 13035 2985
rect 13065 2965 13085 2985
rect 13115 2965 13135 2985
rect 13165 2965 13185 2985
rect 13215 2965 13235 2985
rect 13265 2965 13285 2985
rect 13315 2965 13335 2985
rect 13365 2965 13385 2985
rect 13415 2965 13435 2985
rect 13465 2965 13485 2985
rect 13515 2965 13535 2985
rect 13565 2965 13585 2985
rect 13615 2965 13635 2985
rect 13665 2965 13685 2985
rect 13715 2965 13735 2985
rect 13765 2965 13785 2985
rect 13815 2965 13835 2985
rect 13865 2965 13885 2985
rect 13915 2965 13935 2985
rect 13965 2965 13985 2985
rect 14015 2965 14035 2985
rect 14065 2965 14085 2985
rect 14115 2965 14135 2985
rect 14165 2965 14185 2985
rect 14215 2965 14235 2985
rect 14265 2965 14285 2985
rect 14315 2965 14335 2985
rect 14365 2965 14385 2985
rect 14415 2965 14435 2985
rect 14465 2965 14485 2985
rect 14515 2965 14535 2985
rect 14565 2965 14585 2985
rect 14615 2965 14635 2985
rect 14665 2965 14685 2985
rect 14715 2965 14735 2985
rect 14765 2965 14785 2985
rect 14815 2965 14835 2985
rect 14865 2965 14885 2985
rect 14915 2965 14935 2985
rect 14965 2965 14985 2985
rect 15015 2965 15035 2985
rect 15065 2965 15085 2985
rect 15115 2965 15135 2985
rect 15165 2965 15185 2985
rect 15215 2965 15235 2985
rect 15265 2965 15285 2985
rect 15315 2965 15335 2985
rect 15365 2965 15385 2985
rect 15415 2965 15435 2985
rect 15465 2965 15485 2985
rect 15515 2965 15535 2985
rect 15565 2965 15585 2985
rect 15615 2965 15635 2985
rect 15665 2965 15685 2985
rect 15715 2965 15735 2985
rect 15765 2965 15785 2985
rect 15815 2965 15835 2985
rect 15865 2965 15885 2985
rect 15915 2965 15935 2985
rect 15965 2965 15985 2985
rect 16015 2965 16035 2985
rect 16065 2965 16085 2985
rect 16115 2965 16135 2985
rect 16165 2965 16185 2985
rect 16215 2965 16235 2985
rect 16265 2965 16285 2985
rect 16315 2965 16335 2985
rect 16365 2965 16385 2985
rect 16415 2965 16435 2985
rect 16465 2965 16485 2985
rect 16515 2965 16535 2985
rect 16565 2965 16585 2985
rect 16615 2965 16635 2985
rect 16665 2965 16685 2985
rect 16715 2965 16735 2985
rect 16765 2965 16785 2985
rect 16815 2965 16835 2985
rect 16865 2965 16885 2985
rect 16915 2965 16935 2985
rect 16965 2965 16985 2985
rect 17015 2965 17035 2985
rect 17065 2965 17085 2985
rect 17115 2965 17135 2985
rect 17165 2965 17185 2985
rect 17215 2965 17235 2985
rect 17265 2965 17285 2985
rect 17315 2965 17335 2985
rect 17365 2965 17385 2985
rect 17415 2965 17435 2985
rect 17465 2965 17485 2985
rect 17515 2965 17535 2985
rect 17565 2965 17585 2985
rect 17615 2965 17635 2985
rect 17665 2965 17685 2985
rect 17715 2965 17735 2985
rect 17765 2965 17785 2985
rect 17815 2965 17835 2985
rect 17865 2965 17885 2985
rect 17915 2965 17935 2985
rect 17965 2965 17985 2985
rect 18015 2965 18035 2985
rect 18065 2965 18085 2985
rect 18115 2965 18135 2985
rect 18165 2965 18185 2985
rect 18215 2965 18235 2985
rect 18265 2965 18285 2985
rect 18315 2965 18335 2985
rect 18365 2965 18385 2985
rect 18415 2965 18435 2985
rect 18465 2965 18485 2985
rect 18515 2965 18535 2985
rect 18565 2965 18585 2985
rect 18615 2965 18635 2985
rect 18665 2965 18685 2985
rect 18715 2965 18735 2985
rect 18765 2965 18785 2985
rect 18815 2965 18835 2985
rect 18865 2965 18885 2985
rect 18915 2965 18935 2985
rect 18965 2965 18985 2985
rect 19015 2965 19035 2985
rect 19065 2965 19085 2985
rect 19115 2965 19135 2985
rect 19165 2965 19185 2985
rect 19215 2965 19235 2985
rect 19265 2965 19285 2985
rect 19315 2965 19335 2985
rect 19365 2965 19385 2985
rect 19415 2965 19435 2985
rect 19465 2965 19485 2985
rect 19515 2965 19535 2985
rect 19565 2965 19585 2985
rect 19615 2965 19635 2985
rect 19665 2965 19685 2985
rect 19715 2965 19735 2985
rect 19765 2965 19785 2985
rect 19815 2965 19835 2985
rect 19865 2965 19885 2985
rect 19915 2965 19935 2985
rect 19965 2965 19985 2985
rect 20015 2965 20035 2985
rect 20065 2965 20085 2985
rect 20115 2965 20135 2985
rect 20165 2965 20185 2985
rect 20215 2965 20235 2985
rect 20265 2965 20285 2985
rect 20315 2965 20335 2985
rect 20365 2965 20385 2985
rect 20415 2965 20435 2985
rect 20465 2965 20485 2985
rect 20515 2965 20535 2985
rect 20565 2965 20585 2985
rect 20615 2965 20635 2985
rect 20665 2965 20685 2985
rect 20715 2965 20735 2985
rect 20765 2965 20785 2985
rect 20815 2965 20835 2985
rect 20865 2965 20885 2985
rect 20915 2965 20935 2985
rect 20965 2965 20985 2985
rect 21015 2965 21035 2985
rect 21065 2965 21085 2985
rect 21115 2965 21135 2985
rect 21165 2965 21185 2985
rect 21215 2965 21235 2985
rect 21265 2965 21285 2985
rect 21315 2965 21335 2985
rect 21365 2965 21385 2985
rect 21415 2965 21435 2985
rect 21465 2965 21485 2985
rect 21515 2965 21535 2985
rect 21565 2965 21585 2985
rect 21615 2965 21635 2985
rect 21665 2965 21685 2985
rect 21715 2965 21735 2985
rect 21765 2965 21785 2985
rect 21815 2965 21835 2985
rect 21865 2965 21885 2985
rect 21915 2965 21935 2985
rect 21965 2965 21985 2985
rect 22015 2965 22035 2985
rect 22065 2965 22085 2985
rect 22115 2965 22135 2985
rect 22165 2965 22185 2985
rect 22215 2965 22235 2985
rect 22265 2965 22285 2985
rect 22315 2965 22335 2985
rect 22365 2965 22385 2985
rect 22415 2965 22435 2985
rect 22465 2965 22485 2985
rect 22515 2965 22535 2985
rect 22565 2965 22585 2985
rect 22615 2965 22635 2985
rect 22665 2965 22685 2985
rect 22715 2965 22735 2985
rect 22765 2965 22785 2985
rect 22815 2965 22835 2985
rect 22865 2965 22885 2985
rect 22915 2965 22935 2985
rect 22965 2965 22985 2985
rect 23015 2965 23035 2985
rect 23065 2965 23085 2985
rect 23115 2965 23135 2985
rect 23165 2965 23185 2985
rect 23215 2965 23235 2985
rect 23265 2965 23285 2985
rect 23315 2965 23335 2985
rect 23365 2965 23385 2985
rect 23415 2965 23435 2985
rect 23465 2965 23485 2985
rect 23515 2965 23535 2985
rect 23565 2965 23585 2985
rect 23615 2965 23635 2985
rect 23665 2965 23685 2985
rect 23715 2965 23735 2985
rect 23765 2965 23785 2985
rect 23815 2965 23835 2985
rect 23865 2965 23885 2985
rect 23915 2965 23935 2985
rect 23965 2965 23985 2985
rect 24015 2965 24035 2985
rect 24065 2965 24085 2985
rect 24115 2965 24135 2985
rect 24165 2965 24185 2985
rect 24215 2965 24235 2985
rect 24265 2965 24285 2985
rect 24315 2965 24335 2985
rect 24365 2965 24385 2985
rect 24415 2965 24435 2985
rect 24465 2965 24485 2985
rect 24515 2965 24535 2985
rect 24565 2965 24585 2985
rect 24615 2965 24635 2985
rect 24665 2965 24685 2985
rect 24715 2965 24735 2985
rect 24765 2965 24785 2985
rect 24815 2965 24835 2985
rect 24865 2965 24885 2985
rect 24915 2965 24935 2985
rect 24965 2965 24985 2985
rect 25015 2965 25035 2985
rect 25065 2965 25085 2985
rect 25115 2965 25135 2985
rect 25165 2965 25185 2985
rect 25215 2965 25235 2985
rect 25265 2965 25285 2985
rect 25315 2965 25335 2985
rect 25365 2965 25385 2985
rect 25415 2965 25435 2985
rect 25465 2965 25485 2985
rect 25515 2965 25535 2985
rect 25565 2965 25585 2985
rect 25615 2965 25635 2985
rect 25665 2965 25685 2985
rect 25715 2965 25735 2985
rect 25765 2965 25785 2985
rect 25815 2965 25835 2985
rect 25865 2965 25885 2985
rect 25915 2965 25935 2985
rect 25965 2965 25985 2985
rect 26015 2965 26035 2985
rect 26065 2965 26085 2985
rect 26115 2965 26135 2985
rect 26165 2965 26185 2985
rect 26215 2965 26235 2985
rect 26265 2965 26285 2985
rect 26315 2965 26335 2985
rect 26365 2965 26385 2985
rect 26415 2965 26435 2985
rect 26465 2965 26485 2985
rect 26515 2965 26535 2985
rect 26565 2965 26585 2985
rect 26615 2965 26635 2985
rect 26665 2965 26685 2985
rect 26715 2965 26735 2985
rect 26765 2965 26785 2985
rect 26815 2965 26835 2985
rect 26865 2965 26885 2985
rect 26915 2965 26935 2985
rect 26965 2965 26985 2985
rect 27015 2965 27035 2985
rect 27065 2965 27085 2985
rect 27115 2965 27135 2985
rect 27165 2965 27185 2985
rect 27215 2965 27235 2985
rect 27265 2965 27285 2985
rect 27315 2965 27335 2985
rect 27365 2965 27385 2985
rect 27415 2965 27435 2985
rect 27465 2965 27485 2985
rect 27515 2965 27535 2985
rect 27565 2965 27585 2985
rect 27615 2965 27635 2985
rect 27665 2965 27685 2985
rect 27715 2965 27735 2985
rect 27765 2965 27785 2985
rect 27815 2965 27835 2985
rect 27865 2965 27885 2985
rect 27915 2965 27935 2985
rect 27965 2965 27985 2985
rect 28015 2965 28035 2985
rect 28065 2965 28085 2985
rect 28115 2965 28135 2985
rect 28165 2965 28185 2985
rect 28215 2965 28235 2985
rect 28265 2965 28285 2985
rect 28315 2965 28335 2985
rect 28365 2965 28385 2985
rect 28415 2965 28435 2985
rect 28465 2965 28485 2985
rect 28515 2965 28535 2985
rect 28565 2965 28585 2985
rect 28615 2965 28635 2985
rect 28665 2965 28685 2985
rect 28715 2965 28735 2985
rect 28765 2965 28785 2985
rect 28815 2965 28835 2985
rect 28865 2965 28885 2985
rect 28915 2965 28935 2985
rect 28965 2965 28985 2985
rect 29015 2965 29035 2985
rect 29065 2965 29085 2985
rect 29115 2965 29135 2985
rect 29165 2965 29185 2985
rect 29215 2965 29235 2985
rect 29265 2965 29285 2985
rect 29315 2965 29335 2985
rect 29365 2965 29385 2985
rect 29415 2965 29435 2985
rect 29465 2965 29485 2985
rect 29515 2965 29535 2985
rect 29565 2965 29585 2985
rect 29615 2965 29635 2985
rect 29665 2965 29685 2985
rect 29715 2965 29735 2985
rect 29765 2965 29785 2985
rect 29815 2965 29835 2985
rect 29865 2965 29885 2985
rect 29915 2965 29935 2985
rect 29965 2965 29985 2985
rect 30015 2965 30035 2985
rect 30065 2965 30085 2985
rect 30115 2965 30135 2985
rect 30165 2965 30185 2985
rect 30215 2965 30235 2985
rect 30265 2965 30285 2985
rect 30315 2965 30335 2985
rect 30365 2965 30385 2985
rect 30415 2965 30435 2985
rect 30465 2965 30485 2985
rect 30515 2965 30535 2985
rect 30565 2965 30585 2985
rect 30615 2965 30635 2985
rect 30665 2965 30685 2985
rect 30715 2965 30735 2985
rect 30765 2965 30785 2985
rect 30815 2965 30835 2985
rect 30865 2965 30885 2985
rect 30915 2965 30935 2985
rect 30965 2965 30985 2985
rect 31015 2965 31035 2985
rect 31065 2965 31085 2985
rect 31115 2965 31135 2985
rect 31165 2965 31185 2985
rect 31215 2965 31235 2985
rect 31265 2965 31285 2985
rect 31315 2965 31335 2985
rect 31365 2965 31385 2985
rect 31415 2965 31435 2985
rect 31465 2965 31485 2985
rect 31515 2965 31535 2985
rect 31565 2965 31585 2985
rect 31615 2965 31635 2985
rect 31665 2965 31685 2985
rect 31715 2965 31735 2985
rect 31765 2965 31785 2985
rect 31815 2965 31835 2985
rect 31865 2965 31885 2985
rect 31915 2965 31935 2985
rect 31965 2965 31985 2985
rect 32015 2965 32035 2985
rect 32065 2965 32085 2985
rect -635 1815 -615 1835
rect -585 1815 -565 1835
rect -535 1815 -515 1835
rect -485 1815 -465 1835
rect -435 1815 -415 1835
rect -385 1815 -365 1835
rect -335 1815 -315 1835
rect -285 1815 -265 1835
rect -235 1815 -215 1835
rect -185 1815 -165 1835
rect -135 1815 -115 1835
rect -85 1815 -65 1835
rect -35 1815 -15 1835
rect 15 1815 35 1835
rect 65 1815 85 1835
rect 115 1815 135 1835
rect 165 1815 185 1835
rect 215 1815 235 1835
rect 265 1815 285 1835
rect 315 1815 335 1835
rect 365 1815 385 1835
rect 415 1815 435 1835
rect 465 1815 485 1835
rect 515 1815 535 1835
rect 565 1815 585 1835
rect 615 1815 635 1835
rect 665 1815 685 1835
rect 715 1815 735 1835
rect 765 1815 785 1835
rect 815 1815 835 1835
rect 865 1815 885 1835
rect 915 1815 935 1835
rect 965 1815 985 1835
rect 1015 1815 1035 1835
rect 1065 1815 1085 1835
rect 1115 1815 1135 1835
rect 1165 1815 1185 1835
rect 1215 1815 1235 1835
rect 1265 1815 1285 1835
rect 1315 1815 1335 1835
rect 1365 1815 1385 1835
rect 1415 1815 1435 1835
rect 1465 1815 1485 1835
rect 1515 1815 1535 1835
rect 1565 1815 1585 1835
rect 1615 1815 1635 1835
rect 1665 1815 1685 1835
rect 1715 1815 1735 1835
rect 1765 1815 1785 1835
rect 1815 1815 1835 1835
rect 1865 1815 1885 1835
rect 1915 1815 1935 1835
rect 1965 1815 1985 1835
rect 2015 1815 2035 1835
rect 2065 1815 2085 1835
rect 2115 1815 2135 1835
rect 2165 1815 2185 1835
rect 2215 1815 2235 1835
rect 2265 1815 2285 1835
rect 2315 1815 2335 1835
rect 2365 1815 2385 1835
rect 2415 1815 2435 1835
rect 2465 1815 2485 1835
rect 2515 1815 2535 1835
rect 2565 1815 2585 1835
rect 2615 1815 2635 1835
rect 2665 1815 2685 1835
rect 2715 1815 2735 1835
rect 2765 1815 2785 1835
rect 2815 1815 2835 1835
rect 2865 1815 2885 1835
rect 2915 1815 2935 1835
rect 2965 1815 2985 1835
rect 3015 1815 3035 1835
rect 3065 1815 3085 1835
rect 3115 1815 3135 1835
rect 3165 1815 3185 1835
rect 3215 1815 3235 1835
rect 3265 1815 3285 1835
rect 3315 1815 3335 1835
rect 3365 1815 3385 1835
rect 3415 1815 3435 1835
rect 3465 1815 3485 1835
rect 3515 1815 3535 1835
rect 3565 1815 3585 1835
rect 3615 1815 3635 1835
rect 3665 1815 3685 1835
rect 3715 1815 3735 1835
rect 3765 1815 3785 1835
rect 3815 1815 3835 1835
rect 3865 1815 3885 1835
rect 3915 1815 3935 1835
rect 3965 1815 3985 1835
rect 4015 1815 4035 1835
rect 4065 1815 4085 1835
rect 4115 1815 4135 1835
rect 4165 1815 4185 1835
rect 4215 1815 4235 1835
rect 4265 1815 4285 1835
rect 4315 1815 4335 1835
rect 4365 1815 4385 1835
rect 4415 1815 4435 1835
rect 4465 1815 4485 1835
rect 4515 1815 4535 1835
rect 4565 1815 4585 1835
rect 4615 1815 4635 1835
rect 4665 1815 4685 1835
rect 4715 1815 4735 1835
rect 4765 1815 4785 1835
rect 4815 1815 4835 1835
rect 4865 1815 4885 1835
rect 4915 1815 4935 1835
rect 4965 1815 4985 1835
rect 5015 1815 5035 1835
rect 5065 1815 5085 1835
rect 5115 1815 5135 1835
rect 5165 1815 5185 1835
rect 5215 1815 5235 1835
rect 5265 1815 5285 1835
rect 5315 1815 5335 1835
rect 5365 1815 5385 1835
rect 5415 1815 5435 1835
rect 5465 1815 5485 1835
rect 5515 1815 5535 1835
rect 5565 1815 5585 1835
rect 5615 1815 5635 1835
rect 5665 1815 5685 1835
rect 5715 1815 5735 1835
rect 5765 1815 5785 1835
rect 5815 1815 5835 1835
rect 5865 1815 5885 1835
rect 5915 1815 5935 1835
rect 5965 1815 5985 1835
rect 6015 1815 6035 1835
rect 6065 1815 6085 1835
rect 6115 1815 6135 1835
rect 6165 1815 6185 1835
rect 6215 1815 6235 1835
rect 6265 1815 6285 1835
rect 6315 1815 6335 1835
rect 6365 1815 6385 1835
rect 6415 1815 6435 1835
rect 6465 1815 6485 1835
rect 6515 1815 6535 1835
rect 6565 1815 6585 1835
rect 6615 1815 6635 1835
rect 6665 1815 6685 1835
rect 6715 1815 6735 1835
rect 6765 1815 6785 1835
rect 6815 1815 6835 1835
rect 6865 1815 6885 1835
rect 6915 1815 6935 1835
rect 6965 1815 6985 1835
rect 7015 1815 7035 1835
rect 7065 1815 7085 1835
rect 7115 1815 7135 1835
rect 7165 1815 7185 1835
rect 7215 1815 7235 1835
rect 7265 1815 7285 1835
rect 7315 1815 7335 1835
rect 7365 1815 7385 1835
rect 7415 1815 7435 1835
rect 7465 1815 7485 1835
rect 7515 1815 7535 1835
rect 7565 1815 7585 1835
rect 7615 1815 7635 1835
rect 7665 1815 7685 1835
rect 7715 1815 7735 1835
rect 7765 1815 7785 1835
rect 7815 1815 7835 1835
rect 7865 1815 7885 1835
rect 7915 1815 7935 1835
rect 7965 1815 7985 1835
rect 8015 1815 8035 1835
rect 8065 1815 8085 1835
rect 8115 1815 8135 1835
rect 8165 1815 8185 1835
rect 8215 1815 8235 1835
rect 8265 1815 8285 1835
rect 8315 1815 8335 1835
rect 8365 1815 8385 1835
rect 8415 1815 8435 1835
rect 8465 1815 8485 1835
rect 8515 1815 8535 1835
rect 8565 1815 8585 1835
rect 8615 1815 8635 1835
rect 8665 1815 8685 1835
rect 8715 1815 8735 1835
rect 8765 1815 8785 1835
rect 8815 1815 8835 1835
rect 8865 1815 8885 1835
rect 8915 1815 8935 1835
rect 8965 1815 8985 1835
rect 9015 1815 9035 1835
rect 9065 1815 9085 1835
rect 9115 1815 9135 1835
rect 9165 1815 9185 1835
rect 9215 1815 9235 1835
rect 9265 1815 9285 1835
rect 9315 1815 9335 1835
rect 9365 1815 9385 1835
rect 9415 1815 9435 1835
rect 9465 1815 9485 1835
rect 9515 1815 9535 1835
rect 9565 1815 9585 1835
rect 9615 1815 9635 1835
rect 9665 1815 9685 1835
rect 9715 1815 9735 1835
rect 9765 1815 9785 1835
rect 9815 1815 9835 1835
rect 9865 1815 9885 1835
rect 9915 1815 9935 1835
rect 9965 1815 9985 1835
rect 10015 1815 10035 1835
rect 10065 1815 10085 1835
rect 10115 1815 10135 1835
rect 10165 1815 10185 1835
rect 10215 1815 10235 1835
rect 10265 1815 10285 1835
rect 10315 1815 10335 1835
rect 10365 1815 10385 1835
rect 10415 1815 10435 1835
rect 10465 1815 10485 1835
rect 10515 1815 10535 1835
rect 10565 1815 10585 1835
rect 10615 1815 10635 1835
rect 10665 1815 10685 1835
rect 10715 1815 10735 1835
rect 10765 1815 10785 1835
rect 10815 1815 10835 1835
rect 10865 1815 10885 1835
rect 10915 1815 10935 1835
rect 10965 1815 10985 1835
rect 11015 1815 11035 1835
rect 11065 1815 11085 1835
rect 11115 1815 11135 1835
rect 11165 1815 11185 1835
rect 11215 1815 11235 1835
rect 11265 1815 11285 1835
rect 11315 1815 11335 1835
rect 11365 1815 11385 1835
rect 11415 1815 11435 1835
rect 11465 1815 11485 1835
rect 11515 1815 11535 1835
rect 11565 1815 11585 1835
rect 11615 1815 11635 1835
rect 11665 1815 11685 1835
rect 11715 1815 11735 1835
rect 11765 1815 11785 1835
rect 11815 1815 11835 1835
rect 11865 1815 11885 1835
rect 11915 1815 11935 1835
rect 11965 1815 11985 1835
rect 12015 1815 12035 1835
rect 12065 1815 12085 1835
rect 12115 1815 12135 1835
rect 12165 1815 12185 1835
rect 12215 1815 12235 1835
rect 12265 1815 12285 1835
rect 12315 1815 12335 1835
rect 12365 1815 12385 1835
rect 12415 1815 12435 1835
rect 12465 1815 12485 1835
rect 12515 1815 12535 1835
rect 12565 1815 12585 1835
rect 12615 1815 12635 1835
rect 12665 1815 12685 1835
rect 12715 1815 12735 1835
rect 12765 1815 12785 1835
rect 12815 1815 12835 1835
rect 12865 1815 12885 1835
rect 12915 1815 12935 1835
rect 12965 1815 12985 1835
rect 13015 1815 13035 1835
rect 13065 1815 13085 1835
rect 13115 1815 13135 1835
rect 13165 1815 13185 1835
rect 13215 1815 13235 1835
rect 13265 1815 13285 1835
rect 13315 1815 13335 1835
rect 13365 1815 13385 1835
rect 13415 1815 13435 1835
rect 13465 1815 13485 1835
rect 13515 1815 13535 1835
rect 13565 1815 13585 1835
rect 13615 1815 13635 1835
rect 13665 1815 13685 1835
rect 13715 1815 13735 1835
rect 13765 1815 13785 1835
rect 13815 1815 13835 1835
rect 13865 1815 13885 1835
rect 13915 1815 13935 1835
rect 13965 1815 13985 1835
rect 14015 1815 14035 1835
rect 14065 1815 14085 1835
rect 14115 1815 14135 1835
rect 14165 1815 14185 1835
rect 14215 1815 14235 1835
rect 14265 1815 14285 1835
rect 14315 1815 14335 1835
rect 14365 1815 14385 1835
rect 14415 1815 14435 1835
rect 14465 1815 14485 1835
rect 14515 1815 14535 1835
rect 14565 1815 14585 1835
rect 14615 1815 14635 1835
rect 14665 1815 14685 1835
rect 14715 1815 14735 1835
rect 14765 1815 14785 1835
rect 14815 1815 14835 1835
rect 14865 1815 14885 1835
rect 14915 1815 14935 1835
rect 14965 1815 14985 1835
rect 15015 1815 15035 1835
rect 15065 1815 15085 1835
rect 15115 1815 15135 1835
rect 15165 1815 15185 1835
rect 15215 1815 15235 1835
rect 15265 1815 15285 1835
rect 15315 1815 15335 1835
rect 15365 1815 15385 1835
rect 15415 1815 15435 1835
rect 15465 1815 15485 1835
rect 15515 1815 15535 1835
rect 15565 1815 15585 1835
rect 15615 1815 15635 1835
rect 15665 1815 15685 1835
rect 15715 1815 15735 1835
rect 15765 1815 15785 1835
rect 15815 1815 15835 1835
rect 15865 1815 15885 1835
rect 15915 1815 15935 1835
rect 15965 1815 15985 1835
rect 16015 1815 16035 1835
rect 16065 1815 16085 1835
rect 16115 1815 16135 1835
rect 16165 1815 16185 1835
rect 16215 1815 16235 1835
rect 16265 1815 16285 1835
rect 16315 1815 16335 1835
rect 16365 1815 16385 1835
rect 16415 1815 16435 1835
rect 16465 1815 16485 1835
rect 16515 1815 16535 1835
rect 16565 1815 16585 1835
rect 16615 1815 16635 1835
rect 16665 1815 16685 1835
rect 16715 1815 16735 1835
rect 16765 1815 16785 1835
rect 16815 1815 16835 1835
rect 16865 1815 16885 1835
rect 16915 1815 16935 1835
rect 16965 1815 16985 1835
rect 17015 1815 17035 1835
rect 17065 1815 17085 1835
rect 17115 1815 17135 1835
rect 17165 1815 17185 1835
rect 17215 1815 17235 1835
rect 17265 1815 17285 1835
rect 17315 1815 17335 1835
rect 17365 1815 17385 1835
rect 17415 1815 17435 1835
rect 17465 1815 17485 1835
rect 17515 1815 17535 1835
rect 17565 1815 17585 1835
rect 17615 1815 17635 1835
rect 17665 1815 17685 1835
rect 17715 1815 17735 1835
rect 17765 1815 17785 1835
rect 17815 1815 17835 1835
rect 17865 1815 17885 1835
rect 17915 1815 17935 1835
rect 17965 1815 17985 1835
rect 18015 1815 18035 1835
rect 18065 1815 18085 1835
rect 18115 1815 18135 1835
rect 18165 1815 18185 1835
rect 18215 1815 18235 1835
rect 18265 1815 18285 1835
rect 18315 1815 18335 1835
rect 18365 1815 18385 1835
rect 18415 1815 18435 1835
rect 18465 1815 18485 1835
rect 18515 1815 18535 1835
rect 18565 1815 18585 1835
rect 18615 1815 18635 1835
rect 18665 1815 18685 1835
rect 18715 1815 18735 1835
rect 18765 1815 18785 1835
rect 18815 1815 18835 1835
rect 18865 1815 18885 1835
rect 18915 1815 18935 1835
rect 18965 1815 18985 1835
rect 19015 1815 19035 1835
rect 19065 1815 19085 1835
rect 19115 1815 19135 1835
rect 19165 1815 19185 1835
rect 19215 1815 19235 1835
rect 19265 1815 19285 1835
rect 19315 1815 19335 1835
rect 19365 1815 19385 1835
rect 19415 1815 19435 1835
rect 19465 1815 19485 1835
rect 19515 1815 19535 1835
rect 19565 1815 19585 1835
rect 19615 1815 19635 1835
rect 19665 1815 19685 1835
rect 19715 1815 19735 1835
rect 19765 1815 19785 1835
rect 19815 1815 19835 1835
rect 19865 1815 19885 1835
rect 19915 1815 19935 1835
rect 19965 1815 19985 1835
rect 20015 1815 20035 1835
rect 20065 1815 20085 1835
rect 20115 1815 20135 1835
rect 20165 1815 20185 1835
rect 20215 1815 20235 1835
rect 20265 1815 20285 1835
rect 20315 1815 20335 1835
rect 20365 1815 20385 1835
rect 20415 1815 20435 1835
rect 20465 1815 20485 1835
rect 20515 1815 20535 1835
rect 20565 1815 20585 1835
rect 20615 1815 20635 1835
rect 20665 1815 20685 1835
rect 20715 1815 20735 1835
rect 20765 1815 20785 1835
rect 20815 1815 20835 1835
rect 20865 1815 20885 1835
rect 20915 1815 20935 1835
rect 20965 1815 20985 1835
rect 21015 1815 21035 1835
rect 21065 1815 21085 1835
rect 21115 1815 21135 1835
rect 21165 1815 21185 1835
rect 21215 1815 21235 1835
rect 21265 1815 21285 1835
rect 21315 1815 21335 1835
rect 21365 1815 21385 1835
rect 21415 1815 21435 1835
rect 21465 1815 21485 1835
rect 21515 1815 21535 1835
rect 21565 1815 21585 1835
rect 21615 1815 21635 1835
rect 21665 1815 21685 1835
rect 21715 1815 21735 1835
rect 21765 1815 21785 1835
rect 21815 1815 21835 1835
rect 21865 1815 21885 1835
rect 21915 1815 21935 1835
rect 21965 1815 21985 1835
rect 22015 1815 22035 1835
rect 22065 1815 22085 1835
rect 22115 1815 22135 1835
rect 22165 1815 22185 1835
rect 22215 1815 22235 1835
rect 22265 1815 22285 1835
rect 22315 1815 22335 1835
rect 22365 1815 22385 1835
rect 22415 1815 22435 1835
rect 22465 1815 22485 1835
rect 22515 1815 22535 1835
rect 22565 1815 22585 1835
rect 22615 1815 22635 1835
rect 22665 1815 22685 1835
rect 22715 1815 22735 1835
rect 22765 1815 22785 1835
rect 22815 1815 22835 1835
rect 22865 1815 22885 1835
rect 22915 1815 22935 1835
rect 22965 1815 22985 1835
rect 23015 1815 23035 1835
rect 23065 1815 23085 1835
rect 23115 1815 23135 1835
rect 23165 1815 23185 1835
rect 23215 1815 23235 1835
rect 23265 1815 23285 1835
rect 23315 1815 23335 1835
rect 23365 1815 23385 1835
rect 23415 1815 23435 1835
rect 23465 1815 23485 1835
rect 23515 1815 23535 1835
rect 23565 1815 23585 1835
rect 23615 1815 23635 1835
rect 23665 1815 23685 1835
rect 23715 1815 23735 1835
rect 23765 1815 23785 1835
rect 23815 1815 23835 1835
rect 23865 1815 23885 1835
rect 23915 1815 23935 1835
rect 23965 1815 23985 1835
rect 24015 1815 24035 1835
rect 24065 1815 24085 1835
rect 24115 1815 24135 1835
rect 24165 1815 24185 1835
rect 24215 1815 24235 1835
rect 24265 1815 24285 1835
rect 24315 1815 24335 1835
rect 24365 1815 24385 1835
rect 24415 1815 24435 1835
rect 24465 1815 24485 1835
rect 24515 1815 24535 1835
rect 24565 1815 24585 1835
rect 24615 1815 24635 1835
rect 24665 1815 24685 1835
rect 24715 1815 24735 1835
rect 24765 1815 24785 1835
rect 24815 1815 24835 1835
rect 24865 1815 24885 1835
rect 24915 1815 24935 1835
rect 24965 1815 24985 1835
rect 25015 1815 25035 1835
rect 25065 1815 25085 1835
rect 25115 1815 25135 1835
rect 25165 1815 25185 1835
rect 25215 1815 25235 1835
rect 25265 1815 25285 1835
rect 25315 1815 25335 1835
rect 25365 1815 25385 1835
rect 25415 1815 25435 1835
rect 25465 1815 25485 1835
rect 25515 1815 25535 1835
rect 25565 1815 25585 1835
rect 25615 1815 25635 1835
rect 25665 1815 25685 1835
rect 25715 1815 25735 1835
rect 25765 1815 25785 1835
rect 25815 1815 25835 1835
rect 25865 1815 25885 1835
rect 25915 1815 25935 1835
rect 25965 1815 25985 1835
rect 26015 1815 26035 1835
rect 26065 1815 26085 1835
rect 26115 1815 26135 1835
rect 26165 1815 26185 1835
rect 26215 1815 26235 1835
rect 26265 1815 26285 1835
rect 26315 1815 26335 1835
rect 26365 1815 26385 1835
rect 26415 1815 26435 1835
rect 26465 1815 26485 1835
rect 26515 1815 26535 1835
rect 26565 1815 26585 1835
rect 26615 1815 26635 1835
rect 26665 1815 26685 1835
rect 26715 1815 26735 1835
rect 26765 1815 26785 1835
rect 26815 1815 26835 1835
rect 26865 1815 26885 1835
rect 26915 1815 26935 1835
rect 26965 1815 26985 1835
rect 27015 1815 27035 1835
rect 27065 1815 27085 1835
rect 27115 1815 27135 1835
rect 27165 1815 27185 1835
rect 27215 1815 27235 1835
rect 27265 1815 27285 1835
rect 27315 1815 27335 1835
rect 27365 1815 27385 1835
rect 27415 1815 27435 1835
rect 27465 1815 27485 1835
rect 27515 1815 27535 1835
rect 27565 1815 27585 1835
rect 27615 1815 27635 1835
rect 27665 1815 27685 1835
rect 27715 1815 27735 1835
rect 27765 1815 27785 1835
rect 27815 1815 27835 1835
rect 27865 1815 27885 1835
rect 27915 1815 27935 1835
rect 27965 1815 27985 1835
rect 28015 1815 28035 1835
rect 28065 1815 28085 1835
rect 28115 1815 28135 1835
rect 28165 1815 28185 1835
rect 28215 1815 28235 1835
rect 28265 1815 28285 1835
rect 28315 1815 28335 1835
rect 28365 1815 28385 1835
rect 28415 1815 28435 1835
rect 28465 1815 28485 1835
rect 28515 1815 28535 1835
rect 28565 1815 28585 1835
rect 28615 1815 28635 1835
rect 28665 1815 28685 1835
rect 28715 1815 28735 1835
rect 28765 1815 28785 1835
rect -635 -1885 -615 -1865
rect -585 -1885 -565 -1865
rect -535 -1885 -515 -1865
rect -485 -1885 -465 -1865
rect -435 -1885 -415 -1865
rect -385 -1885 -365 -1865
rect -335 -1885 -315 -1865
rect -285 -1885 -265 -1865
rect -235 -1885 -215 -1865
rect -185 -1885 -165 -1865
rect -135 -1885 -115 -1865
rect -85 -1885 -65 -1865
rect -35 -1885 -15 -1865
rect 15 -1885 35 -1865
rect 65 -1885 85 -1865
rect 115 -1885 135 -1865
rect 165 -1885 185 -1865
rect 215 -1885 235 -1865
rect 265 -1885 285 -1865
rect 315 -1885 335 -1865
rect 365 -1885 385 -1865
rect 415 -1885 435 -1865
rect 465 -1885 485 -1865
rect 515 -1885 535 -1865
rect 565 -1885 585 -1865
rect 615 -1885 635 -1865
rect 665 -1885 685 -1865
rect 715 -1885 735 -1865
rect 765 -1885 785 -1865
rect 815 -1885 835 -1865
rect 865 -1885 885 -1865
rect 915 -1885 935 -1865
rect 965 -1885 985 -1865
rect 1015 -1885 1035 -1865
rect 1065 -1885 1085 -1865
rect 1115 -1885 1135 -1865
rect 1165 -1885 1185 -1865
rect 1215 -1885 1235 -1865
rect 1265 -1885 1285 -1865
rect 1315 -1885 1335 -1865
rect 1365 -1885 1385 -1865
rect 1415 -1885 1435 -1865
rect 1465 -1885 1485 -1865
rect 1515 -1885 1535 -1865
rect 1565 -1885 1585 -1865
rect 1615 -1885 1635 -1865
rect 1665 -1885 1685 -1865
rect 1715 -1885 1735 -1865
rect 1765 -1885 1785 -1865
rect 1815 -1885 1835 -1865
rect 1865 -1885 1885 -1865
rect 1915 -1885 1935 -1865
rect 1965 -1885 1985 -1865
rect 2015 -1885 2035 -1865
rect 2065 -1885 2085 -1865
rect 2115 -1885 2135 -1865
rect 2165 -1885 2185 -1865
rect 2215 -1885 2235 -1865
rect 2265 -1885 2285 -1865
rect 2315 -1885 2335 -1865
rect 2365 -1885 2385 -1865
rect 2415 -1885 2435 -1865
rect 2465 -1885 2485 -1865
rect 2515 -1885 2535 -1865
rect 2565 -1885 2585 -1865
rect 2615 -1885 2635 -1865
rect 2665 -1885 2685 -1865
rect 2715 -1885 2735 -1865
rect 2765 -1885 2785 -1865
rect 2815 -1885 2835 -1865
rect 2865 -1885 2885 -1865
rect 2915 -1885 2935 -1865
rect 2965 -1885 2985 -1865
rect 3015 -1885 3035 -1865
rect 3065 -1885 3085 -1865
rect 3115 -1885 3135 -1865
rect 3165 -1885 3185 -1865
rect 3215 -1885 3235 -1865
rect 3265 -1885 3285 -1865
rect 3315 -1885 3335 -1865
rect 3365 -1885 3385 -1865
rect 3415 -1885 3435 -1865
rect 3465 -1885 3485 -1865
rect 3515 -1885 3535 -1865
rect 3565 -1885 3585 -1865
rect 3615 -1885 3635 -1865
rect 3665 -1885 3685 -1865
rect 3715 -1885 3735 -1865
rect 3765 -1885 3785 -1865
rect 3815 -1885 3835 -1865
rect 3865 -1885 3885 -1865
rect 3915 -1885 3935 -1865
rect 3965 -1885 3985 -1865
rect 4015 -1885 4035 -1865
rect 4065 -1885 4085 -1865
rect 4115 -1885 4135 -1865
rect 4165 -1885 4185 -1865
rect 4215 -1885 4235 -1865
rect 4265 -1885 4285 -1865
rect 4315 -1885 4335 -1865
rect 4365 -1885 4385 -1865
rect 4415 -1885 4435 -1865
rect 4465 -1885 4485 -1865
rect 4515 -1885 4535 -1865
rect 4565 -1885 4585 -1865
rect 4615 -1885 4635 -1865
rect 4665 -1885 4685 -1865
rect 4715 -1885 4735 -1865
rect 4765 -1885 4785 -1865
rect 4815 -1885 4835 -1865
rect 4865 -1885 4885 -1865
rect 4915 -1885 4935 -1865
rect 4965 -1885 4985 -1865
rect 5015 -1885 5035 -1865
rect 5065 -1885 5085 -1865
rect 5115 -1885 5135 -1865
rect 5165 -1885 5185 -1865
rect 5215 -1885 5235 -1865
rect 5265 -1885 5285 -1865
rect 5315 -1885 5335 -1865
rect 5365 -1885 5385 -1865
rect 5415 -1885 5435 -1865
rect 5465 -1885 5485 -1865
rect 5515 -1885 5535 -1865
rect 5565 -1885 5585 -1865
rect 5615 -1885 5635 -1865
rect 5665 -1885 5685 -1865
rect 5715 -1885 5735 -1865
rect 5765 -1885 5785 -1865
rect 5815 -1885 5835 -1865
rect 5865 -1885 5885 -1865
rect 5915 -1885 5935 -1865
rect 5965 -1885 5985 -1865
rect 6015 -1885 6035 -1865
rect 6065 -1885 6085 -1865
rect 6115 -1885 6135 -1865
rect 6165 -1885 6185 -1865
rect 6215 -1885 6235 -1865
rect 6265 -1885 6285 -1865
rect 6315 -1885 6335 -1865
rect 6365 -1885 6385 -1865
rect 6415 -1885 6435 -1865
rect 6465 -1885 6485 -1865
rect 6515 -1885 6535 -1865
rect 6565 -1885 6585 -1865
rect 6615 -1885 6635 -1865
rect 6665 -1885 6685 -1865
rect 6715 -1885 6735 -1865
rect 6765 -1885 6785 -1865
rect 6815 -1885 6835 -1865
rect 6865 -1885 6885 -1865
rect 6915 -1885 6935 -1865
rect 6965 -1885 6985 -1865
rect 7015 -1885 7035 -1865
rect 7065 -1885 7085 -1865
rect 7115 -1885 7135 -1865
rect 7165 -1885 7185 -1865
rect 7215 -1885 7235 -1865
rect 7265 -1885 7285 -1865
rect 7315 -1885 7335 -1865
rect 7365 -1885 7385 -1865
rect 7415 -1885 7435 -1865
rect 7465 -1885 7485 -1865
rect 7515 -1885 7535 -1865
rect 7565 -1885 7585 -1865
rect 7615 -1885 7635 -1865
rect 7665 -1885 7685 -1865
rect 7715 -1885 7735 -1865
rect 7765 -1885 7785 -1865
rect 7815 -1885 7835 -1865
rect 7865 -1885 7885 -1865
rect 7915 -1885 7935 -1865
rect 7965 -1885 7985 -1865
rect 8015 -1885 8035 -1865
rect 8065 -1885 8085 -1865
rect 8115 -1885 8135 -1865
rect 8165 -1885 8185 -1865
rect 8215 -1885 8235 -1865
rect 8265 -1885 8285 -1865
rect 8315 -1885 8335 -1865
rect 8365 -1885 8385 -1865
rect 8415 -1885 8435 -1865
rect 8465 -1885 8485 -1865
rect 8515 -1885 8535 -1865
rect 8565 -1885 8585 -1865
rect 8615 -1885 8635 -1865
rect 8665 -1885 8685 -1865
rect 8715 -1885 8735 -1865
rect 8765 -1885 8785 -1865
rect 8815 -1885 8835 -1865
rect 8865 -1885 8885 -1865
rect 8915 -1885 8935 -1865
rect 8965 -1885 8985 -1865
rect 9015 -1885 9035 -1865
rect 9065 -1885 9085 -1865
rect 9115 -1885 9135 -1865
rect 9165 -1885 9185 -1865
rect 9215 -1885 9235 -1865
rect 9265 -1885 9285 -1865
rect 9315 -1885 9335 -1865
rect 9365 -1885 9385 -1865
rect 9415 -1885 9435 -1865
rect 9465 -1885 9485 -1865
rect 9515 -1885 9535 -1865
rect 9565 -1885 9585 -1865
rect 9615 -1885 9635 -1865
rect 9665 -1885 9685 -1865
rect 9715 -1885 9735 -1865
rect 9765 -1885 9785 -1865
rect 9815 -1885 9835 -1865
rect 9865 -1885 9885 -1865
rect 9915 -1885 9935 -1865
rect 9965 -1885 9985 -1865
rect 10015 -1885 10035 -1865
rect 10065 -1885 10085 -1865
rect 10115 -1885 10135 -1865
rect 10165 -1885 10185 -1865
rect 10215 -1885 10235 -1865
rect 10265 -1885 10285 -1865
rect 10315 -1885 10335 -1865
rect 10365 -1885 10385 -1865
rect 10415 -1885 10435 -1865
rect 10465 -1885 10485 -1865
rect 10515 -1885 10535 -1865
rect 10565 -1885 10585 -1865
rect 10615 -1885 10635 -1865
rect 10665 -1885 10685 -1865
rect 10715 -1885 10735 -1865
rect 10765 -1885 10785 -1865
rect 10815 -1885 10835 -1865
rect 10865 -1885 10885 -1865
rect 10915 -1885 10935 -1865
rect 10965 -1885 10985 -1865
rect 11015 -1885 11035 -1865
rect 11065 -1885 11085 -1865
rect 11115 -1885 11135 -1865
rect 11165 -1885 11185 -1865
rect 11215 -1885 11235 -1865
rect 11265 -1885 11285 -1865
rect 11315 -1885 11335 -1865
rect 11365 -1885 11385 -1865
rect 11415 -1885 11435 -1865
rect 11465 -1885 11485 -1865
rect 11515 -1885 11535 -1865
rect 11565 -1885 11585 -1865
rect 11615 -1885 11635 -1865
rect 11665 -1885 11685 -1865
rect 11715 -1885 11735 -1865
rect 11765 -1885 11785 -1865
rect 11815 -1885 11835 -1865
rect 11865 -1885 11885 -1865
rect 11915 -1885 11935 -1865
rect 11965 -1885 11985 -1865
rect 12015 -1885 12035 -1865
rect 12065 -1885 12085 -1865
rect 12115 -1885 12135 -1865
rect 12165 -1885 12185 -1865
rect 12215 -1885 12235 -1865
rect 12265 -1885 12285 -1865
rect 12315 -1885 12335 -1865
rect 12365 -1885 12385 -1865
rect 12415 -1885 12435 -1865
rect 12465 -1885 12485 -1865
rect 12515 -1885 12535 -1865
rect 12565 -1885 12585 -1865
rect 12615 -1885 12635 -1865
rect 12665 -1885 12685 -1865
rect 12715 -1885 12735 -1865
rect 12765 -1885 12785 -1865
rect 12815 -1885 12835 -1865
rect 12865 -1885 12885 -1865
rect 12915 -1885 12935 -1865
rect 12965 -1885 12985 -1865
rect 13015 -1885 13035 -1865
rect 13065 -1885 13085 -1865
rect 13115 -1885 13135 -1865
rect 13165 -1885 13185 -1865
rect 13215 -1885 13235 -1865
rect 13265 -1885 13285 -1865
rect 13315 -1885 13335 -1865
rect 13365 -1885 13385 -1865
rect 13415 -1885 13435 -1865
rect 13465 -1885 13485 -1865
rect 13515 -1885 13535 -1865
rect 13565 -1885 13585 -1865
rect 13615 -1885 13635 -1865
rect 13665 -1885 13685 -1865
rect 13715 -1885 13735 -1865
rect 13765 -1885 13785 -1865
rect 13815 -1885 13835 -1865
rect 13865 -1885 13885 -1865
rect 13915 -1885 13935 -1865
rect 13965 -1885 13985 -1865
rect 14015 -1885 14035 -1865
rect 14065 -1885 14085 -1865
rect 14115 -1885 14135 -1865
rect 14165 -1885 14185 -1865
rect 14215 -1885 14235 -1865
rect 14265 -1885 14285 -1865
rect 14315 -1885 14335 -1865
rect 14365 -1885 14385 -1865
rect 14415 -1885 14435 -1865
rect 14465 -1885 14485 -1865
rect 14515 -1885 14535 -1865
rect 14565 -1885 14585 -1865
rect 14615 -1885 14635 -1865
rect 14665 -1885 14685 -1865
rect 14715 -1885 14735 -1865
rect 14765 -1885 14785 -1865
rect 14815 -1885 14835 -1865
rect 14865 -1885 14885 -1865
rect 14915 -1885 14935 -1865
rect 14965 -1885 14985 -1865
rect 15015 -1885 15035 -1865
rect 15065 -1885 15085 -1865
rect 15115 -1885 15135 -1865
rect 15165 -1885 15185 -1865
rect 15215 -1885 15235 -1865
rect 15265 -1885 15285 -1865
rect 15315 -1885 15335 -1865
rect 15365 -1885 15385 -1865
rect 15415 -1885 15435 -1865
rect 15465 -1885 15485 -1865
rect 15515 -1885 15535 -1865
rect 15565 -1885 15585 -1865
rect 15615 -1885 15635 -1865
rect 15665 -1885 15685 -1865
rect 15715 -1885 15735 -1865
rect 15765 -1885 15785 -1865
rect 15815 -1885 15835 -1865
rect 15865 -1885 15885 -1865
rect 15915 -1885 15935 -1865
rect 15965 -1885 15985 -1865
rect 16015 -1885 16035 -1865
rect 16065 -1885 16085 -1865
rect 16115 -1885 16135 -1865
rect 16165 -1885 16185 -1865
rect 16215 -1885 16235 -1865
rect 16265 -1885 16285 -1865
rect 16315 -1885 16335 -1865
rect 16365 -1885 16385 -1865
rect 16415 -1885 16435 -1865
rect 16465 -1885 16485 -1865
rect 16515 -1885 16535 -1865
rect 16565 -1885 16585 -1865
rect 16615 -1885 16635 -1865
rect 16665 -1885 16685 -1865
rect 16715 -1885 16735 -1865
rect 16765 -1885 16785 -1865
rect 16815 -1885 16835 -1865
rect 16865 -1885 16885 -1865
rect 16915 -1885 16935 -1865
rect 16965 -1885 16985 -1865
rect 17015 -1885 17035 -1865
rect 17065 -1885 17085 -1865
rect 17115 -1885 17135 -1865
rect 17165 -1885 17185 -1865
rect 17215 -1885 17235 -1865
rect 17265 -1885 17285 -1865
rect 17315 -1885 17335 -1865
rect 17365 -1885 17385 -1865
rect 17415 -1885 17435 -1865
rect 17465 -1885 17485 -1865
rect 17515 -1885 17535 -1865
rect 17565 -1885 17585 -1865
rect 17615 -1885 17635 -1865
rect 17665 -1885 17685 -1865
rect 17715 -1885 17735 -1865
rect 17765 -1885 17785 -1865
rect 17815 -1885 17835 -1865
rect 17865 -1885 17885 -1865
rect 17915 -1885 17935 -1865
rect 17965 -1885 17985 -1865
rect 18015 -1885 18035 -1865
rect 18065 -1885 18085 -1865
rect 18115 -1885 18135 -1865
rect 18165 -1885 18185 -1865
rect 18215 -1885 18235 -1865
rect 18265 -1885 18285 -1865
rect 18315 -1885 18335 -1865
rect 18365 -1885 18385 -1865
rect 18415 -1885 18435 -1865
rect 18465 -1885 18485 -1865
rect 18515 -1885 18535 -1865
rect 18565 -1885 18585 -1865
rect 18615 -1885 18635 -1865
rect 18665 -1885 18685 -1865
rect 18715 -1885 18735 -1865
rect 18765 -1885 18785 -1865
rect 18815 -1885 18835 -1865
rect 18865 -1885 18885 -1865
rect 18915 -1885 18935 -1865
rect 18965 -1885 18985 -1865
rect 19015 -1885 19035 -1865
rect 19065 -1885 19085 -1865
rect 19115 -1885 19135 -1865
rect 19165 -1885 19185 -1865
rect 19215 -1885 19235 -1865
rect 19265 -1885 19285 -1865
rect 19315 -1885 19335 -1865
rect 19365 -1885 19385 -1865
rect 19415 -1885 19435 -1865
rect 19465 -1885 19485 -1865
rect 19515 -1885 19535 -1865
rect 19565 -1885 19585 -1865
rect 19615 -1885 19635 -1865
rect 19665 -1885 19685 -1865
rect 19715 -1885 19735 -1865
rect 19765 -1885 19785 -1865
rect 19815 -1885 19835 -1865
rect 19865 -1885 19885 -1865
rect 19915 -1885 19935 -1865
rect 19965 -1885 19985 -1865
rect 20015 -1885 20035 -1865
rect 20065 -1885 20085 -1865
rect 20115 -1885 20135 -1865
rect 20165 -1885 20185 -1865
rect 20215 -1885 20235 -1865
rect 20265 -1885 20285 -1865
rect 20315 -1885 20335 -1865
rect 20365 -1885 20385 -1865
rect 20415 -1885 20435 -1865
rect 20465 -1885 20485 -1865
rect 20515 -1885 20535 -1865
rect 20565 -1885 20585 -1865
rect 20615 -1885 20635 -1865
rect 20665 -1885 20685 -1865
rect 20715 -1885 20735 -1865
rect 20765 -1885 20785 -1865
rect 20815 -1885 20835 -1865
rect 20865 -1885 20885 -1865
rect 20915 -1885 20935 -1865
rect 20965 -1885 20985 -1865
rect 21015 -1885 21035 -1865
rect 21065 -1885 21085 -1865
rect 21115 -1885 21135 -1865
rect 21165 -1885 21185 -1865
rect 21215 -1885 21235 -1865
rect 21265 -1885 21285 -1865
rect 21315 -1885 21335 -1865
rect 21365 -1885 21385 -1865
rect 21415 -1885 21435 -1865
rect 21465 -1885 21485 -1865
rect 21515 -1885 21535 -1865
rect 21565 -1885 21585 -1865
rect 21615 -1885 21635 -1865
rect 21665 -1885 21685 -1865
rect 21715 -1885 21735 -1865
rect 21765 -1885 21785 -1865
rect 21815 -1885 21835 -1865
rect 21865 -1885 21885 -1865
rect 21915 -1885 21935 -1865
rect 21965 -1885 21985 -1865
rect 22015 -1885 22035 -1865
rect 22065 -1885 22085 -1865
rect 22115 -1885 22135 -1865
rect 22165 -1885 22185 -1865
rect 22215 -1885 22235 -1865
rect 22265 -1885 22285 -1865
rect 22315 -1885 22335 -1865
rect 22365 -1885 22385 -1865
rect 22415 -1885 22435 -1865
rect 22465 -1885 22485 -1865
rect 22515 -1885 22535 -1865
rect 22565 -1885 22585 -1865
rect 22615 -1885 22635 -1865
rect 22665 -1885 22685 -1865
rect 22715 -1885 22735 -1865
rect 22765 -1885 22785 -1865
rect 22815 -1885 22835 -1865
rect 22865 -1885 22885 -1865
rect 22915 -1885 22935 -1865
rect 22965 -1885 22985 -1865
rect 23015 -1885 23035 -1865
rect 23065 -1885 23085 -1865
rect 23115 -1885 23135 -1865
rect 23165 -1885 23185 -1865
rect 23215 -1885 23235 -1865
rect 23265 -1885 23285 -1865
rect 23315 -1885 23335 -1865
rect 23365 -1885 23385 -1865
rect 23415 -1885 23435 -1865
rect 23465 -1885 23485 -1865
rect 23515 -1885 23535 -1865
rect 23565 -1885 23585 -1865
rect 23615 -1885 23635 -1865
rect 23665 -1885 23685 -1865
rect 23715 -1885 23735 -1865
rect 23765 -1885 23785 -1865
rect 23815 -1885 23835 -1865
rect 23865 -1885 23885 -1865
rect 23915 -1885 23935 -1865
rect 23965 -1885 23985 -1865
rect 24015 -1885 24035 -1865
rect 24065 -1885 24085 -1865
rect 24115 -1885 24135 -1865
rect 24165 -1885 24185 -1865
rect 24215 -1885 24235 -1865
rect 24265 -1885 24285 -1865
rect 24315 -1885 24335 -1865
rect 24365 -1885 24385 -1865
rect 24415 -1885 24435 -1865
rect 24465 -1885 24485 -1865
rect 24515 -1885 24535 -1865
rect 24565 -1885 24585 -1865
rect 24615 -1885 24635 -1865
rect 24665 -1885 24685 -1865
rect 24715 -1885 24735 -1865
rect 24765 -1885 24785 -1865
rect 24815 -1885 24835 -1865
rect 24865 -1885 24885 -1865
rect 24915 -1885 24935 -1865
rect 24965 -1885 24985 -1865
rect 25015 -1885 25035 -1865
rect 25065 -1885 25085 -1865
rect 25115 -1885 25135 -1865
rect 25165 -1885 25185 -1865
rect 25215 -1885 25235 -1865
rect 25265 -1885 25285 -1865
rect 25315 -1885 25335 -1865
rect 25365 -1885 25385 -1865
rect 25415 -1885 25435 -1865
rect 25465 -1885 25485 -1865
rect 25515 -1885 25535 -1865
rect 25565 -1885 25585 -1865
rect 25615 -1885 25635 -1865
rect 25665 -1885 25685 -1865
rect 25715 -1885 25735 -1865
rect 25765 -1885 25785 -1865
rect 25815 -1885 25835 -1865
rect 25865 -1885 25885 -1865
rect 25915 -1885 25935 -1865
rect 25965 -1885 25985 -1865
rect 26015 -1885 26035 -1865
rect 26065 -1885 26085 -1865
rect 26115 -1885 26135 -1865
rect 26165 -1885 26185 -1865
rect 26215 -1885 26235 -1865
rect 26265 -1885 26285 -1865
rect 26315 -1885 26335 -1865
rect 26365 -1885 26385 -1865
rect 26415 -1885 26435 -1865
rect 26465 -1885 26485 -1865
rect 26515 -1885 26535 -1865
rect 26565 -1885 26585 -1865
rect 26615 -1885 26635 -1865
rect 26665 -1885 26685 -1865
rect 26715 -1885 26735 -1865
rect 26765 -1885 26785 -1865
rect 26815 -1885 26835 -1865
rect 26865 -1885 26885 -1865
rect 26915 -1885 26935 -1865
rect 26965 -1885 26985 -1865
rect 27015 -1885 27035 -1865
rect 27065 -1885 27085 -1865
rect 27115 -1885 27135 -1865
rect 27165 -1885 27185 -1865
rect 27215 -1885 27235 -1865
rect 27265 -1885 27285 -1865
rect 27315 -1885 27335 -1865
rect 27365 -1885 27385 -1865
rect 27415 -1885 27435 -1865
rect 27465 -1885 27485 -1865
rect 27515 -1885 27535 -1865
rect 27565 -1885 27585 -1865
rect 27615 -1885 27635 -1865
rect 27665 -1885 27685 -1865
rect 27715 -1885 27735 -1865
rect 27765 -1885 27785 -1865
rect 27815 -1885 27835 -1865
rect 27865 -1885 27885 -1865
rect 27915 -1885 27935 -1865
rect 27965 -1885 27985 -1865
rect 28015 -1885 28035 -1865
rect 28065 -1885 28085 -1865
rect 28115 -1885 28135 -1865
rect 28165 -1885 28185 -1865
rect 28215 -1885 28235 -1865
rect 28265 -1885 28285 -1865
rect 28315 -1885 28335 -1865
rect 28365 -1885 28385 -1865
rect 28415 -1885 28435 -1865
rect 28465 -1885 28485 -1865
rect 28515 -1885 28535 -1865
rect 28565 -1885 28585 -1865
rect 28615 -1885 28635 -1865
rect 28665 -1885 28685 -1865
rect 28715 -1885 28735 -1865
rect 28765 -1885 28785 -1865
<< poly >>
rect -600 5500 -500 5515
rect -450 5500 -350 5515
rect -300 5500 -200 5515
rect -150 5500 -50 5515
rect 0 5500 100 5515
rect 150 5500 250 5515
rect 300 5500 400 5515
rect 450 5500 550 5515
rect 600 5500 700 5515
rect 750 5500 850 5515
rect 900 5500 1000 5515
rect 1050 5500 1150 5515
rect 1200 5500 1300 5515
rect 1350 5500 1450 5515
rect 1500 5500 1600 5515
rect 1650 5500 1750 5515
rect 1800 5500 1900 5515
rect 1950 5500 2050 5515
rect 2100 5500 2200 5515
rect 2250 5500 2350 5515
rect 2400 5500 2500 5515
rect 2550 5500 2650 5515
rect 2700 5500 2800 5515
rect 2850 5500 2950 5515
rect 3000 5500 3100 5515
rect 3150 5500 3250 5515
rect 3300 5500 3400 5515
rect 3450 5500 3550 5515
rect 3600 5500 3700 5515
rect 3750 5500 3850 5515
rect 3900 5500 4000 5515
rect 4050 5500 4150 5515
rect 4200 5500 4300 5515
rect 4350 5500 4450 5515
rect 4500 5500 4600 5515
rect 4650 5500 4750 5515
rect 4800 5500 4900 5515
rect 4950 5500 5050 5515
rect 5100 5500 5200 5515
rect 5250 5500 5350 5515
rect 5400 5500 5500 5515
rect 5550 5500 5650 5515
rect 5700 5500 5800 5515
rect 5850 5500 5950 5515
rect 6000 5500 6100 5515
rect 6150 5500 6250 5515
rect 6300 5500 6400 5515
rect 6450 5500 6550 5515
rect 6600 5500 6700 5515
rect 6750 5500 6850 5515
rect 6900 5500 7000 5515
rect 7050 5500 7150 5515
rect 7200 5500 7300 5515
rect 7350 5500 7450 5515
rect 7500 5500 7600 5515
rect 7650 5500 7750 5515
rect 7800 5500 7900 5515
rect 7950 5500 8050 5515
rect 8100 5500 8200 5515
rect 8250 5500 8350 5515
rect 8400 5500 8500 5515
rect 8550 5500 8650 5515
rect 8700 5500 8800 5515
rect 8850 5500 8950 5515
rect 9000 5500 9100 5515
rect 9150 5500 9250 5515
rect 9300 5500 9400 5515
rect 9450 5500 9550 5515
rect 9600 5500 9700 5515
rect 9750 5500 9850 5515
rect 9900 5500 10000 5515
rect 10050 5500 10150 5515
rect 10200 5500 10300 5515
rect 10350 5500 10450 5515
rect 10500 5500 10600 5515
rect 10650 5500 10750 5515
rect 10800 5500 10900 5515
rect 10950 5500 11050 5515
rect 11100 5500 11200 5515
rect 11250 5500 11350 5515
rect 11400 5500 11500 5515
rect 11550 5500 11650 5515
rect 11700 5500 11800 5515
rect 11850 5500 11950 5515
rect 12000 5500 12100 5515
rect 12150 5500 12250 5515
rect 12300 5500 12400 5515
rect 12450 5500 12550 5515
rect 12600 5500 12700 5515
rect 12750 5500 12850 5515
rect 12900 5500 13000 5515
rect 13050 5500 13150 5515
rect 13200 5500 13300 5515
rect 13350 5500 13450 5515
rect 13500 5500 13600 5515
rect 13650 5500 13750 5515
rect 13800 5500 13900 5515
rect 13950 5500 14050 5515
rect 14100 5500 14200 5515
rect 14250 5500 14350 5515
rect 14400 5500 14500 5515
rect 14550 5500 14650 5515
rect 14700 5500 14800 5515
rect 14850 5500 14950 5515
rect 15000 5500 15100 5515
rect 15150 5500 15250 5515
rect 15300 5500 15400 5515
rect 15450 5500 15550 5515
rect 15600 5500 15700 5515
rect 15750 5500 15850 5515
rect 15900 5500 16000 5515
rect 16050 5500 16150 5515
rect 16200 5500 16300 5515
rect 16350 5500 16450 5515
rect 16500 5500 16600 5515
rect 16650 5500 16750 5515
rect 16800 5500 16900 5515
rect 16950 5500 17050 5515
rect 17100 5500 17200 5515
rect 17250 5500 17350 5515
rect 17400 5500 17500 5515
rect 17550 5500 17650 5515
rect 17700 5500 17800 5515
rect 17850 5500 17950 5515
rect 18000 5500 18100 5515
rect 18150 5500 18250 5515
rect 18300 5500 18400 5515
rect 18450 5500 18550 5515
rect 18600 5500 18700 5515
rect 18750 5500 18850 5515
rect 18900 5500 19000 5515
rect 19050 5500 19150 5515
rect 19200 5500 19300 5515
rect 19350 5500 19450 5515
rect 19500 5500 19600 5515
rect 19650 5500 19750 5515
rect 19800 5500 19900 5515
rect 19950 5500 20050 5515
rect 20100 5500 20200 5515
rect 20250 5500 20350 5515
rect 20400 5500 20500 5515
rect 20550 5500 20650 5515
rect 20700 5500 20800 5515
rect 20850 5500 20950 5515
rect 21000 5500 21100 5515
rect 21150 5500 21250 5515
rect 21300 5500 21400 5515
rect 21450 5500 21550 5515
rect 21600 5500 21700 5515
rect 21750 5500 21850 5515
rect 21900 5500 22000 5515
rect 22050 5500 22150 5515
rect 22200 5500 22300 5515
rect 22350 5500 22450 5515
rect 22500 5500 22600 5515
rect 22650 5500 22750 5515
rect 22800 5500 22900 5515
rect 22950 5500 23050 5515
rect 23100 5500 23200 5515
rect 23250 5500 23350 5515
rect 23400 5500 23500 5515
rect 23550 5500 23650 5515
rect 23700 5500 23800 5515
rect 23850 5500 23950 5515
rect 24000 5500 24100 5515
rect 24150 5500 24250 5515
rect 24300 5500 24400 5515
rect 24450 5500 24550 5515
rect 24600 5500 24700 5515
rect 24750 5500 24850 5515
rect 24900 5500 25000 5515
rect 25050 5500 25150 5515
rect 25200 5500 25300 5515
rect 25350 5500 25450 5515
rect 25500 5500 25600 5515
rect 25650 5500 25750 5515
rect 25800 5500 25900 5515
rect 25950 5500 26050 5515
rect 26100 5500 26200 5515
rect 26250 5500 26350 5515
rect 26400 5500 26500 5515
rect 26550 5500 26650 5515
rect 26700 5500 26800 5515
rect 26850 5500 26950 5515
rect 27000 5500 27100 5515
rect 27150 5500 27250 5515
rect 27300 5500 27400 5515
rect 27450 5500 27550 5515
rect 27600 5500 27700 5515
rect 27750 5500 27850 5515
rect 27900 5500 28000 5515
rect 28050 5500 28150 5515
rect 28200 5500 28300 5515
rect 28350 5500 28450 5515
rect 28500 5500 28600 5515
rect 28650 5500 28750 5515
rect 28800 5500 28900 5515
rect 28950 5500 29050 5515
rect 29100 5500 29200 5515
rect 29250 5500 29350 5515
rect 29400 5500 29500 5515
rect 29550 5500 29650 5515
rect 29700 5500 29800 5515
rect 29850 5500 29950 5515
rect 30000 5500 30100 5515
rect 30150 5500 30250 5515
rect 30300 5500 30400 5515
rect 30450 5500 30550 5515
rect 30600 5500 30700 5515
rect 30750 5500 30850 5515
rect 30900 5500 31000 5515
rect 31050 5500 31150 5515
rect 31200 5500 31300 5515
rect 31350 5500 31450 5515
rect 31500 5500 31600 5515
rect 31650 5500 31750 5515
rect 31800 5500 31900 5515
rect 31950 5500 32050 5515
rect -600 4950 -500 5000
rect -450 4950 -350 5000
rect -600 4935 -350 4950
rect -600 4915 -585 4935
rect -565 4915 -535 4935
rect -515 4915 -485 4935
rect -465 4915 -435 4935
rect -415 4915 -385 4935
rect -365 4915 -350 4935
rect -600 4900 -350 4915
rect -600 4850 -500 4900
rect -450 4850 -350 4900
rect -300 4950 -200 5000
rect -150 4950 -50 5000
rect -300 4935 -50 4950
rect -300 4915 -285 4935
rect -265 4915 -235 4935
rect -215 4915 -185 4935
rect -165 4915 -135 4935
rect -115 4915 -85 4935
rect -65 4915 -50 4935
rect -300 4900 -50 4915
rect -300 4850 -200 4900
rect -150 4850 -50 4900
rect 0 4950 100 5000
rect 150 4950 250 5000
rect 0 4935 250 4950
rect 0 4915 15 4935
rect 35 4915 65 4935
rect 85 4915 115 4935
rect 135 4915 165 4935
rect 185 4915 215 4935
rect 235 4915 250 4935
rect 0 4900 250 4915
rect 0 4850 100 4900
rect 150 4850 250 4900
rect 300 4950 400 5000
rect 450 4950 550 5000
rect 300 4935 550 4950
rect 300 4915 315 4935
rect 335 4915 365 4935
rect 385 4915 415 4935
rect 435 4915 465 4935
rect 485 4915 515 4935
rect 535 4915 550 4935
rect 300 4900 550 4915
rect 300 4850 400 4900
rect 450 4850 550 4900
rect 600 4950 700 5000
rect 750 4950 850 5000
rect 600 4935 850 4950
rect 600 4915 615 4935
rect 635 4915 665 4935
rect 685 4915 715 4935
rect 735 4915 765 4935
rect 785 4915 815 4935
rect 835 4915 850 4935
rect 600 4900 850 4915
rect 600 4850 700 4900
rect 750 4850 850 4900
rect 900 4950 1000 5000
rect 1050 4950 1150 5000
rect 900 4935 1150 4950
rect 900 4915 915 4935
rect 935 4915 965 4935
rect 985 4915 1015 4935
rect 1035 4915 1065 4935
rect 1085 4915 1115 4935
rect 1135 4915 1150 4935
rect 900 4900 1150 4915
rect 900 4850 1000 4900
rect 1050 4850 1150 4900
rect 1200 4950 1300 5000
rect 1350 4950 1450 5000
rect 1200 4935 1450 4950
rect 1200 4915 1215 4935
rect 1235 4915 1265 4935
rect 1285 4915 1315 4935
rect 1335 4915 1365 4935
rect 1385 4915 1415 4935
rect 1435 4915 1450 4935
rect 1200 4900 1450 4915
rect 1200 4850 1300 4900
rect 1350 4850 1450 4900
rect 1500 4950 1600 5000
rect 1650 4950 1750 5000
rect 1500 4935 1750 4950
rect 1500 4915 1515 4935
rect 1535 4915 1565 4935
rect 1585 4915 1615 4935
rect 1635 4915 1665 4935
rect 1685 4915 1715 4935
rect 1735 4915 1750 4935
rect 1500 4900 1750 4915
rect 1500 4850 1600 4900
rect 1650 4850 1750 4900
rect 1800 4950 1900 5000
rect 1950 4950 2050 5000
rect 1800 4935 2050 4950
rect 1800 4915 1815 4935
rect 1835 4915 1865 4935
rect 1885 4915 1915 4935
rect 1935 4915 1965 4935
rect 1985 4915 2015 4935
rect 2035 4915 2050 4935
rect 1800 4900 2050 4915
rect 1800 4850 1900 4900
rect 1950 4850 2050 4900
rect 2100 4950 2200 5000
rect 2250 4950 2350 5000
rect 2100 4935 2350 4950
rect 2100 4915 2115 4935
rect 2135 4915 2165 4935
rect 2185 4915 2215 4935
rect 2235 4915 2265 4935
rect 2285 4915 2315 4935
rect 2335 4915 2350 4935
rect 2100 4900 2350 4915
rect 2100 4850 2200 4900
rect 2250 4850 2350 4900
rect 2400 4950 2500 5000
rect 2550 4950 2650 5000
rect 2400 4935 2650 4950
rect 2400 4915 2415 4935
rect 2435 4915 2465 4935
rect 2485 4915 2515 4935
rect 2535 4915 2565 4935
rect 2585 4915 2615 4935
rect 2635 4915 2650 4935
rect 2400 4900 2650 4915
rect 2400 4850 2500 4900
rect 2550 4850 2650 4900
rect 2700 4950 2800 5000
rect 2850 4950 2950 5000
rect 2700 4935 2950 4950
rect 2700 4915 2715 4935
rect 2735 4915 2765 4935
rect 2785 4915 2815 4935
rect 2835 4915 2865 4935
rect 2885 4915 2915 4935
rect 2935 4915 2950 4935
rect 2700 4900 2950 4915
rect 2700 4850 2800 4900
rect 2850 4850 2950 4900
rect 3000 4950 3100 5000
rect 3150 4950 3250 5000
rect 3000 4935 3250 4950
rect 3000 4915 3015 4935
rect 3035 4915 3065 4935
rect 3085 4915 3115 4935
rect 3135 4915 3165 4935
rect 3185 4915 3215 4935
rect 3235 4915 3250 4935
rect 3000 4900 3250 4915
rect 3000 4850 3100 4900
rect 3150 4850 3250 4900
rect 3300 4950 3400 5000
rect 3450 4950 3550 5000
rect 3300 4935 3550 4950
rect 3300 4915 3315 4935
rect 3335 4915 3365 4935
rect 3385 4915 3415 4935
rect 3435 4915 3465 4935
rect 3485 4915 3515 4935
rect 3535 4915 3550 4935
rect 3300 4900 3550 4915
rect 3300 4850 3400 4900
rect 3450 4850 3550 4900
rect 3600 4950 3700 5000
rect 3750 4950 3850 5000
rect 3600 4935 3850 4950
rect 3600 4915 3615 4935
rect 3635 4915 3665 4935
rect 3685 4915 3715 4935
rect 3735 4915 3765 4935
rect 3785 4915 3815 4935
rect 3835 4915 3850 4935
rect 3600 4900 3850 4915
rect 3600 4850 3700 4900
rect 3750 4850 3850 4900
rect 3900 4950 4000 5000
rect 4050 4950 4150 5000
rect 3900 4935 4150 4950
rect 3900 4915 3915 4935
rect 3935 4915 3965 4935
rect 3985 4915 4015 4935
rect 4035 4915 4065 4935
rect 4085 4915 4115 4935
rect 4135 4915 4150 4935
rect 3900 4900 4150 4915
rect 3900 4850 4000 4900
rect 4050 4850 4150 4900
rect 4200 4950 4300 5000
rect 4350 4950 4450 5000
rect 4200 4935 4450 4950
rect 4200 4915 4215 4935
rect 4235 4915 4265 4935
rect 4285 4915 4315 4935
rect 4335 4915 4365 4935
rect 4385 4915 4415 4935
rect 4435 4915 4450 4935
rect 4200 4900 4450 4915
rect 4200 4850 4300 4900
rect 4350 4850 4450 4900
rect 4500 4950 4600 5000
rect 4650 4950 4750 5000
rect 4500 4935 4750 4950
rect 4500 4915 4515 4935
rect 4535 4915 4565 4935
rect 4585 4915 4615 4935
rect 4635 4915 4665 4935
rect 4685 4915 4715 4935
rect 4735 4915 4750 4935
rect 4500 4900 4750 4915
rect 4500 4850 4600 4900
rect 4650 4850 4750 4900
rect 4800 4950 4900 5000
rect 4950 4950 5050 5000
rect 4800 4935 5050 4950
rect 4800 4915 4815 4935
rect 4835 4915 4865 4935
rect 4885 4915 4915 4935
rect 4935 4915 4965 4935
rect 4985 4915 5015 4935
rect 5035 4915 5050 4935
rect 4800 4900 5050 4915
rect 4800 4850 4900 4900
rect 4950 4850 5050 4900
rect 5100 4950 5200 5000
rect 5250 4950 5350 5000
rect 5100 4935 5350 4950
rect 5100 4915 5115 4935
rect 5135 4915 5165 4935
rect 5185 4915 5215 4935
rect 5235 4915 5265 4935
rect 5285 4915 5315 4935
rect 5335 4915 5350 4935
rect 5100 4900 5350 4915
rect 5100 4850 5200 4900
rect 5250 4850 5350 4900
rect 5400 4950 5500 5000
rect 5550 4950 5650 5000
rect 5400 4935 5650 4950
rect 5400 4915 5415 4935
rect 5435 4915 5465 4935
rect 5485 4915 5515 4935
rect 5535 4915 5565 4935
rect 5585 4915 5615 4935
rect 5635 4915 5650 4935
rect 5400 4900 5650 4915
rect 5400 4850 5500 4900
rect 5550 4850 5650 4900
rect 5700 4950 5800 5000
rect 5850 4950 5950 5000
rect 5700 4935 5950 4950
rect 5700 4915 5715 4935
rect 5735 4915 5765 4935
rect 5785 4915 5815 4935
rect 5835 4915 5865 4935
rect 5885 4915 5915 4935
rect 5935 4915 5950 4935
rect 5700 4900 5950 4915
rect 5700 4850 5800 4900
rect 5850 4850 5950 4900
rect 6000 4950 6100 5000
rect 6150 4950 6250 5000
rect 6000 4935 6250 4950
rect 6000 4915 6015 4935
rect 6035 4915 6065 4935
rect 6085 4915 6115 4935
rect 6135 4915 6165 4935
rect 6185 4915 6215 4935
rect 6235 4915 6250 4935
rect 6000 4900 6250 4915
rect 6000 4850 6100 4900
rect 6150 4850 6250 4900
rect 6300 4950 6400 5000
rect 6450 4950 6550 5000
rect 6300 4935 6550 4950
rect 6300 4915 6315 4935
rect 6335 4915 6365 4935
rect 6385 4915 6415 4935
rect 6435 4915 6465 4935
rect 6485 4915 6515 4935
rect 6535 4915 6550 4935
rect 6300 4900 6550 4915
rect 6300 4850 6400 4900
rect 6450 4850 6550 4900
rect 6600 4950 6700 5000
rect 6750 4950 6850 5000
rect 6600 4935 6850 4950
rect 6600 4915 6615 4935
rect 6635 4915 6665 4935
rect 6685 4915 6715 4935
rect 6735 4915 6765 4935
rect 6785 4915 6815 4935
rect 6835 4915 6850 4935
rect 6600 4900 6850 4915
rect 6600 4850 6700 4900
rect 6750 4850 6850 4900
rect 6900 4950 7000 5000
rect 7050 4950 7150 5000
rect 6900 4935 7150 4950
rect 6900 4915 6915 4935
rect 6935 4915 6965 4935
rect 6985 4915 7015 4935
rect 7035 4915 7065 4935
rect 7085 4915 7115 4935
rect 7135 4915 7150 4935
rect 6900 4900 7150 4915
rect 6900 4850 7000 4900
rect 7050 4850 7150 4900
rect 7200 4950 7300 5000
rect 7350 4950 7450 5000
rect 7200 4935 7450 4950
rect 7200 4915 7215 4935
rect 7235 4915 7265 4935
rect 7285 4915 7315 4935
rect 7335 4915 7365 4935
rect 7385 4915 7415 4935
rect 7435 4915 7450 4935
rect 7200 4900 7450 4915
rect 7200 4850 7300 4900
rect 7350 4850 7450 4900
rect 7500 4950 7600 5000
rect 7650 4950 7750 5000
rect 7500 4935 7750 4950
rect 7500 4915 7515 4935
rect 7535 4915 7565 4935
rect 7585 4915 7615 4935
rect 7635 4915 7665 4935
rect 7685 4915 7715 4935
rect 7735 4915 7750 4935
rect 7500 4900 7750 4915
rect 7500 4850 7600 4900
rect 7650 4850 7750 4900
rect 7800 4950 7900 5000
rect 7950 4950 8050 5000
rect 7800 4935 8050 4950
rect 7800 4915 7815 4935
rect 7835 4915 7865 4935
rect 7885 4915 7915 4935
rect 7935 4915 7965 4935
rect 7985 4915 8015 4935
rect 8035 4915 8050 4935
rect 7800 4900 8050 4915
rect 7800 4850 7900 4900
rect 7950 4850 8050 4900
rect 8100 4950 8200 5000
rect 8250 4950 8350 5000
rect 8100 4935 8350 4950
rect 8100 4915 8115 4935
rect 8135 4915 8165 4935
rect 8185 4915 8215 4935
rect 8235 4915 8265 4935
rect 8285 4915 8315 4935
rect 8335 4915 8350 4935
rect 8100 4900 8350 4915
rect 8100 4850 8200 4900
rect 8250 4850 8350 4900
rect 8400 4950 8500 5000
rect 8550 4950 8650 5000
rect 8400 4935 8650 4950
rect 8400 4915 8415 4935
rect 8435 4915 8465 4935
rect 8485 4915 8515 4935
rect 8535 4915 8565 4935
rect 8585 4915 8615 4935
rect 8635 4915 8650 4935
rect 8400 4900 8650 4915
rect 8400 4850 8500 4900
rect 8550 4850 8650 4900
rect 8700 4950 8800 5000
rect 8850 4950 8950 5000
rect 8700 4935 8950 4950
rect 8700 4915 8715 4935
rect 8735 4915 8765 4935
rect 8785 4915 8815 4935
rect 8835 4915 8865 4935
rect 8885 4915 8915 4935
rect 8935 4915 8950 4935
rect 8700 4900 8950 4915
rect 8700 4850 8800 4900
rect 8850 4850 8950 4900
rect 9000 4950 9100 5000
rect 9150 4950 9250 5000
rect 9000 4935 9250 4950
rect 9000 4915 9015 4935
rect 9035 4915 9065 4935
rect 9085 4915 9115 4935
rect 9135 4915 9165 4935
rect 9185 4915 9215 4935
rect 9235 4915 9250 4935
rect 9000 4900 9250 4915
rect 9000 4850 9100 4900
rect 9150 4850 9250 4900
rect 9300 4950 9400 5000
rect 9450 4950 9550 5000
rect 9300 4935 9550 4950
rect 9300 4915 9315 4935
rect 9335 4915 9365 4935
rect 9385 4915 9415 4935
rect 9435 4915 9465 4935
rect 9485 4915 9515 4935
rect 9535 4915 9550 4935
rect 9300 4900 9550 4915
rect 9300 4850 9400 4900
rect 9450 4850 9550 4900
rect 9600 4950 9700 5000
rect 9750 4950 9850 5000
rect 9600 4935 9850 4950
rect 9600 4915 9615 4935
rect 9635 4915 9665 4935
rect 9685 4915 9715 4935
rect 9735 4915 9765 4935
rect 9785 4915 9815 4935
rect 9835 4915 9850 4935
rect 9600 4900 9850 4915
rect 9600 4850 9700 4900
rect 9750 4850 9850 4900
rect 9900 4950 10000 5000
rect 10050 4950 10150 5000
rect 9900 4935 10150 4950
rect 9900 4915 9915 4935
rect 9935 4915 9965 4935
rect 9985 4915 10015 4935
rect 10035 4915 10065 4935
rect 10085 4915 10115 4935
rect 10135 4915 10150 4935
rect 9900 4900 10150 4915
rect 9900 4850 10000 4900
rect 10050 4850 10150 4900
rect 10200 4950 10300 5000
rect 10350 4950 10450 5000
rect 10200 4935 10450 4950
rect 10200 4915 10215 4935
rect 10235 4915 10265 4935
rect 10285 4915 10315 4935
rect 10335 4915 10365 4935
rect 10385 4915 10415 4935
rect 10435 4915 10450 4935
rect 10200 4900 10450 4915
rect 10200 4850 10300 4900
rect 10350 4850 10450 4900
rect 10500 4950 10600 5000
rect 10650 4950 10750 5000
rect 10500 4935 10750 4950
rect 10500 4915 10515 4935
rect 10535 4915 10565 4935
rect 10585 4915 10615 4935
rect 10635 4915 10665 4935
rect 10685 4915 10715 4935
rect 10735 4915 10750 4935
rect 10500 4900 10750 4915
rect 10500 4850 10600 4900
rect 10650 4850 10750 4900
rect 10800 4950 10900 5000
rect 10950 4950 11050 5000
rect 10800 4935 11050 4950
rect 10800 4915 10815 4935
rect 10835 4915 10865 4935
rect 10885 4915 10915 4935
rect 10935 4915 10965 4935
rect 10985 4915 11015 4935
rect 11035 4915 11050 4935
rect 10800 4900 11050 4915
rect 10800 4850 10900 4900
rect 10950 4850 11050 4900
rect 11100 4950 11200 5000
rect 11250 4950 11350 5000
rect 11100 4935 11350 4950
rect 11100 4915 11115 4935
rect 11135 4915 11165 4935
rect 11185 4915 11215 4935
rect 11235 4915 11265 4935
rect 11285 4915 11315 4935
rect 11335 4915 11350 4935
rect 11100 4900 11350 4915
rect 11100 4850 11200 4900
rect 11250 4850 11350 4900
rect 11400 4950 11500 5000
rect 11550 4950 11650 5000
rect 11400 4935 11650 4950
rect 11400 4915 11415 4935
rect 11435 4915 11465 4935
rect 11485 4915 11515 4935
rect 11535 4915 11565 4935
rect 11585 4915 11615 4935
rect 11635 4915 11650 4935
rect 11400 4900 11650 4915
rect 11400 4850 11500 4900
rect 11550 4850 11650 4900
rect 11700 4950 11800 5000
rect 11850 4950 11950 5000
rect 11700 4935 11950 4950
rect 11700 4915 11715 4935
rect 11735 4915 11765 4935
rect 11785 4915 11815 4935
rect 11835 4915 11865 4935
rect 11885 4915 11915 4935
rect 11935 4915 11950 4935
rect 11700 4900 11950 4915
rect 11700 4850 11800 4900
rect 11850 4850 11950 4900
rect 12000 4950 12100 5000
rect 12150 4950 12250 5000
rect 12000 4935 12250 4950
rect 12000 4915 12015 4935
rect 12035 4915 12065 4935
rect 12085 4915 12115 4935
rect 12135 4915 12165 4935
rect 12185 4915 12215 4935
rect 12235 4915 12250 4935
rect 12000 4900 12250 4915
rect 12000 4850 12100 4900
rect 12150 4850 12250 4900
rect 12300 4950 12400 5000
rect 12450 4950 12550 5000
rect 12300 4935 12550 4950
rect 12300 4915 12315 4935
rect 12335 4915 12365 4935
rect 12385 4915 12415 4935
rect 12435 4915 12465 4935
rect 12485 4915 12515 4935
rect 12535 4915 12550 4935
rect 12300 4900 12550 4915
rect 12300 4850 12400 4900
rect 12450 4850 12550 4900
rect 12600 4950 12700 5000
rect 12750 4950 12850 5000
rect 12600 4935 12850 4950
rect 12600 4915 12615 4935
rect 12635 4915 12665 4935
rect 12685 4915 12715 4935
rect 12735 4915 12765 4935
rect 12785 4915 12815 4935
rect 12835 4915 12850 4935
rect 12600 4900 12850 4915
rect 12600 4850 12700 4900
rect 12750 4850 12850 4900
rect 12900 4950 13000 5000
rect 13050 4950 13150 5000
rect 12900 4935 13150 4950
rect 12900 4915 12915 4935
rect 12935 4915 12965 4935
rect 12985 4915 13015 4935
rect 13035 4915 13065 4935
rect 13085 4915 13115 4935
rect 13135 4915 13150 4935
rect 12900 4900 13150 4915
rect 12900 4850 13000 4900
rect 13050 4850 13150 4900
rect 13200 4950 13300 5000
rect 13350 4950 13450 5000
rect 13200 4935 13450 4950
rect 13200 4915 13215 4935
rect 13235 4915 13265 4935
rect 13285 4915 13315 4935
rect 13335 4915 13365 4935
rect 13385 4915 13415 4935
rect 13435 4915 13450 4935
rect 13200 4900 13450 4915
rect 13200 4850 13300 4900
rect 13350 4850 13450 4900
rect 13500 4950 13600 5000
rect 13650 4950 13750 5000
rect 13500 4935 13750 4950
rect 13500 4915 13515 4935
rect 13535 4915 13565 4935
rect 13585 4915 13615 4935
rect 13635 4915 13665 4935
rect 13685 4915 13715 4935
rect 13735 4915 13750 4935
rect 13500 4900 13750 4915
rect 13500 4850 13600 4900
rect 13650 4850 13750 4900
rect 13800 4950 13900 5000
rect 13950 4950 14050 5000
rect 13800 4935 14050 4950
rect 13800 4915 13815 4935
rect 13835 4915 13865 4935
rect 13885 4915 13915 4935
rect 13935 4915 13965 4935
rect 13985 4915 14015 4935
rect 14035 4915 14050 4935
rect 13800 4900 14050 4915
rect 13800 4850 13900 4900
rect 13950 4850 14050 4900
rect 14100 4950 14200 5000
rect 14250 4950 14350 5000
rect 14100 4935 14350 4950
rect 14100 4915 14115 4935
rect 14135 4915 14165 4935
rect 14185 4915 14215 4935
rect 14235 4915 14265 4935
rect 14285 4915 14315 4935
rect 14335 4915 14350 4935
rect 14100 4900 14350 4915
rect 14100 4850 14200 4900
rect 14250 4850 14350 4900
rect 14400 4950 14500 5000
rect 14550 4950 14650 5000
rect 14400 4935 14650 4950
rect 14400 4915 14415 4935
rect 14435 4915 14465 4935
rect 14485 4915 14515 4935
rect 14535 4915 14565 4935
rect 14585 4915 14615 4935
rect 14635 4915 14650 4935
rect 14400 4900 14650 4915
rect 14400 4850 14500 4900
rect 14550 4850 14650 4900
rect 14700 4950 14800 5000
rect 14850 4950 14950 5000
rect 14700 4935 14950 4950
rect 14700 4915 14715 4935
rect 14735 4915 14765 4935
rect 14785 4915 14815 4935
rect 14835 4915 14865 4935
rect 14885 4915 14915 4935
rect 14935 4915 14950 4935
rect 14700 4900 14950 4915
rect 14700 4850 14800 4900
rect 14850 4850 14950 4900
rect 15000 4950 15100 5000
rect 15150 4950 15250 5000
rect 15000 4935 15250 4950
rect 15000 4915 15015 4935
rect 15035 4915 15065 4935
rect 15085 4915 15115 4935
rect 15135 4915 15165 4935
rect 15185 4915 15215 4935
rect 15235 4915 15250 4935
rect 15000 4900 15250 4915
rect 15000 4850 15100 4900
rect 15150 4850 15250 4900
rect 15300 4950 15400 5000
rect 15450 4950 15550 5000
rect 15300 4935 15550 4950
rect 15300 4915 15315 4935
rect 15335 4915 15365 4935
rect 15385 4915 15415 4935
rect 15435 4915 15465 4935
rect 15485 4915 15515 4935
rect 15535 4915 15550 4935
rect 15300 4900 15550 4915
rect 15300 4850 15400 4900
rect 15450 4850 15550 4900
rect 15600 4950 15700 5000
rect 15750 4950 15850 5000
rect 15600 4935 15850 4950
rect 15600 4915 15615 4935
rect 15635 4915 15665 4935
rect 15685 4915 15715 4935
rect 15735 4915 15765 4935
rect 15785 4915 15815 4935
rect 15835 4915 15850 4935
rect 15600 4900 15850 4915
rect 15600 4850 15700 4900
rect 15750 4850 15850 4900
rect 15900 4950 16000 5000
rect 16050 4950 16150 5000
rect 15900 4935 16150 4950
rect 15900 4915 15915 4935
rect 15935 4915 15965 4935
rect 15985 4915 16015 4935
rect 16035 4915 16065 4935
rect 16085 4915 16115 4935
rect 16135 4915 16150 4935
rect 15900 4900 16150 4915
rect 15900 4850 16000 4900
rect 16050 4850 16150 4900
rect 16200 4950 16300 5000
rect 16350 4950 16450 5000
rect 16200 4935 16450 4950
rect 16200 4915 16215 4935
rect 16235 4915 16265 4935
rect 16285 4915 16315 4935
rect 16335 4915 16365 4935
rect 16385 4915 16415 4935
rect 16435 4915 16450 4935
rect 16200 4900 16450 4915
rect 16200 4850 16300 4900
rect 16350 4850 16450 4900
rect 16500 4950 16600 5000
rect 16650 4950 16750 5000
rect 16500 4935 16750 4950
rect 16500 4915 16515 4935
rect 16535 4915 16565 4935
rect 16585 4915 16615 4935
rect 16635 4915 16665 4935
rect 16685 4915 16715 4935
rect 16735 4915 16750 4935
rect 16500 4900 16750 4915
rect 16500 4850 16600 4900
rect 16650 4850 16750 4900
rect 16800 4950 16900 5000
rect 16950 4950 17050 5000
rect 16800 4935 17050 4950
rect 16800 4915 16815 4935
rect 16835 4915 16865 4935
rect 16885 4915 16915 4935
rect 16935 4915 16965 4935
rect 16985 4915 17015 4935
rect 17035 4915 17050 4935
rect 16800 4900 17050 4915
rect 16800 4850 16900 4900
rect 16950 4850 17050 4900
rect 17100 4950 17200 5000
rect 17250 4950 17350 5000
rect 17100 4935 17350 4950
rect 17100 4915 17115 4935
rect 17135 4915 17165 4935
rect 17185 4915 17215 4935
rect 17235 4915 17265 4935
rect 17285 4915 17315 4935
rect 17335 4915 17350 4935
rect 17100 4900 17350 4915
rect 17100 4850 17200 4900
rect 17250 4850 17350 4900
rect 17400 4950 17500 5000
rect 17550 4950 17650 5000
rect 17400 4935 17650 4950
rect 17400 4915 17415 4935
rect 17435 4915 17465 4935
rect 17485 4915 17515 4935
rect 17535 4915 17565 4935
rect 17585 4915 17615 4935
rect 17635 4915 17650 4935
rect 17400 4900 17650 4915
rect 17400 4850 17500 4900
rect 17550 4850 17650 4900
rect 17700 4950 17800 5000
rect 17850 4950 17950 5000
rect 17700 4935 17950 4950
rect 17700 4915 17715 4935
rect 17735 4915 17765 4935
rect 17785 4915 17815 4935
rect 17835 4915 17865 4935
rect 17885 4915 17915 4935
rect 17935 4915 17950 4935
rect 17700 4900 17950 4915
rect 17700 4850 17800 4900
rect 17850 4850 17950 4900
rect 18000 4950 18100 5000
rect 18150 4950 18250 5000
rect 18000 4935 18250 4950
rect 18000 4915 18015 4935
rect 18035 4915 18065 4935
rect 18085 4915 18115 4935
rect 18135 4915 18165 4935
rect 18185 4915 18215 4935
rect 18235 4915 18250 4935
rect 18000 4900 18250 4915
rect 18000 4850 18100 4900
rect 18150 4850 18250 4900
rect 18300 4950 18400 5000
rect 18450 4950 18550 5000
rect 18300 4935 18550 4950
rect 18300 4915 18315 4935
rect 18335 4915 18365 4935
rect 18385 4915 18415 4935
rect 18435 4915 18465 4935
rect 18485 4915 18515 4935
rect 18535 4915 18550 4935
rect 18300 4900 18550 4915
rect 18300 4850 18400 4900
rect 18450 4850 18550 4900
rect 18600 4950 18700 5000
rect 18750 4950 18850 5000
rect 18600 4935 18850 4950
rect 18600 4915 18615 4935
rect 18635 4915 18665 4935
rect 18685 4915 18715 4935
rect 18735 4915 18765 4935
rect 18785 4915 18815 4935
rect 18835 4915 18850 4935
rect 18600 4900 18850 4915
rect 18600 4850 18700 4900
rect 18750 4850 18850 4900
rect 18900 4950 19000 5000
rect 19050 4950 19150 5000
rect 18900 4935 19150 4950
rect 18900 4915 18915 4935
rect 18935 4915 18965 4935
rect 18985 4915 19015 4935
rect 19035 4915 19065 4935
rect 19085 4915 19115 4935
rect 19135 4915 19150 4935
rect 18900 4900 19150 4915
rect 18900 4850 19000 4900
rect 19050 4850 19150 4900
rect 19200 4950 19300 5000
rect 19350 4950 19450 5000
rect 19200 4935 19450 4950
rect 19200 4915 19215 4935
rect 19235 4915 19265 4935
rect 19285 4915 19315 4935
rect 19335 4915 19365 4935
rect 19385 4915 19415 4935
rect 19435 4915 19450 4935
rect 19200 4900 19450 4915
rect 19200 4850 19300 4900
rect 19350 4850 19450 4900
rect 19500 4950 19600 5000
rect 19650 4950 19750 5000
rect 19500 4935 19750 4950
rect 19500 4915 19515 4935
rect 19535 4915 19565 4935
rect 19585 4915 19615 4935
rect 19635 4915 19665 4935
rect 19685 4915 19715 4935
rect 19735 4915 19750 4935
rect 19500 4900 19750 4915
rect 19500 4850 19600 4900
rect 19650 4850 19750 4900
rect 19800 4950 19900 5000
rect 19950 4950 20050 5000
rect 19800 4935 20050 4950
rect 19800 4915 19815 4935
rect 19835 4915 19865 4935
rect 19885 4915 19915 4935
rect 19935 4915 19965 4935
rect 19985 4915 20015 4935
rect 20035 4915 20050 4935
rect 19800 4900 20050 4915
rect 19800 4850 19900 4900
rect 19950 4850 20050 4900
rect 20100 4950 20200 5000
rect 20250 4950 20350 5000
rect 20100 4935 20350 4950
rect 20100 4915 20115 4935
rect 20135 4915 20165 4935
rect 20185 4915 20215 4935
rect 20235 4915 20265 4935
rect 20285 4915 20315 4935
rect 20335 4915 20350 4935
rect 20100 4900 20350 4915
rect 20100 4850 20200 4900
rect 20250 4850 20350 4900
rect 20400 4950 20500 5000
rect 20550 4950 20650 5000
rect 20400 4935 20650 4950
rect 20400 4915 20415 4935
rect 20435 4915 20465 4935
rect 20485 4915 20515 4935
rect 20535 4915 20565 4935
rect 20585 4915 20615 4935
rect 20635 4915 20650 4935
rect 20400 4900 20650 4915
rect 20400 4850 20500 4900
rect 20550 4850 20650 4900
rect 20700 4950 20800 5000
rect 20850 4950 20950 5000
rect 20700 4935 20950 4950
rect 20700 4915 20715 4935
rect 20735 4915 20765 4935
rect 20785 4915 20815 4935
rect 20835 4915 20865 4935
rect 20885 4915 20915 4935
rect 20935 4915 20950 4935
rect 20700 4900 20950 4915
rect 20700 4850 20800 4900
rect 20850 4850 20950 4900
rect 21000 4950 21100 5000
rect 21150 4950 21250 5000
rect 21300 4950 21400 5000
rect 21000 4935 21400 4950
rect 21000 4915 21015 4935
rect 21035 4915 21065 4935
rect 21085 4915 21115 4935
rect 21135 4915 21165 4935
rect 21185 4915 21215 4935
rect 21235 4915 21265 4935
rect 21285 4915 21315 4935
rect 21335 4915 21365 4935
rect 21385 4915 21400 4935
rect 21000 4900 21400 4915
rect 21000 4850 21100 4900
rect 21150 4850 21250 4900
rect 21300 4850 21400 4900
rect 21450 4950 21550 5000
rect 21600 4950 21700 5000
rect 21750 4950 21850 5000
rect 21450 4935 21850 4950
rect 21450 4915 21465 4935
rect 21485 4915 21515 4935
rect 21535 4915 21565 4935
rect 21585 4915 21615 4935
rect 21635 4915 21665 4935
rect 21685 4915 21715 4935
rect 21735 4915 21765 4935
rect 21785 4915 21815 4935
rect 21835 4915 21850 4935
rect 21450 4900 21850 4915
rect 21450 4850 21550 4900
rect 21600 4850 21700 4900
rect 21750 4850 21850 4900
rect 21900 4950 22000 5000
rect 22050 4950 22150 5000
rect 21900 4935 22150 4950
rect 21900 4915 21915 4935
rect 21935 4915 21965 4935
rect 21985 4915 22015 4935
rect 22035 4915 22065 4935
rect 22085 4915 22115 4935
rect 22135 4915 22150 4935
rect 21900 4900 22150 4915
rect 21900 4850 22000 4900
rect 22050 4850 22150 4900
rect 22200 4950 22300 5000
rect 22350 4950 22450 5000
rect 22200 4935 22450 4950
rect 22200 4915 22215 4935
rect 22235 4915 22265 4935
rect 22285 4915 22315 4935
rect 22335 4915 22365 4935
rect 22385 4915 22415 4935
rect 22435 4915 22450 4935
rect 22200 4900 22450 4915
rect 22200 4850 22300 4900
rect 22350 4850 22450 4900
rect 22500 4950 22600 5000
rect 22650 4950 22750 5000
rect 22500 4935 22750 4950
rect 22500 4915 22515 4935
rect 22535 4915 22565 4935
rect 22585 4915 22615 4935
rect 22635 4915 22665 4935
rect 22685 4915 22715 4935
rect 22735 4915 22750 4935
rect 22500 4900 22750 4915
rect 22500 4850 22600 4900
rect 22650 4850 22750 4900
rect 22800 4950 22900 5000
rect 22950 4950 23050 5000
rect 22800 4935 23050 4950
rect 22800 4915 22815 4935
rect 22835 4915 22865 4935
rect 22885 4915 22915 4935
rect 22935 4915 22965 4935
rect 22985 4915 23015 4935
rect 23035 4915 23050 4935
rect 22800 4900 23050 4915
rect 22800 4850 22900 4900
rect 22950 4850 23050 4900
rect 23100 4950 23200 5000
rect 23250 4950 23350 5000
rect 23400 4950 23500 5000
rect 23100 4935 23500 4950
rect 23100 4915 23115 4935
rect 23135 4915 23165 4935
rect 23185 4915 23215 4935
rect 23235 4915 23265 4935
rect 23285 4915 23315 4935
rect 23335 4915 23365 4935
rect 23385 4915 23415 4935
rect 23435 4915 23465 4935
rect 23485 4915 23500 4935
rect 23100 4900 23500 4915
rect 23100 4850 23200 4900
rect 23250 4850 23350 4900
rect 23400 4850 23500 4900
rect 23550 4950 23650 5000
rect 23700 4950 23800 5000
rect 23850 4950 23950 5000
rect 23550 4935 23950 4950
rect 23550 4915 23565 4935
rect 23585 4915 23615 4935
rect 23635 4915 23665 4935
rect 23685 4915 23715 4935
rect 23735 4915 23765 4935
rect 23785 4915 23815 4935
rect 23835 4915 23865 4935
rect 23885 4915 23915 4935
rect 23935 4915 23950 4935
rect 23550 4900 23950 4915
rect 23550 4850 23650 4900
rect 23700 4850 23800 4900
rect 23850 4850 23950 4900
rect 24000 4950 24100 5000
rect 24150 4950 24250 5000
rect 24000 4935 24250 4950
rect 24000 4915 24015 4935
rect 24035 4915 24065 4935
rect 24085 4915 24115 4935
rect 24135 4915 24165 4935
rect 24185 4915 24215 4935
rect 24235 4915 24250 4935
rect 24000 4900 24250 4915
rect 24000 4850 24100 4900
rect 24150 4850 24250 4900
rect 24300 4950 24400 5000
rect 24450 4950 24550 5000
rect 24300 4935 24550 4950
rect 24300 4915 24315 4935
rect 24335 4915 24365 4935
rect 24385 4915 24415 4935
rect 24435 4915 24465 4935
rect 24485 4915 24515 4935
rect 24535 4915 24550 4935
rect 24300 4900 24550 4915
rect 24300 4850 24400 4900
rect 24450 4850 24550 4900
rect 24600 4950 24700 5000
rect 24750 4950 24850 5000
rect 24600 4935 24850 4950
rect 24600 4915 24615 4935
rect 24635 4915 24665 4935
rect 24685 4915 24715 4935
rect 24735 4915 24765 4935
rect 24785 4915 24815 4935
rect 24835 4915 24850 4935
rect 24600 4900 24850 4915
rect 24600 4850 24700 4900
rect 24750 4850 24850 4900
rect 24900 4950 25000 5000
rect 25050 4950 25150 5000
rect 24900 4935 25150 4950
rect 24900 4915 24915 4935
rect 24935 4915 24965 4935
rect 24985 4915 25015 4935
rect 25035 4915 25065 4935
rect 25085 4915 25115 4935
rect 25135 4915 25150 4935
rect 24900 4900 25150 4915
rect 24900 4850 25000 4900
rect 25050 4850 25150 4900
rect 25200 4950 25300 5000
rect 25350 4950 25450 5000
rect 25500 4950 25600 5000
rect 25200 4935 25600 4950
rect 25200 4915 25215 4935
rect 25235 4915 25265 4935
rect 25285 4915 25315 4935
rect 25335 4915 25365 4935
rect 25385 4915 25415 4935
rect 25435 4915 25465 4935
rect 25485 4915 25515 4935
rect 25535 4915 25565 4935
rect 25585 4915 25600 4935
rect 25200 4900 25600 4915
rect 25200 4850 25300 4900
rect 25350 4850 25450 4900
rect 25500 4850 25600 4900
rect 25650 4950 25750 5000
rect 25800 4950 25900 5000
rect 25950 4950 26050 5000
rect 25650 4935 26050 4950
rect 25650 4915 25665 4935
rect 25685 4915 25715 4935
rect 25735 4915 25765 4935
rect 25785 4915 25815 4935
rect 25835 4915 25865 4935
rect 25885 4915 25915 4935
rect 25935 4915 25965 4935
rect 25985 4915 26015 4935
rect 26035 4915 26050 4935
rect 25650 4900 26050 4915
rect 25650 4850 25750 4900
rect 25800 4850 25900 4900
rect 25950 4850 26050 4900
rect 26100 4950 26200 5000
rect 26250 4950 26350 5000
rect 26100 4935 26350 4950
rect 26100 4915 26115 4935
rect 26135 4915 26165 4935
rect 26185 4915 26215 4935
rect 26235 4915 26265 4935
rect 26285 4915 26315 4935
rect 26335 4915 26350 4935
rect 26100 4900 26350 4915
rect 26100 4850 26200 4900
rect 26250 4850 26350 4900
rect 26400 4950 26500 5000
rect 26550 4950 26650 5000
rect 26400 4935 26650 4950
rect 26400 4915 26415 4935
rect 26435 4915 26465 4935
rect 26485 4915 26515 4935
rect 26535 4915 26565 4935
rect 26585 4915 26615 4935
rect 26635 4915 26650 4935
rect 26400 4900 26650 4915
rect 26400 4850 26500 4900
rect 26550 4850 26650 4900
rect 26700 4950 26800 5000
rect 26850 4950 26950 5000
rect 26700 4935 26950 4950
rect 26700 4915 26715 4935
rect 26735 4915 26765 4935
rect 26785 4915 26815 4935
rect 26835 4915 26865 4935
rect 26885 4915 26915 4935
rect 26935 4915 26950 4935
rect 26700 4900 26950 4915
rect 26700 4850 26800 4900
rect 26850 4850 26950 4900
rect 27000 4950 27100 5000
rect 27150 4950 27250 5000
rect 27000 4935 27250 4950
rect 27000 4915 27015 4935
rect 27035 4915 27065 4935
rect 27085 4915 27115 4935
rect 27135 4915 27165 4935
rect 27185 4915 27215 4935
rect 27235 4915 27250 4935
rect 27000 4900 27250 4915
rect 27000 4850 27100 4900
rect 27150 4850 27250 4900
rect 27300 4950 27400 5000
rect 27450 4950 27550 5000
rect 27600 4950 27700 5000
rect 27300 4935 27700 4950
rect 27300 4915 27315 4935
rect 27335 4915 27365 4935
rect 27385 4915 27415 4935
rect 27435 4915 27465 4935
rect 27485 4915 27515 4935
rect 27535 4915 27565 4935
rect 27585 4915 27615 4935
rect 27635 4915 27665 4935
rect 27685 4915 27700 4935
rect 27300 4900 27700 4915
rect 27300 4850 27400 4900
rect 27450 4850 27550 4900
rect 27600 4850 27700 4900
rect 27750 4950 27850 5000
rect 27900 4950 28000 5000
rect 28050 4950 28150 5000
rect 27750 4935 28150 4950
rect 27750 4915 27765 4935
rect 27785 4915 27815 4935
rect 27835 4915 27865 4935
rect 27885 4915 27915 4935
rect 27935 4915 27965 4935
rect 27985 4915 28015 4935
rect 28035 4915 28065 4935
rect 28085 4915 28115 4935
rect 28135 4915 28150 4935
rect 27750 4900 28150 4915
rect 27750 4850 27850 4900
rect 27900 4850 28000 4900
rect 28050 4850 28150 4900
rect 28200 4950 28300 5000
rect 28350 4950 28450 5000
rect 28200 4935 28450 4950
rect 28200 4915 28215 4935
rect 28235 4915 28265 4935
rect 28285 4915 28315 4935
rect 28335 4915 28365 4935
rect 28385 4915 28415 4935
rect 28435 4915 28450 4935
rect 28200 4900 28450 4915
rect 28200 4850 28300 4900
rect 28350 4850 28450 4900
rect 28500 4950 28600 5000
rect 28650 4950 28750 5000
rect 28500 4935 28750 4950
rect 28500 4915 28515 4935
rect 28535 4915 28565 4935
rect 28585 4915 28615 4935
rect 28635 4915 28665 4935
rect 28685 4915 28715 4935
rect 28735 4915 28750 4935
rect 28500 4900 28750 4915
rect 28500 4850 28600 4900
rect 28650 4850 28750 4900
rect 28800 4950 28900 5000
rect 28950 4950 29050 5000
rect 28800 4935 29050 4950
rect 28800 4915 28815 4935
rect 28835 4915 28865 4935
rect 28885 4915 28915 4935
rect 28935 4915 28965 4935
rect 28985 4915 29015 4935
rect 29035 4915 29050 4935
rect 28800 4900 29050 4915
rect 28800 4850 28900 4900
rect 28950 4850 29050 4900
rect 29100 4950 29200 5000
rect 29250 4950 29350 5000
rect 29100 4935 29350 4950
rect 29100 4915 29115 4935
rect 29135 4915 29165 4935
rect 29185 4915 29215 4935
rect 29235 4915 29265 4935
rect 29285 4915 29315 4935
rect 29335 4915 29350 4935
rect 29100 4900 29350 4915
rect 29100 4850 29200 4900
rect 29250 4850 29350 4900
rect 29400 4950 29500 5000
rect 29550 4950 29650 5000
rect 29700 4950 29800 5000
rect 29400 4935 29800 4950
rect 29400 4915 29415 4935
rect 29435 4915 29465 4935
rect 29485 4915 29515 4935
rect 29535 4915 29565 4935
rect 29585 4915 29615 4935
rect 29635 4915 29665 4935
rect 29685 4915 29715 4935
rect 29735 4915 29765 4935
rect 29785 4915 29800 4935
rect 29400 4900 29800 4915
rect 29400 4850 29500 4900
rect 29550 4850 29650 4900
rect 29700 4850 29800 4900
rect 29850 4950 29950 5000
rect 30000 4950 30100 5000
rect 29850 4935 30100 4950
rect 29850 4915 29865 4935
rect 29885 4915 29915 4935
rect 29935 4915 29965 4935
rect 29985 4915 30015 4935
rect 30035 4915 30065 4935
rect 30085 4915 30100 4935
rect 29850 4900 30100 4915
rect 29850 4850 29950 4900
rect 30000 4850 30100 4900
rect 30150 4950 30250 5000
rect 30300 4950 30400 5000
rect 30150 4935 30400 4950
rect 30150 4915 30165 4935
rect 30185 4915 30215 4935
rect 30235 4915 30265 4935
rect 30285 4915 30315 4935
rect 30335 4915 30365 4935
rect 30385 4915 30400 4935
rect 30150 4900 30400 4915
rect 30150 4850 30250 4900
rect 30300 4850 30400 4900
rect 30450 4950 30550 5000
rect 30600 4950 30700 5000
rect 30450 4935 30700 4950
rect 30450 4915 30465 4935
rect 30485 4915 30515 4935
rect 30535 4915 30565 4935
rect 30585 4915 30615 4935
rect 30635 4915 30665 4935
rect 30685 4915 30700 4935
rect 30450 4900 30700 4915
rect 30450 4850 30550 4900
rect 30600 4850 30700 4900
rect 30750 4950 30850 5000
rect 30900 4950 31000 5000
rect 30750 4935 31000 4950
rect 30750 4915 30765 4935
rect 30785 4915 30815 4935
rect 30835 4915 30865 4935
rect 30885 4915 30915 4935
rect 30935 4915 30965 4935
rect 30985 4915 31000 4935
rect 30750 4900 31000 4915
rect 30750 4850 30850 4900
rect 30900 4850 31000 4900
rect 31050 4950 31150 5000
rect 31200 4950 31300 5000
rect 31350 4950 31450 5000
rect 31050 4935 31450 4950
rect 31050 4915 31065 4935
rect 31085 4915 31115 4935
rect 31135 4915 31165 4935
rect 31185 4915 31215 4935
rect 31235 4915 31265 4935
rect 31285 4915 31315 4935
rect 31335 4915 31365 4935
rect 31385 4915 31415 4935
rect 31435 4915 31450 4935
rect 31050 4900 31450 4915
rect 31050 4850 31150 4900
rect 31200 4850 31300 4900
rect 31350 4850 31450 4900
rect 31500 4950 31600 5000
rect 31650 4950 31750 5000
rect 31500 4935 31750 4950
rect 31500 4915 31515 4935
rect 31535 4915 31565 4935
rect 31585 4915 31615 4935
rect 31635 4915 31665 4935
rect 31685 4915 31715 4935
rect 31735 4915 31750 4935
rect 31500 4900 31750 4915
rect 31500 4850 31600 4900
rect 31650 4850 31750 4900
rect 31800 4950 31900 5000
rect 31950 4950 32050 5000
rect 31800 4935 32050 4950
rect 31800 4915 31815 4935
rect 31835 4915 31865 4935
rect 31885 4915 31915 4935
rect 31935 4915 31965 4935
rect 31985 4915 32015 4935
rect 32035 4915 32050 4935
rect 31800 4900 32050 4915
rect 31800 4850 31900 4900
rect 31950 4850 32050 4900
rect -600 4335 -500 4350
rect -450 4335 -350 4350
rect -300 4335 -200 4350
rect -150 4335 -50 4350
rect 0 4335 100 4350
rect 150 4335 250 4350
rect 300 4335 400 4350
rect 450 4335 550 4350
rect 600 4335 700 4350
rect 750 4335 850 4350
rect 900 4335 1000 4350
rect 1050 4335 1150 4350
rect 1200 4335 1300 4350
rect 1350 4335 1450 4350
rect 1500 4335 1600 4350
rect 1650 4335 1750 4350
rect 1800 4335 1900 4350
rect 1950 4335 2050 4350
rect 2100 4335 2200 4350
rect 2250 4335 2350 4350
rect 2400 4335 2500 4350
rect 2550 4335 2650 4350
rect 2700 4335 2800 4350
rect 2850 4335 2950 4350
rect 3000 4335 3100 4350
rect 3150 4335 3250 4350
rect 3300 4335 3400 4350
rect 3450 4335 3550 4350
rect 3600 4335 3700 4350
rect 3750 4335 3850 4350
rect 3900 4335 4000 4350
rect 4050 4335 4150 4350
rect 4200 4335 4300 4350
rect 4350 4335 4450 4350
rect 4500 4335 4600 4350
rect 4650 4335 4750 4350
rect 4800 4335 4900 4350
rect 4950 4335 5050 4350
rect 5100 4335 5200 4350
rect 5250 4335 5350 4350
rect 5400 4335 5500 4350
rect 5550 4335 5650 4350
rect 5700 4335 5800 4350
rect 5850 4335 5950 4350
rect 6000 4335 6100 4350
rect 6150 4335 6250 4350
rect 6300 4335 6400 4350
rect 6450 4335 6550 4350
rect 6600 4335 6700 4350
rect 6750 4335 6850 4350
rect 6900 4335 7000 4350
rect 7050 4335 7150 4350
rect 7200 4335 7300 4350
rect 7350 4335 7450 4350
rect 7500 4335 7600 4350
rect 7650 4335 7750 4350
rect 7800 4335 7900 4350
rect 7950 4335 8050 4350
rect 8100 4335 8200 4350
rect 8250 4335 8350 4350
rect 8400 4335 8500 4350
rect 8550 4335 8650 4350
rect 8700 4335 8800 4350
rect 8850 4335 8950 4350
rect 9000 4335 9100 4350
rect 9150 4335 9250 4350
rect 9300 4335 9400 4350
rect 9450 4335 9550 4350
rect 9600 4335 9700 4350
rect 9750 4335 9850 4350
rect 9900 4335 10000 4350
rect 10050 4335 10150 4350
rect 10200 4335 10300 4350
rect 10350 4335 10450 4350
rect 10500 4335 10600 4350
rect 10650 4335 10750 4350
rect 10800 4335 10900 4350
rect 10950 4335 11050 4350
rect 11100 4335 11200 4350
rect 11250 4335 11350 4350
rect 11400 4335 11500 4350
rect 11550 4335 11650 4350
rect 11700 4335 11800 4350
rect 11850 4335 11950 4350
rect 12000 4335 12100 4350
rect 12150 4335 12250 4350
rect 12300 4335 12400 4350
rect 12450 4335 12550 4350
rect 12600 4335 12700 4350
rect 12750 4335 12850 4350
rect 12900 4335 13000 4350
rect 13050 4335 13150 4350
rect 13200 4335 13300 4350
rect 13350 4335 13450 4350
rect 13500 4335 13600 4350
rect 13650 4335 13750 4350
rect 13800 4335 13900 4350
rect 13950 4335 14050 4350
rect 14100 4335 14200 4350
rect 14250 4335 14350 4350
rect 14400 4335 14500 4350
rect 14550 4335 14650 4350
rect 14700 4335 14800 4350
rect 14850 4335 14950 4350
rect 15000 4335 15100 4350
rect 15150 4335 15250 4350
rect 15300 4335 15400 4350
rect 15450 4335 15550 4350
rect 15600 4335 15700 4350
rect 15750 4335 15850 4350
rect 15900 4335 16000 4350
rect 16050 4335 16150 4350
rect 16200 4335 16300 4350
rect 16350 4335 16450 4350
rect 16500 4335 16600 4350
rect 16650 4335 16750 4350
rect 16800 4335 16900 4350
rect 16950 4335 17050 4350
rect 17100 4335 17200 4350
rect 17250 4335 17350 4350
rect 17400 4335 17500 4350
rect 17550 4335 17650 4350
rect 17700 4335 17800 4350
rect 17850 4335 17950 4350
rect 18000 4335 18100 4350
rect 18150 4335 18250 4350
rect 18300 4335 18400 4350
rect 18450 4335 18550 4350
rect 18600 4335 18700 4350
rect 18750 4335 18850 4350
rect 18900 4335 19000 4350
rect 19050 4335 19150 4350
rect 19200 4335 19300 4350
rect 19350 4335 19450 4350
rect 19500 4335 19600 4350
rect 19650 4335 19750 4350
rect 19800 4335 19900 4350
rect 19950 4335 20050 4350
rect 20100 4335 20200 4350
rect 20250 4335 20350 4350
rect 20400 4335 20500 4350
rect 20550 4335 20650 4350
rect 20700 4335 20800 4350
rect 20850 4335 20950 4350
rect 21000 4335 21100 4350
rect 21150 4335 21250 4350
rect 21300 4335 21400 4350
rect 21450 4335 21550 4350
rect 21600 4335 21700 4350
rect 21750 4335 21850 4350
rect 21900 4335 22000 4350
rect 22050 4335 22150 4350
rect 22200 4335 22300 4350
rect 22350 4335 22450 4350
rect 22500 4335 22600 4350
rect 22650 4335 22750 4350
rect 22800 4335 22900 4350
rect 22950 4335 23050 4350
rect 23100 4335 23200 4350
rect 23250 4335 23350 4350
rect 23400 4335 23500 4350
rect 23550 4335 23650 4350
rect 23700 4335 23800 4350
rect 23850 4335 23950 4350
rect 24000 4335 24100 4350
rect 24150 4335 24250 4350
rect 24300 4335 24400 4350
rect 24450 4335 24550 4350
rect 24600 4335 24700 4350
rect 24750 4335 24850 4350
rect 24900 4335 25000 4350
rect 25050 4335 25150 4350
rect 25200 4335 25300 4350
rect 25350 4335 25450 4350
rect 25500 4335 25600 4350
rect 25650 4335 25750 4350
rect 25800 4335 25900 4350
rect 25950 4335 26050 4350
rect 26100 4335 26200 4350
rect 26250 4335 26350 4350
rect 26400 4335 26500 4350
rect 26550 4335 26650 4350
rect 26700 4335 26800 4350
rect 26850 4335 26950 4350
rect 27000 4335 27100 4350
rect 27150 4335 27250 4350
rect 27300 4335 27400 4350
rect 27450 4335 27550 4350
rect 27600 4335 27700 4350
rect 27750 4335 27850 4350
rect 27900 4335 28000 4350
rect 28050 4335 28150 4350
rect 28200 4335 28300 4350
rect 28350 4335 28450 4350
rect 28500 4335 28600 4350
rect 28650 4335 28750 4350
rect 28800 4335 28900 4350
rect 28950 4335 29050 4350
rect 29100 4335 29200 4350
rect 29250 4335 29350 4350
rect 29400 4335 29500 4350
rect 29550 4335 29650 4350
rect 29700 4335 29800 4350
rect 29850 4335 29950 4350
rect 30000 4335 30100 4350
rect 30150 4335 30250 4350
rect 30300 4335 30400 4350
rect 30450 4335 30550 4350
rect 30600 4335 30700 4350
rect 30750 4335 30850 4350
rect 30900 4335 31000 4350
rect 31050 4335 31150 4350
rect 31200 4335 31300 4350
rect 31350 4335 31450 4350
rect 31500 4335 31600 4350
rect 31650 4335 31750 4350
rect 31800 4335 31900 4350
rect 31950 4335 32050 4350
rect -600 4200 -500 4215
rect -450 4200 -350 4215
rect -300 4200 -200 4215
rect -150 4200 -50 4215
rect 0 4200 100 4215
rect 150 4200 250 4215
rect 300 4200 400 4215
rect 450 4200 550 4215
rect 600 4200 700 4215
rect 750 4200 850 4215
rect 900 4200 1000 4215
rect 1050 4200 1150 4215
rect 1200 4200 1300 4215
rect 1350 4200 1450 4215
rect 1500 4200 1600 4215
rect 1650 4200 1750 4215
rect 1800 4200 1900 4215
rect 1950 4200 2050 4215
rect 2100 4200 2200 4215
rect 2250 4200 2350 4215
rect 2400 4200 2500 4215
rect 2550 4200 2650 4215
rect 2700 4200 2800 4215
rect 2850 4200 2950 4215
rect 3000 4200 3100 4215
rect 3150 4200 3250 4215
rect 3300 4200 3400 4215
rect 3450 4200 3550 4215
rect 3600 4200 3700 4215
rect 3750 4200 3850 4215
rect 3900 4200 4000 4215
rect 4050 4200 4150 4215
rect 4200 4200 4300 4215
rect 4350 4200 4450 4215
rect 4500 4200 4600 4215
rect 4650 4200 4750 4215
rect 4800 4200 4900 4215
rect 4950 4200 5050 4215
rect 5100 4200 5200 4215
rect 5250 4200 5350 4215
rect 5400 4200 5500 4215
rect 5550 4200 5650 4215
rect 5700 4200 5800 4215
rect 5850 4200 5950 4215
rect 6000 4200 6100 4215
rect 6150 4200 6250 4215
rect 6300 4200 6400 4215
rect 6450 4200 6550 4215
rect 6600 4200 6700 4215
rect 6750 4200 6850 4215
rect 6900 4200 7000 4215
rect 7050 4200 7150 4215
rect 7200 4200 7300 4215
rect 7350 4200 7450 4215
rect 7500 4200 7600 4215
rect 7650 4200 7750 4215
rect 7800 4200 7900 4215
rect 7950 4200 8050 4215
rect 8100 4200 8200 4215
rect 8250 4200 8350 4215
rect 8400 4200 8500 4215
rect 8550 4200 8650 4215
rect 8700 4200 8800 4215
rect 8850 4200 8950 4215
rect 9000 4200 9100 4215
rect 9150 4200 9250 4215
rect 9300 4200 9400 4215
rect 9450 4200 9550 4215
rect 9600 4200 9700 4215
rect 9750 4200 9850 4215
rect 9900 4200 10000 4215
rect 10050 4200 10150 4215
rect 10200 4200 10300 4215
rect 10350 4200 10450 4215
rect 10500 4200 10600 4215
rect 10650 4200 10750 4215
rect 10800 4200 10900 4215
rect 10950 4200 11050 4215
rect 11100 4200 11200 4215
rect 11250 4200 11350 4215
rect 11400 4200 11500 4215
rect 11550 4200 11650 4215
rect 11700 4200 11800 4215
rect 11850 4200 11950 4215
rect 12000 4200 12100 4215
rect 12150 4200 12250 4215
rect 12300 4200 12400 4215
rect 12450 4200 12550 4215
rect 12600 4200 12700 4215
rect 12750 4200 12850 4215
rect 12900 4200 13000 4215
rect 13050 4200 13150 4215
rect 13200 4200 13300 4215
rect 13350 4200 13450 4215
rect 13500 4200 13600 4215
rect 13650 4200 13750 4215
rect 13800 4200 13900 4215
rect 13950 4200 14050 4215
rect 14100 4200 14200 4215
rect 14250 4200 14350 4215
rect 14400 4200 14500 4215
rect 14550 4200 14650 4215
rect 14700 4200 14800 4215
rect 14850 4200 14950 4215
rect 15000 4200 15100 4215
rect 15150 4200 15250 4215
rect 15300 4200 15400 4215
rect 15450 4200 15550 4215
rect 15600 4200 15700 4215
rect 15750 4200 15850 4215
rect 15900 4200 16000 4215
rect 16050 4200 16150 4215
rect 16200 4200 16300 4215
rect 16350 4200 16450 4215
rect 16500 4200 16600 4215
rect 16650 4200 16750 4215
rect 16800 4200 16900 4215
rect 16950 4200 17050 4215
rect 17100 4200 17200 4215
rect 17250 4200 17350 4215
rect 17400 4200 17500 4215
rect 17550 4200 17650 4215
rect 17700 4200 17800 4215
rect 17850 4200 17950 4215
rect 18000 4200 18100 4215
rect 18150 4200 18250 4215
rect 18300 4200 18400 4215
rect 18450 4200 18550 4215
rect 18600 4200 18700 4215
rect 18750 4200 18850 4215
rect 18900 4200 19000 4215
rect 19050 4200 19150 4215
rect 19200 4200 19300 4215
rect 19350 4200 19450 4215
rect 19500 4200 19600 4215
rect 19650 4200 19750 4215
rect 19800 4200 19900 4215
rect 19950 4200 20050 4215
rect 20100 4200 20200 4215
rect 20250 4200 20350 4215
rect 20400 4200 20500 4215
rect 20550 4200 20650 4215
rect 20700 4200 20800 4215
rect 20850 4200 20950 4215
rect 21000 4200 21100 4215
rect 21150 4200 21250 4215
rect 21300 4200 21400 4215
rect 21450 4200 21550 4215
rect 21600 4200 21700 4215
rect 21750 4200 21850 4215
rect 21900 4200 22000 4215
rect 22050 4200 22150 4215
rect 22200 4200 22300 4215
rect 22350 4200 22450 4215
rect 22500 4200 22600 4215
rect 22650 4200 22750 4215
rect 22800 4200 22900 4215
rect 22950 4200 23050 4215
rect 23100 4200 23200 4215
rect 23250 4200 23350 4215
rect 23400 4200 23500 4215
rect 23550 4200 23650 4215
rect 23700 4200 23800 4215
rect 23850 4200 23950 4215
rect 24000 4200 24100 4215
rect 24150 4200 24250 4215
rect 24300 4200 24400 4215
rect 24450 4200 24550 4215
rect 24600 4200 24700 4215
rect 24750 4200 24850 4215
rect 24900 4200 25000 4215
rect 25050 4200 25150 4215
rect 25200 4200 25300 4215
rect 25350 4200 25450 4215
rect 25500 4200 25600 4215
rect 25650 4200 25750 4215
rect 25800 4200 25900 4215
rect 25950 4200 26050 4215
rect 26100 4200 26200 4215
rect 26250 4200 26350 4215
rect 26400 4200 26500 4215
rect 26550 4200 26650 4215
rect 26700 4200 26800 4215
rect 26850 4200 26950 4215
rect 27000 4200 27100 4215
rect 27150 4200 27250 4215
rect 27300 4200 27400 4215
rect 27450 4200 27550 4215
rect 27600 4200 27700 4215
rect 27750 4200 27850 4215
rect 27900 4200 28000 4215
rect 28050 4200 28150 4215
rect 28200 4200 28300 4215
rect 28350 4200 28450 4215
rect 28500 4200 28600 4215
rect 28650 4200 28750 4215
rect 28800 4200 28900 4215
rect 28950 4200 29050 4215
rect 29100 4200 29200 4215
rect 29250 4200 29350 4215
rect 29400 4200 29500 4215
rect 29550 4200 29650 4215
rect 29700 4200 29800 4215
rect 29850 4200 29950 4215
rect 30000 4200 30100 4215
rect 30150 4200 30250 4215
rect 30300 4200 30400 4215
rect 30450 4200 30550 4215
rect 30600 4200 30700 4215
rect 30750 4200 30850 4215
rect 30900 4200 31000 4215
rect 31050 4200 31150 4215
rect 31200 4200 31300 4215
rect 31350 4200 31450 4215
rect 31500 4200 31600 4215
rect 31650 4200 31750 4215
rect 31800 4200 31900 4215
rect 31950 4200 32050 4215
rect -600 3650 -500 3700
rect -450 3650 -350 3700
rect -600 3635 -350 3650
rect -600 3615 -585 3635
rect -565 3615 -535 3635
rect -515 3615 -485 3635
rect -465 3615 -435 3635
rect -415 3615 -385 3635
rect -365 3615 -350 3635
rect -600 3600 -350 3615
rect -600 3550 -500 3600
rect -450 3550 -350 3600
rect -300 3650 -200 3700
rect -150 3650 -50 3700
rect -300 3635 -50 3650
rect -300 3615 -285 3635
rect -265 3615 -235 3635
rect -215 3615 -185 3635
rect -165 3615 -135 3635
rect -115 3615 -85 3635
rect -65 3615 -50 3635
rect -300 3600 -50 3615
rect -300 3550 -200 3600
rect -150 3550 -50 3600
rect 0 3650 100 3700
rect 150 3650 250 3700
rect 0 3635 250 3650
rect 0 3615 15 3635
rect 35 3615 65 3635
rect 85 3615 115 3635
rect 135 3615 165 3635
rect 185 3615 215 3635
rect 235 3615 250 3635
rect 0 3600 250 3615
rect 0 3550 100 3600
rect 150 3550 250 3600
rect 300 3650 400 3700
rect 450 3650 550 3700
rect 300 3635 550 3650
rect 300 3615 315 3635
rect 335 3615 365 3635
rect 385 3615 415 3635
rect 435 3615 465 3635
rect 485 3615 515 3635
rect 535 3615 550 3635
rect 300 3600 550 3615
rect 300 3550 400 3600
rect 450 3550 550 3600
rect 600 3650 700 3700
rect 750 3650 850 3700
rect 600 3635 850 3650
rect 600 3615 615 3635
rect 635 3615 665 3635
rect 685 3615 715 3635
rect 735 3615 765 3635
rect 785 3615 815 3635
rect 835 3615 850 3635
rect 600 3600 850 3615
rect 600 3550 700 3600
rect 750 3550 850 3600
rect 900 3650 1000 3700
rect 1050 3650 1150 3700
rect 900 3635 1150 3650
rect 900 3615 915 3635
rect 935 3615 965 3635
rect 985 3615 1015 3635
rect 1035 3615 1065 3635
rect 1085 3615 1115 3635
rect 1135 3615 1150 3635
rect 900 3600 1150 3615
rect 900 3550 1000 3600
rect 1050 3550 1150 3600
rect 1200 3650 1300 3700
rect 1350 3650 1450 3700
rect 1200 3635 1450 3650
rect 1200 3615 1215 3635
rect 1235 3615 1265 3635
rect 1285 3615 1315 3635
rect 1335 3615 1365 3635
rect 1385 3615 1415 3635
rect 1435 3615 1450 3635
rect 1200 3600 1450 3615
rect 1200 3550 1300 3600
rect 1350 3550 1450 3600
rect 1500 3650 1600 3700
rect 1650 3650 1750 3700
rect 1500 3635 1750 3650
rect 1500 3615 1515 3635
rect 1535 3615 1565 3635
rect 1585 3615 1615 3635
rect 1635 3615 1665 3635
rect 1685 3615 1715 3635
rect 1735 3615 1750 3635
rect 1500 3600 1750 3615
rect 1500 3550 1600 3600
rect 1650 3550 1750 3600
rect 1800 3650 1900 3700
rect 1950 3650 2050 3700
rect 1800 3635 2050 3650
rect 1800 3615 1815 3635
rect 1835 3615 1865 3635
rect 1885 3615 1915 3635
rect 1935 3615 1965 3635
rect 1985 3615 2015 3635
rect 2035 3615 2050 3635
rect 1800 3600 2050 3615
rect 1800 3550 1900 3600
rect 1950 3550 2050 3600
rect 2100 3650 2200 3700
rect 2250 3650 2350 3700
rect 2100 3635 2350 3650
rect 2100 3615 2115 3635
rect 2135 3615 2165 3635
rect 2185 3615 2215 3635
rect 2235 3615 2265 3635
rect 2285 3615 2315 3635
rect 2335 3615 2350 3635
rect 2100 3600 2350 3615
rect 2100 3550 2200 3600
rect 2250 3550 2350 3600
rect 2400 3650 2500 3700
rect 2550 3650 2650 3700
rect 2400 3635 2650 3650
rect 2400 3615 2415 3635
rect 2435 3615 2465 3635
rect 2485 3615 2515 3635
rect 2535 3615 2565 3635
rect 2585 3615 2615 3635
rect 2635 3615 2650 3635
rect 2400 3600 2650 3615
rect 2400 3550 2500 3600
rect 2550 3550 2650 3600
rect 2700 3650 2800 3700
rect 2850 3650 2950 3700
rect 2700 3635 2950 3650
rect 2700 3615 2715 3635
rect 2735 3615 2765 3635
rect 2785 3615 2815 3635
rect 2835 3615 2865 3635
rect 2885 3615 2915 3635
rect 2935 3615 2950 3635
rect 2700 3600 2950 3615
rect 2700 3550 2800 3600
rect 2850 3550 2950 3600
rect 3000 3650 3100 3700
rect 3150 3650 3250 3700
rect 3000 3635 3250 3650
rect 3000 3615 3015 3635
rect 3035 3615 3065 3635
rect 3085 3615 3115 3635
rect 3135 3615 3165 3635
rect 3185 3615 3215 3635
rect 3235 3615 3250 3635
rect 3000 3600 3250 3615
rect 3000 3550 3100 3600
rect 3150 3550 3250 3600
rect 3300 3650 3400 3700
rect 3450 3650 3550 3700
rect 3300 3635 3550 3650
rect 3300 3615 3315 3635
rect 3335 3615 3365 3635
rect 3385 3615 3415 3635
rect 3435 3615 3465 3635
rect 3485 3615 3515 3635
rect 3535 3615 3550 3635
rect 3300 3600 3550 3615
rect 3300 3550 3400 3600
rect 3450 3550 3550 3600
rect 3600 3650 3700 3700
rect 3750 3650 3850 3700
rect 3600 3635 3850 3650
rect 3600 3615 3615 3635
rect 3635 3615 3665 3635
rect 3685 3615 3715 3635
rect 3735 3615 3765 3635
rect 3785 3615 3815 3635
rect 3835 3615 3850 3635
rect 3600 3600 3850 3615
rect 3600 3550 3700 3600
rect 3750 3550 3850 3600
rect 3900 3650 4000 3700
rect 4050 3650 4150 3700
rect 3900 3635 4150 3650
rect 3900 3615 3915 3635
rect 3935 3615 3965 3635
rect 3985 3615 4015 3635
rect 4035 3615 4065 3635
rect 4085 3615 4115 3635
rect 4135 3615 4150 3635
rect 3900 3600 4150 3615
rect 3900 3550 4000 3600
rect 4050 3550 4150 3600
rect 4200 3650 4300 3700
rect 4350 3650 4450 3700
rect 4200 3635 4450 3650
rect 4200 3615 4215 3635
rect 4235 3615 4265 3635
rect 4285 3615 4315 3635
rect 4335 3615 4365 3635
rect 4385 3615 4415 3635
rect 4435 3615 4450 3635
rect 4200 3600 4450 3615
rect 4200 3550 4300 3600
rect 4350 3550 4450 3600
rect 4500 3650 4600 3700
rect 4650 3650 4750 3700
rect 4500 3635 4750 3650
rect 4500 3615 4515 3635
rect 4535 3615 4565 3635
rect 4585 3615 4615 3635
rect 4635 3615 4665 3635
rect 4685 3615 4715 3635
rect 4735 3615 4750 3635
rect 4500 3600 4750 3615
rect 4500 3550 4600 3600
rect 4650 3550 4750 3600
rect 4800 3650 4900 3700
rect 4950 3650 5050 3700
rect 4800 3635 5050 3650
rect 4800 3615 4815 3635
rect 4835 3615 4865 3635
rect 4885 3615 4915 3635
rect 4935 3615 4965 3635
rect 4985 3615 5015 3635
rect 5035 3615 5050 3635
rect 4800 3600 5050 3615
rect 4800 3550 4900 3600
rect 4950 3550 5050 3600
rect 5100 3650 5200 3700
rect 5250 3650 5350 3700
rect 5100 3635 5350 3650
rect 5100 3615 5115 3635
rect 5135 3615 5165 3635
rect 5185 3615 5215 3635
rect 5235 3615 5265 3635
rect 5285 3615 5315 3635
rect 5335 3615 5350 3635
rect 5100 3600 5350 3615
rect 5100 3550 5200 3600
rect 5250 3550 5350 3600
rect 5400 3650 5500 3700
rect 5550 3650 5650 3700
rect 5400 3635 5650 3650
rect 5400 3615 5415 3635
rect 5435 3615 5465 3635
rect 5485 3615 5515 3635
rect 5535 3615 5565 3635
rect 5585 3615 5615 3635
rect 5635 3615 5650 3635
rect 5400 3600 5650 3615
rect 5400 3550 5500 3600
rect 5550 3550 5650 3600
rect 5700 3650 5800 3700
rect 5850 3650 5950 3700
rect 5700 3635 5950 3650
rect 5700 3615 5715 3635
rect 5735 3615 5765 3635
rect 5785 3615 5815 3635
rect 5835 3615 5865 3635
rect 5885 3615 5915 3635
rect 5935 3615 5950 3635
rect 5700 3600 5950 3615
rect 5700 3550 5800 3600
rect 5850 3550 5950 3600
rect 6000 3650 6100 3700
rect 6150 3650 6250 3700
rect 6000 3635 6250 3650
rect 6000 3615 6015 3635
rect 6035 3615 6065 3635
rect 6085 3615 6115 3635
rect 6135 3615 6165 3635
rect 6185 3615 6215 3635
rect 6235 3615 6250 3635
rect 6000 3600 6250 3615
rect 6000 3550 6100 3600
rect 6150 3550 6250 3600
rect 6300 3650 6400 3700
rect 6450 3650 6550 3700
rect 6300 3635 6550 3650
rect 6300 3615 6315 3635
rect 6335 3615 6365 3635
rect 6385 3615 6415 3635
rect 6435 3615 6465 3635
rect 6485 3615 6515 3635
rect 6535 3615 6550 3635
rect 6300 3600 6550 3615
rect 6300 3550 6400 3600
rect 6450 3550 6550 3600
rect 6600 3650 6700 3700
rect 6750 3650 6850 3700
rect 6600 3635 6850 3650
rect 6600 3615 6615 3635
rect 6635 3615 6665 3635
rect 6685 3615 6715 3635
rect 6735 3615 6765 3635
rect 6785 3615 6815 3635
rect 6835 3615 6850 3635
rect 6600 3600 6850 3615
rect 6600 3550 6700 3600
rect 6750 3550 6850 3600
rect 6900 3650 7000 3700
rect 7050 3650 7150 3700
rect 6900 3635 7150 3650
rect 6900 3615 6915 3635
rect 6935 3615 6965 3635
rect 6985 3615 7015 3635
rect 7035 3615 7065 3635
rect 7085 3615 7115 3635
rect 7135 3615 7150 3635
rect 6900 3600 7150 3615
rect 6900 3550 7000 3600
rect 7050 3550 7150 3600
rect 7200 3650 7300 3700
rect 7350 3650 7450 3700
rect 7200 3635 7450 3650
rect 7200 3615 7215 3635
rect 7235 3615 7265 3635
rect 7285 3615 7315 3635
rect 7335 3615 7365 3635
rect 7385 3615 7415 3635
rect 7435 3615 7450 3635
rect 7200 3600 7450 3615
rect 7200 3550 7300 3600
rect 7350 3550 7450 3600
rect 7500 3650 7600 3700
rect 7650 3650 7750 3700
rect 7500 3635 7750 3650
rect 7500 3615 7515 3635
rect 7535 3615 7565 3635
rect 7585 3615 7615 3635
rect 7635 3615 7665 3635
rect 7685 3615 7715 3635
rect 7735 3615 7750 3635
rect 7500 3600 7750 3615
rect 7500 3550 7600 3600
rect 7650 3550 7750 3600
rect 7800 3650 7900 3700
rect 7950 3650 8050 3700
rect 7800 3635 8050 3650
rect 7800 3615 7815 3635
rect 7835 3615 7865 3635
rect 7885 3615 7915 3635
rect 7935 3615 7965 3635
rect 7985 3615 8015 3635
rect 8035 3615 8050 3635
rect 7800 3600 8050 3615
rect 7800 3550 7900 3600
rect 7950 3550 8050 3600
rect 8100 3650 8200 3700
rect 8250 3650 8350 3700
rect 8100 3635 8350 3650
rect 8100 3615 8115 3635
rect 8135 3615 8165 3635
rect 8185 3615 8215 3635
rect 8235 3615 8265 3635
rect 8285 3615 8315 3635
rect 8335 3615 8350 3635
rect 8100 3600 8350 3615
rect 8100 3550 8200 3600
rect 8250 3550 8350 3600
rect 8400 3650 8500 3700
rect 8550 3650 8650 3700
rect 8400 3635 8650 3650
rect 8400 3615 8415 3635
rect 8435 3615 8465 3635
rect 8485 3615 8515 3635
rect 8535 3615 8565 3635
rect 8585 3615 8615 3635
rect 8635 3615 8650 3635
rect 8400 3600 8650 3615
rect 8400 3550 8500 3600
rect 8550 3550 8650 3600
rect 8700 3650 8800 3700
rect 8850 3650 8950 3700
rect 8700 3635 8950 3650
rect 8700 3615 8715 3635
rect 8735 3615 8765 3635
rect 8785 3615 8815 3635
rect 8835 3615 8865 3635
rect 8885 3615 8915 3635
rect 8935 3615 8950 3635
rect 8700 3600 8950 3615
rect 8700 3550 8800 3600
rect 8850 3550 8950 3600
rect 9000 3650 9100 3700
rect 9150 3650 9250 3700
rect 9000 3635 9250 3650
rect 9000 3615 9015 3635
rect 9035 3615 9065 3635
rect 9085 3615 9115 3635
rect 9135 3615 9165 3635
rect 9185 3615 9215 3635
rect 9235 3615 9250 3635
rect 9000 3600 9250 3615
rect 9000 3550 9100 3600
rect 9150 3550 9250 3600
rect 9300 3650 9400 3700
rect 9450 3650 9550 3700
rect 9300 3635 9550 3650
rect 9300 3615 9315 3635
rect 9335 3615 9365 3635
rect 9385 3615 9415 3635
rect 9435 3615 9465 3635
rect 9485 3615 9515 3635
rect 9535 3615 9550 3635
rect 9300 3600 9550 3615
rect 9300 3550 9400 3600
rect 9450 3550 9550 3600
rect 9600 3650 9700 3700
rect 9750 3650 9850 3700
rect 9600 3635 9850 3650
rect 9600 3615 9615 3635
rect 9635 3615 9665 3635
rect 9685 3615 9715 3635
rect 9735 3615 9765 3635
rect 9785 3615 9815 3635
rect 9835 3615 9850 3635
rect 9600 3600 9850 3615
rect 9600 3550 9700 3600
rect 9750 3550 9850 3600
rect 9900 3650 10000 3700
rect 10050 3650 10150 3700
rect 9900 3635 10150 3650
rect 9900 3615 9915 3635
rect 9935 3615 9965 3635
rect 9985 3615 10015 3635
rect 10035 3615 10065 3635
rect 10085 3615 10115 3635
rect 10135 3615 10150 3635
rect 9900 3600 10150 3615
rect 9900 3550 10000 3600
rect 10050 3550 10150 3600
rect 10200 3650 10300 3700
rect 10350 3650 10450 3700
rect 10200 3635 10450 3650
rect 10200 3615 10215 3635
rect 10235 3615 10265 3635
rect 10285 3615 10315 3635
rect 10335 3615 10365 3635
rect 10385 3615 10415 3635
rect 10435 3615 10450 3635
rect 10200 3600 10450 3615
rect 10200 3550 10300 3600
rect 10350 3550 10450 3600
rect 10500 3650 10600 3700
rect 10650 3650 10750 3700
rect 10500 3635 10750 3650
rect 10500 3615 10515 3635
rect 10535 3615 10565 3635
rect 10585 3615 10615 3635
rect 10635 3615 10665 3635
rect 10685 3615 10715 3635
rect 10735 3615 10750 3635
rect 10500 3600 10750 3615
rect 10500 3550 10600 3600
rect 10650 3550 10750 3600
rect 10800 3650 10900 3700
rect 10950 3650 11050 3700
rect 10800 3635 11050 3650
rect 10800 3615 10815 3635
rect 10835 3615 10865 3635
rect 10885 3615 10915 3635
rect 10935 3615 10965 3635
rect 10985 3615 11015 3635
rect 11035 3615 11050 3635
rect 10800 3600 11050 3615
rect 10800 3550 10900 3600
rect 10950 3550 11050 3600
rect 11100 3650 11200 3700
rect 11250 3650 11350 3700
rect 11100 3635 11350 3650
rect 11100 3615 11115 3635
rect 11135 3615 11165 3635
rect 11185 3615 11215 3635
rect 11235 3615 11265 3635
rect 11285 3615 11315 3635
rect 11335 3615 11350 3635
rect 11100 3600 11350 3615
rect 11100 3550 11200 3600
rect 11250 3550 11350 3600
rect 11400 3650 11500 3700
rect 11550 3650 11650 3700
rect 11400 3635 11650 3650
rect 11400 3615 11415 3635
rect 11435 3615 11465 3635
rect 11485 3615 11515 3635
rect 11535 3615 11565 3635
rect 11585 3615 11615 3635
rect 11635 3615 11650 3635
rect 11400 3600 11650 3615
rect 11400 3550 11500 3600
rect 11550 3550 11650 3600
rect 11700 3650 11800 3700
rect 11850 3650 11950 3700
rect 11700 3635 11950 3650
rect 11700 3615 11715 3635
rect 11735 3615 11765 3635
rect 11785 3615 11815 3635
rect 11835 3615 11865 3635
rect 11885 3615 11915 3635
rect 11935 3615 11950 3635
rect 11700 3600 11950 3615
rect 11700 3550 11800 3600
rect 11850 3550 11950 3600
rect 12000 3650 12100 3700
rect 12150 3650 12250 3700
rect 12000 3635 12250 3650
rect 12000 3615 12015 3635
rect 12035 3615 12065 3635
rect 12085 3615 12115 3635
rect 12135 3615 12165 3635
rect 12185 3615 12215 3635
rect 12235 3615 12250 3635
rect 12000 3600 12250 3615
rect 12000 3550 12100 3600
rect 12150 3550 12250 3600
rect 12300 3650 12400 3700
rect 12450 3650 12550 3700
rect 12300 3635 12550 3650
rect 12300 3615 12315 3635
rect 12335 3615 12365 3635
rect 12385 3615 12415 3635
rect 12435 3615 12465 3635
rect 12485 3615 12515 3635
rect 12535 3615 12550 3635
rect 12300 3600 12550 3615
rect 12300 3550 12400 3600
rect 12450 3550 12550 3600
rect 12600 3650 12700 3700
rect 12750 3650 12850 3700
rect 12600 3635 12850 3650
rect 12600 3615 12615 3635
rect 12635 3615 12665 3635
rect 12685 3615 12715 3635
rect 12735 3615 12765 3635
rect 12785 3615 12815 3635
rect 12835 3615 12850 3635
rect 12600 3600 12850 3615
rect 12600 3550 12700 3600
rect 12750 3550 12850 3600
rect 12900 3650 13000 3700
rect 13050 3650 13150 3700
rect 12900 3635 13150 3650
rect 12900 3615 12915 3635
rect 12935 3615 12965 3635
rect 12985 3615 13015 3635
rect 13035 3615 13065 3635
rect 13085 3615 13115 3635
rect 13135 3615 13150 3635
rect 12900 3600 13150 3615
rect 12900 3550 13000 3600
rect 13050 3550 13150 3600
rect 13200 3650 13300 3700
rect 13350 3650 13450 3700
rect 13200 3635 13450 3650
rect 13200 3615 13215 3635
rect 13235 3615 13265 3635
rect 13285 3615 13315 3635
rect 13335 3615 13365 3635
rect 13385 3615 13415 3635
rect 13435 3615 13450 3635
rect 13200 3600 13450 3615
rect 13200 3550 13300 3600
rect 13350 3550 13450 3600
rect 13500 3650 13600 3700
rect 13650 3650 13750 3700
rect 13500 3635 13750 3650
rect 13500 3615 13515 3635
rect 13535 3615 13565 3635
rect 13585 3615 13615 3635
rect 13635 3615 13665 3635
rect 13685 3615 13715 3635
rect 13735 3615 13750 3635
rect 13500 3600 13750 3615
rect 13500 3550 13600 3600
rect 13650 3550 13750 3600
rect 13800 3650 13900 3700
rect 13950 3650 14050 3700
rect 13800 3635 14050 3650
rect 13800 3615 13815 3635
rect 13835 3615 13865 3635
rect 13885 3615 13915 3635
rect 13935 3615 13965 3635
rect 13985 3615 14015 3635
rect 14035 3615 14050 3635
rect 13800 3600 14050 3615
rect 13800 3550 13900 3600
rect 13950 3550 14050 3600
rect 14100 3650 14200 3700
rect 14250 3650 14350 3700
rect 14100 3635 14350 3650
rect 14100 3615 14115 3635
rect 14135 3615 14165 3635
rect 14185 3615 14215 3635
rect 14235 3615 14265 3635
rect 14285 3615 14315 3635
rect 14335 3615 14350 3635
rect 14100 3600 14350 3615
rect 14100 3550 14200 3600
rect 14250 3550 14350 3600
rect 14400 3650 14500 3700
rect 14550 3650 14650 3700
rect 14400 3635 14650 3650
rect 14400 3615 14415 3635
rect 14435 3615 14465 3635
rect 14485 3615 14515 3635
rect 14535 3615 14565 3635
rect 14585 3615 14615 3635
rect 14635 3615 14650 3635
rect 14400 3600 14650 3615
rect 14400 3550 14500 3600
rect 14550 3550 14650 3600
rect 14700 3650 14800 3700
rect 14850 3650 14950 3700
rect 14700 3635 14950 3650
rect 14700 3615 14715 3635
rect 14735 3615 14765 3635
rect 14785 3615 14815 3635
rect 14835 3615 14865 3635
rect 14885 3615 14915 3635
rect 14935 3615 14950 3635
rect 14700 3600 14950 3615
rect 14700 3550 14800 3600
rect 14850 3550 14950 3600
rect 15000 3650 15100 3700
rect 15150 3650 15250 3700
rect 15000 3635 15250 3650
rect 15000 3615 15015 3635
rect 15035 3615 15065 3635
rect 15085 3615 15115 3635
rect 15135 3615 15165 3635
rect 15185 3615 15215 3635
rect 15235 3615 15250 3635
rect 15000 3600 15250 3615
rect 15000 3550 15100 3600
rect 15150 3550 15250 3600
rect 15300 3650 15400 3700
rect 15450 3650 15550 3700
rect 15300 3635 15550 3650
rect 15300 3615 15315 3635
rect 15335 3615 15365 3635
rect 15385 3615 15415 3635
rect 15435 3615 15465 3635
rect 15485 3615 15515 3635
rect 15535 3615 15550 3635
rect 15300 3600 15550 3615
rect 15300 3550 15400 3600
rect 15450 3550 15550 3600
rect 15600 3650 15700 3700
rect 15750 3650 15850 3700
rect 15600 3635 15850 3650
rect 15600 3615 15615 3635
rect 15635 3615 15665 3635
rect 15685 3615 15715 3635
rect 15735 3615 15765 3635
rect 15785 3615 15815 3635
rect 15835 3615 15850 3635
rect 15600 3600 15850 3615
rect 15600 3550 15700 3600
rect 15750 3550 15850 3600
rect 15900 3650 16000 3700
rect 16050 3650 16150 3700
rect 15900 3635 16150 3650
rect 15900 3615 15915 3635
rect 15935 3615 15965 3635
rect 15985 3615 16015 3635
rect 16035 3615 16065 3635
rect 16085 3615 16115 3635
rect 16135 3615 16150 3635
rect 15900 3600 16150 3615
rect 15900 3550 16000 3600
rect 16050 3550 16150 3600
rect 16200 3650 16300 3700
rect 16350 3650 16450 3700
rect 16200 3635 16450 3650
rect 16200 3615 16215 3635
rect 16235 3615 16265 3635
rect 16285 3615 16315 3635
rect 16335 3615 16365 3635
rect 16385 3615 16415 3635
rect 16435 3615 16450 3635
rect 16200 3600 16450 3615
rect 16200 3550 16300 3600
rect 16350 3550 16450 3600
rect 16500 3650 16600 3700
rect 16650 3650 16750 3700
rect 16500 3635 16750 3650
rect 16500 3615 16515 3635
rect 16535 3615 16565 3635
rect 16585 3615 16615 3635
rect 16635 3615 16665 3635
rect 16685 3615 16715 3635
rect 16735 3615 16750 3635
rect 16500 3600 16750 3615
rect 16500 3550 16600 3600
rect 16650 3550 16750 3600
rect 16800 3650 16900 3700
rect 16950 3650 17050 3700
rect 16800 3635 17050 3650
rect 16800 3615 16815 3635
rect 16835 3615 16865 3635
rect 16885 3615 16915 3635
rect 16935 3615 16965 3635
rect 16985 3615 17015 3635
rect 17035 3615 17050 3635
rect 16800 3600 17050 3615
rect 16800 3550 16900 3600
rect 16950 3550 17050 3600
rect 17100 3650 17200 3700
rect 17250 3650 17350 3700
rect 17100 3635 17350 3650
rect 17100 3615 17115 3635
rect 17135 3615 17165 3635
rect 17185 3615 17215 3635
rect 17235 3615 17265 3635
rect 17285 3615 17315 3635
rect 17335 3615 17350 3635
rect 17100 3600 17350 3615
rect 17100 3550 17200 3600
rect 17250 3550 17350 3600
rect 17400 3650 17500 3700
rect 17550 3650 17650 3700
rect 17400 3635 17650 3650
rect 17400 3615 17415 3635
rect 17435 3615 17465 3635
rect 17485 3615 17515 3635
rect 17535 3615 17565 3635
rect 17585 3615 17615 3635
rect 17635 3615 17650 3635
rect 17400 3600 17650 3615
rect 17400 3550 17500 3600
rect 17550 3550 17650 3600
rect 17700 3650 17800 3700
rect 17850 3650 17950 3700
rect 17700 3635 17950 3650
rect 17700 3615 17715 3635
rect 17735 3615 17765 3635
rect 17785 3615 17815 3635
rect 17835 3615 17865 3635
rect 17885 3615 17915 3635
rect 17935 3615 17950 3635
rect 17700 3600 17950 3615
rect 17700 3550 17800 3600
rect 17850 3550 17950 3600
rect 18000 3650 18100 3700
rect 18150 3650 18250 3700
rect 18000 3635 18250 3650
rect 18000 3615 18015 3635
rect 18035 3615 18065 3635
rect 18085 3615 18115 3635
rect 18135 3615 18165 3635
rect 18185 3615 18215 3635
rect 18235 3615 18250 3635
rect 18000 3600 18250 3615
rect 18000 3550 18100 3600
rect 18150 3550 18250 3600
rect 18300 3650 18400 3700
rect 18450 3650 18550 3700
rect 18300 3635 18550 3650
rect 18300 3615 18315 3635
rect 18335 3615 18365 3635
rect 18385 3615 18415 3635
rect 18435 3615 18465 3635
rect 18485 3615 18515 3635
rect 18535 3615 18550 3635
rect 18300 3600 18550 3615
rect 18300 3550 18400 3600
rect 18450 3550 18550 3600
rect 18600 3650 18700 3700
rect 18750 3650 18850 3700
rect 18600 3635 18850 3650
rect 18600 3615 18615 3635
rect 18635 3615 18665 3635
rect 18685 3615 18715 3635
rect 18735 3615 18765 3635
rect 18785 3615 18815 3635
rect 18835 3615 18850 3635
rect 18600 3600 18850 3615
rect 18600 3550 18700 3600
rect 18750 3550 18850 3600
rect 18900 3650 19000 3700
rect 19050 3650 19150 3700
rect 18900 3635 19150 3650
rect 18900 3615 18915 3635
rect 18935 3615 18965 3635
rect 18985 3615 19015 3635
rect 19035 3615 19065 3635
rect 19085 3615 19115 3635
rect 19135 3615 19150 3635
rect 18900 3600 19150 3615
rect 18900 3550 19000 3600
rect 19050 3550 19150 3600
rect 19200 3650 19300 3700
rect 19350 3650 19450 3700
rect 19200 3635 19450 3650
rect 19200 3615 19215 3635
rect 19235 3615 19265 3635
rect 19285 3615 19315 3635
rect 19335 3615 19365 3635
rect 19385 3615 19415 3635
rect 19435 3615 19450 3635
rect 19200 3600 19450 3615
rect 19200 3550 19300 3600
rect 19350 3550 19450 3600
rect 19500 3650 19600 3700
rect 19650 3650 19750 3700
rect 19500 3635 19750 3650
rect 19500 3615 19515 3635
rect 19535 3615 19565 3635
rect 19585 3615 19615 3635
rect 19635 3615 19665 3635
rect 19685 3615 19715 3635
rect 19735 3615 19750 3635
rect 19500 3600 19750 3615
rect 19500 3550 19600 3600
rect 19650 3550 19750 3600
rect 19800 3650 19900 3700
rect 19950 3650 20050 3700
rect 19800 3635 20050 3650
rect 19800 3615 19815 3635
rect 19835 3615 19865 3635
rect 19885 3615 19915 3635
rect 19935 3615 19965 3635
rect 19985 3615 20015 3635
rect 20035 3615 20050 3635
rect 19800 3600 20050 3615
rect 19800 3550 19900 3600
rect 19950 3550 20050 3600
rect 20100 3650 20200 3700
rect 20250 3650 20350 3700
rect 20100 3635 20350 3650
rect 20100 3615 20115 3635
rect 20135 3615 20165 3635
rect 20185 3615 20215 3635
rect 20235 3615 20265 3635
rect 20285 3615 20315 3635
rect 20335 3615 20350 3635
rect 20100 3600 20350 3615
rect 20100 3550 20200 3600
rect 20250 3550 20350 3600
rect 20400 3650 20500 3700
rect 20550 3650 20650 3700
rect 20400 3635 20650 3650
rect 20400 3615 20415 3635
rect 20435 3615 20465 3635
rect 20485 3615 20515 3635
rect 20535 3615 20565 3635
rect 20585 3615 20615 3635
rect 20635 3615 20650 3635
rect 20400 3600 20650 3615
rect 20400 3550 20500 3600
rect 20550 3550 20650 3600
rect 20700 3650 20800 3700
rect 20850 3650 20950 3700
rect 20700 3635 20950 3650
rect 20700 3615 20715 3635
rect 20735 3615 20765 3635
rect 20785 3615 20815 3635
rect 20835 3615 20865 3635
rect 20885 3615 20915 3635
rect 20935 3615 20950 3635
rect 20700 3600 20950 3615
rect 20700 3550 20800 3600
rect 20850 3550 20950 3600
rect 21000 3650 21100 3700
rect 21150 3650 21250 3700
rect 21300 3650 21400 3700
rect 21000 3635 21400 3650
rect 21000 3615 21015 3635
rect 21035 3615 21065 3635
rect 21085 3615 21115 3635
rect 21135 3615 21165 3635
rect 21185 3615 21215 3635
rect 21235 3615 21265 3635
rect 21285 3615 21315 3635
rect 21335 3615 21365 3635
rect 21385 3615 21400 3635
rect 21000 3600 21400 3615
rect 21000 3550 21100 3600
rect 21150 3550 21250 3600
rect 21300 3550 21400 3600
rect 21450 3650 21550 3700
rect 21600 3650 21700 3700
rect 21750 3650 21850 3700
rect 21450 3635 21850 3650
rect 21450 3615 21465 3635
rect 21485 3615 21515 3635
rect 21535 3615 21565 3635
rect 21585 3615 21615 3635
rect 21635 3615 21665 3635
rect 21685 3615 21715 3635
rect 21735 3615 21765 3635
rect 21785 3615 21815 3635
rect 21835 3615 21850 3635
rect 21450 3600 21850 3615
rect 21450 3550 21550 3600
rect 21600 3550 21700 3600
rect 21750 3550 21850 3600
rect 21900 3650 22000 3700
rect 22050 3650 22150 3700
rect 21900 3635 22150 3650
rect 21900 3615 21915 3635
rect 21935 3615 21965 3635
rect 21985 3615 22015 3635
rect 22035 3615 22065 3635
rect 22085 3615 22115 3635
rect 22135 3615 22150 3635
rect 21900 3600 22150 3615
rect 21900 3550 22000 3600
rect 22050 3550 22150 3600
rect 22200 3650 22300 3700
rect 22350 3650 22450 3700
rect 22200 3635 22450 3650
rect 22200 3615 22215 3635
rect 22235 3615 22265 3635
rect 22285 3615 22315 3635
rect 22335 3615 22365 3635
rect 22385 3615 22415 3635
rect 22435 3615 22450 3635
rect 22200 3600 22450 3615
rect 22200 3550 22300 3600
rect 22350 3550 22450 3600
rect 22500 3650 22600 3700
rect 22650 3650 22750 3700
rect 22500 3635 22750 3650
rect 22500 3615 22515 3635
rect 22535 3615 22565 3635
rect 22585 3615 22615 3635
rect 22635 3615 22665 3635
rect 22685 3615 22715 3635
rect 22735 3615 22750 3635
rect 22500 3600 22750 3615
rect 22500 3550 22600 3600
rect 22650 3550 22750 3600
rect 22800 3650 22900 3700
rect 22950 3650 23050 3700
rect 22800 3635 23050 3650
rect 22800 3615 22815 3635
rect 22835 3615 22865 3635
rect 22885 3615 22915 3635
rect 22935 3615 22965 3635
rect 22985 3615 23015 3635
rect 23035 3615 23050 3635
rect 22800 3600 23050 3615
rect 22800 3550 22900 3600
rect 22950 3550 23050 3600
rect 23100 3650 23200 3700
rect 23250 3650 23350 3700
rect 23400 3650 23500 3700
rect 23100 3635 23500 3650
rect 23100 3615 23115 3635
rect 23135 3615 23165 3635
rect 23185 3615 23215 3635
rect 23235 3615 23265 3635
rect 23285 3615 23315 3635
rect 23335 3615 23365 3635
rect 23385 3615 23415 3635
rect 23435 3615 23465 3635
rect 23485 3615 23500 3635
rect 23100 3600 23500 3615
rect 23100 3550 23200 3600
rect 23250 3550 23350 3600
rect 23400 3550 23500 3600
rect 23550 3650 23650 3700
rect 23700 3650 23800 3700
rect 23850 3650 23950 3700
rect 23550 3635 23950 3650
rect 23550 3615 23565 3635
rect 23585 3615 23615 3635
rect 23635 3615 23665 3635
rect 23685 3615 23715 3635
rect 23735 3615 23765 3635
rect 23785 3615 23815 3635
rect 23835 3615 23865 3635
rect 23885 3615 23915 3635
rect 23935 3615 23950 3635
rect 23550 3600 23950 3615
rect 23550 3550 23650 3600
rect 23700 3550 23800 3600
rect 23850 3550 23950 3600
rect 24000 3650 24100 3700
rect 24150 3650 24250 3700
rect 24000 3635 24250 3650
rect 24000 3615 24015 3635
rect 24035 3615 24065 3635
rect 24085 3615 24115 3635
rect 24135 3615 24165 3635
rect 24185 3615 24215 3635
rect 24235 3615 24250 3635
rect 24000 3600 24250 3615
rect 24000 3550 24100 3600
rect 24150 3550 24250 3600
rect 24300 3650 24400 3700
rect 24450 3650 24550 3700
rect 24300 3635 24550 3650
rect 24300 3615 24315 3635
rect 24335 3615 24365 3635
rect 24385 3615 24415 3635
rect 24435 3615 24465 3635
rect 24485 3615 24515 3635
rect 24535 3615 24550 3635
rect 24300 3600 24550 3615
rect 24300 3550 24400 3600
rect 24450 3550 24550 3600
rect 24600 3650 24700 3700
rect 24750 3650 24850 3700
rect 24600 3635 24850 3650
rect 24600 3615 24615 3635
rect 24635 3615 24665 3635
rect 24685 3615 24715 3635
rect 24735 3615 24765 3635
rect 24785 3615 24815 3635
rect 24835 3615 24850 3635
rect 24600 3600 24850 3615
rect 24600 3550 24700 3600
rect 24750 3550 24850 3600
rect 24900 3650 25000 3700
rect 25050 3650 25150 3700
rect 24900 3635 25150 3650
rect 24900 3615 24915 3635
rect 24935 3615 24965 3635
rect 24985 3615 25015 3635
rect 25035 3615 25065 3635
rect 25085 3615 25115 3635
rect 25135 3615 25150 3635
rect 24900 3600 25150 3615
rect 24900 3550 25000 3600
rect 25050 3550 25150 3600
rect 25200 3650 25300 3700
rect 25350 3650 25450 3700
rect 25500 3650 25600 3700
rect 25200 3635 25600 3650
rect 25200 3615 25215 3635
rect 25235 3615 25265 3635
rect 25285 3615 25315 3635
rect 25335 3615 25365 3635
rect 25385 3615 25415 3635
rect 25435 3615 25465 3635
rect 25485 3615 25515 3635
rect 25535 3615 25565 3635
rect 25585 3615 25600 3635
rect 25200 3600 25600 3615
rect 25200 3550 25300 3600
rect 25350 3550 25450 3600
rect 25500 3550 25600 3600
rect 25650 3650 25750 3700
rect 25800 3650 25900 3700
rect 25950 3650 26050 3700
rect 25650 3635 26050 3650
rect 25650 3615 25665 3635
rect 25685 3615 25715 3635
rect 25735 3615 25765 3635
rect 25785 3615 25815 3635
rect 25835 3615 25865 3635
rect 25885 3615 25915 3635
rect 25935 3615 25965 3635
rect 25985 3615 26015 3635
rect 26035 3615 26050 3635
rect 25650 3600 26050 3615
rect 25650 3550 25750 3600
rect 25800 3550 25900 3600
rect 25950 3550 26050 3600
rect 26100 3650 26200 3700
rect 26250 3650 26350 3700
rect 26100 3635 26350 3650
rect 26100 3615 26115 3635
rect 26135 3615 26165 3635
rect 26185 3615 26215 3635
rect 26235 3615 26265 3635
rect 26285 3615 26315 3635
rect 26335 3615 26350 3635
rect 26100 3600 26350 3615
rect 26100 3550 26200 3600
rect 26250 3550 26350 3600
rect 26400 3650 26500 3700
rect 26550 3650 26650 3700
rect 26400 3635 26650 3650
rect 26400 3615 26415 3635
rect 26435 3615 26465 3635
rect 26485 3615 26515 3635
rect 26535 3615 26565 3635
rect 26585 3615 26615 3635
rect 26635 3615 26650 3635
rect 26400 3600 26650 3615
rect 26400 3550 26500 3600
rect 26550 3550 26650 3600
rect 26700 3650 26800 3700
rect 26850 3650 26950 3700
rect 26700 3635 26950 3650
rect 26700 3615 26715 3635
rect 26735 3615 26765 3635
rect 26785 3615 26815 3635
rect 26835 3615 26865 3635
rect 26885 3615 26915 3635
rect 26935 3615 26950 3635
rect 26700 3600 26950 3615
rect 26700 3550 26800 3600
rect 26850 3550 26950 3600
rect 27000 3650 27100 3700
rect 27150 3650 27250 3700
rect 27000 3635 27250 3650
rect 27000 3615 27015 3635
rect 27035 3615 27065 3635
rect 27085 3615 27115 3635
rect 27135 3615 27165 3635
rect 27185 3615 27215 3635
rect 27235 3615 27250 3635
rect 27000 3600 27250 3615
rect 27000 3550 27100 3600
rect 27150 3550 27250 3600
rect 27300 3650 27400 3700
rect 27450 3650 27550 3700
rect 27600 3650 27700 3700
rect 27300 3635 27700 3650
rect 27300 3615 27315 3635
rect 27335 3615 27365 3635
rect 27385 3615 27415 3635
rect 27435 3615 27465 3635
rect 27485 3615 27515 3635
rect 27535 3615 27565 3635
rect 27585 3615 27615 3635
rect 27635 3615 27665 3635
rect 27685 3615 27700 3635
rect 27300 3600 27700 3615
rect 27300 3550 27400 3600
rect 27450 3550 27550 3600
rect 27600 3550 27700 3600
rect 27750 3650 27850 3700
rect 27900 3650 28000 3700
rect 28050 3650 28150 3700
rect 27750 3635 28150 3650
rect 27750 3615 27765 3635
rect 27785 3615 27815 3635
rect 27835 3615 27865 3635
rect 27885 3615 27915 3635
rect 27935 3615 27965 3635
rect 27985 3615 28015 3635
rect 28035 3615 28065 3635
rect 28085 3615 28115 3635
rect 28135 3615 28150 3635
rect 27750 3600 28150 3615
rect 27750 3550 27850 3600
rect 27900 3550 28000 3600
rect 28050 3550 28150 3600
rect 28200 3650 28300 3700
rect 28350 3650 28450 3700
rect 28200 3635 28450 3650
rect 28200 3615 28215 3635
rect 28235 3615 28265 3635
rect 28285 3615 28315 3635
rect 28335 3615 28365 3635
rect 28385 3615 28415 3635
rect 28435 3615 28450 3635
rect 28200 3600 28450 3615
rect 28200 3550 28300 3600
rect 28350 3550 28450 3600
rect 28500 3650 28600 3700
rect 28650 3650 28750 3700
rect 28500 3635 28750 3650
rect 28500 3615 28515 3635
rect 28535 3615 28565 3635
rect 28585 3615 28615 3635
rect 28635 3615 28665 3635
rect 28685 3615 28715 3635
rect 28735 3615 28750 3635
rect 28500 3600 28750 3615
rect 28500 3550 28600 3600
rect 28650 3550 28750 3600
rect 28800 3650 28900 3700
rect 28950 3650 29050 3700
rect 28800 3635 29050 3650
rect 28800 3615 28815 3635
rect 28835 3615 28865 3635
rect 28885 3615 28915 3635
rect 28935 3615 28965 3635
rect 28985 3615 29015 3635
rect 29035 3615 29050 3635
rect 28800 3600 29050 3615
rect 28800 3550 28900 3600
rect 28950 3550 29050 3600
rect 29100 3650 29200 3700
rect 29250 3650 29350 3700
rect 29100 3635 29350 3650
rect 29100 3615 29115 3635
rect 29135 3615 29165 3635
rect 29185 3615 29215 3635
rect 29235 3615 29265 3635
rect 29285 3615 29315 3635
rect 29335 3615 29350 3635
rect 29100 3600 29350 3615
rect 29100 3550 29200 3600
rect 29250 3550 29350 3600
rect 29400 3650 29500 3700
rect 29550 3650 29650 3700
rect 29700 3650 29800 3700
rect 29400 3635 29800 3650
rect 29400 3615 29415 3635
rect 29435 3615 29465 3635
rect 29485 3615 29515 3635
rect 29535 3615 29565 3635
rect 29585 3615 29615 3635
rect 29635 3615 29665 3635
rect 29685 3615 29715 3635
rect 29735 3615 29765 3635
rect 29785 3615 29800 3635
rect 29400 3600 29800 3615
rect 29400 3550 29500 3600
rect 29550 3550 29650 3600
rect 29700 3550 29800 3600
rect 29850 3650 29950 3700
rect 30000 3650 30100 3700
rect 29850 3635 30100 3650
rect 29850 3615 29865 3635
rect 29885 3615 29915 3635
rect 29935 3615 29965 3635
rect 29985 3615 30015 3635
rect 30035 3615 30065 3635
rect 30085 3615 30100 3635
rect 29850 3600 30100 3615
rect 29850 3550 29950 3600
rect 30000 3550 30100 3600
rect 30150 3650 30250 3700
rect 30300 3650 30400 3700
rect 30150 3635 30400 3650
rect 30150 3615 30165 3635
rect 30185 3615 30215 3635
rect 30235 3615 30265 3635
rect 30285 3615 30315 3635
rect 30335 3615 30365 3635
rect 30385 3615 30400 3635
rect 30150 3600 30400 3615
rect 30150 3550 30250 3600
rect 30300 3550 30400 3600
rect 30450 3650 30550 3700
rect 30600 3650 30700 3700
rect 30450 3635 30700 3650
rect 30450 3615 30465 3635
rect 30485 3615 30515 3635
rect 30535 3615 30565 3635
rect 30585 3615 30615 3635
rect 30635 3615 30665 3635
rect 30685 3615 30700 3635
rect 30450 3600 30700 3615
rect 30450 3550 30550 3600
rect 30600 3550 30700 3600
rect 30750 3650 30850 3700
rect 30900 3650 31000 3700
rect 30750 3635 31000 3650
rect 30750 3615 30765 3635
rect 30785 3615 30815 3635
rect 30835 3615 30865 3635
rect 30885 3615 30915 3635
rect 30935 3615 30965 3635
rect 30985 3615 31000 3635
rect 30750 3600 31000 3615
rect 30750 3550 30850 3600
rect 30900 3550 31000 3600
rect 31050 3650 31150 3700
rect 31200 3650 31300 3700
rect 31350 3650 31450 3700
rect 31050 3635 31450 3650
rect 31050 3615 31065 3635
rect 31085 3615 31115 3635
rect 31135 3615 31165 3635
rect 31185 3615 31215 3635
rect 31235 3615 31265 3635
rect 31285 3615 31315 3635
rect 31335 3615 31365 3635
rect 31385 3615 31415 3635
rect 31435 3615 31450 3635
rect 31050 3600 31450 3615
rect 31050 3550 31150 3600
rect 31200 3550 31300 3600
rect 31350 3550 31450 3600
rect 31500 3650 31600 3700
rect 31650 3650 31750 3700
rect 31500 3635 31750 3650
rect 31500 3615 31515 3635
rect 31535 3615 31565 3635
rect 31585 3615 31615 3635
rect 31635 3615 31665 3635
rect 31685 3615 31715 3635
rect 31735 3615 31750 3635
rect 31500 3600 31750 3615
rect 31500 3550 31600 3600
rect 31650 3550 31750 3600
rect 31800 3650 31900 3700
rect 31950 3650 32050 3700
rect 31800 3635 32050 3650
rect 31800 3615 31815 3635
rect 31835 3615 31865 3635
rect 31885 3615 31915 3635
rect 31935 3615 31965 3635
rect 31985 3615 32015 3635
rect 32035 3615 32050 3635
rect 31800 3600 32050 3615
rect 31800 3550 31900 3600
rect 31950 3550 32050 3600
rect -600 3035 -500 3050
rect -450 3035 -350 3050
rect -300 3035 -200 3050
rect -150 3035 -50 3050
rect 0 3035 100 3050
rect 150 3035 250 3050
rect 300 3035 400 3050
rect 450 3035 550 3050
rect 600 3035 700 3050
rect 750 3035 850 3050
rect 900 3035 1000 3050
rect 1050 3035 1150 3050
rect 1200 3035 1300 3050
rect 1350 3035 1450 3050
rect 1500 3035 1600 3050
rect 1650 3035 1750 3050
rect 1800 3035 1900 3050
rect 1950 3035 2050 3050
rect 2100 3035 2200 3050
rect 2250 3035 2350 3050
rect 2400 3035 2500 3050
rect 2550 3035 2650 3050
rect 2700 3035 2800 3050
rect 2850 3035 2950 3050
rect 3000 3035 3100 3050
rect 3150 3035 3250 3050
rect 3300 3035 3400 3050
rect 3450 3035 3550 3050
rect 3600 3035 3700 3050
rect 3750 3035 3850 3050
rect 3900 3035 4000 3050
rect 4050 3035 4150 3050
rect 4200 3035 4300 3050
rect 4350 3035 4450 3050
rect 4500 3035 4600 3050
rect 4650 3035 4750 3050
rect 4800 3035 4900 3050
rect 4950 3035 5050 3050
rect 5100 3035 5200 3050
rect 5250 3035 5350 3050
rect 5400 3035 5500 3050
rect 5550 3035 5650 3050
rect 5700 3035 5800 3050
rect 5850 3035 5950 3050
rect 6000 3035 6100 3050
rect 6150 3035 6250 3050
rect 6300 3035 6400 3050
rect 6450 3035 6550 3050
rect 6600 3035 6700 3050
rect 6750 3035 6850 3050
rect 6900 3035 7000 3050
rect 7050 3035 7150 3050
rect 7200 3035 7300 3050
rect 7350 3035 7450 3050
rect 7500 3035 7600 3050
rect 7650 3035 7750 3050
rect 7800 3035 7900 3050
rect 7950 3035 8050 3050
rect 8100 3035 8200 3050
rect 8250 3035 8350 3050
rect 8400 3035 8500 3050
rect 8550 3035 8650 3050
rect 8700 3035 8800 3050
rect 8850 3035 8950 3050
rect 9000 3035 9100 3050
rect 9150 3035 9250 3050
rect 9300 3035 9400 3050
rect 9450 3035 9550 3050
rect 9600 3035 9700 3050
rect 9750 3035 9850 3050
rect 9900 3035 10000 3050
rect 10050 3035 10150 3050
rect 10200 3035 10300 3050
rect 10350 3035 10450 3050
rect 10500 3035 10600 3050
rect 10650 3035 10750 3050
rect 10800 3035 10900 3050
rect 10950 3035 11050 3050
rect 11100 3035 11200 3050
rect 11250 3035 11350 3050
rect 11400 3035 11500 3050
rect 11550 3035 11650 3050
rect 11700 3035 11800 3050
rect 11850 3035 11950 3050
rect 12000 3035 12100 3050
rect 12150 3035 12250 3050
rect 12300 3035 12400 3050
rect 12450 3035 12550 3050
rect 12600 3035 12700 3050
rect 12750 3035 12850 3050
rect 12900 3035 13000 3050
rect 13050 3035 13150 3050
rect 13200 3035 13300 3050
rect 13350 3035 13450 3050
rect 13500 3035 13600 3050
rect 13650 3035 13750 3050
rect 13800 3035 13900 3050
rect 13950 3035 14050 3050
rect 14100 3035 14200 3050
rect 14250 3035 14350 3050
rect 14400 3035 14500 3050
rect 14550 3035 14650 3050
rect 14700 3035 14800 3050
rect 14850 3035 14950 3050
rect 15000 3035 15100 3050
rect 15150 3035 15250 3050
rect 15300 3035 15400 3050
rect 15450 3035 15550 3050
rect 15600 3035 15700 3050
rect 15750 3035 15850 3050
rect 15900 3035 16000 3050
rect 16050 3035 16150 3050
rect 16200 3035 16300 3050
rect 16350 3035 16450 3050
rect 16500 3035 16600 3050
rect 16650 3035 16750 3050
rect 16800 3035 16900 3050
rect 16950 3035 17050 3050
rect 17100 3035 17200 3050
rect 17250 3035 17350 3050
rect 17400 3035 17500 3050
rect 17550 3035 17650 3050
rect 17700 3035 17800 3050
rect 17850 3035 17950 3050
rect 18000 3035 18100 3050
rect 18150 3035 18250 3050
rect 18300 3035 18400 3050
rect 18450 3035 18550 3050
rect 18600 3035 18700 3050
rect 18750 3035 18850 3050
rect 18900 3035 19000 3050
rect 19050 3035 19150 3050
rect 19200 3035 19300 3050
rect 19350 3035 19450 3050
rect 19500 3035 19600 3050
rect 19650 3035 19750 3050
rect 19800 3035 19900 3050
rect 19950 3035 20050 3050
rect 20100 3035 20200 3050
rect 20250 3035 20350 3050
rect 20400 3035 20500 3050
rect 20550 3035 20650 3050
rect 20700 3035 20800 3050
rect 20850 3035 20950 3050
rect 21000 3035 21100 3050
rect 21150 3035 21250 3050
rect 21300 3035 21400 3050
rect 21450 3035 21550 3050
rect 21600 3035 21700 3050
rect 21750 3035 21850 3050
rect 21900 3035 22000 3050
rect 22050 3035 22150 3050
rect 22200 3035 22300 3050
rect 22350 3035 22450 3050
rect 22500 3035 22600 3050
rect 22650 3035 22750 3050
rect 22800 3035 22900 3050
rect 22950 3035 23050 3050
rect 23100 3035 23200 3050
rect 23250 3035 23350 3050
rect 23400 3035 23500 3050
rect 23550 3035 23650 3050
rect 23700 3035 23800 3050
rect 23850 3035 23950 3050
rect 24000 3035 24100 3050
rect 24150 3035 24250 3050
rect 24300 3035 24400 3050
rect 24450 3035 24550 3050
rect 24600 3035 24700 3050
rect 24750 3035 24850 3050
rect 24900 3035 25000 3050
rect 25050 3035 25150 3050
rect 25200 3035 25300 3050
rect 25350 3035 25450 3050
rect 25500 3035 25600 3050
rect 25650 3035 25750 3050
rect 25800 3035 25900 3050
rect 25950 3035 26050 3050
rect 26100 3035 26200 3050
rect 26250 3035 26350 3050
rect 26400 3035 26500 3050
rect 26550 3035 26650 3050
rect 26700 3035 26800 3050
rect 26850 3035 26950 3050
rect 27000 3035 27100 3050
rect 27150 3035 27250 3050
rect 27300 3035 27400 3050
rect 27450 3035 27550 3050
rect 27600 3035 27700 3050
rect 27750 3035 27850 3050
rect 27900 3035 28000 3050
rect 28050 3035 28150 3050
rect 28200 3035 28300 3050
rect 28350 3035 28450 3050
rect 28500 3035 28600 3050
rect 28650 3035 28750 3050
rect 28800 3035 28900 3050
rect 28950 3035 29050 3050
rect 29100 3035 29200 3050
rect 29250 3035 29350 3050
rect 29400 3035 29500 3050
rect 29550 3035 29650 3050
rect 29700 3035 29800 3050
rect 29850 3035 29950 3050
rect 30000 3035 30100 3050
rect 30150 3035 30250 3050
rect 30300 3035 30400 3050
rect 30450 3035 30550 3050
rect 30600 3035 30700 3050
rect 30750 3035 30850 3050
rect 30900 3035 31000 3050
rect 31050 3035 31150 3050
rect 31200 3035 31300 3050
rect 31350 3035 31450 3050
rect 31500 3035 31600 3050
rect 31650 3035 31750 3050
rect 31800 3035 31900 3050
rect 31950 3035 32050 3050
rect -600 1600 -500 1615
rect -450 1600 -350 1615
rect -300 1600 -200 1615
rect -150 1600 -50 1615
rect 0 1600 100 1615
rect 150 1600 250 1615
rect 300 1600 400 1615
rect 450 1600 550 1615
rect 600 1600 700 1615
rect 750 1600 850 1615
rect 900 1600 1000 1615
rect 1050 1600 1150 1615
rect 1200 1600 1300 1615
rect 1350 1600 1450 1615
rect 1500 1600 1600 1615
rect 1650 1600 1750 1615
rect 1800 1600 1900 1615
rect 1950 1600 2050 1615
rect 2100 1600 2200 1615
rect 2250 1600 2350 1615
rect 2400 1600 2500 1615
rect 2550 1600 2650 1615
rect 2700 1600 2800 1615
rect 2850 1600 2950 1615
rect 3000 1600 3100 1615
rect 3150 1600 3250 1615
rect 3300 1600 3400 1615
rect 3450 1600 3550 1615
rect 3600 1600 3700 1615
rect 3750 1600 3850 1615
rect 3900 1600 4000 1615
rect 4050 1600 4150 1615
rect 4200 1600 4300 1615
rect 4350 1600 4450 1615
rect 4500 1600 4600 1615
rect 4650 1600 4750 1615
rect 4800 1600 4900 1615
rect 4950 1600 5050 1615
rect 5100 1600 5200 1615
rect 5250 1600 5350 1615
rect 5400 1600 5500 1615
rect 5550 1600 5650 1615
rect 5700 1600 5800 1615
rect 5850 1600 5950 1615
rect 6000 1600 6100 1615
rect 6150 1600 6250 1615
rect 6300 1600 6400 1615
rect 6450 1600 6550 1615
rect 6600 1600 6700 1615
rect 6750 1600 6850 1615
rect 6900 1600 7000 1615
rect 7050 1600 7150 1615
rect 7200 1600 7300 1615
rect 7350 1600 7450 1615
rect 7500 1600 7600 1615
rect 7650 1600 7750 1615
rect 7800 1600 7900 1615
rect 7950 1600 8050 1615
rect 8100 1600 8200 1615
rect 8250 1600 8350 1615
rect 8400 1600 8500 1615
rect 8550 1600 8650 1615
rect 8700 1600 8800 1615
rect 8850 1600 8950 1615
rect 9000 1600 9100 1615
rect 9150 1600 9250 1615
rect 9300 1600 9400 1615
rect 9450 1600 9550 1615
rect 9600 1600 9700 1615
rect 9750 1600 9850 1615
rect 9900 1600 10000 1615
rect 10050 1600 10150 1615
rect 10200 1600 10300 1615
rect 10350 1600 10450 1615
rect 10500 1600 10600 1615
rect 10650 1600 10750 1615
rect 10800 1600 10900 1615
rect 10950 1600 11050 1615
rect 11100 1600 11200 1615
rect 11250 1600 11350 1615
rect 11400 1600 11500 1615
rect 11550 1600 11650 1615
rect 11700 1600 11800 1615
rect 11850 1600 11950 1615
rect 12000 1600 12100 1615
rect 12150 1600 12250 1615
rect 12300 1600 12400 1615
rect 12450 1600 12550 1615
rect 12600 1600 12700 1615
rect 12750 1600 12850 1615
rect 12900 1600 13000 1615
rect 13050 1600 13150 1615
rect 13200 1600 13300 1615
rect 13350 1600 13450 1615
rect 13500 1600 13600 1615
rect 13650 1600 13750 1615
rect 13800 1600 13900 1615
rect 13950 1600 14050 1615
rect 14100 1600 14200 1615
rect 14250 1600 14350 1615
rect 14400 1600 14500 1615
rect 14550 1600 14650 1615
rect 14700 1600 14800 1615
rect 14850 1600 14950 1615
rect 15000 1600 15100 1615
rect 15150 1600 15250 1615
rect 15300 1600 15400 1615
rect 15450 1600 15550 1615
rect 15600 1600 15700 1615
rect 15750 1600 15850 1615
rect 15900 1600 16000 1615
rect 16050 1600 16150 1615
rect 16200 1600 16300 1615
rect 16350 1600 16450 1615
rect 16500 1600 16600 1615
rect 16650 1600 16750 1615
rect 16800 1600 16900 1615
rect 16950 1600 17050 1615
rect 17100 1600 17200 1615
rect 17250 1600 17350 1615
rect 17400 1600 17500 1615
rect 17550 1600 17650 1615
rect 17700 1600 17800 1615
rect 17850 1600 17950 1615
rect 18000 1600 18100 1615
rect 18150 1600 18250 1615
rect 18300 1600 18400 1615
rect 18450 1600 18550 1615
rect 18600 1600 18700 1615
rect 18750 1600 18850 1615
rect 18900 1600 19000 1615
rect 19050 1600 19150 1615
rect 19200 1600 19300 1615
rect 19350 1600 19450 1615
rect 19500 1600 19600 1615
rect 19650 1600 19750 1615
rect 19800 1600 19900 1615
rect 19950 1600 20050 1615
rect 20100 1600 20200 1615
rect 20250 1600 20350 1615
rect 20400 1600 20500 1615
rect 20550 1600 20650 1615
rect 20700 1600 20800 1615
rect 20850 1600 20950 1615
rect 21000 1600 21100 1615
rect 21150 1600 21250 1615
rect 21300 1600 21400 1615
rect 21450 1600 21550 1615
rect 21600 1600 21700 1615
rect 21750 1600 21850 1615
rect 21900 1600 22000 1615
rect 22050 1600 22150 1615
rect 22200 1600 22300 1615
rect 22350 1600 22450 1615
rect 22500 1600 22600 1615
rect 22650 1600 22750 1615
rect 22800 1600 22900 1615
rect 22950 1600 23050 1615
rect 23100 1600 23200 1615
rect 23250 1600 23350 1615
rect 23400 1600 23500 1615
rect 23550 1600 23650 1615
rect 23700 1600 23800 1615
rect 23850 1600 23950 1615
rect 24000 1600 24100 1615
rect 24150 1600 24250 1615
rect 24300 1600 24400 1615
rect 24450 1600 24550 1615
rect 24600 1600 24700 1615
rect 24750 1600 24850 1615
rect 24900 1600 25000 1615
rect 25050 1600 25150 1615
rect 25200 1600 25300 1615
rect 25350 1600 25450 1615
rect 25500 1600 25600 1615
rect 25650 1600 25750 1615
rect 25800 1600 25900 1615
rect 25950 1600 26050 1615
rect 26100 1600 26200 1615
rect 26250 1600 26350 1615
rect 26400 1600 26500 1615
rect 26550 1600 26650 1615
rect 26700 1600 26800 1615
rect 26850 1600 26950 1615
rect 27000 1600 27100 1615
rect 27150 1600 27250 1615
rect 27300 1600 27400 1615
rect 27450 1600 27550 1615
rect 27600 1600 27700 1615
rect 27750 1600 27850 1615
rect 27900 1600 28000 1615
rect 28050 1600 28150 1615
rect 28200 1600 28300 1615
rect 28350 1600 28450 1615
rect 28500 1600 28600 1615
rect 28650 1600 28750 1615
rect -600 850 -500 900
rect -450 850 -350 900
rect -600 835 -350 850
rect -600 815 -585 835
rect -565 815 -535 835
rect -515 815 -485 835
rect -465 815 -435 835
rect -415 815 -385 835
rect -365 815 -350 835
rect -600 800 -350 815
rect -600 750 -500 800
rect -450 750 -350 800
rect -300 850 -200 900
rect -150 850 -50 900
rect -300 835 -50 850
rect -300 815 -285 835
rect -265 815 -235 835
rect -215 815 -185 835
rect -165 815 -135 835
rect -115 815 -85 835
rect -65 815 -50 835
rect -300 800 -50 815
rect -300 750 -200 800
rect -150 750 -50 800
rect 0 850 100 900
rect 150 850 250 900
rect 0 835 250 850
rect 0 815 15 835
rect 35 815 65 835
rect 85 815 115 835
rect 135 815 165 835
rect 185 815 215 835
rect 235 815 250 835
rect 0 800 250 815
rect 0 750 100 800
rect 150 750 250 800
rect 300 850 400 900
rect 450 850 550 900
rect 300 835 550 850
rect 300 815 315 835
rect 335 815 365 835
rect 385 815 415 835
rect 435 815 465 835
rect 485 815 515 835
rect 535 815 550 835
rect 300 800 550 815
rect 300 750 400 800
rect 450 750 550 800
rect 600 850 700 900
rect 750 850 850 900
rect 600 835 850 850
rect 600 815 615 835
rect 635 815 665 835
rect 685 815 715 835
rect 735 815 765 835
rect 785 815 815 835
rect 835 815 850 835
rect 600 800 850 815
rect 600 750 700 800
rect 750 750 850 800
rect 900 850 1000 900
rect 1050 850 1150 900
rect 900 835 1150 850
rect 900 815 915 835
rect 935 815 965 835
rect 985 815 1015 835
rect 1035 815 1065 835
rect 1085 815 1115 835
rect 1135 815 1150 835
rect 900 800 1150 815
rect 900 750 1000 800
rect 1050 750 1150 800
rect 1200 850 1300 900
rect 1350 850 1450 900
rect 1200 835 1450 850
rect 1200 815 1215 835
rect 1235 815 1265 835
rect 1285 815 1315 835
rect 1335 815 1365 835
rect 1385 815 1415 835
rect 1435 815 1450 835
rect 1200 800 1450 815
rect 1200 750 1300 800
rect 1350 750 1450 800
rect 1500 850 1600 900
rect 1650 850 1750 900
rect 1500 835 1750 850
rect 1500 815 1515 835
rect 1535 815 1565 835
rect 1585 815 1615 835
rect 1635 815 1665 835
rect 1685 815 1715 835
rect 1735 815 1750 835
rect 1500 800 1750 815
rect 1500 750 1600 800
rect 1650 750 1750 800
rect 1800 850 1900 900
rect 1950 850 2050 900
rect 1800 835 2050 850
rect 1800 815 1815 835
rect 1835 815 1865 835
rect 1885 815 1915 835
rect 1935 815 1965 835
rect 1985 815 2015 835
rect 2035 815 2050 835
rect 1800 800 2050 815
rect 1800 750 1900 800
rect 1950 750 2050 800
rect 2100 850 2200 900
rect 2250 850 2350 900
rect 2100 835 2350 850
rect 2100 815 2115 835
rect 2135 815 2165 835
rect 2185 815 2215 835
rect 2235 815 2265 835
rect 2285 815 2315 835
rect 2335 815 2350 835
rect 2100 800 2350 815
rect 2100 750 2200 800
rect 2250 750 2350 800
rect 2400 850 2500 900
rect 2550 850 2650 900
rect 2400 835 2650 850
rect 2400 815 2415 835
rect 2435 815 2465 835
rect 2485 815 2515 835
rect 2535 815 2565 835
rect 2585 815 2615 835
rect 2635 815 2650 835
rect 2400 800 2650 815
rect 2400 750 2500 800
rect 2550 750 2650 800
rect 2700 850 2800 900
rect 2850 850 2950 900
rect 2700 835 2950 850
rect 2700 815 2715 835
rect 2735 815 2765 835
rect 2785 815 2815 835
rect 2835 815 2865 835
rect 2885 815 2915 835
rect 2935 815 2950 835
rect 2700 800 2950 815
rect 2700 750 2800 800
rect 2850 750 2950 800
rect 3000 850 3100 900
rect 3150 850 3250 900
rect 3000 835 3250 850
rect 3000 815 3015 835
rect 3035 815 3065 835
rect 3085 815 3115 835
rect 3135 815 3165 835
rect 3185 815 3215 835
rect 3235 815 3250 835
rect 3000 800 3250 815
rect 3000 750 3100 800
rect 3150 750 3250 800
rect 3300 850 3400 900
rect 3450 850 3550 900
rect 3300 835 3550 850
rect 3300 815 3315 835
rect 3335 815 3365 835
rect 3385 815 3415 835
rect 3435 815 3465 835
rect 3485 815 3515 835
rect 3535 815 3550 835
rect 3300 800 3550 815
rect 3300 750 3400 800
rect 3450 750 3550 800
rect 3600 850 3700 900
rect 3750 850 3850 900
rect 3600 835 3850 850
rect 3600 815 3615 835
rect 3635 815 3665 835
rect 3685 815 3715 835
rect 3735 815 3765 835
rect 3785 815 3815 835
rect 3835 815 3850 835
rect 3600 800 3850 815
rect 3600 750 3700 800
rect 3750 750 3850 800
rect 3900 850 4000 900
rect 4050 850 4150 900
rect 3900 835 4150 850
rect 3900 815 3915 835
rect 3935 815 3965 835
rect 3985 815 4015 835
rect 4035 815 4065 835
rect 4085 815 4115 835
rect 4135 815 4150 835
rect 3900 800 4150 815
rect 3900 750 4000 800
rect 4050 750 4150 800
rect 4200 850 4300 900
rect 4350 850 4450 900
rect 4200 835 4450 850
rect 4200 815 4215 835
rect 4235 815 4265 835
rect 4285 815 4315 835
rect 4335 815 4365 835
rect 4385 815 4415 835
rect 4435 815 4450 835
rect 4200 800 4450 815
rect 4200 750 4300 800
rect 4350 750 4450 800
rect 4500 850 4600 900
rect 4650 850 4750 900
rect 4500 835 4750 850
rect 4500 815 4515 835
rect 4535 815 4565 835
rect 4585 815 4615 835
rect 4635 815 4665 835
rect 4685 815 4715 835
rect 4735 815 4750 835
rect 4500 800 4750 815
rect 4500 750 4600 800
rect 4650 750 4750 800
rect 4800 850 4900 900
rect 4950 850 5050 900
rect 4800 835 5050 850
rect 4800 815 4815 835
rect 4835 815 4865 835
rect 4885 815 4915 835
rect 4935 815 4965 835
rect 4985 815 5015 835
rect 5035 815 5050 835
rect 4800 800 5050 815
rect 4800 750 4900 800
rect 4950 750 5050 800
rect 5100 850 5200 900
rect 5250 850 5350 900
rect 5100 835 5350 850
rect 5100 815 5115 835
rect 5135 815 5165 835
rect 5185 815 5215 835
rect 5235 815 5265 835
rect 5285 815 5315 835
rect 5335 815 5350 835
rect 5100 800 5350 815
rect 5100 750 5200 800
rect 5250 750 5350 800
rect 5400 850 5500 900
rect 5550 850 5650 900
rect 5400 835 5650 850
rect 5400 815 5415 835
rect 5435 815 5465 835
rect 5485 815 5515 835
rect 5535 815 5565 835
rect 5585 815 5615 835
rect 5635 815 5650 835
rect 5400 800 5650 815
rect 5400 750 5500 800
rect 5550 750 5650 800
rect 5700 850 5800 900
rect 5850 850 5950 900
rect 5700 835 5950 850
rect 5700 815 5715 835
rect 5735 815 5765 835
rect 5785 815 5815 835
rect 5835 815 5865 835
rect 5885 815 5915 835
rect 5935 815 5950 835
rect 5700 800 5950 815
rect 5700 750 5800 800
rect 5850 750 5950 800
rect 6000 850 6100 900
rect 6150 850 6250 900
rect 6000 835 6250 850
rect 6000 815 6015 835
rect 6035 815 6065 835
rect 6085 815 6115 835
rect 6135 815 6165 835
rect 6185 815 6215 835
rect 6235 815 6250 835
rect 6000 800 6250 815
rect 6000 750 6100 800
rect 6150 750 6250 800
rect 6300 850 6400 900
rect 6450 850 6550 900
rect 6300 835 6550 850
rect 6300 815 6315 835
rect 6335 815 6365 835
rect 6385 815 6415 835
rect 6435 815 6465 835
rect 6485 815 6515 835
rect 6535 815 6550 835
rect 6300 800 6550 815
rect 6300 750 6400 800
rect 6450 750 6550 800
rect 6600 850 6700 900
rect 6750 850 6850 900
rect 6600 835 6850 850
rect 6600 815 6615 835
rect 6635 815 6665 835
rect 6685 815 6715 835
rect 6735 815 6765 835
rect 6785 815 6815 835
rect 6835 815 6850 835
rect 6600 800 6850 815
rect 6600 750 6700 800
rect 6750 750 6850 800
rect 6900 850 7000 900
rect 7050 850 7150 900
rect 6900 835 7150 850
rect 6900 815 6915 835
rect 6935 815 6965 835
rect 6985 815 7015 835
rect 7035 815 7065 835
rect 7085 815 7115 835
rect 7135 815 7150 835
rect 6900 800 7150 815
rect 6900 750 7000 800
rect 7050 750 7150 800
rect 7200 850 7300 900
rect 7350 850 7450 900
rect 7200 835 7450 850
rect 7200 815 7215 835
rect 7235 815 7265 835
rect 7285 815 7315 835
rect 7335 815 7365 835
rect 7385 815 7415 835
rect 7435 815 7450 835
rect 7200 800 7450 815
rect 7200 750 7300 800
rect 7350 750 7450 800
rect 7500 850 7600 900
rect 7650 850 7750 900
rect 7500 835 7750 850
rect 7500 815 7515 835
rect 7535 815 7565 835
rect 7585 815 7615 835
rect 7635 815 7665 835
rect 7685 815 7715 835
rect 7735 815 7750 835
rect 7500 800 7750 815
rect 7500 750 7600 800
rect 7650 750 7750 800
rect 7800 850 7900 900
rect 7950 850 8050 900
rect 7800 835 8050 850
rect 7800 815 7815 835
rect 7835 815 7865 835
rect 7885 815 7915 835
rect 7935 815 7965 835
rect 7985 815 8015 835
rect 8035 815 8050 835
rect 7800 800 8050 815
rect 7800 750 7900 800
rect 7950 750 8050 800
rect 8100 850 8200 900
rect 8250 850 8350 900
rect 8100 835 8350 850
rect 8100 815 8115 835
rect 8135 815 8165 835
rect 8185 815 8215 835
rect 8235 815 8265 835
rect 8285 815 8315 835
rect 8335 815 8350 835
rect 8100 800 8350 815
rect 8100 750 8200 800
rect 8250 750 8350 800
rect 8400 850 8500 900
rect 8550 850 8650 900
rect 8400 835 8650 850
rect 8400 815 8415 835
rect 8435 815 8465 835
rect 8485 815 8515 835
rect 8535 815 8565 835
rect 8585 815 8615 835
rect 8635 815 8650 835
rect 8400 800 8650 815
rect 8400 750 8500 800
rect 8550 750 8650 800
rect 8700 850 8800 900
rect 8850 850 8950 900
rect 8700 835 8950 850
rect 8700 815 8715 835
rect 8735 815 8765 835
rect 8785 815 8815 835
rect 8835 815 8865 835
rect 8885 815 8915 835
rect 8935 815 8950 835
rect 8700 800 8950 815
rect 8700 750 8800 800
rect 8850 750 8950 800
rect 9000 850 9100 900
rect 9150 850 9250 900
rect 9000 835 9250 850
rect 9000 815 9015 835
rect 9035 815 9065 835
rect 9085 815 9115 835
rect 9135 815 9165 835
rect 9185 815 9215 835
rect 9235 815 9250 835
rect 9000 800 9250 815
rect 9000 750 9100 800
rect 9150 750 9250 800
rect 9300 850 9400 900
rect 9450 850 9550 900
rect 9300 835 9550 850
rect 9300 815 9315 835
rect 9335 815 9365 835
rect 9385 815 9415 835
rect 9435 815 9465 835
rect 9485 815 9515 835
rect 9535 815 9550 835
rect 9300 800 9550 815
rect 9300 750 9400 800
rect 9450 750 9550 800
rect 9600 850 9700 900
rect 9750 850 9850 900
rect 9600 835 9850 850
rect 9600 815 9615 835
rect 9635 815 9665 835
rect 9685 815 9715 835
rect 9735 815 9765 835
rect 9785 815 9815 835
rect 9835 815 9850 835
rect 9600 800 9850 815
rect 9600 750 9700 800
rect 9750 750 9850 800
rect 9900 850 10000 900
rect 10050 850 10150 900
rect 9900 835 10150 850
rect 9900 815 9915 835
rect 9935 815 9965 835
rect 9985 815 10015 835
rect 10035 815 10065 835
rect 10085 815 10115 835
rect 10135 815 10150 835
rect 9900 800 10150 815
rect 9900 750 10000 800
rect 10050 750 10150 800
rect 10200 850 10300 900
rect 10350 850 10450 900
rect 10200 835 10450 850
rect 10200 815 10215 835
rect 10235 815 10265 835
rect 10285 815 10315 835
rect 10335 815 10365 835
rect 10385 815 10415 835
rect 10435 815 10450 835
rect 10200 800 10450 815
rect 10200 750 10300 800
rect 10350 750 10450 800
rect 10500 850 10600 900
rect 10650 850 10750 900
rect 10500 835 10750 850
rect 10500 815 10515 835
rect 10535 815 10565 835
rect 10585 815 10615 835
rect 10635 815 10665 835
rect 10685 815 10715 835
rect 10735 815 10750 835
rect 10500 800 10750 815
rect 10500 750 10600 800
rect 10650 750 10750 800
rect 10800 850 10900 900
rect 10950 850 11050 900
rect 10800 835 11050 850
rect 10800 815 10815 835
rect 10835 815 10865 835
rect 10885 815 10915 835
rect 10935 815 10965 835
rect 10985 815 11015 835
rect 11035 815 11050 835
rect 10800 800 11050 815
rect 10800 750 10900 800
rect 10950 750 11050 800
rect 11100 850 11200 900
rect 11250 850 11350 900
rect 11100 835 11350 850
rect 11100 815 11115 835
rect 11135 815 11165 835
rect 11185 815 11215 835
rect 11235 815 11265 835
rect 11285 815 11315 835
rect 11335 815 11350 835
rect 11100 800 11350 815
rect 11100 750 11200 800
rect 11250 750 11350 800
rect 11400 850 11500 900
rect 11550 850 11650 900
rect 11400 835 11650 850
rect 11400 815 11415 835
rect 11435 815 11465 835
rect 11485 815 11515 835
rect 11535 815 11565 835
rect 11585 815 11615 835
rect 11635 815 11650 835
rect 11400 800 11650 815
rect 11400 750 11500 800
rect 11550 750 11650 800
rect 11700 850 11800 900
rect 11850 850 11950 900
rect 11700 835 11950 850
rect 11700 815 11715 835
rect 11735 815 11765 835
rect 11785 815 11815 835
rect 11835 815 11865 835
rect 11885 815 11915 835
rect 11935 815 11950 835
rect 11700 800 11950 815
rect 11700 750 11800 800
rect 11850 750 11950 800
rect 12000 850 12100 900
rect 12150 850 12250 900
rect 12000 835 12250 850
rect 12000 815 12015 835
rect 12035 815 12065 835
rect 12085 815 12115 835
rect 12135 815 12165 835
rect 12185 815 12215 835
rect 12235 815 12250 835
rect 12000 800 12250 815
rect 12000 750 12100 800
rect 12150 750 12250 800
rect 12300 850 12400 900
rect 12450 850 12550 900
rect 12300 835 12550 850
rect 12300 815 12315 835
rect 12335 815 12365 835
rect 12385 815 12415 835
rect 12435 815 12465 835
rect 12485 815 12515 835
rect 12535 815 12550 835
rect 12300 800 12550 815
rect 12300 750 12400 800
rect 12450 750 12550 800
rect 12600 850 12700 900
rect 12750 850 12850 900
rect 12600 835 12850 850
rect 12600 815 12615 835
rect 12635 815 12665 835
rect 12685 815 12715 835
rect 12735 815 12765 835
rect 12785 815 12815 835
rect 12835 815 12850 835
rect 12600 800 12850 815
rect 12600 750 12700 800
rect 12750 750 12850 800
rect 12900 850 13000 900
rect 13050 850 13150 900
rect 12900 835 13150 850
rect 12900 815 12915 835
rect 12935 815 12965 835
rect 12985 815 13015 835
rect 13035 815 13065 835
rect 13085 815 13115 835
rect 13135 815 13150 835
rect 12900 800 13150 815
rect 12900 750 13000 800
rect 13050 750 13150 800
rect 13200 850 13300 900
rect 13350 850 13450 900
rect 13200 835 13450 850
rect 13200 815 13215 835
rect 13235 815 13265 835
rect 13285 815 13315 835
rect 13335 815 13365 835
rect 13385 815 13415 835
rect 13435 815 13450 835
rect 13200 800 13450 815
rect 13200 750 13300 800
rect 13350 750 13450 800
rect 13500 850 13600 900
rect 13650 850 13750 900
rect 13500 835 13750 850
rect 13500 815 13515 835
rect 13535 815 13565 835
rect 13585 815 13615 835
rect 13635 815 13665 835
rect 13685 815 13715 835
rect 13735 815 13750 835
rect 13500 800 13750 815
rect 13500 750 13600 800
rect 13650 750 13750 800
rect 13800 850 13900 900
rect 13950 850 14050 900
rect 13800 835 14050 850
rect 13800 815 13815 835
rect 13835 815 13865 835
rect 13885 815 13915 835
rect 13935 815 13965 835
rect 13985 815 14015 835
rect 14035 815 14050 835
rect 13800 800 14050 815
rect 13800 750 13900 800
rect 13950 750 14050 800
rect 14100 850 14200 900
rect 14250 850 14350 900
rect 14100 835 14350 850
rect 14100 815 14115 835
rect 14135 815 14165 835
rect 14185 815 14215 835
rect 14235 815 14265 835
rect 14285 815 14315 835
rect 14335 815 14350 835
rect 14100 800 14350 815
rect 14100 750 14200 800
rect 14250 750 14350 800
rect 14400 850 14500 900
rect 14550 850 14650 900
rect 14400 835 14650 850
rect 14400 815 14415 835
rect 14435 815 14465 835
rect 14485 815 14515 835
rect 14535 815 14565 835
rect 14585 815 14615 835
rect 14635 815 14650 835
rect 14400 800 14650 815
rect 14400 750 14500 800
rect 14550 750 14650 800
rect 14700 850 14800 900
rect 14850 850 14950 900
rect 14700 835 14950 850
rect 14700 815 14715 835
rect 14735 815 14765 835
rect 14785 815 14815 835
rect 14835 815 14865 835
rect 14885 815 14915 835
rect 14935 815 14950 835
rect 14700 800 14950 815
rect 14700 750 14800 800
rect 14850 750 14950 800
rect 15000 850 15100 900
rect 15150 850 15250 900
rect 15000 835 15250 850
rect 15000 815 15015 835
rect 15035 815 15065 835
rect 15085 815 15115 835
rect 15135 815 15165 835
rect 15185 815 15215 835
rect 15235 815 15250 835
rect 15000 800 15250 815
rect 15000 750 15100 800
rect 15150 750 15250 800
rect 15300 850 15400 900
rect 15450 850 15550 900
rect 15300 835 15550 850
rect 15300 815 15315 835
rect 15335 815 15365 835
rect 15385 815 15415 835
rect 15435 815 15465 835
rect 15485 815 15515 835
rect 15535 815 15550 835
rect 15300 800 15550 815
rect 15300 750 15400 800
rect 15450 750 15550 800
rect 15600 850 15700 900
rect 15750 850 15850 900
rect 15600 835 15850 850
rect 15600 815 15615 835
rect 15635 815 15665 835
rect 15685 815 15715 835
rect 15735 815 15765 835
rect 15785 815 15815 835
rect 15835 815 15850 835
rect 15600 800 15850 815
rect 15600 750 15700 800
rect 15750 750 15850 800
rect 15900 850 16000 900
rect 16050 850 16150 900
rect 15900 835 16150 850
rect 15900 815 15915 835
rect 15935 815 15965 835
rect 15985 815 16015 835
rect 16035 815 16065 835
rect 16085 815 16115 835
rect 16135 815 16150 835
rect 15900 800 16150 815
rect 15900 750 16000 800
rect 16050 750 16150 800
rect 16200 850 16300 900
rect 16350 850 16450 900
rect 16200 835 16450 850
rect 16200 815 16215 835
rect 16235 815 16265 835
rect 16285 815 16315 835
rect 16335 815 16365 835
rect 16385 815 16415 835
rect 16435 815 16450 835
rect 16200 800 16450 815
rect 16200 750 16300 800
rect 16350 750 16450 800
rect 16500 850 16600 900
rect 16650 850 16750 900
rect 16500 835 16750 850
rect 16500 815 16515 835
rect 16535 815 16565 835
rect 16585 815 16615 835
rect 16635 815 16665 835
rect 16685 815 16715 835
rect 16735 815 16750 835
rect 16500 800 16750 815
rect 16500 750 16600 800
rect 16650 750 16750 800
rect 16800 850 16900 900
rect 16950 850 17050 900
rect 16800 835 17050 850
rect 16800 815 16815 835
rect 16835 815 16865 835
rect 16885 815 16915 835
rect 16935 815 16965 835
rect 16985 815 17015 835
rect 17035 815 17050 835
rect 16800 800 17050 815
rect 16800 750 16900 800
rect 16950 750 17050 800
rect 17100 850 17200 900
rect 17250 850 17350 900
rect 17100 835 17350 850
rect 17100 815 17115 835
rect 17135 815 17165 835
rect 17185 815 17215 835
rect 17235 815 17265 835
rect 17285 815 17315 835
rect 17335 815 17350 835
rect 17100 800 17350 815
rect 17100 750 17200 800
rect 17250 750 17350 800
rect 17400 850 17500 900
rect 17550 850 17650 900
rect 17400 835 17650 850
rect 17400 815 17415 835
rect 17435 815 17465 835
rect 17485 815 17515 835
rect 17535 815 17565 835
rect 17585 815 17615 835
rect 17635 815 17650 835
rect 17400 800 17650 815
rect 17400 750 17500 800
rect 17550 750 17650 800
rect 17700 850 17800 900
rect 17850 850 17950 900
rect 17700 835 17950 850
rect 17700 815 17715 835
rect 17735 815 17765 835
rect 17785 815 17815 835
rect 17835 815 17865 835
rect 17885 815 17915 835
rect 17935 815 17950 835
rect 17700 800 17950 815
rect 17700 750 17800 800
rect 17850 750 17950 800
rect 18000 850 18100 900
rect 18150 850 18250 900
rect 18000 835 18250 850
rect 18000 815 18015 835
rect 18035 815 18065 835
rect 18085 815 18115 835
rect 18135 815 18165 835
rect 18185 815 18215 835
rect 18235 815 18250 835
rect 18000 800 18250 815
rect 18000 750 18100 800
rect 18150 750 18250 800
rect 18300 850 18400 900
rect 18450 850 18550 900
rect 18300 835 18550 850
rect 18300 815 18315 835
rect 18335 815 18365 835
rect 18385 815 18415 835
rect 18435 815 18465 835
rect 18485 815 18515 835
rect 18535 815 18550 835
rect 18300 800 18550 815
rect 18300 750 18400 800
rect 18450 750 18550 800
rect 18600 850 18700 900
rect 18750 850 18850 900
rect 18600 835 18850 850
rect 18600 815 18615 835
rect 18635 815 18665 835
rect 18685 815 18715 835
rect 18735 815 18765 835
rect 18785 815 18815 835
rect 18835 815 18850 835
rect 18600 800 18850 815
rect 18600 750 18700 800
rect 18750 750 18850 800
rect 18900 850 19000 900
rect 19050 850 19150 900
rect 18900 835 19150 850
rect 18900 815 18915 835
rect 18935 815 18965 835
rect 18985 815 19015 835
rect 19035 815 19065 835
rect 19085 815 19115 835
rect 19135 815 19150 835
rect 18900 800 19150 815
rect 18900 750 19000 800
rect 19050 750 19150 800
rect 19200 850 19300 900
rect 19350 850 19450 900
rect 19200 835 19450 850
rect 19200 815 19215 835
rect 19235 815 19265 835
rect 19285 815 19315 835
rect 19335 815 19365 835
rect 19385 815 19415 835
rect 19435 815 19450 835
rect 19200 800 19450 815
rect 19200 750 19300 800
rect 19350 750 19450 800
rect 19500 850 19600 900
rect 19650 850 19750 900
rect 19500 835 19750 850
rect 19500 815 19515 835
rect 19535 815 19565 835
rect 19585 815 19615 835
rect 19635 815 19665 835
rect 19685 815 19715 835
rect 19735 815 19750 835
rect 19500 800 19750 815
rect 19500 750 19600 800
rect 19650 750 19750 800
rect 19800 850 19900 900
rect 19950 850 20050 900
rect 19800 835 20050 850
rect 19800 815 19815 835
rect 19835 815 19865 835
rect 19885 815 19915 835
rect 19935 815 19965 835
rect 19985 815 20015 835
rect 20035 815 20050 835
rect 19800 800 20050 815
rect 19800 750 19900 800
rect 19950 750 20050 800
rect 20100 850 20200 900
rect 20250 850 20350 900
rect 20100 835 20350 850
rect 20100 815 20115 835
rect 20135 815 20165 835
rect 20185 815 20215 835
rect 20235 815 20265 835
rect 20285 815 20315 835
rect 20335 815 20350 835
rect 20100 800 20350 815
rect 20100 750 20200 800
rect 20250 750 20350 800
rect 20400 850 20500 900
rect 20550 850 20650 900
rect 20400 835 20650 850
rect 20400 815 20415 835
rect 20435 815 20465 835
rect 20485 815 20515 835
rect 20535 815 20565 835
rect 20585 815 20615 835
rect 20635 815 20650 835
rect 20400 800 20650 815
rect 20400 750 20500 800
rect 20550 750 20650 800
rect 20700 850 20800 900
rect 20850 850 20950 900
rect 20700 835 20950 850
rect 20700 815 20715 835
rect 20735 815 20765 835
rect 20785 815 20815 835
rect 20835 815 20865 835
rect 20885 815 20915 835
rect 20935 815 20950 835
rect 20700 800 20950 815
rect 20700 750 20800 800
rect 20850 750 20950 800
rect 21000 850 21100 900
rect 21150 850 21250 900
rect 21000 835 21250 850
rect 21000 815 21015 835
rect 21035 815 21065 835
rect 21085 815 21115 835
rect 21135 815 21165 835
rect 21185 815 21215 835
rect 21235 815 21250 835
rect 21000 800 21250 815
rect 21000 750 21100 800
rect 21150 750 21250 800
rect 21300 850 21400 900
rect 21450 850 21550 900
rect 21300 835 21550 850
rect 21300 815 21315 835
rect 21335 815 21365 835
rect 21385 815 21415 835
rect 21435 815 21465 835
rect 21485 815 21515 835
rect 21535 815 21550 835
rect 21300 800 21550 815
rect 21300 750 21400 800
rect 21450 750 21550 800
rect 21600 850 21700 900
rect 21750 850 21850 900
rect 21600 835 21850 850
rect 21600 815 21615 835
rect 21635 815 21665 835
rect 21685 815 21715 835
rect 21735 815 21765 835
rect 21785 815 21815 835
rect 21835 815 21850 835
rect 21600 800 21850 815
rect 21600 750 21700 800
rect 21750 750 21850 800
rect 21900 850 22000 900
rect 22050 850 22150 900
rect 21900 835 22150 850
rect 21900 815 21915 835
rect 21935 815 21965 835
rect 21985 815 22015 835
rect 22035 815 22065 835
rect 22085 815 22115 835
rect 22135 815 22150 835
rect 21900 800 22150 815
rect 21900 750 22000 800
rect 22050 750 22150 800
rect 22200 850 22300 900
rect 22350 850 22450 900
rect 22200 835 22450 850
rect 22200 815 22215 835
rect 22235 815 22265 835
rect 22285 815 22315 835
rect 22335 815 22365 835
rect 22385 815 22415 835
rect 22435 815 22450 835
rect 22200 800 22450 815
rect 22200 750 22300 800
rect 22350 750 22450 800
rect 22500 850 22600 900
rect 22650 850 22750 900
rect 22500 835 22750 850
rect 22500 815 22515 835
rect 22535 815 22565 835
rect 22585 815 22615 835
rect 22635 815 22665 835
rect 22685 815 22715 835
rect 22735 815 22750 835
rect 22500 800 22750 815
rect 22500 750 22600 800
rect 22650 750 22750 800
rect 22800 850 22900 900
rect 22950 850 23050 900
rect 22800 835 23050 850
rect 22800 815 22815 835
rect 22835 815 22865 835
rect 22885 815 22915 835
rect 22935 815 22965 835
rect 22985 815 23015 835
rect 23035 815 23050 835
rect 22800 800 23050 815
rect 22800 750 22900 800
rect 22950 750 23050 800
rect 23100 850 23200 900
rect 23250 850 23350 900
rect 23100 835 23350 850
rect 23100 815 23115 835
rect 23135 815 23165 835
rect 23185 815 23215 835
rect 23235 815 23265 835
rect 23285 815 23315 835
rect 23335 815 23350 835
rect 23100 800 23350 815
rect 23100 750 23200 800
rect 23250 750 23350 800
rect 23400 850 23500 900
rect 23550 850 23650 900
rect 23400 835 23650 850
rect 23400 815 23415 835
rect 23435 815 23465 835
rect 23485 815 23515 835
rect 23535 815 23565 835
rect 23585 815 23615 835
rect 23635 815 23650 835
rect 23400 800 23650 815
rect 23400 750 23500 800
rect 23550 750 23650 800
rect 23700 850 23800 900
rect 23850 850 23950 900
rect 23700 835 23950 850
rect 23700 815 23715 835
rect 23735 815 23765 835
rect 23785 815 23815 835
rect 23835 815 23865 835
rect 23885 815 23915 835
rect 23935 815 23950 835
rect 23700 800 23950 815
rect 23700 750 23800 800
rect 23850 750 23950 800
rect 24000 850 24100 900
rect 24150 850 24250 900
rect 24000 835 24250 850
rect 24000 815 24015 835
rect 24035 815 24065 835
rect 24085 815 24115 835
rect 24135 815 24165 835
rect 24185 815 24215 835
rect 24235 815 24250 835
rect 24000 800 24250 815
rect 24000 750 24100 800
rect 24150 750 24250 800
rect 24300 850 24400 900
rect 24450 850 24550 900
rect 24300 835 24550 850
rect 24300 815 24315 835
rect 24335 815 24365 835
rect 24385 815 24415 835
rect 24435 815 24465 835
rect 24485 815 24515 835
rect 24535 815 24550 835
rect 24300 800 24550 815
rect 24300 750 24400 800
rect 24450 750 24550 800
rect 24600 850 24700 900
rect 24750 850 24850 900
rect 24600 835 24850 850
rect 24600 815 24615 835
rect 24635 815 24665 835
rect 24685 815 24715 835
rect 24735 815 24765 835
rect 24785 815 24815 835
rect 24835 815 24850 835
rect 24600 800 24850 815
rect 24600 750 24700 800
rect 24750 750 24850 800
rect 24900 850 25000 900
rect 25050 850 25150 900
rect 24900 835 25150 850
rect 24900 815 24915 835
rect 24935 815 24965 835
rect 24985 815 25015 835
rect 25035 815 25065 835
rect 25085 815 25115 835
rect 25135 815 25150 835
rect 24900 800 25150 815
rect 24900 750 25000 800
rect 25050 750 25150 800
rect 25200 850 25300 900
rect 25350 850 25450 900
rect 25200 835 25450 850
rect 25200 815 25215 835
rect 25235 815 25265 835
rect 25285 815 25315 835
rect 25335 815 25365 835
rect 25385 815 25415 835
rect 25435 815 25450 835
rect 25200 800 25450 815
rect 25200 750 25300 800
rect 25350 750 25450 800
rect 25500 850 25600 900
rect 25650 850 25750 900
rect 25500 835 25750 850
rect 25500 815 25515 835
rect 25535 815 25565 835
rect 25585 815 25615 835
rect 25635 815 25665 835
rect 25685 815 25715 835
rect 25735 815 25750 835
rect 25500 800 25750 815
rect 25500 750 25600 800
rect 25650 750 25750 800
rect 25800 850 25900 900
rect 25950 850 26050 900
rect 25800 835 26050 850
rect 25800 815 25815 835
rect 25835 815 25865 835
rect 25885 815 25915 835
rect 25935 815 25965 835
rect 25985 815 26015 835
rect 26035 815 26050 835
rect 25800 800 26050 815
rect 25800 750 25900 800
rect 25950 750 26050 800
rect 26100 850 26200 900
rect 26250 850 26350 900
rect 26100 835 26350 850
rect 26100 815 26115 835
rect 26135 815 26165 835
rect 26185 815 26215 835
rect 26235 815 26265 835
rect 26285 815 26315 835
rect 26335 815 26350 835
rect 26100 800 26350 815
rect 26100 750 26200 800
rect 26250 750 26350 800
rect 26400 850 26500 900
rect 26550 850 26650 900
rect 26400 835 26650 850
rect 26400 815 26415 835
rect 26435 815 26465 835
rect 26485 815 26515 835
rect 26535 815 26565 835
rect 26585 815 26615 835
rect 26635 815 26650 835
rect 26400 800 26650 815
rect 26400 750 26500 800
rect 26550 750 26650 800
rect 26700 850 26800 900
rect 26850 850 26950 900
rect 26700 835 26950 850
rect 26700 815 26715 835
rect 26735 815 26765 835
rect 26785 815 26815 835
rect 26835 815 26865 835
rect 26885 815 26915 835
rect 26935 815 26950 835
rect 26700 800 26950 815
rect 26700 750 26800 800
rect 26850 750 26950 800
rect 27000 850 27100 900
rect 27150 850 27250 900
rect 27000 835 27250 850
rect 27000 815 27015 835
rect 27035 815 27065 835
rect 27085 815 27115 835
rect 27135 815 27165 835
rect 27185 815 27215 835
rect 27235 815 27250 835
rect 27000 800 27250 815
rect 27000 750 27100 800
rect 27150 750 27250 800
rect 27300 850 27400 900
rect 27450 850 27550 900
rect 27300 835 27550 850
rect 27300 815 27315 835
rect 27335 815 27365 835
rect 27385 815 27415 835
rect 27435 815 27465 835
rect 27485 815 27515 835
rect 27535 815 27550 835
rect 27300 800 27550 815
rect 27300 750 27400 800
rect 27450 750 27550 800
rect 27600 850 27700 900
rect 27750 850 27850 900
rect 27600 835 27850 850
rect 27600 815 27615 835
rect 27635 815 27665 835
rect 27685 815 27715 835
rect 27735 815 27765 835
rect 27785 815 27815 835
rect 27835 815 27850 835
rect 27600 800 27850 815
rect 27600 750 27700 800
rect 27750 750 27850 800
rect 27900 850 28000 900
rect 28050 850 28150 900
rect 27900 835 28150 850
rect 27900 815 27915 835
rect 27935 815 27965 835
rect 27985 815 28015 835
rect 28035 815 28065 835
rect 28085 815 28115 835
rect 28135 815 28150 835
rect 27900 800 28150 815
rect 27900 750 28000 800
rect 28050 750 28150 800
rect 28200 850 28300 900
rect 28350 850 28450 900
rect 28200 835 28450 850
rect 28200 815 28215 835
rect 28235 815 28265 835
rect 28285 815 28315 835
rect 28335 815 28365 835
rect 28385 815 28415 835
rect 28435 815 28450 835
rect 28200 800 28450 815
rect 28200 750 28300 800
rect 28350 750 28450 800
rect 28500 850 28600 900
rect 28650 850 28750 900
rect 28500 835 28750 850
rect 28500 815 28515 835
rect 28535 815 28565 835
rect 28585 815 28615 835
rect 28635 815 28665 835
rect 28685 815 28715 835
rect 28735 815 28750 835
rect 28500 800 28750 815
rect 28500 750 28600 800
rect 28650 750 28750 800
rect -600 35 -500 50
rect -450 35 -350 50
rect -300 35 -200 50
rect -150 35 -50 50
rect 0 35 100 50
rect 150 35 250 50
rect 300 35 400 50
rect 450 35 550 50
rect 600 35 700 50
rect 750 35 850 50
rect 900 35 1000 50
rect 1050 35 1150 50
rect 1200 35 1300 50
rect 1350 35 1450 50
rect 1500 35 1600 50
rect 1650 35 1750 50
rect 1800 35 1900 50
rect 1950 35 2050 50
rect 2100 35 2200 50
rect 2250 35 2350 50
rect 2400 35 2500 50
rect 2550 35 2650 50
rect 2700 35 2800 50
rect 2850 35 2950 50
rect 3000 35 3100 50
rect 3150 35 3250 50
rect 3300 35 3400 50
rect 3450 35 3550 50
rect 3600 35 3700 50
rect 3750 35 3850 50
rect 3900 35 4000 50
rect 4050 35 4150 50
rect 4200 35 4300 50
rect 4350 35 4450 50
rect 4500 35 4600 50
rect 4650 35 4750 50
rect 4800 35 4900 50
rect 4950 35 5050 50
rect 5100 35 5200 50
rect 5250 35 5350 50
rect 5400 35 5500 50
rect 5550 35 5650 50
rect 5700 35 5800 50
rect 5850 35 5950 50
rect 6000 35 6100 50
rect 6150 35 6250 50
rect 6300 35 6400 50
rect 6450 35 6550 50
rect 6600 35 6700 50
rect 6750 35 6850 50
rect 6900 35 7000 50
rect 7050 35 7150 50
rect 7200 35 7300 50
rect 7350 35 7450 50
rect 7500 35 7600 50
rect 7650 35 7750 50
rect 7800 35 7900 50
rect 7950 35 8050 50
rect 8100 35 8200 50
rect 8250 35 8350 50
rect 8400 35 8500 50
rect 8550 35 8650 50
rect 8700 35 8800 50
rect 8850 35 8950 50
rect 9000 35 9100 50
rect 9150 35 9250 50
rect 9300 35 9400 50
rect 9450 35 9550 50
rect 9600 35 9700 50
rect 9750 35 9850 50
rect 9900 35 10000 50
rect 10050 35 10150 50
rect 10200 35 10300 50
rect 10350 35 10450 50
rect 10500 35 10600 50
rect 10650 35 10750 50
rect 10800 35 10900 50
rect 10950 35 11050 50
rect 11100 35 11200 50
rect 11250 35 11350 50
rect 11400 35 11500 50
rect 11550 35 11650 50
rect 11700 35 11800 50
rect 11850 35 11950 50
rect 12000 35 12100 50
rect 12150 35 12250 50
rect 12300 35 12400 50
rect 12450 35 12550 50
rect 12600 35 12700 50
rect 12750 35 12850 50
rect 12900 35 13000 50
rect 13050 35 13150 50
rect 13200 35 13300 50
rect 13350 35 13450 50
rect 13500 35 13600 50
rect 13650 35 13750 50
rect 13800 35 13900 50
rect 13950 35 14050 50
rect 14100 35 14200 50
rect 14250 35 14350 50
rect 14400 35 14500 50
rect 14550 35 14650 50
rect 14700 35 14800 50
rect 14850 35 14950 50
rect 15000 35 15100 50
rect 15150 35 15250 50
rect 15300 35 15400 50
rect 15450 35 15550 50
rect 15600 35 15700 50
rect 15750 35 15850 50
rect 15900 35 16000 50
rect 16050 35 16150 50
rect 16200 35 16300 50
rect 16350 35 16450 50
rect 16500 35 16600 50
rect 16650 35 16750 50
rect 16800 35 16900 50
rect 16950 35 17050 50
rect 17100 35 17200 50
rect 17250 35 17350 50
rect 17400 35 17500 50
rect 17550 35 17650 50
rect 17700 35 17800 50
rect 17850 35 17950 50
rect 18000 35 18100 50
rect 18150 35 18250 50
rect 18300 35 18400 50
rect 18450 35 18550 50
rect 18600 35 18700 50
rect 18750 35 18850 50
rect 18900 35 19000 50
rect 19050 35 19150 50
rect 19200 35 19300 50
rect 19350 35 19450 50
rect 19500 35 19600 50
rect 19650 35 19750 50
rect 19800 35 19900 50
rect 19950 35 20050 50
rect 20100 35 20200 50
rect 20250 35 20350 50
rect 20400 35 20500 50
rect 20550 35 20650 50
rect 20700 35 20800 50
rect 20850 35 20950 50
rect 21000 35 21100 50
rect 21150 35 21250 50
rect 21300 35 21400 50
rect 21450 35 21550 50
rect 21600 35 21700 50
rect 21750 35 21850 50
rect 21900 35 22000 50
rect 22050 35 22150 50
rect 22200 35 22300 50
rect 22350 35 22450 50
rect 22500 35 22600 50
rect 22650 35 22750 50
rect 22800 35 22900 50
rect 22950 35 23050 50
rect 23100 35 23200 50
rect 23250 35 23350 50
rect 23400 35 23500 50
rect 23550 35 23650 50
rect 23700 35 23800 50
rect 23850 35 23950 50
rect 24000 35 24100 50
rect 24150 35 24250 50
rect 24300 35 24400 50
rect 24450 35 24550 50
rect 24600 35 24700 50
rect 24750 35 24850 50
rect 24900 35 25000 50
rect 25050 35 25150 50
rect 25200 35 25300 50
rect 25350 35 25450 50
rect 25500 35 25600 50
rect 25650 35 25750 50
rect 25800 35 25900 50
rect 25950 35 26050 50
rect 26100 35 26200 50
rect 26250 35 26350 50
rect 26400 35 26500 50
rect 26550 35 26650 50
rect 26700 35 26800 50
rect 26850 35 26950 50
rect 27000 35 27100 50
rect 27150 35 27250 50
rect 27300 35 27400 50
rect 27450 35 27550 50
rect 27600 35 27700 50
rect 27750 35 27850 50
rect 27900 35 28000 50
rect 28050 35 28150 50
rect 28200 35 28300 50
rect 28350 35 28450 50
rect 28500 35 28600 50
rect 28650 35 28750 50
rect -600 -100 -500 -85
rect -450 -100 -350 -85
rect -300 -100 -200 -85
rect -150 -100 -50 -85
rect 0 -100 100 -85
rect 150 -100 250 -85
rect 300 -100 400 -85
rect 450 -100 550 -85
rect 600 -100 700 -85
rect 750 -100 850 -85
rect 900 -100 1000 -85
rect 1050 -100 1150 -85
rect 1200 -100 1300 -85
rect 1350 -100 1450 -85
rect 1500 -100 1600 -85
rect 1650 -100 1750 -85
rect 1800 -100 1900 -85
rect 1950 -100 2050 -85
rect 2100 -100 2200 -85
rect 2250 -100 2350 -85
rect 2400 -100 2500 -85
rect 2550 -100 2650 -85
rect 2700 -100 2800 -85
rect 2850 -100 2950 -85
rect 3000 -100 3100 -85
rect 3150 -100 3250 -85
rect 3300 -100 3400 -85
rect 3450 -100 3550 -85
rect 3600 -100 3700 -85
rect 3750 -100 3850 -85
rect 3900 -100 4000 -85
rect 4050 -100 4150 -85
rect 4200 -100 4300 -85
rect 4350 -100 4450 -85
rect 4500 -100 4600 -85
rect 4650 -100 4750 -85
rect 4800 -100 4900 -85
rect 4950 -100 5050 -85
rect 5100 -100 5200 -85
rect 5250 -100 5350 -85
rect 5400 -100 5500 -85
rect 5550 -100 5650 -85
rect 5700 -100 5800 -85
rect 5850 -100 5950 -85
rect 6000 -100 6100 -85
rect 6150 -100 6250 -85
rect 6300 -100 6400 -85
rect 6450 -100 6550 -85
rect 6600 -100 6700 -85
rect 6750 -100 6850 -85
rect 6900 -100 7000 -85
rect 7050 -100 7150 -85
rect 7200 -100 7300 -85
rect 7350 -100 7450 -85
rect 7500 -100 7600 -85
rect 7650 -100 7750 -85
rect 7800 -100 7900 -85
rect 7950 -100 8050 -85
rect 8100 -100 8200 -85
rect 8250 -100 8350 -85
rect 8400 -100 8500 -85
rect 8550 -100 8650 -85
rect 8700 -100 8800 -85
rect 8850 -100 8950 -85
rect 9000 -100 9100 -85
rect 9150 -100 9250 -85
rect 9300 -100 9400 -85
rect 9450 -100 9550 -85
rect 9600 -100 9700 -85
rect 9750 -100 9850 -85
rect 9900 -100 10000 -85
rect 10050 -100 10150 -85
rect 10200 -100 10300 -85
rect 10350 -100 10450 -85
rect 10500 -100 10600 -85
rect 10650 -100 10750 -85
rect 10800 -100 10900 -85
rect 10950 -100 11050 -85
rect 11100 -100 11200 -85
rect 11250 -100 11350 -85
rect 11400 -100 11500 -85
rect 11550 -100 11650 -85
rect 11700 -100 11800 -85
rect 11850 -100 11950 -85
rect 12000 -100 12100 -85
rect 12150 -100 12250 -85
rect 12300 -100 12400 -85
rect 12450 -100 12550 -85
rect 12600 -100 12700 -85
rect 12750 -100 12850 -85
rect 12900 -100 13000 -85
rect 13050 -100 13150 -85
rect 13200 -100 13300 -85
rect 13350 -100 13450 -85
rect 13500 -100 13600 -85
rect 13650 -100 13750 -85
rect 13800 -100 13900 -85
rect 13950 -100 14050 -85
rect 14100 -100 14200 -85
rect 14250 -100 14350 -85
rect 14400 -100 14500 -85
rect 14550 -100 14650 -85
rect 14700 -100 14800 -85
rect 14850 -100 14950 -85
rect 15000 -100 15100 -85
rect 15150 -100 15250 -85
rect 15300 -100 15400 -85
rect 15450 -100 15550 -85
rect 15600 -100 15700 -85
rect 15750 -100 15850 -85
rect 15900 -100 16000 -85
rect 16050 -100 16150 -85
rect 16200 -100 16300 -85
rect 16350 -100 16450 -85
rect 16500 -100 16600 -85
rect 16650 -100 16750 -85
rect 16800 -100 16900 -85
rect 16950 -100 17050 -85
rect 17100 -100 17200 -85
rect 17250 -100 17350 -85
rect 17400 -100 17500 -85
rect 17550 -100 17650 -85
rect 17700 -100 17800 -85
rect 17850 -100 17950 -85
rect 18000 -100 18100 -85
rect 18150 -100 18250 -85
rect 18300 -100 18400 -85
rect 18450 -100 18550 -85
rect 18600 -100 18700 -85
rect 18750 -100 18850 -85
rect 18900 -100 19000 -85
rect 19050 -100 19150 -85
rect 19200 -100 19300 -85
rect 19350 -100 19450 -85
rect 19500 -100 19600 -85
rect 19650 -100 19750 -85
rect 19800 -100 19900 -85
rect 19950 -100 20050 -85
rect 20100 -100 20200 -85
rect 20250 -100 20350 -85
rect 20400 -100 20500 -85
rect 20550 -100 20650 -85
rect 20700 -100 20800 -85
rect 20850 -100 20950 -85
rect 21000 -100 21100 -85
rect 21150 -100 21250 -85
rect 21300 -100 21400 -85
rect 21450 -100 21550 -85
rect 21600 -100 21700 -85
rect 21750 -100 21850 -85
rect 21900 -100 22000 -85
rect 22050 -100 22150 -85
rect 22200 -100 22300 -85
rect 22350 -100 22450 -85
rect 22500 -100 22600 -85
rect 22650 -100 22750 -85
rect 22800 -100 22900 -85
rect 22950 -100 23050 -85
rect 23100 -100 23200 -85
rect 23250 -100 23350 -85
rect 23400 -100 23500 -85
rect 23550 -100 23650 -85
rect 23700 -100 23800 -85
rect 23850 -100 23950 -85
rect 24000 -100 24100 -85
rect 24150 -100 24250 -85
rect 24300 -100 24400 -85
rect 24450 -100 24550 -85
rect 24600 -100 24700 -85
rect 24750 -100 24850 -85
rect 24900 -100 25000 -85
rect 25050 -100 25150 -85
rect 25200 -100 25300 -85
rect 25350 -100 25450 -85
rect 25500 -100 25600 -85
rect 25650 -100 25750 -85
rect 25800 -100 25900 -85
rect 25950 -100 26050 -85
rect 26100 -100 26200 -85
rect 26250 -100 26350 -85
rect 26400 -100 26500 -85
rect 26550 -100 26650 -85
rect 26700 -100 26800 -85
rect 26850 -100 26950 -85
rect 27000 -100 27100 -85
rect 27150 -100 27250 -85
rect 27300 -100 27400 -85
rect 27450 -100 27550 -85
rect 27600 -100 27700 -85
rect 27750 -100 27850 -85
rect 27900 -100 28000 -85
rect 28050 -100 28150 -85
rect 28200 -100 28300 -85
rect 28350 -100 28450 -85
rect 28500 -100 28600 -85
rect 28650 -100 28750 -85
rect -600 -850 -500 -800
rect -450 -850 -350 -800
rect -600 -865 -350 -850
rect -600 -885 -585 -865
rect -565 -885 -535 -865
rect -515 -885 -485 -865
rect -465 -885 -435 -865
rect -415 -885 -385 -865
rect -365 -885 -350 -865
rect -600 -900 -350 -885
rect -600 -950 -500 -900
rect -450 -950 -350 -900
rect -300 -850 -200 -800
rect -150 -850 -50 -800
rect -300 -865 -50 -850
rect -300 -885 -285 -865
rect -265 -885 -235 -865
rect -215 -885 -185 -865
rect -165 -885 -135 -865
rect -115 -885 -85 -865
rect -65 -885 -50 -865
rect -300 -900 -50 -885
rect -300 -950 -200 -900
rect -150 -950 -50 -900
rect 0 -850 100 -800
rect 150 -850 250 -800
rect 0 -865 250 -850
rect 0 -885 15 -865
rect 35 -885 65 -865
rect 85 -885 115 -865
rect 135 -885 165 -865
rect 185 -885 215 -865
rect 235 -885 250 -865
rect 0 -900 250 -885
rect 0 -950 100 -900
rect 150 -950 250 -900
rect 300 -850 400 -800
rect 450 -850 550 -800
rect 300 -865 550 -850
rect 300 -885 315 -865
rect 335 -885 365 -865
rect 385 -885 415 -865
rect 435 -885 465 -865
rect 485 -885 515 -865
rect 535 -885 550 -865
rect 300 -900 550 -885
rect 300 -950 400 -900
rect 450 -950 550 -900
rect 600 -850 700 -800
rect 750 -850 850 -800
rect 600 -865 850 -850
rect 600 -885 615 -865
rect 635 -885 665 -865
rect 685 -885 715 -865
rect 735 -885 765 -865
rect 785 -885 815 -865
rect 835 -885 850 -865
rect 600 -900 850 -885
rect 600 -950 700 -900
rect 750 -950 850 -900
rect 900 -850 1000 -800
rect 1050 -850 1150 -800
rect 900 -865 1150 -850
rect 900 -885 915 -865
rect 935 -885 965 -865
rect 985 -885 1015 -865
rect 1035 -885 1065 -865
rect 1085 -885 1115 -865
rect 1135 -885 1150 -865
rect 900 -900 1150 -885
rect 900 -950 1000 -900
rect 1050 -950 1150 -900
rect 1200 -850 1300 -800
rect 1350 -850 1450 -800
rect 1200 -865 1450 -850
rect 1200 -885 1215 -865
rect 1235 -885 1265 -865
rect 1285 -885 1315 -865
rect 1335 -885 1365 -865
rect 1385 -885 1415 -865
rect 1435 -885 1450 -865
rect 1200 -900 1450 -885
rect 1200 -950 1300 -900
rect 1350 -950 1450 -900
rect 1500 -850 1600 -800
rect 1650 -850 1750 -800
rect 1500 -865 1750 -850
rect 1500 -885 1515 -865
rect 1535 -885 1565 -865
rect 1585 -885 1615 -865
rect 1635 -885 1665 -865
rect 1685 -885 1715 -865
rect 1735 -885 1750 -865
rect 1500 -900 1750 -885
rect 1500 -950 1600 -900
rect 1650 -950 1750 -900
rect 1800 -850 1900 -800
rect 1950 -850 2050 -800
rect 1800 -865 2050 -850
rect 1800 -885 1815 -865
rect 1835 -885 1865 -865
rect 1885 -885 1915 -865
rect 1935 -885 1965 -865
rect 1985 -885 2015 -865
rect 2035 -885 2050 -865
rect 1800 -900 2050 -885
rect 1800 -950 1900 -900
rect 1950 -950 2050 -900
rect 2100 -850 2200 -800
rect 2250 -850 2350 -800
rect 2100 -865 2350 -850
rect 2100 -885 2115 -865
rect 2135 -885 2165 -865
rect 2185 -885 2215 -865
rect 2235 -885 2265 -865
rect 2285 -885 2315 -865
rect 2335 -885 2350 -865
rect 2100 -900 2350 -885
rect 2100 -950 2200 -900
rect 2250 -950 2350 -900
rect 2400 -850 2500 -800
rect 2550 -850 2650 -800
rect 2400 -865 2650 -850
rect 2400 -885 2415 -865
rect 2435 -885 2465 -865
rect 2485 -885 2515 -865
rect 2535 -885 2565 -865
rect 2585 -885 2615 -865
rect 2635 -885 2650 -865
rect 2400 -900 2650 -885
rect 2400 -950 2500 -900
rect 2550 -950 2650 -900
rect 2700 -850 2800 -800
rect 2850 -850 2950 -800
rect 2700 -865 2950 -850
rect 2700 -885 2715 -865
rect 2735 -885 2765 -865
rect 2785 -885 2815 -865
rect 2835 -885 2865 -865
rect 2885 -885 2915 -865
rect 2935 -885 2950 -865
rect 2700 -900 2950 -885
rect 2700 -950 2800 -900
rect 2850 -950 2950 -900
rect 3000 -850 3100 -800
rect 3150 -850 3250 -800
rect 3000 -865 3250 -850
rect 3000 -885 3015 -865
rect 3035 -885 3065 -865
rect 3085 -885 3115 -865
rect 3135 -885 3165 -865
rect 3185 -885 3215 -865
rect 3235 -885 3250 -865
rect 3000 -900 3250 -885
rect 3000 -950 3100 -900
rect 3150 -950 3250 -900
rect 3300 -850 3400 -800
rect 3450 -850 3550 -800
rect 3300 -865 3550 -850
rect 3300 -885 3315 -865
rect 3335 -885 3365 -865
rect 3385 -885 3415 -865
rect 3435 -885 3465 -865
rect 3485 -885 3515 -865
rect 3535 -885 3550 -865
rect 3300 -900 3550 -885
rect 3300 -950 3400 -900
rect 3450 -950 3550 -900
rect 3600 -850 3700 -800
rect 3750 -850 3850 -800
rect 3600 -865 3850 -850
rect 3600 -885 3615 -865
rect 3635 -885 3665 -865
rect 3685 -885 3715 -865
rect 3735 -885 3765 -865
rect 3785 -885 3815 -865
rect 3835 -885 3850 -865
rect 3600 -900 3850 -885
rect 3600 -950 3700 -900
rect 3750 -950 3850 -900
rect 3900 -850 4000 -800
rect 4050 -850 4150 -800
rect 3900 -865 4150 -850
rect 3900 -885 3915 -865
rect 3935 -885 3965 -865
rect 3985 -885 4015 -865
rect 4035 -885 4065 -865
rect 4085 -885 4115 -865
rect 4135 -885 4150 -865
rect 3900 -900 4150 -885
rect 3900 -950 4000 -900
rect 4050 -950 4150 -900
rect 4200 -850 4300 -800
rect 4350 -850 4450 -800
rect 4200 -865 4450 -850
rect 4200 -885 4215 -865
rect 4235 -885 4265 -865
rect 4285 -885 4315 -865
rect 4335 -885 4365 -865
rect 4385 -885 4415 -865
rect 4435 -885 4450 -865
rect 4200 -900 4450 -885
rect 4200 -950 4300 -900
rect 4350 -950 4450 -900
rect 4500 -850 4600 -800
rect 4650 -850 4750 -800
rect 4500 -865 4750 -850
rect 4500 -885 4515 -865
rect 4535 -885 4565 -865
rect 4585 -885 4615 -865
rect 4635 -885 4665 -865
rect 4685 -885 4715 -865
rect 4735 -885 4750 -865
rect 4500 -900 4750 -885
rect 4500 -950 4600 -900
rect 4650 -950 4750 -900
rect 4800 -850 4900 -800
rect 4950 -850 5050 -800
rect 4800 -865 5050 -850
rect 4800 -885 4815 -865
rect 4835 -885 4865 -865
rect 4885 -885 4915 -865
rect 4935 -885 4965 -865
rect 4985 -885 5015 -865
rect 5035 -885 5050 -865
rect 4800 -900 5050 -885
rect 4800 -950 4900 -900
rect 4950 -950 5050 -900
rect 5100 -850 5200 -800
rect 5250 -850 5350 -800
rect 5100 -865 5350 -850
rect 5100 -885 5115 -865
rect 5135 -885 5165 -865
rect 5185 -885 5215 -865
rect 5235 -885 5265 -865
rect 5285 -885 5315 -865
rect 5335 -885 5350 -865
rect 5100 -900 5350 -885
rect 5100 -950 5200 -900
rect 5250 -950 5350 -900
rect 5400 -850 5500 -800
rect 5550 -850 5650 -800
rect 5400 -865 5650 -850
rect 5400 -885 5415 -865
rect 5435 -885 5465 -865
rect 5485 -885 5515 -865
rect 5535 -885 5565 -865
rect 5585 -885 5615 -865
rect 5635 -885 5650 -865
rect 5400 -900 5650 -885
rect 5400 -950 5500 -900
rect 5550 -950 5650 -900
rect 5700 -850 5800 -800
rect 5850 -850 5950 -800
rect 5700 -865 5950 -850
rect 5700 -885 5715 -865
rect 5735 -885 5765 -865
rect 5785 -885 5815 -865
rect 5835 -885 5865 -865
rect 5885 -885 5915 -865
rect 5935 -885 5950 -865
rect 5700 -900 5950 -885
rect 5700 -950 5800 -900
rect 5850 -950 5950 -900
rect 6000 -850 6100 -800
rect 6150 -850 6250 -800
rect 6000 -865 6250 -850
rect 6000 -885 6015 -865
rect 6035 -885 6065 -865
rect 6085 -885 6115 -865
rect 6135 -885 6165 -865
rect 6185 -885 6215 -865
rect 6235 -885 6250 -865
rect 6000 -900 6250 -885
rect 6000 -950 6100 -900
rect 6150 -950 6250 -900
rect 6300 -850 6400 -800
rect 6450 -850 6550 -800
rect 6300 -865 6550 -850
rect 6300 -885 6315 -865
rect 6335 -885 6365 -865
rect 6385 -885 6415 -865
rect 6435 -885 6465 -865
rect 6485 -885 6515 -865
rect 6535 -885 6550 -865
rect 6300 -900 6550 -885
rect 6300 -950 6400 -900
rect 6450 -950 6550 -900
rect 6600 -850 6700 -800
rect 6750 -850 6850 -800
rect 6600 -865 6850 -850
rect 6600 -885 6615 -865
rect 6635 -885 6665 -865
rect 6685 -885 6715 -865
rect 6735 -885 6765 -865
rect 6785 -885 6815 -865
rect 6835 -885 6850 -865
rect 6600 -900 6850 -885
rect 6600 -950 6700 -900
rect 6750 -950 6850 -900
rect 6900 -850 7000 -800
rect 7050 -850 7150 -800
rect 6900 -865 7150 -850
rect 6900 -885 6915 -865
rect 6935 -885 6965 -865
rect 6985 -885 7015 -865
rect 7035 -885 7065 -865
rect 7085 -885 7115 -865
rect 7135 -885 7150 -865
rect 6900 -900 7150 -885
rect 6900 -950 7000 -900
rect 7050 -950 7150 -900
rect 7200 -850 7300 -800
rect 7350 -850 7450 -800
rect 7200 -865 7450 -850
rect 7200 -885 7215 -865
rect 7235 -885 7265 -865
rect 7285 -885 7315 -865
rect 7335 -885 7365 -865
rect 7385 -885 7415 -865
rect 7435 -885 7450 -865
rect 7200 -900 7450 -885
rect 7200 -950 7300 -900
rect 7350 -950 7450 -900
rect 7500 -850 7600 -800
rect 7650 -850 7750 -800
rect 7500 -865 7750 -850
rect 7500 -885 7515 -865
rect 7535 -885 7565 -865
rect 7585 -885 7615 -865
rect 7635 -885 7665 -865
rect 7685 -885 7715 -865
rect 7735 -885 7750 -865
rect 7500 -900 7750 -885
rect 7500 -950 7600 -900
rect 7650 -950 7750 -900
rect 7800 -850 7900 -800
rect 7950 -850 8050 -800
rect 7800 -865 8050 -850
rect 7800 -885 7815 -865
rect 7835 -885 7865 -865
rect 7885 -885 7915 -865
rect 7935 -885 7965 -865
rect 7985 -885 8015 -865
rect 8035 -885 8050 -865
rect 7800 -900 8050 -885
rect 7800 -950 7900 -900
rect 7950 -950 8050 -900
rect 8100 -850 8200 -800
rect 8250 -850 8350 -800
rect 8100 -865 8350 -850
rect 8100 -885 8115 -865
rect 8135 -885 8165 -865
rect 8185 -885 8215 -865
rect 8235 -885 8265 -865
rect 8285 -885 8315 -865
rect 8335 -885 8350 -865
rect 8100 -900 8350 -885
rect 8100 -950 8200 -900
rect 8250 -950 8350 -900
rect 8400 -850 8500 -800
rect 8550 -850 8650 -800
rect 8400 -865 8650 -850
rect 8400 -885 8415 -865
rect 8435 -885 8465 -865
rect 8485 -885 8515 -865
rect 8535 -885 8565 -865
rect 8585 -885 8615 -865
rect 8635 -885 8650 -865
rect 8400 -900 8650 -885
rect 8400 -950 8500 -900
rect 8550 -950 8650 -900
rect 8700 -850 8800 -800
rect 8850 -850 8950 -800
rect 8700 -865 8950 -850
rect 8700 -885 8715 -865
rect 8735 -885 8765 -865
rect 8785 -885 8815 -865
rect 8835 -885 8865 -865
rect 8885 -885 8915 -865
rect 8935 -885 8950 -865
rect 8700 -900 8950 -885
rect 8700 -950 8800 -900
rect 8850 -950 8950 -900
rect 9000 -850 9100 -800
rect 9150 -850 9250 -800
rect 9000 -865 9250 -850
rect 9000 -885 9015 -865
rect 9035 -885 9065 -865
rect 9085 -885 9115 -865
rect 9135 -885 9165 -865
rect 9185 -885 9215 -865
rect 9235 -885 9250 -865
rect 9000 -900 9250 -885
rect 9000 -950 9100 -900
rect 9150 -950 9250 -900
rect 9300 -850 9400 -800
rect 9450 -850 9550 -800
rect 9300 -865 9550 -850
rect 9300 -885 9315 -865
rect 9335 -885 9365 -865
rect 9385 -885 9415 -865
rect 9435 -885 9465 -865
rect 9485 -885 9515 -865
rect 9535 -885 9550 -865
rect 9300 -900 9550 -885
rect 9300 -950 9400 -900
rect 9450 -950 9550 -900
rect 9600 -850 9700 -800
rect 9750 -850 9850 -800
rect 9600 -865 9850 -850
rect 9600 -885 9615 -865
rect 9635 -885 9665 -865
rect 9685 -885 9715 -865
rect 9735 -885 9765 -865
rect 9785 -885 9815 -865
rect 9835 -885 9850 -865
rect 9600 -900 9850 -885
rect 9600 -950 9700 -900
rect 9750 -950 9850 -900
rect 9900 -850 10000 -800
rect 10050 -850 10150 -800
rect 9900 -865 10150 -850
rect 9900 -885 9915 -865
rect 9935 -885 9965 -865
rect 9985 -885 10015 -865
rect 10035 -885 10065 -865
rect 10085 -885 10115 -865
rect 10135 -885 10150 -865
rect 9900 -900 10150 -885
rect 9900 -950 10000 -900
rect 10050 -950 10150 -900
rect 10200 -850 10300 -800
rect 10350 -850 10450 -800
rect 10200 -865 10450 -850
rect 10200 -885 10215 -865
rect 10235 -885 10265 -865
rect 10285 -885 10315 -865
rect 10335 -885 10365 -865
rect 10385 -885 10415 -865
rect 10435 -885 10450 -865
rect 10200 -900 10450 -885
rect 10200 -950 10300 -900
rect 10350 -950 10450 -900
rect 10500 -850 10600 -800
rect 10650 -850 10750 -800
rect 10500 -865 10750 -850
rect 10500 -885 10515 -865
rect 10535 -885 10565 -865
rect 10585 -885 10615 -865
rect 10635 -885 10665 -865
rect 10685 -885 10715 -865
rect 10735 -885 10750 -865
rect 10500 -900 10750 -885
rect 10500 -950 10600 -900
rect 10650 -950 10750 -900
rect 10800 -850 10900 -800
rect 10950 -850 11050 -800
rect 10800 -865 11050 -850
rect 10800 -885 10815 -865
rect 10835 -885 10865 -865
rect 10885 -885 10915 -865
rect 10935 -885 10965 -865
rect 10985 -885 11015 -865
rect 11035 -885 11050 -865
rect 10800 -900 11050 -885
rect 10800 -950 10900 -900
rect 10950 -950 11050 -900
rect 11100 -850 11200 -800
rect 11250 -850 11350 -800
rect 11100 -865 11350 -850
rect 11100 -885 11115 -865
rect 11135 -885 11165 -865
rect 11185 -885 11215 -865
rect 11235 -885 11265 -865
rect 11285 -885 11315 -865
rect 11335 -885 11350 -865
rect 11100 -900 11350 -885
rect 11100 -950 11200 -900
rect 11250 -950 11350 -900
rect 11400 -850 11500 -800
rect 11550 -850 11650 -800
rect 11400 -865 11650 -850
rect 11400 -885 11415 -865
rect 11435 -885 11465 -865
rect 11485 -885 11515 -865
rect 11535 -885 11565 -865
rect 11585 -885 11615 -865
rect 11635 -885 11650 -865
rect 11400 -900 11650 -885
rect 11400 -950 11500 -900
rect 11550 -950 11650 -900
rect 11700 -850 11800 -800
rect 11850 -850 11950 -800
rect 11700 -865 11950 -850
rect 11700 -885 11715 -865
rect 11735 -885 11765 -865
rect 11785 -885 11815 -865
rect 11835 -885 11865 -865
rect 11885 -885 11915 -865
rect 11935 -885 11950 -865
rect 11700 -900 11950 -885
rect 11700 -950 11800 -900
rect 11850 -950 11950 -900
rect 12000 -850 12100 -800
rect 12150 -850 12250 -800
rect 12000 -865 12250 -850
rect 12000 -885 12015 -865
rect 12035 -885 12065 -865
rect 12085 -885 12115 -865
rect 12135 -885 12165 -865
rect 12185 -885 12215 -865
rect 12235 -885 12250 -865
rect 12000 -900 12250 -885
rect 12000 -950 12100 -900
rect 12150 -950 12250 -900
rect 12300 -850 12400 -800
rect 12450 -850 12550 -800
rect 12300 -865 12550 -850
rect 12300 -885 12315 -865
rect 12335 -885 12365 -865
rect 12385 -885 12415 -865
rect 12435 -885 12465 -865
rect 12485 -885 12515 -865
rect 12535 -885 12550 -865
rect 12300 -900 12550 -885
rect 12300 -950 12400 -900
rect 12450 -950 12550 -900
rect 12600 -850 12700 -800
rect 12750 -850 12850 -800
rect 12600 -865 12850 -850
rect 12600 -885 12615 -865
rect 12635 -885 12665 -865
rect 12685 -885 12715 -865
rect 12735 -885 12765 -865
rect 12785 -885 12815 -865
rect 12835 -885 12850 -865
rect 12600 -900 12850 -885
rect 12600 -950 12700 -900
rect 12750 -950 12850 -900
rect 12900 -850 13000 -800
rect 13050 -850 13150 -800
rect 12900 -865 13150 -850
rect 12900 -885 12915 -865
rect 12935 -885 12965 -865
rect 12985 -885 13015 -865
rect 13035 -885 13065 -865
rect 13085 -885 13115 -865
rect 13135 -885 13150 -865
rect 12900 -900 13150 -885
rect 12900 -950 13000 -900
rect 13050 -950 13150 -900
rect 13200 -850 13300 -800
rect 13350 -850 13450 -800
rect 13200 -865 13450 -850
rect 13200 -885 13215 -865
rect 13235 -885 13265 -865
rect 13285 -885 13315 -865
rect 13335 -885 13365 -865
rect 13385 -885 13415 -865
rect 13435 -885 13450 -865
rect 13200 -900 13450 -885
rect 13200 -950 13300 -900
rect 13350 -950 13450 -900
rect 13500 -850 13600 -800
rect 13650 -850 13750 -800
rect 13500 -865 13750 -850
rect 13500 -885 13515 -865
rect 13535 -885 13565 -865
rect 13585 -885 13615 -865
rect 13635 -885 13665 -865
rect 13685 -885 13715 -865
rect 13735 -885 13750 -865
rect 13500 -900 13750 -885
rect 13500 -950 13600 -900
rect 13650 -950 13750 -900
rect 13800 -850 13900 -800
rect 13950 -850 14050 -800
rect 13800 -865 14050 -850
rect 13800 -885 13815 -865
rect 13835 -885 13865 -865
rect 13885 -885 13915 -865
rect 13935 -885 13965 -865
rect 13985 -885 14015 -865
rect 14035 -885 14050 -865
rect 13800 -900 14050 -885
rect 13800 -950 13900 -900
rect 13950 -950 14050 -900
rect 14100 -850 14200 -800
rect 14250 -850 14350 -800
rect 14100 -865 14350 -850
rect 14100 -885 14115 -865
rect 14135 -885 14165 -865
rect 14185 -885 14215 -865
rect 14235 -885 14265 -865
rect 14285 -885 14315 -865
rect 14335 -885 14350 -865
rect 14100 -900 14350 -885
rect 14100 -950 14200 -900
rect 14250 -950 14350 -900
rect 14400 -850 14500 -800
rect 14550 -850 14650 -800
rect 14400 -865 14650 -850
rect 14400 -885 14415 -865
rect 14435 -885 14465 -865
rect 14485 -885 14515 -865
rect 14535 -885 14565 -865
rect 14585 -885 14615 -865
rect 14635 -885 14650 -865
rect 14400 -900 14650 -885
rect 14400 -950 14500 -900
rect 14550 -950 14650 -900
rect 14700 -850 14800 -800
rect 14850 -850 14950 -800
rect 14700 -865 14950 -850
rect 14700 -885 14715 -865
rect 14735 -885 14765 -865
rect 14785 -885 14815 -865
rect 14835 -885 14865 -865
rect 14885 -885 14915 -865
rect 14935 -885 14950 -865
rect 14700 -900 14950 -885
rect 14700 -950 14800 -900
rect 14850 -950 14950 -900
rect 15000 -850 15100 -800
rect 15150 -850 15250 -800
rect 15000 -865 15250 -850
rect 15000 -885 15015 -865
rect 15035 -885 15065 -865
rect 15085 -885 15115 -865
rect 15135 -885 15165 -865
rect 15185 -885 15215 -865
rect 15235 -885 15250 -865
rect 15000 -900 15250 -885
rect 15000 -950 15100 -900
rect 15150 -950 15250 -900
rect 15300 -850 15400 -800
rect 15450 -850 15550 -800
rect 15300 -865 15550 -850
rect 15300 -885 15315 -865
rect 15335 -885 15365 -865
rect 15385 -885 15415 -865
rect 15435 -885 15465 -865
rect 15485 -885 15515 -865
rect 15535 -885 15550 -865
rect 15300 -900 15550 -885
rect 15300 -950 15400 -900
rect 15450 -950 15550 -900
rect 15600 -850 15700 -800
rect 15750 -850 15850 -800
rect 15600 -865 15850 -850
rect 15600 -885 15615 -865
rect 15635 -885 15665 -865
rect 15685 -885 15715 -865
rect 15735 -885 15765 -865
rect 15785 -885 15815 -865
rect 15835 -885 15850 -865
rect 15600 -900 15850 -885
rect 15600 -950 15700 -900
rect 15750 -950 15850 -900
rect 15900 -850 16000 -800
rect 16050 -850 16150 -800
rect 15900 -865 16150 -850
rect 15900 -885 15915 -865
rect 15935 -885 15965 -865
rect 15985 -885 16015 -865
rect 16035 -885 16065 -865
rect 16085 -885 16115 -865
rect 16135 -885 16150 -865
rect 15900 -900 16150 -885
rect 15900 -950 16000 -900
rect 16050 -950 16150 -900
rect 16200 -850 16300 -800
rect 16350 -850 16450 -800
rect 16200 -865 16450 -850
rect 16200 -885 16215 -865
rect 16235 -885 16265 -865
rect 16285 -885 16315 -865
rect 16335 -885 16365 -865
rect 16385 -885 16415 -865
rect 16435 -885 16450 -865
rect 16200 -900 16450 -885
rect 16200 -950 16300 -900
rect 16350 -950 16450 -900
rect 16500 -850 16600 -800
rect 16650 -850 16750 -800
rect 16500 -865 16750 -850
rect 16500 -885 16515 -865
rect 16535 -885 16565 -865
rect 16585 -885 16615 -865
rect 16635 -885 16665 -865
rect 16685 -885 16715 -865
rect 16735 -885 16750 -865
rect 16500 -900 16750 -885
rect 16500 -950 16600 -900
rect 16650 -950 16750 -900
rect 16800 -850 16900 -800
rect 16950 -850 17050 -800
rect 16800 -865 17050 -850
rect 16800 -885 16815 -865
rect 16835 -885 16865 -865
rect 16885 -885 16915 -865
rect 16935 -885 16965 -865
rect 16985 -885 17015 -865
rect 17035 -885 17050 -865
rect 16800 -900 17050 -885
rect 16800 -950 16900 -900
rect 16950 -950 17050 -900
rect 17100 -850 17200 -800
rect 17250 -850 17350 -800
rect 17100 -865 17350 -850
rect 17100 -885 17115 -865
rect 17135 -885 17165 -865
rect 17185 -885 17215 -865
rect 17235 -885 17265 -865
rect 17285 -885 17315 -865
rect 17335 -885 17350 -865
rect 17100 -900 17350 -885
rect 17100 -950 17200 -900
rect 17250 -950 17350 -900
rect 17400 -850 17500 -800
rect 17550 -850 17650 -800
rect 17400 -865 17650 -850
rect 17400 -885 17415 -865
rect 17435 -885 17465 -865
rect 17485 -885 17515 -865
rect 17535 -885 17565 -865
rect 17585 -885 17615 -865
rect 17635 -885 17650 -865
rect 17400 -900 17650 -885
rect 17400 -950 17500 -900
rect 17550 -950 17650 -900
rect 17700 -850 17800 -800
rect 17850 -850 17950 -800
rect 17700 -865 17950 -850
rect 17700 -885 17715 -865
rect 17735 -885 17765 -865
rect 17785 -885 17815 -865
rect 17835 -885 17865 -865
rect 17885 -885 17915 -865
rect 17935 -885 17950 -865
rect 17700 -900 17950 -885
rect 17700 -950 17800 -900
rect 17850 -950 17950 -900
rect 18000 -850 18100 -800
rect 18150 -850 18250 -800
rect 18000 -865 18250 -850
rect 18000 -885 18015 -865
rect 18035 -885 18065 -865
rect 18085 -885 18115 -865
rect 18135 -885 18165 -865
rect 18185 -885 18215 -865
rect 18235 -885 18250 -865
rect 18000 -900 18250 -885
rect 18000 -950 18100 -900
rect 18150 -950 18250 -900
rect 18300 -850 18400 -800
rect 18450 -850 18550 -800
rect 18300 -865 18550 -850
rect 18300 -885 18315 -865
rect 18335 -885 18365 -865
rect 18385 -885 18415 -865
rect 18435 -885 18465 -865
rect 18485 -885 18515 -865
rect 18535 -885 18550 -865
rect 18300 -900 18550 -885
rect 18300 -950 18400 -900
rect 18450 -950 18550 -900
rect 18600 -850 18700 -800
rect 18750 -850 18850 -800
rect 18600 -865 18850 -850
rect 18600 -885 18615 -865
rect 18635 -885 18665 -865
rect 18685 -885 18715 -865
rect 18735 -885 18765 -865
rect 18785 -885 18815 -865
rect 18835 -885 18850 -865
rect 18600 -900 18850 -885
rect 18600 -950 18700 -900
rect 18750 -950 18850 -900
rect 18900 -850 19000 -800
rect 19050 -850 19150 -800
rect 18900 -865 19150 -850
rect 18900 -885 18915 -865
rect 18935 -885 18965 -865
rect 18985 -885 19015 -865
rect 19035 -885 19065 -865
rect 19085 -885 19115 -865
rect 19135 -885 19150 -865
rect 18900 -900 19150 -885
rect 18900 -950 19000 -900
rect 19050 -950 19150 -900
rect 19200 -850 19300 -800
rect 19350 -850 19450 -800
rect 19200 -865 19450 -850
rect 19200 -885 19215 -865
rect 19235 -885 19265 -865
rect 19285 -885 19315 -865
rect 19335 -885 19365 -865
rect 19385 -885 19415 -865
rect 19435 -885 19450 -865
rect 19200 -900 19450 -885
rect 19200 -950 19300 -900
rect 19350 -950 19450 -900
rect 19500 -850 19600 -800
rect 19650 -850 19750 -800
rect 19500 -865 19750 -850
rect 19500 -885 19515 -865
rect 19535 -885 19565 -865
rect 19585 -885 19615 -865
rect 19635 -885 19665 -865
rect 19685 -885 19715 -865
rect 19735 -885 19750 -865
rect 19500 -900 19750 -885
rect 19500 -950 19600 -900
rect 19650 -950 19750 -900
rect 19800 -850 19900 -800
rect 19950 -850 20050 -800
rect 19800 -865 20050 -850
rect 19800 -885 19815 -865
rect 19835 -885 19865 -865
rect 19885 -885 19915 -865
rect 19935 -885 19965 -865
rect 19985 -885 20015 -865
rect 20035 -885 20050 -865
rect 19800 -900 20050 -885
rect 19800 -950 19900 -900
rect 19950 -950 20050 -900
rect 20100 -850 20200 -800
rect 20250 -850 20350 -800
rect 20100 -865 20350 -850
rect 20100 -885 20115 -865
rect 20135 -885 20165 -865
rect 20185 -885 20215 -865
rect 20235 -885 20265 -865
rect 20285 -885 20315 -865
rect 20335 -885 20350 -865
rect 20100 -900 20350 -885
rect 20100 -950 20200 -900
rect 20250 -950 20350 -900
rect 20400 -850 20500 -800
rect 20550 -850 20650 -800
rect 20400 -865 20650 -850
rect 20400 -885 20415 -865
rect 20435 -885 20465 -865
rect 20485 -885 20515 -865
rect 20535 -885 20565 -865
rect 20585 -885 20615 -865
rect 20635 -885 20650 -865
rect 20400 -900 20650 -885
rect 20400 -950 20500 -900
rect 20550 -950 20650 -900
rect 20700 -850 20800 -800
rect 20850 -850 20950 -800
rect 20700 -865 20950 -850
rect 20700 -885 20715 -865
rect 20735 -885 20765 -865
rect 20785 -885 20815 -865
rect 20835 -885 20865 -865
rect 20885 -885 20915 -865
rect 20935 -885 20950 -865
rect 20700 -900 20950 -885
rect 20700 -950 20800 -900
rect 20850 -950 20950 -900
rect 21000 -850 21100 -800
rect 21150 -850 21250 -800
rect 21000 -865 21250 -850
rect 21000 -885 21015 -865
rect 21035 -885 21065 -865
rect 21085 -885 21115 -865
rect 21135 -885 21165 -865
rect 21185 -885 21215 -865
rect 21235 -885 21250 -865
rect 21000 -900 21250 -885
rect 21000 -950 21100 -900
rect 21150 -950 21250 -900
rect 21300 -850 21400 -800
rect 21450 -850 21550 -800
rect 21300 -865 21550 -850
rect 21300 -885 21315 -865
rect 21335 -885 21365 -865
rect 21385 -885 21415 -865
rect 21435 -885 21465 -865
rect 21485 -885 21515 -865
rect 21535 -885 21550 -865
rect 21300 -900 21550 -885
rect 21300 -950 21400 -900
rect 21450 -950 21550 -900
rect 21600 -850 21700 -800
rect 21750 -850 21850 -800
rect 21600 -865 21850 -850
rect 21600 -885 21615 -865
rect 21635 -885 21665 -865
rect 21685 -885 21715 -865
rect 21735 -885 21765 -865
rect 21785 -885 21815 -865
rect 21835 -885 21850 -865
rect 21600 -900 21850 -885
rect 21600 -950 21700 -900
rect 21750 -950 21850 -900
rect 21900 -850 22000 -800
rect 22050 -850 22150 -800
rect 21900 -865 22150 -850
rect 21900 -885 21915 -865
rect 21935 -885 21965 -865
rect 21985 -885 22015 -865
rect 22035 -885 22065 -865
rect 22085 -885 22115 -865
rect 22135 -885 22150 -865
rect 21900 -900 22150 -885
rect 21900 -950 22000 -900
rect 22050 -950 22150 -900
rect 22200 -850 22300 -800
rect 22350 -850 22450 -800
rect 22200 -865 22450 -850
rect 22200 -885 22215 -865
rect 22235 -885 22265 -865
rect 22285 -885 22315 -865
rect 22335 -885 22365 -865
rect 22385 -885 22415 -865
rect 22435 -885 22450 -865
rect 22200 -900 22450 -885
rect 22200 -950 22300 -900
rect 22350 -950 22450 -900
rect 22500 -850 22600 -800
rect 22650 -850 22750 -800
rect 22500 -865 22750 -850
rect 22500 -885 22515 -865
rect 22535 -885 22565 -865
rect 22585 -885 22615 -865
rect 22635 -885 22665 -865
rect 22685 -885 22715 -865
rect 22735 -885 22750 -865
rect 22500 -900 22750 -885
rect 22500 -950 22600 -900
rect 22650 -950 22750 -900
rect 22800 -850 22900 -800
rect 22950 -850 23050 -800
rect 22800 -865 23050 -850
rect 22800 -885 22815 -865
rect 22835 -885 22865 -865
rect 22885 -885 22915 -865
rect 22935 -885 22965 -865
rect 22985 -885 23015 -865
rect 23035 -885 23050 -865
rect 22800 -900 23050 -885
rect 22800 -950 22900 -900
rect 22950 -950 23050 -900
rect 23100 -850 23200 -800
rect 23250 -850 23350 -800
rect 23100 -865 23350 -850
rect 23100 -885 23115 -865
rect 23135 -885 23165 -865
rect 23185 -885 23215 -865
rect 23235 -885 23265 -865
rect 23285 -885 23315 -865
rect 23335 -885 23350 -865
rect 23100 -900 23350 -885
rect 23100 -950 23200 -900
rect 23250 -950 23350 -900
rect 23400 -850 23500 -800
rect 23550 -850 23650 -800
rect 23400 -865 23650 -850
rect 23400 -885 23415 -865
rect 23435 -885 23465 -865
rect 23485 -885 23515 -865
rect 23535 -885 23565 -865
rect 23585 -885 23615 -865
rect 23635 -885 23650 -865
rect 23400 -900 23650 -885
rect 23400 -950 23500 -900
rect 23550 -950 23650 -900
rect 23700 -850 23800 -800
rect 23850 -850 23950 -800
rect 23700 -865 23950 -850
rect 23700 -885 23715 -865
rect 23735 -885 23765 -865
rect 23785 -885 23815 -865
rect 23835 -885 23865 -865
rect 23885 -885 23915 -865
rect 23935 -885 23950 -865
rect 23700 -900 23950 -885
rect 23700 -950 23800 -900
rect 23850 -950 23950 -900
rect 24000 -850 24100 -800
rect 24150 -850 24250 -800
rect 24000 -865 24250 -850
rect 24000 -885 24015 -865
rect 24035 -885 24065 -865
rect 24085 -885 24115 -865
rect 24135 -885 24165 -865
rect 24185 -885 24215 -865
rect 24235 -885 24250 -865
rect 24000 -900 24250 -885
rect 24000 -950 24100 -900
rect 24150 -950 24250 -900
rect 24300 -850 24400 -800
rect 24450 -850 24550 -800
rect 24300 -865 24550 -850
rect 24300 -885 24315 -865
rect 24335 -885 24365 -865
rect 24385 -885 24415 -865
rect 24435 -885 24465 -865
rect 24485 -885 24515 -865
rect 24535 -885 24550 -865
rect 24300 -900 24550 -885
rect 24300 -950 24400 -900
rect 24450 -950 24550 -900
rect 24600 -850 24700 -800
rect 24750 -850 24850 -800
rect 24600 -865 24850 -850
rect 24600 -885 24615 -865
rect 24635 -885 24665 -865
rect 24685 -885 24715 -865
rect 24735 -885 24765 -865
rect 24785 -885 24815 -865
rect 24835 -885 24850 -865
rect 24600 -900 24850 -885
rect 24600 -950 24700 -900
rect 24750 -950 24850 -900
rect 24900 -850 25000 -800
rect 25050 -850 25150 -800
rect 24900 -865 25150 -850
rect 24900 -885 24915 -865
rect 24935 -885 24965 -865
rect 24985 -885 25015 -865
rect 25035 -885 25065 -865
rect 25085 -885 25115 -865
rect 25135 -885 25150 -865
rect 24900 -900 25150 -885
rect 24900 -950 25000 -900
rect 25050 -950 25150 -900
rect 25200 -850 25300 -800
rect 25350 -850 25450 -800
rect 25200 -865 25450 -850
rect 25200 -885 25215 -865
rect 25235 -885 25265 -865
rect 25285 -885 25315 -865
rect 25335 -885 25365 -865
rect 25385 -885 25415 -865
rect 25435 -885 25450 -865
rect 25200 -900 25450 -885
rect 25200 -950 25300 -900
rect 25350 -950 25450 -900
rect 25500 -850 25600 -800
rect 25650 -850 25750 -800
rect 25500 -865 25750 -850
rect 25500 -885 25515 -865
rect 25535 -885 25565 -865
rect 25585 -885 25615 -865
rect 25635 -885 25665 -865
rect 25685 -885 25715 -865
rect 25735 -885 25750 -865
rect 25500 -900 25750 -885
rect 25500 -950 25600 -900
rect 25650 -950 25750 -900
rect 25800 -850 25900 -800
rect 25950 -850 26050 -800
rect 25800 -865 26050 -850
rect 25800 -885 25815 -865
rect 25835 -885 25865 -865
rect 25885 -885 25915 -865
rect 25935 -885 25965 -865
rect 25985 -885 26015 -865
rect 26035 -885 26050 -865
rect 25800 -900 26050 -885
rect 25800 -950 25900 -900
rect 25950 -950 26050 -900
rect 26100 -850 26200 -800
rect 26250 -850 26350 -800
rect 26100 -865 26350 -850
rect 26100 -885 26115 -865
rect 26135 -885 26165 -865
rect 26185 -885 26215 -865
rect 26235 -885 26265 -865
rect 26285 -885 26315 -865
rect 26335 -885 26350 -865
rect 26100 -900 26350 -885
rect 26100 -950 26200 -900
rect 26250 -950 26350 -900
rect 26400 -850 26500 -800
rect 26550 -850 26650 -800
rect 26400 -865 26650 -850
rect 26400 -885 26415 -865
rect 26435 -885 26465 -865
rect 26485 -885 26515 -865
rect 26535 -885 26565 -865
rect 26585 -885 26615 -865
rect 26635 -885 26650 -865
rect 26400 -900 26650 -885
rect 26400 -950 26500 -900
rect 26550 -950 26650 -900
rect 26700 -850 26800 -800
rect 26850 -850 26950 -800
rect 26700 -865 26950 -850
rect 26700 -885 26715 -865
rect 26735 -885 26765 -865
rect 26785 -885 26815 -865
rect 26835 -885 26865 -865
rect 26885 -885 26915 -865
rect 26935 -885 26950 -865
rect 26700 -900 26950 -885
rect 26700 -950 26800 -900
rect 26850 -950 26950 -900
rect 27000 -850 27100 -800
rect 27150 -850 27250 -800
rect 27000 -865 27250 -850
rect 27000 -885 27015 -865
rect 27035 -885 27065 -865
rect 27085 -885 27115 -865
rect 27135 -885 27165 -865
rect 27185 -885 27215 -865
rect 27235 -885 27250 -865
rect 27000 -900 27250 -885
rect 27000 -950 27100 -900
rect 27150 -950 27250 -900
rect 27300 -850 27400 -800
rect 27450 -850 27550 -800
rect 27300 -865 27550 -850
rect 27300 -885 27315 -865
rect 27335 -885 27365 -865
rect 27385 -885 27415 -865
rect 27435 -885 27465 -865
rect 27485 -885 27515 -865
rect 27535 -885 27550 -865
rect 27300 -900 27550 -885
rect 27300 -950 27400 -900
rect 27450 -950 27550 -900
rect 27600 -850 27700 -800
rect 27750 -850 27850 -800
rect 27600 -865 27850 -850
rect 27600 -885 27615 -865
rect 27635 -885 27665 -865
rect 27685 -885 27715 -865
rect 27735 -885 27765 -865
rect 27785 -885 27815 -865
rect 27835 -885 27850 -865
rect 27600 -900 27850 -885
rect 27600 -950 27700 -900
rect 27750 -950 27850 -900
rect 27900 -850 28000 -800
rect 28050 -850 28150 -800
rect 27900 -865 28150 -850
rect 27900 -885 27915 -865
rect 27935 -885 27965 -865
rect 27985 -885 28015 -865
rect 28035 -885 28065 -865
rect 28085 -885 28115 -865
rect 28135 -885 28150 -865
rect 27900 -900 28150 -885
rect 27900 -950 28000 -900
rect 28050 -950 28150 -900
rect 28200 -850 28300 -800
rect 28350 -850 28450 -800
rect 28200 -865 28450 -850
rect 28200 -885 28215 -865
rect 28235 -885 28265 -865
rect 28285 -885 28315 -865
rect 28335 -885 28365 -865
rect 28385 -885 28415 -865
rect 28435 -885 28450 -865
rect 28200 -900 28450 -885
rect 28200 -950 28300 -900
rect 28350 -950 28450 -900
rect 28500 -850 28600 -800
rect 28650 -850 28750 -800
rect 28500 -865 28750 -850
rect 28500 -885 28515 -865
rect 28535 -885 28565 -865
rect 28585 -885 28615 -865
rect 28635 -885 28665 -865
rect 28685 -885 28715 -865
rect 28735 -885 28750 -865
rect 28500 -900 28750 -885
rect 28500 -950 28600 -900
rect 28650 -950 28750 -900
rect -600 -1665 -500 -1650
rect -450 -1665 -350 -1650
rect -300 -1665 -200 -1650
rect -150 -1665 -50 -1650
rect 0 -1665 100 -1650
rect 150 -1665 250 -1650
rect 300 -1665 400 -1650
rect 450 -1665 550 -1650
rect 600 -1665 700 -1650
rect 750 -1665 850 -1650
rect 900 -1665 1000 -1650
rect 1050 -1665 1150 -1650
rect 1200 -1665 1300 -1650
rect 1350 -1665 1450 -1650
rect 1500 -1665 1600 -1650
rect 1650 -1665 1750 -1650
rect 1800 -1665 1900 -1650
rect 1950 -1665 2050 -1650
rect 2100 -1665 2200 -1650
rect 2250 -1665 2350 -1650
rect 2400 -1665 2500 -1650
rect 2550 -1665 2650 -1650
rect 2700 -1665 2800 -1650
rect 2850 -1665 2950 -1650
rect 3000 -1665 3100 -1650
rect 3150 -1665 3250 -1650
rect 3300 -1665 3400 -1650
rect 3450 -1665 3550 -1650
rect 3600 -1665 3700 -1650
rect 3750 -1665 3850 -1650
rect 3900 -1665 4000 -1650
rect 4050 -1665 4150 -1650
rect 4200 -1665 4300 -1650
rect 4350 -1665 4450 -1650
rect 4500 -1665 4600 -1650
rect 4650 -1665 4750 -1650
rect 4800 -1665 4900 -1650
rect 4950 -1665 5050 -1650
rect 5100 -1665 5200 -1650
rect 5250 -1665 5350 -1650
rect 5400 -1665 5500 -1650
rect 5550 -1665 5650 -1650
rect 5700 -1665 5800 -1650
rect 5850 -1665 5950 -1650
rect 6000 -1665 6100 -1650
rect 6150 -1665 6250 -1650
rect 6300 -1665 6400 -1650
rect 6450 -1665 6550 -1650
rect 6600 -1665 6700 -1650
rect 6750 -1665 6850 -1650
rect 6900 -1665 7000 -1650
rect 7050 -1665 7150 -1650
rect 7200 -1665 7300 -1650
rect 7350 -1665 7450 -1650
rect 7500 -1665 7600 -1650
rect 7650 -1665 7750 -1650
rect 7800 -1665 7900 -1650
rect 7950 -1665 8050 -1650
rect 8100 -1665 8200 -1650
rect 8250 -1665 8350 -1650
rect 8400 -1665 8500 -1650
rect 8550 -1665 8650 -1650
rect 8700 -1665 8800 -1650
rect 8850 -1665 8950 -1650
rect 9000 -1665 9100 -1650
rect 9150 -1665 9250 -1650
rect 9300 -1665 9400 -1650
rect 9450 -1665 9550 -1650
rect 9600 -1665 9700 -1650
rect 9750 -1665 9850 -1650
rect 9900 -1665 10000 -1650
rect 10050 -1665 10150 -1650
rect 10200 -1665 10300 -1650
rect 10350 -1665 10450 -1650
rect 10500 -1665 10600 -1650
rect 10650 -1665 10750 -1650
rect 10800 -1665 10900 -1650
rect 10950 -1665 11050 -1650
rect 11100 -1665 11200 -1650
rect 11250 -1665 11350 -1650
rect 11400 -1665 11500 -1650
rect 11550 -1665 11650 -1650
rect 11700 -1665 11800 -1650
rect 11850 -1665 11950 -1650
rect 12000 -1665 12100 -1650
rect 12150 -1665 12250 -1650
rect 12300 -1665 12400 -1650
rect 12450 -1665 12550 -1650
rect 12600 -1665 12700 -1650
rect 12750 -1665 12850 -1650
rect 12900 -1665 13000 -1650
rect 13050 -1665 13150 -1650
rect 13200 -1665 13300 -1650
rect 13350 -1665 13450 -1650
rect 13500 -1665 13600 -1650
rect 13650 -1665 13750 -1650
rect 13800 -1665 13900 -1650
rect 13950 -1665 14050 -1650
rect 14100 -1665 14200 -1650
rect 14250 -1665 14350 -1650
rect 14400 -1665 14500 -1650
rect 14550 -1665 14650 -1650
rect 14700 -1665 14800 -1650
rect 14850 -1665 14950 -1650
rect 15000 -1665 15100 -1650
rect 15150 -1665 15250 -1650
rect 15300 -1665 15400 -1650
rect 15450 -1665 15550 -1650
rect 15600 -1665 15700 -1650
rect 15750 -1665 15850 -1650
rect 15900 -1665 16000 -1650
rect 16050 -1665 16150 -1650
rect 16200 -1665 16300 -1650
rect 16350 -1665 16450 -1650
rect 16500 -1665 16600 -1650
rect 16650 -1665 16750 -1650
rect 16800 -1665 16900 -1650
rect 16950 -1665 17050 -1650
rect 17100 -1665 17200 -1650
rect 17250 -1665 17350 -1650
rect 17400 -1665 17500 -1650
rect 17550 -1665 17650 -1650
rect 17700 -1665 17800 -1650
rect 17850 -1665 17950 -1650
rect 18000 -1665 18100 -1650
rect 18150 -1665 18250 -1650
rect 18300 -1665 18400 -1650
rect 18450 -1665 18550 -1650
rect 18600 -1665 18700 -1650
rect 18750 -1665 18850 -1650
rect 18900 -1665 19000 -1650
rect 19050 -1665 19150 -1650
rect 19200 -1665 19300 -1650
rect 19350 -1665 19450 -1650
rect 19500 -1665 19600 -1650
rect 19650 -1665 19750 -1650
rect 19800 -1665 19900 -1650
rect 19950 -1665 20050 -1650
rect 20100 -1665 20200 -1650
rect 20250 -1665 20350 -1650
rect 20400 -1665 20500 -1650
rect 20550 -1665 20650 -1650
rect 20700 -1665 20800 -1650
rect 20850 -1665 20950 -1650
rect 21000 -1665 21100 -1650
rect 21150 -1665 21250 -1650
rect 21300 -1665 21400 -1650
rect 21450 -1665 21550 -1650
rect 21600 -1665 21700 -1650
rect 21750 -1665 21850 -1650
rect 21900 -1665 22000 -1650
rect 22050 -1665 22150 -1650
rect 22200 -1665 22300 -1650
rect 22350 -1665 22450 -1650
rect 22500 -1665 22600 -1650
rect 22650 -1665 22750 -1650
rect 22800 -1665 22900 -1650
rect 22950 -1665 23050 -1650
rect 23100 -1665 23200 -1650
rect 23250 -1665 23350 -1650
rect 23400 -1665 23500 -1650
rect 23550 -1665 23650 -1650
rect 23700 -1665 23800 -1650
rect 23850 -1665 23950 -1650
rect 24000 -1665 24100 -1650
rect 24150 -1665 24250 -1650
rect 24300 -1665 24400 -1650
rect 24450 -1665 24550 -1650
rect 24600 -1665 24700 -1650
rect 24750 -1665 24850 -1650
rect 24900 -1665 25000 -1650
rect 25050 -1665 25150 -1650
rect 25200 -1665 25300 -1650
rect 25350 -1665 25450 -1650
rect 25500 -1665 25600 -1650
rect 25650 -1665 25750 -1650
rect 25800 -1665 25900 -1650
rect 25950 -1665 26050 -1650
rect 26100 -1665 26200 -1650
rect 26250 -1665 26350 -1650
rect 26400 -1665 26500 -1650
rect 26550 -1665 26650 -1650
rect 26700 -1665 26800 -1650
rect 26850 -1665 26950 -1650
rect 27000 -1665 27100 -1650
rect 27150 -1665 27250 -1650
rect 27300 -1665 27400 -1650
rect 27450 -1665 27550 -1650
rect 27600 -1665 27700 -1650
rect 27750 -1665 27850 -1650
rect 27900 -1665 28000 -1650
rect 28050 -1665 28150 -1650
rect 28200 -1665 28300 -1650
rect 28350 -1665 28450 -1650
rect 28500 -1665 28600 -1650
rect 28650 -1665 28750 -1650
<< polycont >>
rect -585 4915 -565 4935
rect -535 4915 -515 4935
rect -485 4915 -465 4935
rect -435 4915 -415 4935
rect -385 4915 -365 4935
rect -285 4915 -265 4935
rect -235 4915 -215 4935
rect -185 4915 -165 4935
rect -135 4915 -115 4935
rect -85 4915 -65 4935
rect 15 4915 35 4935
rect 65 4915 85 4935
rect 115 4915 135 4935
rect 165 4915 185 4935
rect 215 4915 235 4935
rect 315 4915 335 4935
rect 365 4915 385 4935
rect 415 4915 435 4935
rect 465 4915 485 4935
rect 515 4915 535 4935
rect 615 4915 635 4935
rect 665 4915 685 4935
rect 715 4915 735 4935
rect 765 4915 785 4935
rect 815 4915 835 4935
rect 915 4915 935 4935
rect 965 4915 985 4935
rect 1015 4915 1035 4935
rect 1065 4915 1085 4935
rect 1115 4915 1135 4935
rect 1215 4915 1235 4935
rect 1265 4915 1285 4935
rect 1315 4915 1335 4935
rect 1365 4915 1385 4935
rect 1415 4915 1435 4935
rect 1515 4915 1535 4935
rect 1565 4915 1585 4935
rect 1615 4915 1635 4935
rect 1665 4915 1685 4935
rect 1715 4915 1735 4935
rect 1815 4915 1835 4935
rect 1865 4915 1885 4935
rect 1915 4915 1935 4935
rect 1965 4915 1985 4935
rect 2015 4915 2035 4935
rect 2115 4915 2135 4935
rect 2165 4915 2185 4935
rect 2215 4915 2235 4935
rect 2265 4915 2285 4935
rect 2315 4915 2335 4935
rect 2415 4915 2435 4935
rect 2465 4915 2485 4935
rect 2515 4915 2535 4935
rect 2565 4915 2585 4935
rect 2615 4915 2635 4935
rect 2715 4915 2735 4935
rect 2765 4915 2785 4935
rect 2815 4915 2835 4935
rect 2865 4915 2885 4935
rect 2915 4915 2935 4935
rect 3015 4915 3035 4935
rect 3065 4915 3085 4935
rect 3115 4915 3135 4935
rect 3165 4915 3185 4935
rect 3215 4915 3235 4935
rect 3315 4915 3335 4935
rect 3365 4915 3385 4935
rect 3415 4915 3435 4935
rect 3465 4915 3485 4935
rect 3515 4915 3535 4935
rect 3615 4915 3635 4935
rect 3665 4915 3685 4935
rect 3715 4915 3735 4935
rect 3765 4915 3785 4935
rect 3815 4915 3835 4935
rect 3915 4915 3935 4935
rect 3965 4915 3985 4935
rect 4015 4915 4035 4935
rect 4065 4915 4085 4935
rect 4115 4915 4135 4935
rect 4215 4915 4235 4935
rect 4265 4915 4285 4935
rect 4315 4915 4335 4935
rect 4365 4915 4385 4935
rect 4415 4915 4435 4935
rect 4515 4915 4535 4935
rect 4565 4915 4585 4935
rect 4615 4915 4635 4935
rect 4665 4915 4685 4935
rect 4715 4915 4735 4935
rect 4815 4915 4835 4935
rect 4865 4915 4885 4935
rect 4915 4915 4935 4935
rect 4965 4915 4985 4935
rect 5015 4915 5035 4935
rect 5115 4915 5135 4935
rect 5165 4915 5185 4935
rect 5215 4915 5235 4935
rect 5265 4915 5285 4935
rect 5315 4915 5335 4935
rect 5415 4915 5435 4935
rect 5465 4915 5485 4935
rect 5515 4915 5535 4935
rect 5565 4915 5585 4935
rect 5615 4915 5635 4935
rect 5715 4915 5735 4935
rect 5765 4915 5785 4935
rect 5815 4915 5835 4935
rect 5865 4915 5885 4935
rect 5915 4915 5935 4935
rect 6015 4915 6035 4935
rect 6065 4915 6085 4935
rect 6115 4915 6135 4935
rect 6165 4915 6185 4935
rect 6215 4915 6235 4935
rect 6315 4915 6335 4935
rect 6365 4915 6385 4935
rect 6415 4915 6435 4935
rect 6465 4915 6485 4935
rect 6515 4915 6535 4935
rect 6615 4915 6635 4935
rect 6665 4915 6685 4935
rect 6715 4915 6735 4935
rect 6765 4915 6785 4935
rect 6815 4915 6835 4935
rect 6915 4915 6935 4935
rect 6965 4915 6985 4935
rect 7015 4915 7035 4935
rect 7065 4915 7085 4935
rect 7115 4915 7135 4935
rect 7215 4915 7235 4935
rect 7265 4915 7285 4935
rect 7315 4915 7335 4935
rect 7365 4915 7385 4935
rect 7415 4915 7435 4935
rect 7515 4915 7535 4935
rect 7565 4915 7585 4935
rect 7615 4915 7635 4935
rect 7665 4915 7685 4935
rect 7715 4915 7735 4935
rect 7815 4915 7835 4935
rect 7865 4915 7885 4935
rect 7915 4915 7935 4935
rect 7965 4915 7985 4935
rect 8015 4915 8035 4935
rect 8115 4915 8135 4935
rect 8165 4915 8185 4935
rect 8215 4915 8235 4935
rect 8265 4915 8285 4935
rect 8315 4915 8335 4935
rect 8415 4915 8435 4935
rect 8465 4915 8485 4935
rect 8515 4915 8535 4935
rect 8565 4915 8585 4935
rect 8615 4915 8635 4935
rect 8715 4915 8735 4935
rect 8765 4915 8785 4935
rect 8815 4915 8835 4935
rect 8865 4915 8885 4935
rect 8915 4915 8935 4935
rect 9015 4915 9035 4935
rect 9065 4915 9085 4935
rect 9115 4915 9135 4935
rect 9165 4915 9185 4935
rect 9215 4915 9235 4935
rect 9315 4915 9335 4935
rect 9365 4915 9385 4935
rect 9415 4915 9435 4935
rect 9465 4915 9485 4935
rect 9515 4915 9535 4935
rect 9615 4915 9635 4935
rect 9665 4915 9685 4935
rect 9715 4915 9735 4935
rect 9765 4915 9785 4935
rect 9815 4915 9835 4935
rect 9915 4915 9935 4935
rect 9965 4915 9985 4935
rect 10015 4915 10035 4935
rect 10065 4915 10085 4935
rect 10115 4915 10135 4935
rect 10215 4915 10235 4935
rect 10265 4915 10285 4935
rect 10315 4915 10335 4935
rect 10365 4915 10385 4935
rect 10415 4915 10435 4935
rect 10515 4915 10535 4935
rect 10565 4915 10585 4935
rect 10615 4915 10635 4935
rect 10665 4915 10685 4935
rect 10715 4915 10735 4935
rect 10815 4915 10835 4935
rect 10865 4915 10885 4935
rect 10915 4915 10935 4935
rect 10965 4915 10985 4935
rect 11015 4915 11035 4935
rect 11115 4915 11135 4935
rect 11165 4915 11185 4935
rect 11215 4915 11235 4935
rect 11265 4915 11285 4935
rect 11315 4915 11335 4935
rect 11415 4915 11435 4935
rect 11465 4915 11485 4935
rect 11515 4915 11535 4935
rect 11565 4915 11585 4935
rect 11615 4915 11635 4935
rect 11715 4915 11735 4935
rect 11765 4915 11785 4935
rect 11815 4915 11835 4935
rect 11865 4915 11885 4935
rect 11915 4915 11935 4935
rect 12015 4915 12035 4935
rect 12065 4915 12085 4935
rect 12115 4915 12135 4935
rect 12165 4915 12185 4935
rect 12215 4915 12235 4935
rect 12315 4915 12335 4935
rect 12365 4915 12385 4935
rect 12415 4915 12435 4935
rect 12465 4915 12485 4935
rect 12515 4915 12535 4935
rect 12615 4915 12635 4935
rect 12665 4915 12685 4935
rect 12715 4915 12735 4935
rect 12765 4915 12785 4935
rect 12815 4915 12835 4935
rect 12915 4915 12935 4935
rect 12965 4915 12985 4935
rect 13015 4915 13035 4935
rect 13065 4915 13085 4935
rect 13115 4915 13135 4935
rect 13215 4915 13235 4935
rect 13265 4915 13285 4935
rect 13315 4915 13335 4935
rect 13365 4915 13385 4935
rect 13415 4915 13435 4935
rect 13515 4915 13535 4935
rect 13565 4915 13585 4935
rect 13615 4915 13635 4935
rect 13665 4915 13685 4935
rect 13715 4915 13735 4935
rect 13815 4915 13835 4935
rect 13865 4915 13885 4935
rect 13915 4915 13935 4935
rect 13965 4915 13985 4935
rect 14015 4915 14035 4935
rect 14115 4915 14135 4935
rect 14165 4915 14185 4935
rect 14215 4915 14235 4935
rect 14265 4915 14285 4935
rect 14315 4915 14335 4935
rect 14415 4915 14435 4935
rect 14465 4915 14485 4935
rect 14515 4915 14535 4935
rect 14565 4915 14585 4935
rect 14615 4915 14635 4935
rect 14715 4915 14735 4935
rect 14765 4915 14785 4935
rect 14815 4915 14835 4935
rect 14865 4915 14885 4935
rect 14915 4915 14935 4935
rect 15015 4915 15035 4935
rect 15065 4915 15085 4935
rect 15115 4915 15135 4935
rect 15165 4915 15185 4935
rect 15215 4915 15235 4935
rect 15315 4915 15335 4935
rect 15365 4915 15385 4935
rect 15415 4915 15435 4935
rect 15465 4915 15485 4935
rect 15515 4915 15535 4935
rect 15615 4915 15635 4935
rect 15665 4915 15685 4935
rect 15715 4915 15735 4935
rect 15765 4915 15785 4935
rect 15815 4915 15835 4935
rect 15915 4915 15935 4935
rect 15965 4915 15985 4935
rect 16015 4915 16035 4935
rect 16065 4915 16085 4935
rect 16115 4915 16135 4935
rect 16215 4915 16235 4935
rect 16265 4915 16285 4935
rect 16315 4915 16335 4935
rect 16365 4915 16385 4935
rect 16415 4915 16435 4935
rect 16515 4915 16535 4935
rect 16565 4915 16585 4935
rect 16615 4915 16635 4935
rect 16665 4915 16685 4935
rect 16715 4915 16735 4935
rect 16815 4915 16835 4935
rect 16865 4915 16885 4935
rect 16915 4915 16935 4935
rect 16965 4915 16985 4935
rect 17015 4915 17035 4935
rect 17115 4915 17135 4935
rect 17165 4915 17185 4935
rect 17215 4915 17235 4935
rect 17265 4915 17285 4935
rect 17315 4915 17335 4935
rect 17415 4915 17435 4935
rect 17465 4915 17485 4935
rect 17515 4915 17535 4935
rect 17565 4915 17585 4935
rect 17615 4915 17635 4935
rect 17715 4915 17735 4935
rect 17765 4915 17785 4935
rect 17815 4915 17835 4935
rect 17865 4915 17885 4935
rect 17915 4915 17935 4935
rect 18015 4915 18035 4935
rect 18065 4915 18085 4935
rect 18115 4915 18135 4935
rect 18165 4915 18185 4935
rect 18215 4915 18235 4935
rect 18315 4915 18335 4935
rect 18365 4915 18385 4935
rect 18415 4915 18435 4935
rect 18465 4915 18485 4935
rect 18515 4915 18535 4935
rect 18615 4915 18635 4935
rect 18665 4915 18685 4935
rect 18715 4915 18735 4935
rect 18765 4915 18785 4935
rect 18815 4915 18835 4935
rect 18915 4915 18935 4935
rect 18965 4915 18985 4935
rect 19015 4915 19035 4935
rect 19065 4915 19085 4935
rect 19115 4915 19135 4935
rect 19215 4915 19235 4935
rect 19265 4915 19285 4935
rect 19315 4915 19335 4935
rect 19365 4915 19385 4935
rect 19415 4915 19435 4935
rect 19515 4915 19535 4935
rect 19565 4915 19585 4935
rect 19615 4915 19635 4935
rect 19665 4915 19685 4935
rect 19715 4915 19735 4935
rect 19815 4915 19835 4935
rect 19865 4915 19885 4935
rect 19915 4915 19935 4935
rect 19965 4915 19985 4935
rect 20015 4915 20035 4935
rect 20115 4915 20135 4935
rect 20165 4915 20185 4935
rect 20215 4915 20235 4935
rect 20265 4915 20285 4935
rect 20315 4915 20335 4935
rect 20415 4915 20435 4935
rect 20465 4915 20485 4935
rect 20515 4915 20535 4935
rect 20565 4915 20585 4935
rect 20615 4915 20635 4935
rect 20715 4915 20735 4935
rect 20765 4915 20785 4935
rect 20815 4915 20835 4935
rect 20865 4915 20885 4935
rect 20915 4915 20935 4935
rect 21015 4915 21035 4935
rect 21065 4915 21085 4935
rect 21115 4915 21135 4935
rect 21165 4915 21185 4935
rect 21215 4915 21235 4935
rect 21265 4915 21285 4935
rect 21315 4915 21335 4935
rect 21365 4915 21385 4935
rect 21465 4915 21485 4935
rect 21515 4915 21535 4935
rect 21565 4915 21585 4935
rect 21615 4915 21635 4935
rect 21665 4915 21685 4935
rect 21715 4915 21735 4935
rect 21765 4915 21785 4935
rect 21815 4915 21835 4935
rect 21915 4915 21935 4935
rect 21965 4915 21985 4935
rect 22015 4915 22035 4935
rect 22065 4915 22085 4935
rect 22115 4915 22135 4935
rect 22215 4915 22235 4935
rect 22265 4915 22285 4935
rect 22315 4915 22335 4935
rect 22365 4915 22385 4935
rect 22415 4915 22435 4935
rect 22515 4915 22535 4935
rect 22565 4915 22585 4935
rect 22615 4915 22635 4935
rect 22665 4915 22685 4935
rect 22715 4915 22735 4935
rect 22815 4915 22835 4935
rect 22865 4915 22885 4935
rect 22915 4915 22935 4935
rect 22965 4915 22985 4935
rect 23015 4915 23035 4935
rect 23115 4915 23135 4935
rect 23165 4915 23185 4935
rect 23215 4915 23235 4935
rect 23265 4915 23285 4935
rect 23315 4915 23335 4935
rect 23365 4915 23385 4935
rect 23415 4915 23435 4935
rect 23465 4915 23485 4935
rect 23565 4915 23585 4935
rect 23615 4915 23635 4935
rect 23665 4915 23685 4935
rect 23715 4915 23735 4935
rect 23765 4915 23785 4935
rect 23815 4915 23835 4935
rect 23865 4915 23885 4935
rect 23915 4915 23935 4935
rect 24015 4915 24035 4935
rect 24065 4915 24085 4935
rect 24115 4915 24135 4935
rect 24165 4915 24185 4935
rect 24215 4915 24235 4935
rect 24315 4915 24335 4935
rect 24365 4915 24385 4935
rect 24415 4915 24435 4935
rect 24465 4915 24485 4935
rect 24515 4915 24535 4935
rect 24615 4915 24635 4935
rect 24665 4915 24685 4935
rect 24715 4915 24735 4935
rect 24765 4915 24785 4935
rect 24815 4915 24835 4935
rect 24915 4915 24935 4935
rect 24965 4915 24985 4935
rect 25015 4915 25035 4935
rect 25065 4915 25085 4935
rect 25115 4915 25135 4935
rect 25215 4915 25235 4935
rect 25265 4915 25285 4935
rect 25315 4915 25335 4935
rect 25365 4915 25385 4935
rect 25415 4915 25435 4935
rect 25465 4915 25485 4935
rect 25515 4915 25535 4935
rect 25565 4915 25585 4935
rect 25665 4915 25685 4935
rect 25715 4915 25735 4935
rect 25765 4915 25785 4935
rect 25815 4915 25835 4935
rect 25865 4915 25885 4935
rect 25915 4915 25935 4935
rect 25965 4915 25985 4935
rect 26015 4915 26035 4935
rect 26115 4915 26135 4935
rect 26165 4915 26185 4935
rect 26215 4915 26235 4935
rect 26265 4915 26285 4935
rect 26315 4915 26335 4935
rect 26415 4915 26435 4935
rect 26465 4915 26485 4935
rect 26515 4915 26535 4935
rect 26565 4915 26585 4935
rect 26615 4915 26635 4935
rect 26715 4915 26735 4935
rect 26765 4915 26785 4935
rect 26815 4915 26835 4935
rect 26865 4915 26885 4935
rect 26915 4915 26935 4935
rect 27015 4915 27035 4935
rect 27065 4915 27085 4935
rect 27115 4915 27135 4935
rect 27165 4915 27185 4935
rect 27215 4915 27235 4935
rect 27315 4915 27335 4935
rect 27365 4915 27385 4935
rect 27415 4915 27435 4935
rect 27465 4915 27485 4935
rect 27515 4915 27535 4935
rect 27565 4915 27585 4935
rect 27615 4915 27635 4935
rect 27665 4915 27685 4935
rect 27765 4915 27785 4935
rect 27815 4915 27835 4935
rect 27865 4915 27885 4935
rect 27915 4915 27935 4935
rect 27965 4915 27985 4935
rect 28015 4915 28035 4935
rect 28065 4915 28085 4935
rect 28115 4915 28135 4935
rect 28215 4915 28235 4935
rect 28265 4915 28285 4935
rect 28315 4915 28335 4935
rect 28365 4915 28385 4935
rect 28415 4915 28435 4935
rect 28515 4915 28535 4935
rect 28565 4915 28585 4935
rect 28615 4915 28635 4935
rect 28665 4915 28685 4935
rect 28715 4915 28735 4935
rect 28815 4915 28835 4935
rect 28865 4915 28885 4935
rect 28915 4915 28935 4935
rect 28965 4915 28985 4935
rect 29015 4915 29035 4935
rect 29115 4915 29135 4935
rect 29165 4915 29185 4935
rect 29215 4915 29235 4935
rect 29265 4915 29285 4935
rect 29315 4915 29335 4935
rect 29415 4915 29435 4935
rect 29465 4915 29485 4935
rect 29515 4915 29535 4935
rect 29565 4915 29585 4935
rect 29615 4915 29635 4935
rect 29665 4915 29685 4935
rect 29715 4915 29735 4935
rect 29765 4915 29785 4935
rect 29865 4915 29885 4935
rect 29915 4915 29935 4935
rect 29965 4915 29985 4935
rect 30015 4915 30035 4935
rect 30065 4915 30085 4935
rect 30165 4915 30185 4935
rect 30215 4915 30235 4935
rect 30265 4915 30285 4935
rect 30315 4915 30335 4935
rect 30365 4915 30385 4935
rect 30465 4915 30485 4935
rect 30515 4915 30535 4935
rect 30565 4915 30585 4935
rect 30615 4915 30635 4935
rect 30665 4915 30685 4935
rect 30765 4915 30785 4935
rect 30815 4915 30835 4935
rect 30865 4915 30885 4935
rect 30915 4915 30935 4935
rect 30965 4915 30985 4935
rect 31065 4915 31085 4935
rect 31115 4915 31135 4935
rect 31165 4915 31185 4935
rect 31215 4915 31235 4935
rect 31265 4915 31285 4935
rect 31315 4915 31335 4935
rect 31365 4915 31385 4935
rect 31415 4915 31435 4935
rect 31515 4915 31535 4935
rect 31565 4915 31585 4935
rect 31615 4915 31635 4935
rect 31665 4915 31685 4935
rect 31715 4915 31735 4935
rect 31815 4915 31835 4935
rect 31865 4915 31885 4935
rect 31915 4915 31935 4935
rect 31965 4915 31985 4935
rect 32015 4915 32035 4935
rect -585 3615 -565 3635
rect -535 3615 -515 3635
rect -485 3615 -465 3635
rect -435 3615 -415 3635
rect -385 3615 -365 3635
rect -285 3615 -265 3635
rect -235 3615 -215 3635
rect -185 3615 -165 3635
rect -135 3615 -115 3635
rect -85 3615 -65 3635
rect 15 3615 35 3635
rect 65 3615 85 3635
rect 115 3615 135 3635
rect 165 3615 185 3635
rect 215 3615 235 3635
rect 315 3615 335 3635
rect 365 3615 385 3635
rect 415 3615 435 3635
rect 465 3615 485 3635
rect 515 3615 535 3635
rect 615 3615 635 3635
rect 665 3615 685 3635
rect 715 3615 735 3635
rect 765 3615 785 3635
rect 815 3615 835 3635
rect 915 3615 935 3635
rect 965 3615 985 3635
rect 1015 3615 1035 3635
rect 1065 3615 1085 3635
rect 1115 3615 1135 3635
rect 1215 3615 1235 3635
rect 1265 3615 1285 3635
rect 1315 3615 1335 3635
rect 1365 3615 1385 3635
rect 1415 3615 1435 3635
rect 1515 3615 1535 3635
rect 1565 3615 1585 3635
rect 1615 3615 1635 3635
rect 1665 3615 1685 3635
rect 1715 3615 1735 3635
rect 1815 3615 1835 3635
rect 1865 3615 1885 3635
rect 1915 3615 1935 3635
rect 1965 3615 1985 3635
rect 2015 3615 2035 3635
rect 2115 3615 2135 3635
rect 2165 3615 2185 3635
rect 2215 3615 2235 3635
rect 2265 3615 2285 3635
rect 2315 3615 2335 3635
rect 2415 3615 2435 3635
rect 2465 3615 2485 3635
rect 2515 3615 2535 3635
rect 2565 3615 2585 3635
rect 2615 3615 2635 3635
rect 2715 3615 2735 3635
rect 2765 3615 2785 3635
rect 2815 3615 2835 3635
rect 2865 3615 2885 3635
rect 2915 3615 2935 3635
rect 3015 3615 3035 3635
rect 3065 3615 3085 3635
rect 3115 3615 3135 3635
rect 3165 3615 3185 3635
rect 3215 3615 3235 3635
rect 3315 3615 3335 3635
rect 3365 3615 3385 3635
rect 3415 3615 3435 3635
rect 3465 3615 3485 3635
rect 3515 3615 3535 3635
rect 3615 3615 3635 3635
rect 3665 3615 3685 3635
rect 3715 3615 3735 3635
rect 3765 3615 3785 3635
rect 3815 3615 3835 3635
rect 3915 3615 3935 3635
rect 3965 3615 3985 3635
rect 4015 3615 4035 3635
rect 4065 3615 4085 3635
rect 4115 3615 4135 3635
rect 4215 3615 4235 3635
rect 4265 3615 4285 3635
rect 4315 3615 4335 3635
rect 4365 3615 4385 3635
rect 4415 3615 4435 3635
rect 4515 3615 4535 3635
rect 4565 3615 4585 3635
rect 4615 3615 4635 3635
rect 4665 3615 4685 3635
rect 4715 3615 4735 3635
rect 4815 3615 4835 3635
rect 4865 3615 4885 3635
rect 4915 3615 4935 3635
rect 4965 3615 4985 3635
rect 5015 3615 5035 3635
rect 5115 3615 5135 3635
rect 5165 3615 5185 3635
rect 5215 3615 5235 3635
rect 5265 3615 5285 3635
rect 5315 3615 5335 3635
rect 5415 3615 5435 3635
rect 5465 3615 5485 3635
rect 5515 3615 5535 3635
rect 5565 3615 5585 3635
rect 5615 3615 5635 3635
rect 5715 3615 5735 3635
rect 5765 3615 5785 3635
rect 5815 3615 5835 3635
rect 5865 3615 5885 3635
rect 5915 3615 5935 3635
rect 6015 3615 6035 3635
rect 6065 3615 6085 3635
rect 6115 3615 6135 3635
rect 6165 3615 6185 3635
rect 6215 3615 6235 3635
rect 6315 3615 6335 3635
rect 6365 3615 6385 3635
rect 6415 3615 6435 3635
rect 6465 3615 6485 3635
rect 6515 3615 6535 3635
rect 6615 3615 6635 3635
rect 6665 3615 6685 3635
rect 6715 3615 6735 3635
rect 6765 3615 6785 3635
rect 6815 3615 6835 3635
rect 6915 3615 6935 3635
rect 6965 3615 6985 3635
rect 7015 3615 7035 3635
rect 7065 3615 7085 3635
rect 7115 3615 7135 3635
rect 7215 3615 7235 3635
rect 7265 3615 7285 3635
rect 7315 3615 7335 3635
rect 7365 3615 7385 3635
rect 7415 3615 7435 3635
rect 7515 3615 7535 3635
rect 7565 3615 7585 3635
rect 7615 3615 7635 3635
rect 7665 3615 7685 3635
rect 7715 3615 7735 3635
rect 7815 3615 7835 3635
rect 7865 3615 7885 3635
rect 7915 3615 7935 3635
rect 7965 3615 7985 3635
rect 8015 3615 8035 3635
rect 8115 3615 8135 3635
rect 8165 3615 8185 3635
rect 8215 3615 8235 3635
rect 8265 3615 8285 3635
rect 8315 3615 8335 3635
rect 8415 3615 8435 3635
rect 8465 3615 8485 3635
rect 8515 3615 8535 3635
rect 8565 3615 8585 3635
rect 8615 3615 8635 3635
rect 8715 3615 8735 3635
rect 8765 3615 8785 3635
rect 8815 3615 8835 3635
rect 8865 3615 8885 3635
rect 8915 3615 8935 3635
rect 9015 3615 9035 3635
rect 9065 3615 9085 3635
rect 9115 3615 9135 3635
rect 9165 3615 9185 3635
rect 9215 3615 9235 3635
rect 9315 3615 9335 3635
rect 9365 3615 9385 3635
rect 9415 3615 9435 3635
rect 9465 3615 9485 3635
rect 9515 3615 9535 3635
rect 9615 3615 9635 3635
rect 9665 3615 9685 3635
rect 9715 3615 9735 3635
rect 9765 3615 9785 3635
rect 9815 3615 9835 3635
rect 9915 3615 9935 3635
rect 9965 3615 9985 3635
rect 10015 3615 10035 3635
rect 10065 3615 10085 3635
rect 10115 3615 10135 3635
rect 10215 3615 10235 3635
rect 10265 3615 10285 3635
rect 10315 3615 10335 3635
rect 10365 3615 10385 3635
rect 10415 3615 10435 3635
rect 10515 3615 10535 3635
rect 10565 3615 10585 3635
rect 10615 3615 10635 3635
rect 10665 3615 10685 3635
rect 10715 3615 10735 3635
rect 10815 3615 10835 3635
rect 10865 3615 10885 3635
rect 10915 3615 10935 3635
rect 10965 3615 10985 3635
rect 11015 3615 11035 3635
rect 11115 3615 11135 3635
rect 11165 3615 11185 3635
rect 11215 3615 11235 3635
rect 11265 3615 11285 3635
rect 11315 3615 11335 3635
rect 11415 3615 11435 3635
rect 11465 3615 11485 3635
rect 11515 3615 11535 3635
rect 11565 3615 11585 3635
rect 11615 3615 11635 3635
rect 11715 3615 11735 3635
rect 11765 3615 11785 3635
rect 11815 3615 11835 3635
rect 11865 3615 11885 3635
rect 11915 3615 11935 3635
rect 12015 3615 12035 3635
rect 12065 3615 12085 3635
rect 12115 3615 12135 3635
rect 12165 3615 12185 3635
rect 12215 3615 12235 3635
rect 12315 3615 12335 3635
rect 12365 3615 12385 3635
rect 12415 3615 12435 3635
rect 12465 3615 12485 3635
rect 12515 3615 12535 3635
rect 12615 3615 12635 3635
rect 12665 3615 12685 3635
rect 12715 3615 12735 3635
rect 12765 3615 12785 3635
rect 12815 3615 12835 3635
rect 12915 3615 12935 3635
rect 12965 3615 12985 3635
rect 13015 3615 13035 3635
rect 13065 3615 13085 3635
rect 13115 3615 13135 3635
rect 13215 3615 13235 3635
rect 13265 3615 13285 3635
rect 13315 3615 13335 3635
rect 13365 3615 13385 3635
rect 13415 3615 13435 3635
rect 13515 3615 13535 3635
rect 13565 3615 13585 3635
rect 13615 3615 13635 3635
rect 13665 3615 13685 3635
rect 13715 3615 13735 3635
rect 13815 3615 13835 3635
rect 13865 3615 13885 3635
rect 13915 3615 13935 3635
rect 13965 3615 13985 3635
rect 14015 3615 14035 3635
rect 14115 3615 14135 3635
rect 14165 3615 14185 3635
rect 14215 3615 14235 3635
rect 14265 3615 14285 3635
rect 14315 3615 14335 3635
rect 14415 3615 14435 3635
rect 14465 3615 14485 3635
rect 14515 3615 14535 3635
rect 14565 3615 14585 3635
rect 14615 3615 14635 3635
rect 14715 3615 14735 3635
rect 14765 3615 14785 3635
rect 14815 3615 14835 3635
rect 14865 3615 14885 3635
rect 14915 3615 14935 3635
rect 15015 3615 15035 3635
rect 15065 3615 15085 3635
rect 15115 3615 15135 3635
rect 15165 3615 15185 3635
rect 15215 3615 15235 3635
rect 15315 3615 15335 3635
rect 15365 3615 15385 3635
rect 15415 3615 15435 3635
rect 15465 3615 15485 3635
rect 15515 3615 15535 3635
rect 15615 3615 15635 3635
rect 15665 3615 15685 3635
rect 15715 3615 15735 3635
rect 15765 3615 15785 3635
rect 15815 3615 15835 3635
rect 15915 3615 15935 3635
rect 15965 3615 15985 3635
rect 16015 3615 16035 3635
rect 16065 3615 16085 3635
rect 16115 3615 16135 3635
rect 16215 3615 16235 3635
rect 16265 3615 16285 3635
rect 16315 3615 16335 3635
rect 16365 3615 16385 3635
rect 16415 3615 16435 3635
rect 16515 3615 16535 3635
rect 16565 3615 16585 3635
rect 16615 3615 16635 3635
rect 16665 3615 16685 3635
rect 16715 3615 16735 3635
rect 16815 3615 16835 3635
rect 16865 3615 16885 3635
rect 16915 3615 16935 3635
rect 16965 3615 16985 3635
rect 17015 3615 17035 3635
rect 17115 3615 17135 3635
rect 17165 3615 17185 3635
rect 17215 3615 17235 3635
rect 17265 3615 17285 3635
rect 17315 3615 17335 3635
rect 17415 3615 17435 3635
rect 17465 3615 17485 3635
rect 17515 3615 17535 3635
rect 17565 3615 17585 3635
rect 17615 3615 17635 3635
rect 17715 3615 17735 3635
rect 17765 3615 17785 3635
rect 17815 3615 17835 3635
rect 17865 3615 17885 3635
rect 17915 3615 17935 3635
rect 18015 3615 18035 3635
rect 18065 3615 18085 3635
rect 18115 3615 18135 3635
rect 18165 3615 18185 3635
rect 18215 3615 18235 3635
rect 18315 3615 18335 3635
rect 18365 3615 18385 3635
rect 18415 3615 18435 3635
rect 18465 3615 18485 3635
rect 18515 3615 18535 3635
rect 18615 3615 18635 3635
rect 18665 3615 18685 3635
rect 18715 3615 18735 3635
rect 18765 3615 18785 3635
rect 18815 3615 18835 3635
rect 18915 3615 18935 3635
rect 18965 3615 18985 3635
rect 19015 3615 19035 3635
rect 19065 3615 19085 3635
rect 19115 3615 19135 3635
rect 19215 3615 19235 3635
rect 19265 3615 19285 3635
rect 19315 3615 19335 3635
rect 19365 3615 19385 3635
rect 19415 3615 19435 3635
rect 19515 3615 19535 3635
rect 19565 3615 19585 3635
rect 19615 3615 19635 3635
rect 19665 3615 19685 3635
rect 19715 3615 19735 3635
rect 19815 3615 19835 3635
rect 19865 3615 19885 3635
rect 19915 3615 19935 3635
rect 19965 3615 19985 3635
rect 20015 3615 20035 3635
rect 20115 3615 20135 3635
rect 20165 3615 20185 3635
rect 20215 3615 20235 3635
rect 20265 3615 20285 3635
rect 20315 3615 20335 3635
rect 20415 3615 20435 3635
rect 20465 3615 20485 3635
rect 20515 3615 20535 3635
rect 20565 3615 20585 3635
rect 20615 3615 20635 3635
rect 20715 3615 20735 3635
rect 20765 3615 20785 3635
rect 20815 3615 20835 3635
rect 20865 3615 20885 3635
rect 20915 3615 20935 3635
rect 21015 3615 21035 3635
rect 21065 3615 21085 3635
rect 21115 3615 21135 3635
rect 21165 3615 21185 3635
rect 21215 3615 21235 3635
rect 21265 3615 21285 3635
rect 21315 3615 21335 3635
rect 21365 3615 21385 3635
rect 21465 3615 21485 3635
rect 21515 3615 21535 3635
rect 21565 3615 21585 3635
rect 21615 3615 21635 3635
rect 21665 3615 21685 3635
rect 21715 3615 21735 3635
rect 21765 3615 21785 3635
rect 21815 3615 21835 3635
rect 21915 3615 21935 3635
rect 21965 3615 21985 3635
rect 22015 3615 22035 3635
rect 22065 3615 22085 3635
rect 22115 3615 22135 3635
rect 22215 3615 22235 3635
rect 22265 3615 22285 3635
rect 22315 3615 22335 3635
rect 22365 3615 22385 3635
rect 22415 3615 22435 3635
rect 22515 3615 22535 3635
rect 22565 3615 22585 3635
rect 22615 3615 22635 3635
rect 22665 3615 22685 3635
rect 22715 3615 22735 3635
rect 22815 3615 22835 3635
rect 22865 3615 22885 3635
rect 22915 3615 22935 3635
rect 22965 3615 22985 3635
rect 23015 3615 23035 3635
rect 23115 3615 23135 3635
rect 23165 3615 23185 3635
rect 23215 3615 23235 3635
rect 23265 3615 23285 3635
rect 23315 3615 23335 3635
rect 23365 3615 23385 3635
rect 23415 3615 23435 3635
rect 23465 3615 23485 3635
rect 23565 3615 23585 3635
rect 23615 3615 23635 3635
rect 23665 3615 23685 3635
rect 23715 3615 23735 3635
rect 23765 3615 23785 3635
rect 23815 3615 23835 3635
rect 23865 3615 23885 3635
rect 23915 3615 23935 3635
rect 24015 3615 24035 3635
rect 24065 3615 24085 3635
rect 24115 3615 24135 3635
rect 24165 3615 24185 3635
rect 24215 3615 24235 3635
rect 24315 3615 24335 3635
rect 24365 3615 24385 3635
rect 24415 3615 24435 3635
rect 24465 3615 24485 3635
rect 24515 3615 24535 3635
rect 24615 3615 24635 3635
rect 24665 3615 24685 3635
rect 24715 3615 24735 3635
rect 24765 3615 24785 3635
rect 24815 3615 24835 3635
rect 24915 3615 24935 3635
rect 24965 3615 24985 3635
rect 25015 3615 25035 3635
rect 25065 3615 25085 3635
rect 25115 3615 25135 3635
rect 25215 3615 25235 3635
rect 25265 3615 25285 3635
rect 25315 3615 25335 3635
rect 25365 3615 25385 3635
rect 25415 3615 25435 3635
rect 25465 3615 25485 3635
rect 25515 3615 25535 3635
rect 25565 3615 25585 3635
rect 25665 3615 25685 3635
rect 25715 3615 25735 3635
rect 25765 3615 25785 3635
rect 25815 3615 25835 3635
rect 25865 3615 25885 3635
rect 25915 3615 25935 3635
rect 25965 3615 25985 3635
rect 26015 3615 26035 3635
rect 26115 3615 26135 3635
rect 26165 3615 26185 3635
rect 26215 3615 26235 3635
rect 26265 3615 26285 3635
rect 26315 3615 26335 3635
rect 26415 3615 26435 3635
rect 26465 3615 26485 3635
rect 26515 3615 26535 3635
rect 26565 3615 26585 3635
rect 26615 3615 26635 3635
rect 26715 3615 26735 3635
rect 26765 3615 26785 3635
rect 26815 3615 26835 3635
rect 26865 3615 26885 3635
rect 26915 3615 26935 3635
rect 27015 3615 27035 3635
rect 27065 3615 27085 3635
rect 27115 3615 27135 3635
rect 27165 3615 27185 3635
rect 27215 3615 27235 3635
rect 27315 3615 27335 3635
rect 27365 3615 27385 3635
rect 27415 3615 27435 3635
rect 27465 3615 27485 3635
rect 27515 3615 27535 3635
rect 27565 3615 27585 3635
rect 27615 3615 27635 3635
rect 27665 3615 27685 3635
rect 27765 3615 27785 3635
rect 27815 3615 27835 3635
rect 27865 3615 27885 3635
rect 27915 3615 27935 3635
rect 27965 3615 27985 3635
rect 28015 3615 28035 3635
rect 28065 3615 28085 3635
rect 28115 3615 28135 3635
rect 28215 3615 28235 3635
rect 28265 3615 28285 3635
rect 28315 3615 28335 3635
rect 28365 3615 28385 3635
rect 28415 3615 28435 3635
rect 28515 3615 28535 3635
rect 28565 3615 28585 3635
rect 28615 3615 28635 3635
rect 28665 3615 28685 3635
rect 28715 3615 28735 3635
rect 28815 3615 28835 3635
rect 28865 3615 28885 3635
rect 28915 3615 28935 3635
rect 28965 3615 28985 3635
rect 29015 3615 29035 3635
rect 29115 3615 29135 3635
rect 29165 3615 29185 3635
rect 29215 3615 29235 3635
rect 29265 3615 29285 3635
rect 29315 3615 29335 3635
rect 29415 3615 29435 3635
rect 29465 3615 29485 3635
rect 29515 3615 29535 3635
rect 29565 3615 29585 3635
rect 29615 3615 29635 3635
rect 29665 3615 29685 3635
rect 29715 3615 29735 3635
rect 29765 3615 29785 3635
rect 29865 3615 29885 3635
rect 29915 3615 29935 3635
rect 29965 3615 29985 3635
rect 30015 3615 30035 3635
rect 30065 3615 30085 3635
rect 30165 3615 30185 3635
rect 30215 3615 30235 3635
rect 30265 3615 30285 3635
rect 30315 3615 30335 3635
rect 30365 3615 30385 3635
rect 30465 3615 30485 3635
rect 30515 3615 30535 3635
rect 30565 3615 30585 3635
rect 30615 3615 30635 3635
rect 30665 3615 30685 3635
rect 30765 3615 30785 3635
rect 30815 3615 30835 3635
rect 30865 3615 30885 3635
rect 30915 3615 30935 3635
rect 30965 3615 30985 3635
rect 31065 3615 31085 3635
rect 31115 3615 31135 3635
rect 31165 3615 31185 3635
rect 31215 3615 31235 3635
rect 31265 3615 31285 3635
rect 31315 3615 31335 3635
rect 31365 3615 31385 3635
rect 31415 3615 31435 3635
rect 31515 3615 31535 3635
rect 31565 3615 31585 3635
rect 31615 3615 31635 3635
rect 31665 3615 31685 3635
rect 31715 3615 31735 3635
rect 31815 3615 31835 3635
rect 31865 3615 31885 3635
rect 31915 3615 31935 3635
rect 31965 3615 31985 3635
rect 32015 3615 32035 3635
rect -585 815 -565 835
rect -535 815 -515 835
rect -485 815 -465 835
rect -435 815 -415 835
rect -385 815 -365 835
rect -285 815 -265 835
rect -235 815 -215 835
rect -185 815 -165 835
rect -135 815 -115 835
rect -85 815 -65 835
rect 15 815 35 835
rect 65 815 85 835
rect 115 815 135 835
rect 165 815 185 835
rect 215 815 235 835
rect 315 815 335 835
rect 365 815 385 835
rect 415 815 435 835
rect 465 815 485 835
rect 515 815 535 835
rect 615 815 635 835
rect 665 815 685 835
rect 715 815 735 835
rect 765 815 785 835
rect 815 815 835 835
rect 915 815 935 835
rect 965 815 985 835
rect 1015 815 1035 835
rect 1065 815 1085 835
rect 1115 815 1135 835
rect 1215 815 1235 835
rect 1265 815 1285 835
rect 1315 815 1335 835
rect 1365 815 1385 835
rect 1415 815 1435 835
rect 1515 815 1535 835
rect 1565 815 1585 835
rect 1615 815 1635 835
rect 1665 815 1685 835
rect 1715 815 1735 835
rect 1815 815 1835 835
rect 1865 815 1885 835
rect 1915 815 1935 835
rect 1965 815 1985 835
rect 2015 815 2035 835
rect 2115 815 2135 835
rect 2165 815 2185 835
rect 2215 815 2235 835
rect 2265 815 2285 835
rect 2315 815 2335 835
rect 2415 815 2435 835
rect 2465 815 2485 835
rect 2515 815 2535 835
rect 2565 815 2585 835
rect 2615 815 2635 835
rect 2715 815 2735 835
rect 2765 815 2785 835
rect 2815 815 2835 835
rect 2865 815 2885 835
rect 2915 815 2935 835
rect 3015 815 3035 835
rect 3065 815 3085 835
rect 3115 815 3135 835
rect 3165 815 3185 835
rect 3215 815 3235 835
rect 3315 815 3335 835
rect 3365 815 3385 835
rect 3415 815 3435 835
rect 3465 815 3485 835
rect 3515 815 3535 835
rect 3615 815 3635 835
rect 3665 815 3685 835
rect 3715 815 3735 835
rect 3765 815 3785 835
rect 3815 815 3835 835
rect 3915 815 3935 835
rect 3965 815 3985 835
rect 4015 815 4035 835
rect 4065 815 4085 835
rect 4115 815 4135 835
rect 4215 815 4235 835
rect 4265 815 4285 835
rect 4315 815 4335 835
rect 4365 815 4385 835
rect 4415 815 4435 835
rect 4515 815 4535 835
rect 4565 815 4585 835
rect 4615 815 4635 835
rect 4665 815 4685 835
rect 4715 815 4735 835
rect 4815 815 4835 835
rect 4865 815 4885 835
rect 4915 815 4935 835
rect 4965 815 4985 835
rect 5015 815 5035 835
rect 5115 815 5135 835
rect 5165 815 5185 835
rect 5215 815 5235 835
rect 5265 815 5285 835
rect 5315 815 5335 835
rect 5415 815 5435 835
rect 5465 815 5485 835
rect 5515 815 5535 835
rect 5565 815 5585 835
rect 5615 815 5635 835
rect 5715 815 5735 835
rect 5765 815 5785 835
rect 5815 815 5835 835
rect 5865 815 5885 835
rect 5915 815 5935 835
rect 6015 815 6035 835
rect 6065 815 6085 835
rect 6115 815 6135 835
rect 6165 815 6185 835
rect 6215 815 6235 835
rect 6315 815 6335 835
rect 6365 815 6385 835
rect 6415 815 6435 835
rect 6465 815 6485 835
rect 6515 815 6535 835
rect 6615 815 6635 835
rect 6665 815 6685 835
rect 6715 815 6735 835
rect 6765 815 6785 835
rect 6815 815 6835 835
rect 6915 815 6935 835
rect 6965 815 6985 835
rect 7015 815 7035 835
rect 7065 815 7085 835
rect 7115 815 7135 835
rect 7215 815 7235 835
rect 7265 815 7285 835
rect 7315 815 7335 835
rect 7365 815 7385 835
rect 7415 815 7435 835
rect 7515 815 7535 835
rect 7565 815 7585 835
rect 7615 815 7635 835
rect 7665 815 7685 835
rect 7715 815 7735 835
rect 7815 815 7835 835
rect 7865 815 7885 835
rect 7915 815 7935 835
rect 7965 815 7985 835
rect 8015 815 8035 835
rect 8115 815 8135 835
rect 8165 815 8185 835
rect 8215 815 8235 835
rect 8265 815 8285 835
rect 8315 815 8335 835
rect 8415 815 8435 835
rect 8465 815 8485 835
rect 8515 815 8535 835
rect 8565 815 8585 835
rect 8615 815 8635 835
rect 8715 815 8735 835
rect 8765 815 8785 835
rect 8815 815 8835 835
rect 8865 815 8885 835
rect 8915 815 8935 835
rect 9015 815 9035 835
rect 9065 815 9085 835
rect 9115 815 9135 835
rect 9165 815 9185 835
rect 9215 815 9235 835
rect 9315 815 9335 835
rect 9365 815 9385 835
rect 9415 815 9435 835
rect 9465 815 9485 835
rect 9515 815 9535 835
rect 9615 815 9635 835
rect 9665 815 9685 835
rect 9715 815 9735 835
rect 9765 815 9785 835
rect 9815 815 9835 835
rect 9915 815 9935 835
rect 9965 815 9985 835
rect 10015 815 10035 835
rect 10065 815 10085 835
rect 10115 815 10135 835
rect 10215 815 10235 835
rect 10265 815 10285 835
rect 10315 815 10335 835
rect 10365 815 10385 835
rect 10415 815 10435 835
rect 10515 815 10535 835
rect 10565 815 10585 835
rect 10615 815 10635 835
rect 10665 815 10685 835
rect 10715 815 10735 835
rect 10815 815 10835 835
rect 10865 815 10885 835
rect 10915 815 10935 835
rect 10965 815 10985 835
rect 11015 815 11035 835
rect 11115 815 11135 835
rect 11165 815 11185 835
rect 11215 815 11235 835
rect 11265 815 11285 835
rect 11315 815 11335 835
rect 11415 815 11435 835
rect 11465 815 11485 835
rect 11515 815 11535 835
rect 11565 815 11585 835
rect 11615 815 11635 835
rect 11715 815 11735 835
rect 11765 815 11785 835
rect 11815 815 11835 835
rect 11865 815 11885 835
rect 11915 815 11935 835
rect 12015 815 12035 835
rect 12065 815 12085 835
rect 12115 815 12135 835
rect 12165 815 12185 835
rect 12215 815 12235 835
rect 12315 815 12335 835
rect 12365 815 12385 835
rect 12415 815 12435 835
rect 12465 815 12485 835
rect 12515 815 12535 835
rect 12615 815 12635 835
rect 12665 815 12685 835
rect 12715 815 12735 835
rect 12765 815 12785 835
rect 12815 815 12835 835
rect 12915 815 12935 835
rect 12965 815 12985 835
rect 13015 815 13035 835
rect 13065 815 13085 835
rect 13115 815 13135 835
rect 13215 815 13235 835
rect 13265 815 13285 835
rect 13315 815 13335 835
rect 13365 815 13385 835
rect 13415 815 13435 835
rect 13515 815 13535 835
rect 13565 815 13585 835
rect 13615 815 13635 835
rect 13665 815 13685 835
rect 13715 815 13735 835
rect 13815 815 13835 835
rect 13865 815 13885 835
rect 13915 815 13935 835
rect 13965 815 13985 835
rect 14015 815 14035 835
rect 14115 815 14135 835
rect 14165 815 14185 835
rect 14215 815 14235 835
rect 14265 815 14285 835
rect 14315 815 14335 835
rect 14415 815 14435 835
rect 14465 815 14485 835
rect 14515 815 14535 835
rect 14565 815 14585 835
rect 14615 815 14635 835
rect 14715 815 14735 835
rect 14765 815 14785 835
rect 14815 815 14835 835
rect 14865 815 14885 835
rect 14915 815 14935 835
rect 15015 815 15035 835
rect 15065 815 15085 835
rect 15115 815 15135 835
rect 15165 815 15185 835
rect 15215 815 15235 835
rect 15315 815 15335 835
rect 15365 815 15385 835
rect 15415 815 15435 835
rect 15465 815 15485 835
rect 15515 815 15535 835
rect 15615 815 15635 835
rect 15665 815 15685 835
rect 15715 815 15735 835
rect 15765 815 15785 835
rect 15815 815 15835 835
rect 15915 815 15935 835
rect 15965 815 15985 835
rect 16015 815 16035 835
rect 16065 815 16085 835
rect 16115 815 16135 835
rect 16215 815 16235 835
rect 16265 815 16285 835
rect 16315 815 16335 835
rect 16365 815 16385 835
rect 16415 815 16435 835
rect 16515 815 16535 835
rect 16565 815 16585 835
rect 16615 815 16635 835
rect 16665 815 16685 835
rect 16715 815 16735 835
rect 16815 815 16835 835
rect 16865 815 16885 835
rect 16915 815 16935 835
rect 16965 815 16985 835
rect 17015 815 17035 835
rect 17115 815 17135 835
rect 17165 815 17185 835
rect 17215 815 17235 835
rect 17265 815 17285 835
rect 17315 815 17335 835
rect 17415 815 17435 835
rect 17465 815 17485 835
rect 17515 815 17535 835
rect 17565 815 17585 835
rect 17615 815 17635 835
rect 17715 815 17735 835
rect 17765 815 17785 835
rect 17815 815 17835 835
rect 17865 815 17885 835
rect 17915 815 17935 835
rect 18015 815 18035 835
rect 18065 815 18085 835
rect 18115 815 18135 835
rect 18165 815 18185 835
rect 18215 815 18235 835
rect 18315 815 18335 835
rect 18365 815 18385 835
rect 18415 815 18435 835
rect 18465 815 18485 835
rect 18515 815 18535 835
rect 18615 815 18635 835
rect 18665 815 18685 835
rect 18715 815 18735 835
rect 18765 815 18785 835
rect 18815 815 18835 835
rect 18915 815 18935 835
rect 18965 815 18985 835
rect 19015 815 19035 835
rect 19065 815 19085 835
rect 19115 815 19135 835
rect 19215 815 19235 835
rect 19265 815 19285 835
rect 19315 815 19335 835
rect 19365 815 19385 835
rect 19415 815 19435 835
rect 19515 815 19535 835
rect 19565 815 19585 835
rect 19615 815 19635 835
rect 19665 815 19685 835
rect 19715 815 19735 835
rect 19815 815 19835 835
rect 19865 815 19885 835
rect 19915 815 19935 835
rect 19965 815 19985 835
rect 20015 815 20035 835
rect 20115 815 20135 835
rect 20165 815 20185 835
rect 20215 815 20235 835
rect 20265 815 20285 835
rect 20315 815 20335 835
rect 20415 815 20435 835
rect 20465 815 20485 835
rect 20515 815 20535 835
rect 20565 815 20585 835
rect 20615 815 20635 835
rect 20715 815 20735 835
rect 20765 815 20785 835
rect 20815 815 20835 835
rect 20865 815 20885 835
rect 20915 815 20935 835
rect 21015 815 21035 835
rect 21065 815 21085 835
rect 21115 815 21135 835
rect 21165 815 21185 835
rect 21215 815 21235 835
rect 21315 815 21335 835
rect 21365 815 21385 835
rect 21415 815 21435 835
rect 21465 815 21485 835
rect 21515 815 21535 835
rect 21615 815 21635 835
rect 21665 815 21685 835
rect 21715 815 21735 835
rect 21765 815 21785 835
rect 21815 815 21835 835
rect 21915 815 21935 835
rect 21965 815 21985 835
rect 22015 815 22035 835
rect 22065 815 22085 835
rect 22115 815 22135 835
rect 22215 815 22235 835
rect 22265 815 22285 835
rect 22315 815 22335 835
rect 22365 815 22385 835
rect 22415 815 22435 835
rect 22515 815 22535 835
rect 22565 815 22585 835
rect 22615 815 22635 835
rect 22665 815 22685 835
rect 22715 815 22735 835
rect 22815 815 22835 835
rect 22865 815 22885 835
rect 22915 815 22935 835
rect 22965 815 22985 835
rect 23015 815 23035 835
rect 23115 815 23135 835
rect 23165 815 23185 835
rect 23215 815 23235 835
rect 23265 815 23285 835
rect 23315 815 23335 835
rect 23415 815 23435 835
rect 23465 815 23485 835
rect 23515 815 23535 835
rect 23565 815 23585 835
rect 23615 815 23635 835
rect 23715 815 23735 835
rect 23765 815 23785 835
rect 23815 815 23835 835
rect 23865 815 23885 835
rect 23915 815 23935 835
rect 24015 815 24035 835
rect 24065 815 24085 835
rect 24115 815 24135 835
rect 24165 815 24185 835
rect 24215 815 24235 835
rect 24315 815 24335 835
rect 24365 815 24385 835
rect 24415 815 24435 835
rect 24465 815 24485 835
rect 24515 815 24535 835
rect 24615 815 24635 835
rect 24665 815 24685 835
rect 24715 815 24735 835
rect 24765 815 24785 835
rect 24815 815 24835 835
rect 24915 815 24935 835
rect 24965 815 24985 835
rect 25015 815 25035 835
rect 25065 815 25085 835
rect 25115 815 25135 835
rect 25215 815 25235 835
rect 25265 815 25285 835
rect 25315 815 25335 835
rect 25365 815 25385 835
rect 25415 815 25435 835
rect 25515 815 25535 835
rect 25565 815 25585 835
rect 25615 815 25635 835
rect 25665 815 25685 835
rect 25715 815 25735 835
rect 25815 815 25835 835
rect 25865 815 25885 835
rect 25915 815 25935 835
rect 25965 815 25985 835
rect 26015 815 26035 835
rect 26115 815 26135 835
rect 26165 815 26185 835
rect 26215 815 26235 835
rect 26265 815 26285 835
rect 26315 815 26335 835
rect 26415 815 26435 835
rect 26465 815 26485 835
rect 26515 815 26535 835
rect 26565 815 26585 835
rect 26615 815 26635 835
rect 26715 815 26735 835
rect 26765 815 26785 835
rect 26815 815 26835 835
rect 26865 815 26885 835
rect 26915 815 26935 835
rect 27015 815 27035 835
rect 27065 815 27085 835
rect 27115 815 27135 835
rect 27165 815 27185 835
rect 27215 815 27235 835
rect 27315 815 27335 835
rect 27365 815 27385 835
rect 27415 815 27435 835
rect 27465 815 27485 835
rect 27515 815 27535 835
rect 27615 815 27635 835
rect 27665 815 27685 835
rect 27715 815 27735 835
rect 27765 815 27785 835
rect 27815 815 27835 835
rect 27915 815 27935 835
rect 27965 815 27985 835
rect 28015 815 28035 835
rect 28065 815 28085 835
rect 28115 815 28135 835
rect 28215 815 28235 835
rect 28265 815 28285 835
rect 28315 815 28335 835
rect 28365 815 28385 835
rect 28415 815 28435 835
rect 28515 815 28535 835
rect 28565 815 28585 835
rect 28615 815 28635 835
rect 28665 815 28685 835
rect 28715 815 28735 835
rect -585 -885 -565 -865
rect -535 -885 -515 -865
rect -485 -885 -465 -865
rect -435 -885 -415 -865
rect -385 -885 -365 -865
rect -285 -885 -265 -865
rect -235 -885 -215 -865
rect -185 -885 -165 -865
rect -135 -885 -115 -865
rect -85 -885 -65 -865
rect 15 -885 35 -865
rect 65 -885 85 -865
rect 115 -885 135 -865
rect 165 -885 185 -865
rect 215 -885 235 -865
rect 315 -885 335 -865
rect 365 -885 385 -865
rect 415 -885 435 -865
rect 465 -885 485 -865
rect 515 -885 535 -865
rect 615 -885 635 -865
rect 665 -885 685 -865
rect 715 -885 735 -865
rect 765 -885 785 -865
rect 815 -885 835 -865
rect 915 -885 935 -865
rect 965 -885 985 -865
rect 1015 -885 1035 -865
rect 1065 -885 1085 -865
rect 1115 -885 1135 -865
rect 1215 -885 1235 -865
rect 1265 -885 1285 -865
rect 1315 -885 1335 -865
rect 1365 -885 1385 -865
rect 1415 -885 1435 -865
rect 1515 -885 1535 -865
rect 1565 -885 1585 -865
rect 1615 -885 1635 -865
rect 1665 -885 1685 -865
rect 1715 -885 1735 -865
rect 1815 -885 1835 -865
rect 1865 -885 1885 -865
rect 1915 -885 1935 -865
rect 1965 -885 1985 -865
rect 2015 -885 2035 -865
rect 2115 -885 2135 -865
rect 2165 -885 2185 -865
rect 2215 -885 2235 -865
rect 2265 -885 2285 -865
rect 2315 -885 2335 -865
rect 2415 -885 2435 -865
rect 2465 -885 2485 -865
rect 2515 -885 2535 -865
rect 2565 -885 2585 -865
rect 2615 -885 2635 -865
rect 2715 -885 2735 -865
rect 2765 -885 2785 -865
rect 2815 -885 2835 -865
rect 2865 -885 2885 -865
rect 2915 -885 2935 -865
rect 3015 -885 3035 -865
rect 3065 -885 3085 -865
rect 3115 -885 3135 -865
rect 3165 -885 3185 -865
rect 3215 -885 3235 -865
rect 3315 -885 3335 -865
rect 3365 -885 3385 -865
rect 3415 -885 3435 -865
rect 3465 -885 3485 -865
rect 3515 -885 3535 -865
rect 3615 -885 3635 -865
rect 3665 -885 3685 -865
rect 3715 -885 3735 -865
rect 3765 -885 3785 -865
rect 3815 -885 3835 -865
rect 3915 -885 3935 -865
rect 3965 -885 3985 -865
rect 4015 -885 4035 -865
rect 4065 -885 4085 -865
rect 4115 -885 4135 -865
rect 4215 -885 4235 -865
rect 4265 -885 4285 -865
rect 4315 -885 4335 -865
rect 4365 -885 4385 -865
rect 4415 -885 4435 -865
rect 4515 -885 4535 -865
rect 4565 -885 4585 -865
rect 4615 -885 4635 -865
rect 4665 -885 4685 -865
rect 4715 -885 4735 -865
rect 4815 -885 4835 -865
rect 4865 -885 4885 -865
rect 4915 -885 4935 -865
rect 4965 -885 4985 -865
rect 5015 -885 5035 -865
rect 5115 -885 5135 -865
rect 5165 -885 5185 -865
rect 5215 -885 5235 -865
rect 5265 -885 5285 -865
rect 5315 -885 5335 -865
rect 5415 -885 5435 -865
rect 5465 -885 5485 -865
rect 5515 -885 5535 -865
rect 5565 -885 5585 -865
rect 5615 -885 5635 -865
rect 5715 -885 5735 -865
rect 5765 -885 5785 -865
rect 5815 -885 5835 -865
rect 5865 -885 5885 -865
rect 5915 -885 5935 -865
rect 6015 -885 6035 -865
rect 6065 -885 6085 -865
rect 6115 -885 6135 -865
rect 6165 -885 6185 -865
rect 6215 -885 6235 -865
rect 6315 -885 6335 -865
rect 6365 -885 6385 -865
rect 6415 -885 6435 -865
rect 6465 -885 6485 -865
rect 6515 -885 6535 -865
rect 6615 -885 6635 -865
rect 6665 -885 6685 -865
rect 6715 -885 6735 -865
rect 6765 -885 6785 -865
rect 6815 -885 6835 -865
rect 6915 -885 6935 -865
rect 6965 -885 6985 -865
rect 7015 -885 7035 -865
rect 7065 -885 7085 -865
rect 7115 -885 7135 -865
rect 7215 -885 7235 -865
rect 7265 -885 7285 -865
rect 7315 -885 7335 -865
rect 7365 -885 7385 -865
rect 7415 -885 7435 -865
rect 7515 -885 7535 -865
rect 7565 -885 7585 -865
rect 7615 -885 7635 -865
rect 7665 -885 7685 -865
rect 7715 -885 7735 -865
rect 7815 -885 7835 -865
rect 7865 -885 7885 -865
rect 7915 -885 7935 -865
rect 7965 -885 7985 -865
rect 8015 -885 8035 -865
rect 8115 -885 8135 -865
rect 8165 -885 8185 -865
rect 8215 -885 8235 -865
rect 8265 -885 8285 -865
rect 8315 -885 8335 -865
rect 8415 -885 8435 -865
rect 8465 -885 8485 -865
rect 8515 -885 8535 -865
rect 8565 -885 8585 -865
rect 8615 -885 8635 -865
rect 8715 -885 8735 -865
rect 8765 -885 8785 -865
rect 8815 -885 8835 -865
rect 8865 -885 8885 -865
rect 8915 -885 8935 -865
rect 9015 -885 9035 -865
rect 9065 -885 9085 -865
rect 9115 -885 9135 -865
rect 9165 -885 9185 -865
rect 9215 -885 9235 -865
rect 9315 -885 9335 -865
rect 9365 -885 9385 -865
rect 9415 -885 9435 -865
rect 9465 -885 9485 -865
rect 9515 -885 9535 -865
rect 9615 -885 9635 -865
rect 9665 -885 9685 -865
rect 9715 -885 9735 -865
rect 9765 -885 9785 -865
rect 9815 -885 9835 -865
rect 9915 -885 9935 -865
rect 9965 -885 9985 -865
rect 10015 -885 10035 -865
rect 10065 -885 10085 -865
rect 10115 -885 10135 -865
rect 10215 -885 10235 -865
rect 10265 -885 10285 -865
rect 10315 -885 10335 -865
rect 10365 -885 10385 -865
rect 10415 -885 10435 -865
rect 10515 -885 10535 -865
rect 10565 -885 10585 -865
rect 10615 -885 10635 -865
rect 10665 -885 10685 -865
rect 10715 -885 10735 -865
rect 10815 -885 10835 -865
rect 10865 -885 10885 -865
rect 10915 -885 10935 -865
rect 10965 -885 10985 -865
rect 11015 -885 11035 -865
rect 11115 -885 11135 -865
rect 11165 -885 11185 -865
rect 11215 -885 11235 -865
rect 11265 -885 11285 -865
rect 11315 -885 11335 -865
rect 11415 -885 11435 -865
rect 11465 -885 11485 -865
rect 11515 -885 11535 -865
rect 11565 -885 11585 -865
rect 11615 -885 11635 -865
rect 11715 -885 11735 -865
rect 11765 -885 11785 -865
rect 11815 -885 11835 -865
rect 11865 -885 11885 -865
rect 11915 -885 11935 -865
rect 12015 -885 12035 -865
rect 12065 -885 12085 -865
rect 12115 -885 12135 -865
rect 12165 -885 12185 -865
rect 12215 -885 12235 -865
rect 12315 -885 12335 -865
rect 12365 -885 12385 -865
rect 12415 -885 12435 -865
rect 12465 -885 12485 -865
rect 12515 -885 12535 -865
rect 12615 -885 12635 -865
rect 12665 -885 12685 -865
rect 12715 -885 12735 -865
rect 12765 -885 12785 -865
rect 12815 -885 12835 -865
rect 12915 -885 12935 -865
rect 12965 -885 12985 -865
rect 13015 -885 13035 -865
rect 13065 -885 13085 -865
rect 13115 -885 13135 -865
rect 13215 -885 13235 -865
rect 13265 -885 13285 -865
rect 13315 -885 13335 -865
rect 13365 -885 13385 -865
rect 13415 -885 13435 -865
rect 13515 -885 13535 -865
rect 13565 -885 13585 -865
rect 13615 -885 13635 -865
rect 13665 -885 13685 -865
rect 13715 -885 13735 -865
rect 13815 -885 13835 -865
rect 13865 -885 13885 -865
rect 13915 -885 13935 -865
rect 13965 -885 13985 -865
rect 14015 -885 14035 -865
rect 14115 -885 14135 -865
rect 14165 -885 14185 -865
rect 14215 -885 14235 -865
rect 14265 -885 14285 -865
rect 14315 -885 14335 -865
rect 14415 -885 14435 -865
rect 14465 -885 14485 -865
rect 14515 -885 14535 -865
rect 14565 -885 14585 -865
rect 14615 -885 14635 -865
rect 14715 -885 14735 -865
rect 14765 -885 14785 -865
rect 14815 -885 14835 -865
rect 14865 -885 14885 -865
rect 14915 -885 14935 -865
rect 15015 -885 15035 -865
rect 15065 -885 15085 -865
rect 15115 -885 15135 -865
rect 15165 -885 15185 -865
rect 15215 -885 15235 -865
rect 15315 -885 15335 -865
rect 15365 -885 15385 -865
rect 15415 -885 15435 -865
rect 15465 -885 15485 -865
rect 15515 -885 15535 -865
rect 15615 -885 15635 -865
rect 15665 -885 15685 -865
rect 15715 -885 15735 -865
rect 15765 -885 15785 -865
rect 15815 -885 15835 -865
rect 15915 -885 15935 -865
rect 15965 -885 15985 -865
rect 16015 -885 16035 -865
rect 16065 -885 16085 -865
rect 16115 -885 16135 -865
rect 16215 -885 16235 -865
rect 16265 -885 16285 -865
rect 16315 -885 16335 -865
rect 16365 -885 16385 -865
rect 16415 -885 16435 -865
rect 16515 -885 16535 -865
rect 16565 -885 16585 -865
rect 16615 -885 16635 -865
rect 16665 -885 16685 -865
rect 16715 -885 16735 -865
rect 16815 -885 16835 -865
rect 16865 -885 16885 -865
rect 16915 -885 16935 -865
rect 16965 -885 16985 -865
rect 17015 -885 17035 -865
rect 17115 -885 17135 -865
rect 17165 -885 17185 -865
rect 17215 -885 17235 -865
rect 17265 -885 17285 -865
rect 17315 -885 17335 -865
rect 17415 -885 17435 -865
rect 17465 -885 17485 -865
rect 17515 -885 17535 -865
rect 17565 -885 17585 -865
rect 17615 -885 17635 -865
rect 17715 -885 17735 -865
rect 17765 -885 17785 -865
rect 17815 -885 17835 -865
rect 17865 -885 17885 -865
rect 17915 -885 17935 -865
rect 18015 -885 18035 -865
rect 18065 -885 18085 -865
rect 18115 -885 18135 -865
rect 18165 -885 18185 -865
rect 18215 -885 18235 -865
rect 18315 -885 18335 -865
rect 18365 -885 18385 -865
rect 18415 -885 18435 -865
rect 18465 -885 18485 -865
rect 18515 -885 18535 -865
rect 18615 -885 18635 -865
rect 18665 -885 18685 -865
rect 18715 -885 18735 -865
rect 18765 -885 18785 -865
rect 18815 -885 18835 -865
rect 18915 -885 18935 -865
rect 18965 -885 18985 -865
rect 19015 -885 19035 -865
rect 19065 -885 19085 -865
rect 19115 -885 19135 -865
rect 19215 -885 19235 -865
rect 19265 -885 19285 -865
rect 19315 -885 19335 -865
rect 19365 -885 19385 -865
rect 19415 -885 19435 -865
rect 19515 -885 19535 -865
rect 19565 -885 19585 -865
rect 19615 -885 19635 -865
rect 19665 -885 19685 -865
rect 19715 -885 19735 -865
rect 19815 -885 19835 -865
rect 19865 -885 19885 -865
rect 19915 -885 19935 -865
rect 19965 -885 19985 -865
rect 20015 -885 20035 -865
rect 20115 -885 20135 -865
rect 20165 -885 20185 -865
rect 20215 -885 20235 -865
rect 20265 -885 20285 -865
rect 20315 -885 20335 -865
rect 20415 -885 20435 -865
rect 20465 -885 20485 -865
rect 20515 -885 20535 -865
rect 20565 -885 20585 -865
rect 20615 -885 20635 -865
rect 20715 -885 20735 -865
rect 20765 -885 20785 -865
rect 20815 -885 20835 -865
rect 20865 -885 20885 -865
rect 20915 -885 20935 -865
rect 21015 -885 21035 -865
rect 21065 -885 21085 -865
rect 21115 -885 21135 -865
rect 21165 -885 21185 -865
rect 21215 -885 21235 -865
rect 21315 -885 21335 -865
rect 21365 -885 21385 -865
rect 21415 -885 21435 -865
rect 21465 -885 21485 -865
rect 21515 -885 21535 -865
rect 21615 -885 21635 -865
rect 21665 -885 21685 -865
rect 21715 -885 21735 -865
rect 21765 -885 21785 -865
rect 21815 -885 21835 -865
rect 21915 -885 21935 -865
rect 21965 -885 21985 -865
rect 22015 -885 22035 -865
rect 22065 -885 22085 -865
rect 22115 -885 22135 -865
rect 22215 -885 22235 -865
rect 22265 -885 22285 -865
rect 22315 -885 22335 -865
rect 22365 -885 22385 -865
rect 22415 -885 22435 -865
rect 22515 -885 22535 -865
rect 22565 -885 22585 -865
rect 22615 -885 22635 -865
rect 22665 -885 22685 -865
rect 22715 -885 22735 -865
rect 22815 -885 22835 -865
rect 22865 -885 22885 -865
rect 22915 -885 22935 -865
rect 22965 -885 22985 -865
rect 23015 -885 23035 -865
rect 23115 -885 23135 -865
rect 23165 -885 23185 -865
rect 23215 -885 23235 -865
rect 23265 -885 23285 -865
rect 23315 -885 23335 -865
rect 23415 -885 23435 -865
rect 23465 -885 23485 -865
rect 23515 -885 23535 -865
rect 23565 -885 23585 -865
rect 23615 -885 23635 -865
rect 23715 -885 23735 -865
rect 23765 -885 23785 -865
rect 23815 -885 23835 -865
rect 23865 -885 23885 -865
rect 23915 -885 23935 -865
rect 24015 -885 24035 -865
rect 24065 -885 24085 -865
rect 24115 -885 24135 -865
rect 24165 -885 24185 -865
rect 24215 -885 24235 -865
rect 24315 -885 24335 -865
rect 24365 -885 24385 -865
rect 24415 -885 24435 -865
rect 24465 -885 24485 -865
rect 24515 -885 24535 -865
rect 24615 -885 24635 -865
rect 24665 -885 24685 -865
rect 24715 -885 24735 -865
rect 24765 -885 24785 -865
rect 24815 -885 24835 -865
rect 24915 -885 24935 -865
rect 24965 -885 24985 -865
rect 25015 -885 25035 -865
rect 25065 -885 25085 -865
rect 25115 -885 25135 -865
rect 25215 -885 25235 -865
rect 25265 -885 25285 -865
rect 25315 -885 25335 -865
rect 25365 -885 25385 -865
rect 25415 -885 25435 -865
rect 25515 -885 25535 -865
rect 25565 -885 25585 -865
rect 25615 -885 25635 -865
rect 25665 -885 25685 -865
rect 25715 -885 25735 -865
rect 25815 -885 25835 -865
rect 25865 -885 25885 -865
rect 25915 -885 25935 -865
rect 25965 -885 25985 -865
rect 26015 -885 26035 -865
rect 26115 -885 26135 -865
rect 26165 -885 26185 -865
rect 26215 -885 26235 -865
rect 26265 -885 26285 -865
rect 26315 -885 26335 -865
rect 26415 -885 26435 -865
rect 26465 -885 26485 -865
rect 26515 -885 26535 -865
rect 26565 -885 26585 -865
rect 26615 -885 26635 -865
rect 26715 -885 26735 -865
rect 26765 -885 26785 -865
rect 26815 -885 26835 -865
rect 26865 -885 26885 -865
rect 26915 -885 26935 -865
rect 27015 -885 27035 -865
rect 27065 -885 27085 -865
rect 27115 -885 27135 -865
rect 27165 -885 27185 -865
rect 27215 -885 27235 -865
rect 27315 -885 27335 -865
rect 27365 -885 27385 -865
rect 27415 -885 27435 -865
rect 27465 -885 27485 -865
rect 27515 -885 27535 -865
rect 27615 -885 27635 -865
rect 27665 -885 27685 -865
rect 27715 -885 27735 -865
rect 27765 -885 27785 -865
rect 27815 -885 27835 -865
rect 27915 -885 27935 -865
rect 27965 -885 27985 -865
rect 28015 -885 28035 -865
rect 28065 -885 28085 -865
rect 28115 -885 28135 -865
rect 28215 -885 28235 -865
rect 28265 -885 28285 -865
rect 28315 -885 28335 -865
rect 28365 -885 28385 -865
rect 28415 -885 28435 -865
rect 28515 -885 28535 -865
rect 28565 -885 28585 -865
rect 28615 -885 28635 -865
rect 28665 -885 28685 -865
rect 28715 -885 28735 -865
<< locali >>
rect -650 5585 32100 5600
rect -650 5565 -635 5585
rect -615 5565 -585 5585
rect -565 5565 -535 5585
rect -515 5565 -485 5585
rect -465 5565 -435 5585
rect -415 5565 -385 5585
rect -365 5565 -335 5585
rect -315 5565 -285 5585
rect -265 5565 -235 5585
rect -215 5565 -185 5585
rect -165 5565 -135 5585
rect -115 5565 -85 5585
rect -65 5565 -35 5585
rect -15 5565 15 5585
rect 35 5565 65 5585
rect 85 5565 115 5585
rect 135 5565 165 5585
rect 185 5565 215 5585
rect 235 5565 265 5585
rect 285 5565 315 5585
rect 335 5565 365 5585
rect 385 5565 415 5585
rect 435 5565 465 5585
rect 485 5565 515 5585
rect 535 5565 565 5585
rect 585 5565 615 5585
rect 635 5565 665 5585
rect 685 5565 715 5585
rect 735 5565 765 5585
rect 785 5565 815 5585
rect 835 5565 865 5585
rect 885 5565 915 5585
rect 935 5565 965 5585
rect 985 5565 1015 5585
rect 1035 5565 1065 5585
rect 1085 5565 1115 5585
rect 1135 5565 1165 5585
rect 1185 5565 1215 5585
rect 1235 5565 1265 5585
rect 1285 5565 1315 5585
rect 1335 5565 1365 5585
rect 1385 5565 1415 5585
rect 1435 5565 1465 5585
rect 1485 5565 1515 5585
rect 1535 5565 1565 5585
rect 1585 5565 1615 5585
rect 1635 5565 1665 5585
rect 1685 5565 1715 5585
rect 1735 5565 1765 5585
rect 1785 5565 1815 5585
rect 1835 5565 1865 5585
rect 1885 5565 1915 5585
rect 1935 5565 1965 5585
rect 1985 5565 2015 5585
rect 2035 5565 2065 5585
rect 2085 5565 2115 5585
rect 2135 5565 2165 5585
rect 2185 5565 2215 5585
rect 2235 5565 2265 5585
rect 2285 5565 2315 5585
rect 2335 5565 2365 5585
rect 2385 5565 2415 5585
rect 2435 5565 2465 5585
rect 2485 5565 2515 5585
rect 2535 5565 2565 5585
rect 2585 5565 2615 5585
rect 2635 5565 2665 5585
rect 2685 5565 2715 5585
rect 2735 5565 2765 5585
rect 2785 5565 2815 5585
rect 2835 5565 2865 5585
rect 2885 5565 2915 5585
rect 2935 5565 2965 5585
rect 2985 5565 3015 5585
rect 3035 5565 3065 5585
rect 3085 5565 3115 5585
rect 3135 5565 3165 5585
rect 3185 5565 3215 5585
rect 3235 5565 3265 5585
rect 3285 5565 3315 5585
rect 3335 5565 3365 5585
rect 3385 5565 3415 5585
rect 3435 5565 3465 5585
rect 3485 5565 3515 5585
rect 3535 5565 3565 5585
rect 3585 5565 3615 5585
rect 3635 5565 3665 5585
rect 3685 5565 3715 5585
rect 3735 5565 3765 5585
rect 3785 5565 3815 5585
rect 3835 5565 3865 5585
rect 3885 5565 3915 5585
rect 3935 5565 3965 5585
rect 3985 5565 4015 5585
rect 4035 5565 4065 5585
rect 4085 5565 4115 5585
rect 4135 5565 4165 5585
rect 4185 5565 4215 5585
rect 4235 5565 4265 5585
rect 4285 5565 4315 5585
rect 4335 5565 4365 5585
rect 4385 5565 4415 5585
rect 4435 5565 4465 5585
rect 4485 5565 4515 5585
rect 4535 5565 4565 5585
rect 4585 5565 4615 5585
rect 4635 5565 4665 5585
rect 4685 5565 4715 5585
rect 4735 5565 4765 5585
rect 4785 5565 4815 5585
rect 4835 5565 4865 5585
rect 4885 5565 4915 5585
rect 4935 5565 4965 5585
rect 4985 5565 5015 5585
rect 5035 5565 5065 5585
rect 5085 5565 5115 5585
rect 5135 5565 5165 5585
rect 5185 5565 5215 5585
rect 5235 5565 5265 5585
rect 5285 5565 5315 5585
rect 5335 5565 5365 5585
rect 5385 5565 5415 5585
rect 5435 5565 5465 5585
rect 5485 5565 5515 5585
rect 5535 5565 5565 5585
rect 5585 5565 5615 5585
rect 5635 5565 5665 5585
rect 5685 5565 5715 5585
rect 5735 5565 5765 5585
rect 5785 5565 5815 5585
rect 5835 5565 5865 5585
rect 5885 5565 5915 5585
rect 5935 5565 5965 5585
rect 5985 5565 6015 5585
rect 6035 5565 6065 5585
rect 6085 5565 6115 5585
rect 6135 5565 6165 5585
rect 6185 5565 6215 5585
rect 6235 5565 6265 5585
rect 6285 5565 6315 5585
rect 6335 5565 6365 5585
rect 6385 5565 6415 5585
rect 6435 5565 6465 5585
rect 6485 5565 6515 5585
rect 6535 5565 6565 5585
rect 6585 5565 6615 5585
rect 6635 5565 6665 5585
rect 6685 5565 6715 5585
rect 6735 5565 6765 5585
rect 6785 5565 6815 5585
rect 6835 5565 6865 5585
rect 6885 5565 6915 5585
rect 6935 5565 6965 5585
rect 6985 5565 7015 5585
rect 7035 5565 7065 5585
rect 7085 5565 7115 5585
rect 7135 5565 7165 5585
rect 7185 5565 7215 5585
rect 7235 5565 7265 5585
rect 7285 5565 7315 5585
rect 7335 5565 7365 5585
rect 7385 5565 7415 5585
rect 7435 5565 7465 5585
rect 7485 5565 7515 5585
rect 7535 5565 7565 5585
rect 7585 5565 7615 5585
rect 7635 5565 7665 5585
rect 7685 5565 7715 5585
rect 7735 5565 7765 5585
rect 7785 5565 7815 5585
rect 7835 5565 7865 5585
rect 7885 5565 7915 5585
rect 7935 5565 7965 5585
rect 7985 5565 8015 5585
rect 8035 5565 8065 5585
rect 8085 5565 8115 5585
rect 8135 5565 8165 5585
rect 8185 5565 8215 5585
rect 8235 5565 8265 5585
rect 8285 5565 8315 5585
rect 8335 5565 8365 5585
rect 8385 5565 8415 5585
rect 8435 5565 8465 5585
rect 8485 5565 8515 5585
rect 8535 5565 8565 5585
rect 8585 5565 8615 5585
rect 8635 5565 8665 5585
rect 8685 5565 8715 5585
rect 8735 5565 8765 5585
rect 8785 5565 8815 5585
rect 8835 5565 8865 5585
rect 8885 5565 8915 5585
rect 8935 5565 8965 5585
rect 8985 5565 9015 5585
rect 9035 5565 9065 5585
rect 9085 5565 9115 5585
rect 9135 5565 9165 5585
rect 9185 5565 9215 5585
rect 9235 5565 9265 5585
rect 9285 5565 9315 5585
rect 9335 5565 9365 5585
rect 9385 5565 9415 5585
rect 9435 5565 9465 5585
rect 9485 5565 9515 5585
rect 9535 5565 9565 5585
rect 9585 5565 9615 5585
rect 9635 5565 9665 5585
rect 9685 5565 9715 5585
rect 9735 5565 9765 5585
rect 9785 5565 9815 5585
rect 9835 5565 9865 5585
rect 9885 5565 9915 5585
rect 9935 5565 9965 5585
rect 9985 5565 10015 5585
rect 10035 5565 10065 5585
rect 10085 5565 10115 5585
rect 10135 5565 10165 5585
rect 10185 5565 10215 5585
rect 10235 5565 10265 5585
rect 10285 5565 10315 5585
rect 10335 5565 10365 5585
rect 10385 5565 10415 5585
rect 10435 5565 10465 5585
rect 10485 5565 10515 5585
rect 10535 5565 10565 5585
rect 10585 5565 10615 5585
rect 10635 5565 10665 5585
rect 10685 5565 10715 5585
rect 10735 5565 10765 5585
rect 10785 5565 10815 5585
rect 10835 5565 10865 5585
rect 10885 5565 10915 5585
rect 10935 5565 10965 5585
rect 10985 5565 11015 5585
rect 11035 5565 11065 5585
rect 11085 5565 11115 5585
rect 11135 5565 11165 5585
rect 11185 5565 11215 5585
rect 11235 5565 11265 5585
rect 11285 5565 11315 5585
rect 11335 5565 11365 5585
rect 11385 5565 11415 5585
rect 11435 5565 11465 5585
rect 11485 5565 11515 5585
rect 11535 5565 11565 5585
rect 11585 5565 11615 5585
rect 11635 5565 11665 5585
rect 11685 5565 11715 5585
rect 11735 5565 11765 5585
rect 11785 5565 11815 5585
rect 11835 5565 11865 5585
rect 11885 5565 11915 5585
rect 11935 5565 11965 5585
rect 11985 5565 12015 5585
rect 12035 5565 12065 5585
rect 12085 5565 12115 5585
rect 12135 5565 12165 5585
rect 12185 5565 12215 5585
rect 12235 5565 12265 5585
rect 12285 5565 12315 5585
rect 12335 5565 12365 5585
rect 12385 5565 12415 5585
rect 12435 5565 12465 5585
rect 12485 5565 12515 5585
rect 12535 5565 12565 5585
rect 12585 5565 12615 5585
rect 12635 5565 12665 5585
rect 12685 5565 12715 5585
rect 12735 5565 12765 5585
rect 12785 5565 12815 5585
rect 12835 5565 12865 5585
rect 12885 5565 12915 5585
rect 12935 5565 12965 5585
rect 12985 5565 13015 5585
rect 13035 5565 13065 5585
rect 13085 5565 13115 5585
rect 13135 5565 13165 5585
rect 13185 5565 13215 5585
rect 13235 5565 13265 5585
rect 13285 5565 13315 5585
rect 13335 5565 13365 5585
rect 13385 5565 13415 5585
rect 13435 5565 13465 5585
rect 13485 5565 13515 5585
rect 13535 5565 13565 5585
rect 13585 5565 13615 5585
rect 13635 5565 13665 5585
rect 13685 5565 13715 5585
rect 13735 5565 13765 5585
rect 13785 5565 13815 5585
rect 13835 5565 13865 5585
rect 13885 5565 13915 5585
rect 13935 5565 13965 5585
rect 13985 5565 14015 5585
rect 14035 5565 14065 5585
rect 14085 5565 14115 5585
rect 14135 5565 14165 5585
rect 14185 5565 14215 5585
rect 14235 5565 14265 5585
rect 14285 5565 14315 5585
rect 14335 5565 14365 5585
rect 14385 5565 14415 5585
rect 14435 5565 14465 5585
rect 14485 5565 14515 5585
rect 14535 5565 14565 5585
rect 14585 5565 14615 5585
rect 14635 5565 14665 5585
rect 14685 5565 14715 5585
rect 14735 5565 14765 5585
rect 14785 5565 14815 5585
rect 14835 5565 14865 5585
rect 14885 5565 14915 5585
rect 14935 5565 14965 5585
rect 14985 5565 15015 5585
rect 15035 5565 15065 5585
rect 15085 5565 15115 5585
rect 15135 5565 15165 5585
rect 15185 5565 15215 5585
rect 15235 5565 15265 5585
rect 15285 5565 15315 5585
rect 15335 5565 15365 5585
rect 15385 5565 15415 5585
rect 15435 5565 15465 5585
rect 15485 5565 15515 5585
rect 15535 5565 15565 5585
rect 15585 5565 15615 5585
rect 15635 5565 15665 5585
rect 15685 5565 15715 5585
rect 15735 5565 15765 5585
rect 15785 5565 15815 5585
rect 15835 5565 15865 5585
rect 15885 5565 15915 5585
rect 15935 5565 15965 5585
rect 15985 5565 16015 5585
rect 16035 5565 16065 5585
rect 16085 5565 16115 5585
rect 16135 5565 16165 5585
rect 16185 5565 16215 5585
rect 16235 5565 16265 5585
rect 16285 5565 16315 5585
rect 16335 5565 16365 5585
rect 16385 5565 16415 5585
rect 16435 5565 16465 5585
rect 16485 5565 16515 5585
rect 16535 5565 16565 5585
rect 16585 5565 16615 5585
rect 16635 5565 16665 5585
rect 16685 5565 16715 5585
rect 16735 5565 16765 5585
rect 16785 5565 16815 5585
rect 16835 5565 16865 5585
rect 16885 5565 16915 5585
rect 16935 5565 16965 5585
rect 16985 5565 17015 5585
rect 17035 5565 17065 5585
rect 17085 5565 17115 5585
rect 17135 5565 17165 5585
rect 17185 5565 17215 5585
rect 17235 5565 17265 5585
rect 17285 5565 17315 5585
rect 17335 5565 17365 5585
rect 17385 5565 17415 5585
rect 17435 5565 17465 5585
rect 17485 5565 17515 5585
rect 17535 5565 17565 5585
rect 17585 5565 17615 5585
rect 17635 5565 17665 5585
rect 17685 5565 17715 5585
rect 17735 5565 17765 5585
rect 17785 5565 17815 5585
rect 17835 5565 17865 5585
rect 17885 5565 17915 5585
rect 17935 5565 17965 5585
rect 17985 5565 18015 5585
rect 18035 5565 18065 5585
rect 18085 5565 18115 5585
rect 18135 5565 18165 5585
rect 18185 5565 18215 5585
rect 18235 5565 18265 5585
rect 18285 5565 18315 5585
rect 18335 5565 18365 5585
rect 18385 5565 18415 5585
rect 18435 5565 18465 5585
rect 18485 5565 18515 5585
rect 18535 5565 18565 5585
rect 18585 5565 18615 5585
rect 18635 5565 18665 5585
rect 18685 5565 18715 5585
rect 18735 5565 18765 5585
rect 18785 5565 18815 5585
rect 18835 5565 18865 5585
rect 18885 5565 18915 5585
rect 18935 5565 18965 5585
rect 18985 5565 19015 5585
rect 19035 5565 19065 5585
rect 19085 5565 19115 5585
rect 19135 5565 19165 5585
rect 19185 5565 19215 5585
rect 19235 5565 19265 5585
rect 19285 5565 19315 5585
rect 19335 5565 19365 5585
rect 19385 5565 19415 5585
rect 19435 5565 19465 5585
rect 19485 5565 19515 5585
rect 19535 5565 19565 5585
rect 19585 5565 19615 5585
rect 19635 5565 19665 5585
rect 19685 5565 19715 5585
rect 19735 5565 19765 5585
rect 19785 5565 19815 5585
rect 19835 5565 19865 5585
rect 19885 5565 19915 5585
rect 19935 5565 19965 5585
rect 19985 5565 20015 5585
rect 20035 5565 20065 5585
rect 20085 5565 20115 5585
rect 20135 5565 20165 5585
rect 20185 5565 20215 5585
rect 20235 5565 20265 5585
rect 20285 5565 20315 5585
rect 20335 5565 20365 5585
rect 20385 5565 20415 5585
rect 20435 5565 20465 5585
rect 20485 5565 20515 5585
rect 20535 5565 20565 5585
rect 20585 5565 20615 5585
rect 20635 5565 20665 5585
rect 20685 5565 20715 5585
rect 20735 5565 20765 5585
rect 20785 5565 20815 5585
rect 20835 5565 20865 5585
rect 20885 5565 20915 5585
rect 20935 5565 20965 5585
rect 20985 5565 21015 5585
rect 21035 5565 21065 5585
rect 21085 5565 21115 5585
rect 21135 5565 21165 5585
rect 21185 5565 21215 5585
rect 21235 5565 21265 5585
rect 21285 5565 21315 5585
rect 21335 5565 21365 5585
rect 21385 5565 21415 5585
rect 21435 5565 21465 5585
rect 21485 5565 21515 5585
rect 21535 5565 21565 5585
rect 21585 5565 21615 5585
rect 21635 5565 21665 5585
rect 21685 5565 21715 5585
rect 21735 5565 21765 5585
rect 21785 5565 21815 5585
rect 21835 5565 21865 5585
rect 21885 5565 21915 5585
rect 21935 5565 21965 5585
rect 21985 5565 22015 5585
rect 22035 5565 22065 5585
rect 22085 5565 22115 5585
rect 22135 5565 22165 5585
rect 22185 5565 22215 5585
rect 22235 5565 22265 5585
rect 22285 5565 22315 5585
rect 22335 5565 22365 5585
rect 22385 5565 22415 5585
rect 22435 5565 22465 5585
rect 22485 5565 22515 5585
rect 22535 5565 22565 5585
rect 22585 5565 22615 5585
rect 22635 5565 22665 5585
rect 22685 5565 22715 5585
rect 22735 5565 22765 5585
rect 22785 5565 22815 5585
rect 22835 5565 22865 5585
rect 22885 5565 22915 5585
rect 22935 5565 22965 5585
rect 22985 5565 23015 5585
rect 23035 5565 23065 5585
rect 23085 5565 23115 5585
rect 23135 5565 23165 5585
rect 23185 5565 23215 5585
rect 23235 5565 23265 5585
rect 23285 5565 23315 5585
rect 23335 5565 23365 5585
rect 23385 5565 23415 5585
rect 23435 5565 23465 5585
rect 23485 5565 23515 5585
rect 23535 5565 23565 5585
rect 23585 5565 23615 5585
rect 23635 5565 23665 5585
rect 23685 5565 23715 5585
rect 23735 5565 23765 5585
rect 23785 5565 23815 5585
rect 23835 5565 23865 5585
rect 23885 5565 23915 5585
rect 23935 5565 23965 5585
rect 23985 5565 24015 5585
rect 24035 5565 24065 5585
rect 24085 5565 24115 5585
rect 24135 5565 24165 5585
rect 24185 5565 24215 5585
rect 24235 5565 24265 5585
rect 24285 5565 24315 5585
rect 24335 5565 24365 5585
rect 24385 5565 24415 5585
rect 24435 5565 24465 5585
rect 24485 5565 24515 5585
rect 24535 5565 24565 5585
rect 24585 5565 24615 5585
rect 24635 5565 24665 5585
rect 24685 5565 24715 5585
rect 24735 5565 24765 5585
rect 24785 5565 24815 5585
rect 24835 5565 24865 5585
rect 24885 5565 24915 5585
rect 24935 5565 24965 5585
rect 24985 5565 25015 5585
rect 25035 5565 25065 5585
rect 25085 5565 25115 5585
rect 25135 5565 25165 5585
rect 25185 5565 25215 5585
rect 25235 5565 25265 5585
rect 25285 5565 25315 5585
rect 25335 5565 25365 5585
rect 25385 5565 25415 5585
rect 25435 5565 25465 5585
rect 25485 5565 25515 5585
rect 25535 5565 25565 5585
rect 25585 5565 25615 5585
rect 25635 5565 25665 5585
rect 25685 5565 25715 5585
rect 25735 5565 25765 5585
rect 25785 5565 25815 5585
rect 25835 5565 25865 5585
rect 25885 5565 25915 5585
rect 25935 5565 25965 5585
rect 25985 5565 26015 5585
rect 26035 5565 26065 5585
rect 26085 5565 26115 5585
rect 26135 5565 26165 5585
rect 26185 5565 26215 5585
rect 26235 5565 26265 5585
rect 26285 5565 26315 5585
rect 26335 5565 26365 5585
rect 26385 5565 26415 5585
rect 26435 5565 26465 5585
rect 26485 5565 26515 5585
rect 26535 5565 26565 5585
rect 26585 5565 26615 5585
rect 26635 5565 26665 5585
rect 26685 5565 26715 5585
rect 26735 5565 26765 5585
rect 26785 5565 26815 5585
rect 26835 5565 26865 5585
rect 26885 5565 26915 5585
rect 26935 5565 26965 5585
rect 26985 5565 27015 5585
rect 27035 5565 27065 5585
rect 27085 5565 27115 5585
rect 27135 5565 27165 5585
rect 27185 5565 27215 5585
rect 27235 5565 27265 5585
rect 27285 5565 27315 5585
rect 27335 5565 27365 5585
rect 27385 5565 27415 5585
rect 27435 5565 27465 5585
rect 27485 5565 27515 5585
rect 27535 5565 27565 5585
rect 27585 5565 27615 5585
rect 27635 5565 27665 5585
rect 27685 5565 27715 5585
rect 27735 5565 27765 5585
rect 27785 5565 27815 5585
rect 27835 5565 27865 5585
rect 27885 5565 27915 5585
rect 27935 5565 27965 5585
rect 27985 5565 28015 5585
rect 28035 5565 28065 5585
rect 28085 5565 28115 5585
rect 28135 5565 28165 5585
rect 28185 5565 28215 5585
rect 28235 5565 28265 5585
rect 28285 5565 28315 5585
rect 28335 5565 28365 5585
rect 28385 5565 28415 5585
rect 28435 5565 28465 5585
rect 28485 5565 28515 5585
rect 28535 5565 28565 5585
rect 28585 5565 28615 5585
rect 28635 5565 28665 5585
rect 28685 5565 28715 5585
rect 28735 5565 28765 5585
rect 28785 5565 28815 5585
rect 28835 5565 28865 5585
rect 28885 5565 28915 5585
rect 28935 5565 28965 5585
rect 28985 5565 29015 5585
rect 29035 5565 29065 5585
rect 29085 5565 29115 5585
rect 29135 5565 29165 5585
rect 29185 5565 29215 5585
rect 29235 5565 29265 5585
rect 29285 5565 29315 5585
rect 29335 5565 29365 5585
rect 29385 5565 29415 5585
rect 29435 5565 29465 5585
rect 29485 5565 29515 5585
rect 29535 5565 29565 5585
rect 29585 5565 29615 5585
rect 29635 5565 29665 5585
rect 29685 5565 29715 5585
rect 29735 5565 29765 5585
rect 29785 5565 29815 5585
rect 29835 5565 29865 5585
rect 29885 5565 29915 5585
rect 29935 5565 29965 5585
rect 29985 5565 30015 5585
rect 30035 5565 30065 5585
rect 30085 5565 30115 5585
rect 30135 5565 30165 5585
rect 30185 5565 30215 5585
rect 30235 5565 30265 5585
rect 30285 5565 30315 5585
rect 30335 5565 30365 5585
rect 30385 5565 30415 5585
rect 30435 5565 30465 5585
rect 30485 5565 30515 5585
rect 30535 5565 30565 5585
rect 30585 5565 30615 5585
rect 30635 5565 30665 5585
rect 30685 5565 30715 5585
rect 30735 5565 30765 5585
rect 30785 5565 30815 5585
rect 30835 5565 30865 5585
rect 30885 5565 30915 5585
rect 30935 5565 30965 5585
rect 30985 5565 31015 5585
rect 31035 5565 31065 5585
rect 31085 5565 31115 5585
rect 31135 5565 31165 5585
rect 31185 5565 31215 5585
rect 31235 5565 31265 5585
rect 31285 5565 31315 5585
rect 31335 5565 31365 5585
rect 31385 5565 31415 5585
rect 31435 5565 31465 5585
rect 31485 5565 31515 5585
rect 31535 5565 31565 5585
rect 31585 5565 31615 5585
rect 31635 5565 31665 5585
rect 31685 5565 31715 5585
rect 31735 5565 31765 5585
rect 31785 5565 31815 5585
rect 31835 5565 31865 5585
rect 31885 5565 31915 5585
rect 31935 5565 31965 5585
rect 31985 5565 32015 5585
rect 32035 5565 32065 5585
rect 32085 5565 32100 5585
rect -650 5550 32100 5565
rect -650 5485 -600 5500
rect -650 5465 -635 5485
rect -615 5465 -600 5485
rect -650 5435 -600 5465
rect -650 5415 -635 5435
rect -615 5415 -600 5435
rect -650 5385 -600 5415
rect -650 5365 -635 5385
rect -615 5365 -600 5385
rect -650 5335 -600 5365
rect -650 5315 -635 5335
rect -615 5315 -600 5335
rect -650 5285 -600 5315
rect -650 5265 -635 5285
rect -615 5265 -600 5285
rect -650 5235 -600 5265
rect -650 5215 -635 5235
rect -615 5215 -600 5235
rect -650 5185 -600 5215
rect -650 5165 -635 5185
rect -615 5165 -600 5185
rect -650 5135 -600 5165
rect -650 5115 -635 5135
rect -615 5115 -600 5135
rect -650 5085 -600 5115
rect -650 5065 -635 5085
rect -615 5065 -600 5085
rect -650 5035 -600 5065
rect -650 5015 -635 5035
rect -615 5015 -600 5035
rect -650 5000 -600 5015
rect -500 5485 -450 5500
rect -500 5465 -485 5485
rect -465 5465 -450 5485
rect -500 5435 -450 5465
rect -500 5415 -485 5435
rect -465 5415 -450 5435
rect -500 5385 -450 5415
rect -500 5365 -485 5385
rect -465 5365 -450 5385
rect -500 5335 -450 5365
rect -500 5315 -485 5335
rect -465 5315 -450 5335
rect -500 5285 -450 5315
rect -500 5265 -485 5285
rect -465 5265 -450 5285
rect -500 5235 -450 5265
rect -500 5215 -485 5235
rect -465 5215 -450 5235
rect -500 5185 -450 5215
rect -500 5165 -485 5185
rect -465 5165 -450 5185
rect -500 5135 -450 5165
rect -500 5115 -485 5135
rect -465 5115 -450 5135
rect -500 5085 -450 5115
rect -500 5065 -485 5085
rect -465 5065 -450 5085
rect -500 5035 -450 5065
rect -500 5015 -485 5035
rect -465 5015 -450 5035
rect -500 5000 -450 5015
rect -350 5485 -300 5500
rect -350 5465 -335 5485
rect -315 5465 -300 5485
rect -350 5435 -300 5465
rect -350 5415 -335 5435
rect -315 5415 -300 5435
rect -350 5385 -300 5415
rect -350 5365 -335 5385
rect -315 5365 -300 5385
rect -350 5335 -300 5365
rect -350 5315 -335 5335
rect -315 5315 -300 5335
rect -350 5285 -300 5315
rect -350 5265 -335 5285
rect -315 5265 -300 5285
rect -350 5235 -300 5265
rect -350 5215 -335 5235
rect -315 5215 -300 5235
rect -350 5185 -300 5215
rect -350 5165 -335 5185
rect -315 5165 -300 5185
rect -350 5135 -300 5165
rect -350 5115 -335 5135
rect -315 5115 -300 5135
rect -350 5085 -300 5115
rect -350 5065 -335 5085
rect -315 5065 -300 5085
rect -350 5035 -300 5065
rect -350 5015 -335 5035
rect -315 5015 -300 5035
rect -350 5000 -300 5015
rect -200 5485 -150 5500
rect -200 5465 -185 5485
rect -165 5465 -150 5485
rect -200 5435 -150 5465
rect -200 5415 -185 5435
rect -165 5415 -150 5435
rect -200 5385 -150 5415
rect -200 5365 -185 5385
rect -165 5365 -150 5385
rect -200 5335 -150 5365
rect -200 5315 -185 5335
rect -165 5315 -150 5335
rect -200 5285 -150 5315
rect -200 5265 -185 5285
rect -165 5265 -150 5285
rect -200 5235 -150 5265
rect -200 5215 -185 5235
rect -165 5215 -150 5235
rect -200 5185 -150 5215
rect -200 5165 -185 5185
rect -165 5165 -150 5185
rect -200 5135 -150 5165
rect -200 5115 -185 5135
rect -165 5115 -150 5135
rect -200 5085 -150 5115
rect -200 5065 -185 5085
rect -165 5065 -150 5085
rect -200 5035 -150 5065
rect -200 5015 -185 5035
rect -165 5015 -150 5035
rect -200 5000 -150 5015
rect -50 5485 0 5500
rect -50 5465 -35 5485
rect -15 5465 0 5485
rect -50 5435 0 5465
rect -50 5415 -35 5435
rect -15 5415 0 5435
rect -50 5385 0 5415
rect -50 5365 -35 5385
rect -15 5365 0 5385
rect -50 5335 0 5365
rect -50 5315 -35 5335
rect -15 5315 0 5335
rect -50 5285 0 5315
rect -50 5265 -35 5285
rect -15 5265 0 5285
rect -50 5235 0 5265
rect -50 5215 -35 5235
rect -15 5215 0 5235
rect -50 5185 0 5215
rect -50 5165 -35 5185
rect -15 5165 0 5185
rect -50 5135 0 5165
rect -50 5115 -35 5135
rect -15 5115 0 5135
rect -50 5085 0 5115
rect -50 5065 -35 5085
rect -15 5065 0 5085
rect -50 5035 0 5065
rect -50 5015 -35 5035
rect -15 5015 0 5035
rect -50 5000 0 5015
rect 550 5485 600 5500
rect 550 5465 565 5485
rect 585 5465 600 5485
rect 550 5435 600 5465
rect 550 5415 565 5435
rect 585 5415 600 5435
rect 550 5385 600 5415
rect 550 5365 565 5385
rect 585 5365 600 5385
rect 550 5335 600 5365
rect 550 5315 565 5335
rect 585 5315 600 5335
rect 550 5285 600 5315
rect 550 5265 565 5285
rect 585 5265 600 5285
rect 550 5235 600 5265
rect 550 5215 565 5235
rect 585 5215 600 5235
rect 550 5185 600 5215
rect 550 5165 565 5185
rect 585 5165 600 5185
rect 550 5135 600 5165
rect 550 5115 565 5135
rect 585 5115 600 5135
rect 550 5085 600 5115
rect 550 5065 565 5085
rect 585 5065 600 5085
rect 550 5035 600 5065
rect 550 5015 565 5035
rect 585 5015 600 5035
rect 550 5000 600 5015
rect 700 5485 750 5500
rect 700 5465 715 5485
rect 735 5465 750 5485
rect 700 5435 750 5465
rect 700 5415 715 5435
rect 735 5415 750 5435
rect 700 5385 750 5415
rect 700 5365 715 5385
rect 735 5365 750 5385
rect 700 5335 750 5365
rect 700 5315 715 5335
rect 735 5315 750 5335
rect 700 5285 750 5315
rect 700 5265 715 5285
rect 735 5265 750 5285
rect 700 5235 750 5265
rect 700 5215 715 5235
rect 735 5215 750 5235
rect 700 5185 750 5215
rect 700 5165 715 5185
rect 735 5165 750 5185
rect 700 5135 750 5165
rect 700 5115 715 5135
rect 735 5115 750 5135
rect 700 5085 750 5115
rect 700 5065 715 5085
rect 735 5065 750 5085
rect 700 5035 750 5065
rect 700 5015 715 5035
rect 735 5015 750 5035
rect 700 5000 750 5015
rect 850 5485 900 5500
rect 850 5465 865 5485
rect 885 5465 900 5485
rect 850 5435 900 5465
rect 850 5415 865 5435
rect 885 5415 900 5435
rect 850 5385 900 5415
rect 850 5365 865 5385
rect 885 5365 900 5385
rect 850 5335 900 5365
rect 850 5315 865 5335
rect 885 5315 900 5335
rect 850 5285 900 5315
rect 850 5265 865 5285
rect 885 5265 900 5285
rect 850 5235 900 5265
rect 850 5215 865 5235
rect 885 5215 900 5235
rect 850 5185 900 5215
rect 850 5165 865 5185
rect 885 5165 900 5185
rect 850 5135 900 5165
rect 850 5115 865 5135
rect 885 5115 900 5135
rect 850 5085 900 5115
rect 850 5065 865 5085
rect 885 5065 900 5085
rect 850 5035 900 5065
rect 850 5015 865 5035
rect 885 5015 900 5035
rect 850 5000 900 5015
rect 1000 5485 1050 5500
rect 1000 5465 1015 5485
rect 1035 5465 1050 5485
rect 1000 5435 1050 5465
rect 1000 5415 1015 5435
rect 1035 5415 1050 5435
rect 1000 5385 1050 5415
rect 1000 5365 1015 5385
rect 1035 5365 1050 5385
rect 1000 5335 1050 5365
rect 1000 5315 1015 5335
rect 1035 5315 1050 5335
rect 1000 5285 1050 5315
rect 1000 5265 1015 5285
rect 1035 5265 1050 5285
rect 1000 5235 1050 5265
rect 1000 5215 1015 5235
rect 1035 5215 1050 5235
rect 1000 5185 1050 5215
rect 1000 5165 1015 5185
rect 1035 5165 1050 5185
rect 1000 5135 1050 5165
rect 1000 5115 1015 5135
rect 1035 5115 1050 5135
rect 1000 5085 1050 5115
rect 1000 5065 1015 5085
rect 1035 5065 1050 5085
rect 1000 5035 1050 5065
rect 1000 5015 1015 5035
rect 1035 5015 1050 5035
rect 1000 5000 1050 5015
rect 1150 5485 1200 5500
rect 1150 5465 1165 5485
rect 1185 5465 1200 5485
rect 1150 5435 1200 5465
rect 1150 5415 1165 5435
rect 1185 5415 1200 5435
rect 1150 5385 1200 5415
rect 1150 5365 1165 5385
rect 1185 5365 1200 5385
rect 1150 5335 1200 5365
rect 1150 5315 1165 5335
rect 1185 5315 1200 5335
rect 1150 5285 1200 5315
rect 1150 5265 1165 5285
rect 1185 5265 1200 5285
rect 1150 5235 1200 5265
rect 1150 5215 1165 5235
rect 1185 5215 1200 5235
rect 1150 5185 1200 5215
rect 1150 5165 1165 5185
rect 1185 5165 1200 5185
rect 1150 5135 1200 5165
rect 1150 5115 1165 5135
rect 1185 5115 1200 5135
rect 1150 5085 1200 5115
rect 1150 5065 1165 5085
rect 1185 5065 1200 5085
rect 1150 5035 1200 5065
rect 1150 5015 1165 5035
rect 1185 5015 1200 5035
rect 1150 5000 1200 5015
rect 1300 5485 1350 5500
rect 1300 5465 1315 5485
rect 1335 5465 1350 5485
rect 1300 5435 1350 5465
rect 1300 5415 1315 5435
rect 1335 5415 1350 5435
rect 1300 5385 1350 5415
rect 1300 5365 1315 5385
rect 1335 5365 1350 5385
rect 1300 5335 1350 5365
rect 1300 5315 1315 5335
rect 1335 5315 1350 5335
rect 1300 5285 1350 5315
rect 1300 5265 1315 5285
rect 1335 5265 1350 5285
rect 1300 5235 1350 5265
rect 1300 5215 1315 5235
rect 1335 5215 1350 5235
rect 1300 5185 1350 5215
rect 1300 5165 1315 5185
rect 1335 5165 1350 5185
rect 1300 5135 1350 5165
rect 1300 5115 1315 5135
rect 1335 5115 1350 5135
rect 1300 5085 1350 5115
rect 1300 5065 1315 5085
rect 1335 5065 1350 5085
rect 1300 5035 1350 5065
rect 1300 5015 1315 5035
rect 1335 5015 1350 5035
rect 1300 5000 1350 5015
rect 1450 5485 1500 5500
rect 1450 5465 1465 5485
rect 1485 5465 1500 5485
rect 1450 5435 1500 5465
rect 1450 5415 1465 5435
rect 1485 5415 1500 5435
rect 1450 5385 1500 5415
rect 1450 5365 1465 5385
rect 1485 5365 1500 5385
rect 1450 5335 1500 5365
rect 1450 5315 1465 5335
rect 1485 5315 1500 5335
rect 1450 5285 1500 5315
rect 1450 5265 1465 5285
rect 1485 5265 1500 5285
rect 1450 5235 1500 5265
rect 1450 5215 1465 5235
rect 1485 5215 1500 5235
rect 1450 5185 1500 5215
rect 1450 5165 1465 5185
rect 1485 5165 1500 5185
rect 1450 5135 1500 5165
rect 1450 5115 1465 5135
rect 1485 5115 1500 5135
rect 1450 5085 1500 5115
rect 1450 5065 1465 5085
rect 1485 5065 1500 5085
rect 1450 5035 1500 5065
rect 1450 5015 1465 5035
rect 1485 5015 1500 5035
rect 1450 5000 1500 5015
rect 1600 5485 1650 5500
rect 1600 5465 1615 5485
rect 1635 5465 1650 5485
rect 1600 5435 1650 5465
rect 1600 5415 1615 5435
rect 1635 5415 1650 5435
rect 1600 5385 1650 5415
rect 1600 5365 1615 5385
rect 1635 5365 1650 5385
rect 1600 5335 1650 5365
rect 1600 5315 1615 5335
rect 1635 5315 1650 5335
rect 1600 5285 1650 5315
rect 1600 5265 1615 5285
rect 1635 5265 1650 5285
rect 1600 5235 1650 5265
rect 1600 5215 1615 5235
rect 1635 5215 1650 5235
rect 1600 5185 1650 5215
rect 1600 5165 1615 5185
rect 1635 5165 1650 5185
rect 1600 5135 1650 5165
rect 1600 5115 1615 5135
rect 1635 5115 1650 5135
rect 1600 5085 1650 5115
rect 1600 5065 1615 5085
rect 1635 5065 1650 5085
rect 1600 5035 1650 5065
rect 1600 5015 1615 5035
rect 1635 5015 1650 5035
rect 1600 5000 1650 5015
rect 1750 5485 1800 5500
rect 1750 5465 1765 5485
rect 1785 5465 1800 5485
rect 1750 5435 1800 5465
rect 1750 5415 1765 5435
rect 1785 5415 1800 5435
rect 1750 5385 1800 5415
rect 1750 5365 1765 5385
rect 1785 5365 1800 5385
rect 1750 5335 1800 5365
rect 1750 5315 1765 5335
rect 1785 5315 1800 5335
rect 1750 5285 1800 5315
rect 1750 5265 1765 5285
rect 1785 5265 1800 5285
rect 1750 5235 1800 5265
rect 1750 5215 1765 5235
rect 1785 5215 1800 5235
rect 1750 5185 1800 5215
rect 1750 5165 1765 5185
rect 1785 5165 1800 5185
rect 1750 5135 1800 5165
rect 1750 5115 1765 5135
rect 1785 5115 1800 5135
rect 1750 5085 1800 5115
rect 1750 5065 1765 5085
rect 1785 5065 1800 5085
rect 1750 5035 1800 5065
rect 1750 5015 1765 5035
rect 1785 5015 1800 5035
rect 1750 5000 1800 5015
rect 1900 5485 1950 5500
rect 1900 5465 1915 5485
rect 1935 5465 1950 5485
rect 1900 5435 1950 5465
rect 1900 5415 1915 5435
rect 1935 5415 1950 5435
rect 1900 5385 1950 5415
rect 1900 5365 1915 5385
rect 1935 5365 1950 5385
rect 1900 5335 1950 5365
rect 1900 5315 1915 5335
rect 1935 5315 1950 5335
rect 1900 5285 1950 5315
rect 1900 5265 1915 5285
rect 1935 5265 1950 5285
rect 1900 5235 1950 5265
rect 1900 5215 1915 5235
rect 1935 5215 1950 5235
rect 1900 5185 1950 5215
rect 1900 5165 1915 5185
rect 1935 5165 1950 5185
rect 1900 5135 1950 5165
rect 1900 5115 1915 5135
rect 1935 5115 1950 5135
rect 1900 5085 1950 5115
rect 1900 5065 1915 5085
rect 1935 5065 1950 5085
rect 1900 5035 1950 5065
rect 1900 5015 1915 5035
rect 1935 5015 1950 5035
rect 1900 5000 1950 5015
rect 2050 5485 2100 5500
rect 2050 5465 2065 5485
rect 2085 5465 2100 5485
rect 2050 5435 2100 5465
rect 2050 5415 2065 5435
rect 2085 5415 2100 5435
rect 2050 5385 2100 5415
rect 2050 5365 2065 5385
rect 2085 5365 2100 5385
rect 2050 5335 2100 5365
rect 2050 5315 2065 5335
rect 2085 5315 2100 5335
rect 2050 5285 2100 5315
rect 2050 5265 2065 5285
rect 2085 5265 2100 5285
rect 2050 5235 2100 5265
rect 2050 5215 2065 5235
rect 2085 5215 2100 5235
rect 2050 5185 2100 5215
rect 2050 5165 2065 5185
rect 2085 5165 2100 5185
rect 2050 5135 2100 5165
rect 2050 5115 2065 5135
rect 2085 5115 2100 5135
rect 2050 5085 2100 5115
rect 2050 5065 2065 5085
rect 2085 5065 2100 5085
rect 2050 5035 2100 5065
rect 2050 5015 2065 5035
rect 2085 5015 2100 5035
rect 2050 5000 2100 5015
rect 2200 5485 2250 5500
rect 2200 5465 2215 5485
rect 2235 5465 2250 5485
rect 2200 5435 2250 5465
rect 2200 5415 2215 5435
rect 2235 5415 2250 5435
rect 2200 5385 2250 5415
rect 2200 5365 2215 5385
rect 2235 5365 2250 5385
rect 2200 5335 2250 5365
rect 2200 5315 2215 5335
rect 2235 5315 2250 5335
rect 2200 5285 2250 5315
rect 2200 5265 2215 5285
rect 2235 5265 2250 5285
rect 2200 5235 2250 5265
rect 2200 5215 2215 5235
rect 2235 5215 2250 5235
rect 2200 5185 2250 5215
rect 2200 5165 2215 5185
rect 2235 5165 2250 5185
rect 2200 5135 2250 5165
rect 2200 5115 2215 5135
rect 2235 5115 2250 5135
rect 2200 5085 2250 5115
rect 2200 5065 2215 5085
rect 2235 5065 2250 5085
rect 2200 5035 2250 5065
rect 2200 5015 2215 5035
rect 2235 5015 2250 5035
rect 2200 5000 2250 5015
rect 2350 5485 2400 5500
rect 2350 5465 2365 5485
rect 2385 5465 2400 5485
rect 2350 5435 2400 5465
rect 2350 5415 2365 5435
rect 2385 5415 2400 5435
rect 2350 5385 2400 5415
rect 2350 5365 2365 5385
rect 2385 5365 2400 5385
rect 2350 5335 2400 5365
rect 2350 5315 2365 5335
rect 2385 5315 2400 5335
rect 2350 5285 2400 5315
rect 2350 5265 2365 5285
rect 2385 5265 2400 5285
rect 2350 5235 2400 5265
rect 2350 5215 2365 5235
rect 2385 5215 2400 5235
rect 2350 5185 2400 5215
rect 2350 5165 2365 5185
rect 2385 5165 2400 5185
rect 2350 5135 2400 5165
rect 2350 5115 2365 5135
rect 2385 5115 2400 5135
rect 2350 5085 2400 5115
rect 2350 5065 2365 5085
rect 2385 5065 2400 5085
rect 2350 5035 2400 5065
rect 2350 5015 2365 5035
rect 2385 5015 2400 5035
rect 2350 5000 2400 5015
rect 2500 5485 2550 5500
rect 2500 5465 2515 5485
rect 2535 5465 2550 5485
rect 2500 5435 2550 5465
rect 2500 5415 2515 5435
rect 2535 5415 2550 5435
rect 2500 5385 2550 5415
rect 2500 5365 2515 5385
rect 2535 5365 2550 5385
rect 2500 5335 2550 5365
rect 2500 5315 2515 5335
rect 2535 5315 2550 5335
rect 2500 5285 2550 5315
rect 2500 5265 2515 5285
rect 2535 5265 2550 5285
rect 2500 5235 2550 5265
rect 2500 5215 2515 5235
rect 2535 5215 2550 5235
rect 2500 5185 2550 5215
rect 2500 5165 2515 5185
rect 2535 5165 2550 5185
rect 2500 5135 2550 5165
rect 2500 5115 2515 5135
rect 2535 5115 2550 5135
rect 2500 5085 2550 5115
rect 2500 5065 2515 5085
rect 2535 5065 2550 5085
rect 2500 5035 2550 5065
rect 2500 5015 2515 5035
rect 2535 5015 2550 5035
rect 2500 5000 2550 5015
rect 2650 5485 2700 5500
rect 2650 5465 2665 5485
rect 2685 5465 2700 5485
rect 2650 5435 2700 5465
rect 2650 5415 2665 5435
rect 2685 5415 2700 5435
rect 2650 5385 2700 5415
rect 2650 5365 2665 5385
rect 2685 5365 2700 5385
rect 2650 5335 2700 5365
rect 2650 5315 2665 5335
rect 2685 5315 2700 5335
rect 2650 5285 2700 5315
rect 2650 5265 2665 5285
rect 2685 5265 2700 5285
rect 2650 5235 2700 5265
rect 2650 5215 2665 5235
rect 2685 5215 2700 5235
rect 2650 5185 2700 5215
rect 2650 5165 2665 5185
rect 2685 5165 2700 5185
rect 2650 5135 2700 5165
rect 2650 5115 2665 5135
rect 2685 5115 2700 5135
rect 2650 5085 2700 5115
rect 2650 5065 2665 5085
rect 2685 5065 2700 5085
rect 2650 5035 2700 5065
rect 2650 5015 2665 5035
rect 2685 5015 2700 5035
rect 2650 5000 2700 5015
rect 2800 5485 2850 5500
rect 2800 5465 2815 5485
rect 2835 5465 2850 5485
rect 2800 5435 2850 5465
rect 2800 5415 2815 5435
rect 2835 5415 2850 5435
rect 2800 5385 2850 5415
rect 2800 5365 2815 5385
rect 2835 5365 2850 5385
rect 2800 5335 2850 5365
rect 2800 5315 2815 5335
rect 2835 5315 2850 5335
rect 2800 5285 2850 5315
rect 2800 5265 2815 5285
rect 2835 5265 2850 5285
rect 2800 5235 2850 5265
rect 2800 5215 2815 5235
rect 2835 5215 2850 5235
rect 2800 5185 2850 5215
rect 2800 5165 2815 5185
rect 2835 5165 2850 5185
rect 2800 5135 2850 5165
rect 2800 5115 2815 5135
rect 2835 5115 2850 5135
rect 2800 5085 2850 5115
rect 2800 5065 2815 5085
rect 2835 5065 2850 5085
rect 2800 5035 2850 5065
rect 2800 5015 2815 5035
rect 2835 5015 2850 5035
rect 2800 5000 2850 5015
rect 2950 5485 3000 5500
rect 2950 5465 2965 5485
rect 2985 5465 3000 5485
rect 2950 5435 3000 5465
rect 2950 5415 2965 5435
rect 2985 5415 3000 5435
rect 2950 5385 3000 5415
rect 2950 5365 2965 5385
rect 2985 5365 3000 5385
rect 2950 5335 3000 5365
rect 2950 5315 2965 5335
rect 2985 5315 3000 5335
rect 2950 5285 3000 5315
rect 2950 5265 2965 5285
rect 2985 5265 3000 5285
rect 2950 5235 3000 5265
rect 2950 5215 2965 5235
rect 2985 5215 3000 5235
rect 2950 5185 3000 5215
rect 2950 5165 2965 5185
rect 2985 5165 3000 5185
rect 2950 5135 3000 5165
rect 2950 5115 2965 5135
rect 2985 5115 3000 5135
rect 2950 5085 3000 5115
rect 2950 5065 2965 5085
rect 2985 5065 3000 5085
rect 2950 5035 3000 5065
rect 2950 5015 2965 5035
rect 2985 5015 3000 5035
rect 2950 5000 3000 5015
rect 3100 5485 3150 5500
rect 3100 5465 3115 5485
rect 3135 5465 3150 5485
rect 3100 5435 3150 5465
rect 3100 5415 3115 5435
rect 3135 5415 3150 5435
rect 3100 5385 3150 5415
rect 3100 5365 3115 5385
rect 3135 5365 3150 5385
rect 3100 5335 3150 5365
rect 3100 5315 3115 5335
rect 3135 5315 3150 5335
rect 3100 5285 3150 5315
rect 3100 5265 3115 5285
rect 3135 5265 3150 5285
rect 3100 5235 3150 5265
rect 3100 5215 3115 5235
rect 3135 5215 3150 5235
rect 3100 5185 3150 5215
rect 3100 5165 3115 5185
rect 3135 5165 3150 5185
rect 3100 5135 3150 5165
rect 3100 5115 3115 5135
rect 3135 5115 3150 5135
rect 3100 5085 3150 5115
rect 3100 5065 3115 5085
rect 3135 5065 3150 5085
rect 3100 5035 3150 5065
rect 3100 5015 3115 5035
rect 3135 5015 3150 5035
rect 3100 5000 3150 5015
rect 3250 5485 3300 5500
rect 3250 5465 3265 5485
rect 3285 5465 3300 5485
rect 3250 5435 3300 5465
rect 3250 5415 3265 5435
rect 3285 5415 3300 5435
rect 3250 5385 3300 5415
rect 3250 5365 3265 5385
rect 3285 5365 3300 5385
rect 3250 5335 3300 5365
rect 3250 5315 3265 5335
rect 3285 5315 3300 5335
rect 3250 5285 3300 5315
rect 3250 5265 3265 5285
rect 3285 5265 3300 5285
rect 3250 5235 3300 5265
rect 3250 5215 3265 5235
rect 3285 5215 3300 5235
rect 3250 5185 3300 5215
rect 3250 5165 3265 5185
rect 3285 5165 3300 5185
rect 3250 5135 3300 5165
rect 3250 5115 3265 5135
rect 3285 5115 3300 5135
rect 3250 5085 3300 5115
rect 3250 5065 3265 5085
rect 3285 5065 3300 5085
rect 3250 5035 3300 5065
rect 3250 5015 3265 5035
rect 3285 5015 3300 5035
rect 3250 5000 3300 5015
rect 3400 5485 3450 5500
rect 3400 5465 3415 5485
rect 3435 5465 3450 5485
rect 3400 5435 3450 5465
rect 3400 5415 3415 5435
rect 3435 5415 3450 5435
rect 3400 5385 3450 5415
rect 3400 5365 3415 5385
rect 3435 5365 3450 5385
rect 3400 5335 3450 5365
rect 3400 5315 3415 5335
rect 3435 5315 3450 5335
rect 3400 5285 3450 5315
rect 3400 5265 3415 5285
rect 3435 5265 3450 5285
rect 3400 5235 3450 5265
rect 3400 5215 3415 5235
rect 3435 5215 3450 5235
rect 3400 5185 3450 5215
rect 3400 5165 3415 5185
rect 3435 5165 3450 5185
rect 3400 5135 3450 5165
rect 3400 5115 3415 5135
rect 3435 5115 3450 5135
rect 3400 5085 3450 5115
rect 3400 5065 3415 5085
rect 3435 5065 3450 5085
rect 3400 5035 3450 5065
rect 3400 5015 3415 5035
rect 3435 5015 3450 5035
rect 3400 5000 3450 5015
rect 3550 5485 3600 5500
rect 3550 5465 3565 5485
rect 3585 5465 3600 5485
rect 3550 5435 3600 5465
rect 3550 5415 3565 5435
rect 3585 5415 3600 5435
rect 3550 5385 3600 5415
rect 3550 5365 3565 5385
rect 3585 5365 3600 5385
rect 3550 5335 3600 5365
rect 3550 5315 3565 5335
rect 3585 5315 3600 5335
rect 3550 5285 3600 5315
rect 3550 5265 3565 5285
rect 3585 5265 3600 5285
rect 3550 5235 3600 5265
rect 3550 5215 3565 5235
rect 3585 5215 3600 5235
rect 3550 5185 3600 5215
rect 3550 5165 3565 5185
rect 3585 5165 3600 5185
rect 3550 5135 3600 5165
rect 3550 5115 3565 5135
rect 3585 5115 3600 5135
rect 3550 5085 3600 5115
rect 3550 5065 3565 5085
rect 3585 5065 3600 5085
rect 3550 5035 3600 5065
rect 3550 5015 3565 5035
rect 3585 5015 3600 5035
rect 3550 5000 3600 5015
rect 4150 5485 4200 5500
rect 4150 5465 4165 5485
rect 4185 5465 4200 5485
rect 4150 5435 4200 5465
rect 4150 5415 4165 5435
rect 4185 5415 4200 5435
rect 4150 5385 4200 5415
rect 4150 5365 4165 5385
rect 4185 5365 4200 5385
rect 4150 5335 4200 5365
rect 4150 5315 4165 5335
rect 4185 5315 4200 5335
rect 4150 5285 4200 5315
rect 4150 5265 4165 5285
rect 4185 5265 4200 5285
rect 4150 5235 4200 5265
rect 4150 5215 4165 5235
rect 4185 5215 4200 5235
rect 4150 5185 4200 5215
rect 4150 5165 4165 5185
rect 4185 5165 4200 5185
rect 4150 5135 4200 5165
rect 4150 5115 4165 5135
rect 4185 5115 4200 5135
rect 4150 5085 4200 5115
rect 4150 5065 4165 5085
rect 4185 5065 4200 5085
rect 4150 5035 4200 5065
rect 4150 5015 4165 5035
rect 4185 5015 4200 5035
rect 4150 5000 4200 5015
rect 4750 5485 4800 5500
rect 4750 5465 4765 5485
rect 4785 5465 4800 5485
rect 4750 5435 4800 5465
rect 4750 5415 4765 5435
rect 4785 5415 4800 5435
rect 4750 5385 4800 5415
rect 4750 5365 4765 5385
rect 4785 5365 4800 5385
rect 4750 5335 4800 5365
rect 4750 5315 4765 5335
rect 4785 5315 4800 5335
rect 4750 5285 4800 5315
rect 4750 5265 4765 5285
rect 4785 5265 4800 5285
rect 4750 5235 4800 5265
rect 4750 5215 4765 5235
rect 4785 5215 4800 5235
rect 4750 5185 4800 5215
rect 4750 5165 4765 5185
rect 4785 5165 4800 5185
rect 4750 5135 4800 5165
rect 4750 5115 4765 5135
rect 4785 5115 4800 5135
rect 4750 5085 4800 5115
rect 4750 5065 4765 5085
rect 4785 5065 4800 5085
rect 4750 5035 4800 5065
rect 4750 5015 4765 5035
rect 4785 5015 4800 5035
rect 4750 5000 4800 5015
rect 4900 5485 4950 5500
rect 4900 5465 4915 5485
rect 4935 5465 4950 5485
rect 4900 5435 4950 5465
rect 4900 5415 4915 5435
rect 4935 5415 4950 5435
rect 4900 5385 4950 5415
rect 4900 5365 4915 5385
rect 4935 5365 4950 5385
rect 4900 5335 4950 5365
rect 4900 5315 4915 5335
rect 4935 5315 4950 5335
rect 4900 5285 4950 5315
rect 4900 5265 4915 5285
rect 4935 5265 4950 5285
rect 4900 5235 4950 5265
rect 4900 5215 4915 5235
rect 4935 5215 4950 5235
rect 4900 5185 4950 5215
rect 4900 5165 4915 5185
rect 4935 5165 4950 5185
rect 4900 5135 4950 5165
rect 4900 5115 4915 5135
rect 4935 5115 4950 5135
rect 4900 5085 4950 5115
rect 4900 5065 4915 5085
rect 4935 5065 4950 5085
rect 4900 5035 4950 5065
rect 4900 5015 4915 5035
rect 4935 5015 4950 5035
rect 4900 5000 4950 5015
rect 5050 5485 5100 5500
rect 5050 5465 5065 5485
rect 5085 5465 5100 5485
rect 5050 5435 5100 5465
rect 5050 5415 5065 5435
rect 5085 5415 5100 5435
rect 5050 5385 5100 5415
rect 5050 5365 5065 5385
rect 5085 5365 5100 5385
rect 5050 5335 5100 5365
rect 5050 5315 5065 5335
rect 5085 5315 5100 5335
rect 5050 5285 5100 5315
rect 5050 5265 5065 5285
rect 5085 5265 5100 5285
rect 5050 5235 5100 5265
rect 5050 5215 5065 5235
rect 5085 5215 5100 5235
rect 5050 5185 5100 5215
rect 5050 5165 5065 5185
rect 5085 5165 5100 5185
rect 5050 5135 5100 5165
rect 5050 5115 5065 5135
rect 5085 5115 5100 5135
rect 5050 5085 5100 5115
rect 5050 5065 5065 5085
rect 5085 5065 5100 5085
rect 5050 5035 5100 5065
rect 5050 5015 5065 5035
rect 5085 5015 5100 5035
rect 5050 5000 5100 5015
rect 5200 5485 5250 5500
rect 5200 5465 5215 5485
rect 5235 5465 5250 5485
rect 5200 5435 5250 5465
rect 5200 5415 5215 5435
rect 5235 5415 5250 5435
rect 5200 5385 5250 5415
rect 5200 5365 5215 5385
rect 5235 5365 5250 5385
rect 5200 5335 5250 5365
rect 5200 5315 5215 5335
rect 5235 5315 5250 5335
rect 5200 5285 5250 5315
rect 5200 5265 5215 5285
rect 5235 5265 5250 5285
rect 5200 5235 5250 5265
rect 5200 5215 5215 5235
rect 5235 5215 5250 5235
rect 5200 5185 5250 5215
rect 5200 5165 5215 5185
rect 5235 5165 5250 5185
rect 5200 5135 5250 5165
rect 5200 5115 5215 5135
rect 5235 5115 5250 5135
rect 5200 5085 5250 5115
rect 5200 5065 5215 5085
rect 5235 5065 5250 5085
rect 5200 5035 5250 5065
rect 5200 5015 5215 5035
rect 5235 5015 5250 5035
rect 5200 5000 5250 5015
rect 5350 5485 5400 5500
rect 5350 5465 5365 5485
rect 5385 5465 5400 5485
rect 5350 5435 5400 5465
rect 5350 5415 5365 5435
rect 5385 5415 5400 5435
rect 5350 5385 5400 5415
rect 5350 5365 5365 5385
rect 5385 5365 5400 5385
rect 5350 5335 5400 5365
rect 5350 5315 5365 5335
rect 5385 5315 5400 5335
rect 5350 5285 5400 5315
rect 5350 5265 5365 5285
rect 5385 5265 5400 5285
rect 5350 5235 5400 5265
rect 5350 5215 5365 5235
rect 5385 5215 5400 5235
rect 5350 5185 5400 5215
rect 5350 5165 5365 5185
rect 5385 5165 5400 5185
rect 5350 5135 5400 5165
rect 5350 5115 5365 5135
rect 5385 5115 5400 5135
rect 5350 5085 5400 5115
rect 5350 5065 5365 5085
rect 5385 5065 5400 5085
rect 5350 5035 5400 5065
rect 5350 5015 5365 5035
rect 5385 5015 5400 5035
rect 5350 5000 5400 5015
rect 5500 5485 5550 5500
rect 5500 5465 5515 5485
rect 5535 5465 5550 5485
rect 5500 5435 5550 5465
rect 5500 5415 5515 5435
rect 5535 5415 5550 5435
rect 5500 5385 5550 5415
rect 5500 5365 5515 5385
rect 5535 5365 5550 5385
rect 5500 5335 5550 5365
rect 5500 5315 5515 5335
rect 5535 5315 5550 5335
rect 5500 5285 5550 5315
rect 5500 5265 5515 5285
rect 5535 5265 5550 5285
rect 5500 5235 5550 5265
rect 5500 5215 5515 5235
rect 5535 5215 5550 5235
rect 5500 5185 5550 5215
rect 5500 5165 5515 5185
rect 5535 5165 5550 5185
rect 5500 5135 5550 5165
rect 5500 5115 5515 5135
rect 5535 5115 5550 5135
rect 5500 5085 5550 5115
rect 5500 5065 5515 5085
rect 5535 5065 5550 5085
rect 5500 5035 5550 5065
rect 5500 5015 5515 5035
rect 5535 5015 5550 5035
rect 5500 5000 5550 5015
rect 5650 5485 5700 5500
rect 5650 5465 5665 5485
rect 5685 5465 5700 5485
rect 5650 5435 5700 5465
rect 5650 5415 5665 5435
rect 5685 5415 5700 5435
rect 5650 5385 5700 5415
rect 5650 5365 5665 5385
rect 5685 5365 5700 5385
rect 5650 5335 5700 5365
rect 5650 5315 5665 5335
rect 5685 5315 5700 5335
rect 5650 5285 5700 5315
rect 5650 5265 5665 5285
rect 5685 5265 5700 5285
rect 5650 5235 5700 5265
rect 5650 5215 5665 5235
rect 5685 5215 5700 5235
rect 5650 5185 5700 5215
rect 5650 5165 5665 5185
rect 5685 5165 5700 5185
rect 5650 5135 5700 5165
rect 5650 5115 5665 5135
rect 5685 5115 5700 5135
rect 5650 5085 5700 5115
rect 5650 5065 5665 5085
rect 5685 5065 5700 5085
rect 5650 5035 5700 5065
rect 5650 5015 5665 5035
rect 5685 5015 5700 5035
rect 5650 5000 5700 5015
rect 5800 5485 5850 5500
rect 5800 5465 5815 5485
rect 5835 5465 5850 5485
rect 5800 5435 5850 5465
rect 5800 5415 5815 5435
rect 5835 5415 5850 5435
rect 5800 5385 5850 5415
rect 5800 5365 5815 5385
rect 5835 5365 5850 5385
rect 5800 5335 5850 5365
rect 5800 5315 5815 5335
rect 5835 5315 5850 5335
rect 5800 5285 5850 5315
rect 5800 5265 5815 5285
rect 5835 5265 5850 5285
rect 5800 5235 5850 5265
rect 5800 5215 5815 5235
rect 5835 5215 5850 5235
rect 5800 5185 5850 5215
rect 5800 5165 5815 5185
rect 5835 5165 5850 5185
rect 5800 5135 5850 5165
rect 5800 5115 5815 5135
rect 5835 5115 5850 5135
rect 5800 5085 5850 5115
rect 5800 5065 5815 5085
rect 5835 5065 5850 5085
rect 5800 5035 5850 5065
rect 5800 5015 5815 5035
rect 5835 5015 5850 5035
rect 5800 5000 5850 5015
rect 5950 5485 6000 5500
rect 5950 5465 5965 5485
rect 5985 5465 6000 5485
rect 5950 5435 6000 5465
rect 5950 5415 5965 5435
rect 5985 5415 6000 5435
rect 5950 5385 6000 5415
rect 5950 5365 5965 5385
rect 5985 5365 6000 5385
rect 5950 5335 6000 5365
rect 5950 5315 5965 5335
rect 5985 5315 6000 5335
rect 5950 5285 6000 5315
rect 5950 5265 5965 5285
rect 5985 5265 6000 5285
rect 5950 5235 6000 5265
rect 5950 5215 5965 5235
rect 5985 5215 6000 5235
rect 5950 5185 6000 5215
rect 5950 5165 5965 5185
rect 5985 5165 6000 5185
rect 5950 5135 6000 5165
rect 5950 5115 5965 5135
rect 5985 5115 6000 5135
rect 5950 5085 6000 5115
rect 5950 5065 5965 5085
rect 5985 5065 6000 5085
rect 5950 5035 6000 5065
rect 5950 5015 5965 5035
rect 5985 5015 6000 5035
rect 5950 5000 6000 5015
rect 6100 5485 6150 5500
rect 6100 5465 6115 5485
rect 6135 5465 6150 5485
rect 6100 5435 6150 5465
rect 6100 5415 6115 5435
rect 6135 5415 6150 5435
rect 6100 5385 6150 5415
rect 6100 5365 6115 5385
rect 6135 5365 6150 5385
rect 6100 5335 6150 5365
rect 6100 5315 6115 5335
rect 6135 5315 6150 5335
rect 6100 5285 6150 5315
rect 6100 5265 6115 5285
rect 6135 5265 6150 5285
rect 6100 5235 6150 5265
rect 6100 5215 6115 5235
rect 6135 5215 6150 5235
rect 6100 5185 6150 5215
rect 6100 5165 6115 5185
rect 6135 5165 6150 5185
rect 6100 5135 6150 5165
rect 6100 5115 6115 5135
rect 6135 5115 6150 5135
rect 6100 5085 6150 5115
rect 6100 5065 6115 5085
rect 6135 5065 6150 5085
rect 6100 5035 6150 5065
rect 6100 5015 6115 5035
rect 6135 5015 6150 5035
rect 6100 5000 6150 5015
rect 6250 5485 6300 5500
rect 6250 5465 6265 5485
rect 6285 5465 6300 5485
rect 6250 5435 6300 5465
rect 6250 5415 6265 5435
rect 6285 5415 6300 5435
rect 6250 5385 6300 5415
rect 6250 5365 6265 5385
rect 6285 5365 6300 5385
rect 6250 5335 6300 5365
rect 6250 5315 6265 5335
rect 6285 5315 6300 5335
rect 6250 5285 6300 5315
rect 6250 5265 6265 5285
rect 6285 5265 6300 5285
rect 6250 5235 6300 5265
rect 6250 5215 6265 5235
rect 6285 5215 6300 5235
rect 6250 5185 6300 5215
rect 6250 5165 6265 5185
rect 6285 5165 6300 5185
rect 6250 5135 6300 5165
rect 6250 5115 6265 5135
rect 6285 5115 6300 5135
rect 6250 5085 6300 5115
rect 6250 5065 6265 5085
rect 6285 5065 6300 5085
rect 6250 5035 6300 5065
rect 6250 5015 6265 5035
rect 6285 5015 6300 5035
rect 6250 5000 6300 5015
rect 6400 5485 6450 5500
rect 6400 5465 6415 5485
rect 6435 5465 6450 5485
rect 6400 5435 6450 5465
rect 6400 5415 6415 5435
rect 6435 5415 6450 5435
rect 6400 5385 6450 5415
rect 6400 5365 6415 5385
rect 6435 5365 6450 5385
rect 6400 5335 6450 5365
rect 6400 5315 6415 5335
rect 6435 5315 6450 5335
rect 6400 5285 6450 5315
rect 6400 5265 6415 5285
rect 6435 5265 6450 5285
rect 6400 5235 6450 5265
rect 6400 5215 6415 5235
rect 6435 5215 6450 5235
rect 6400 5185 6450 5215
rect 6400 5165 6415 5185
rect 6435 5165 6450 5185
rect 6400 5135 6450 5165
rect 6400 5115 6415 5135
rect 6435 5115 6450 5135
rect 6400 5085 6450 5115
rect 6400 5065 6415 5085
rect 6435 5065 6450 5085
rect 6400 5035 6450 5065
rect 6400 5015 6415 5035
rect 6435 5015 6450 5035
rect 6400 5000 6450 5015
rect 6550 5485 6600 5500
rect 6550 5465 6565 5485
rect 6585 5465 6600 5485
rect 6550 5435 6600 5465
rect 6550 5415 6565 5435
rect 6585 5415 6600 5435
rect 6550 5385 6600 5415
rect 6550 5365 6565 5385
rect 6585 5365 6600 5385
rect 6550 5335 6600 5365
rect 6550 5315 6565 5335
rect 6585 5315 6600 5335
rect 6550 5285 6600 5315
rect 6550 5265 6565 5285
rect 6585 5265 6600 5285
rect 6550 5235 6600 5265
rect 6550 5215 6565 5235
rect 6585 5215 6600 5235
rect 6550 5185 6600 5215
rect 6550 5165 6565 5185
rect 6585 5165 6600 5185
rect 6550 5135 6600 5165
rect 6550 5115 6565 5135
rect 6585 5115 6600 5135
rect 6550 5085 6600 5115
rect 6550 5065 6565 5085
rect 6585 5065 6600 5085
rect 6550 5035 6600 5065
rect 6550 5015 6565 5035
rect 6585 5015 6600 5035
rect 6550 5000 6600 5015
rect 6700 5485 6750 5500
rect 6700 5465 6715 5485
rect 6735 5465 6750 5485
rect 6700 5435 6750 5465
rect 6700 5415 6715 5435
rect 6735 5415 6750 5435
rect 6700 5385 6750 5415
rect 6700 5365 6715 5385
rect 6735 5365 6750 5385
rect 6700 5335 6750 5365
rect 6700 5315 6715 5335
rect 6735 5315 6750 5335
rect 6700 5285 6750 5315
rect 6700 5265 6715 5285
rect 6735 5265 6750 5285
rect 6700 5235 6750 5265
rect 6700 5215 6715 5235
rect 6735 5215 6750 5235
rect 6700 5185 6750 5215
rect 6700 5165 6715 5185
rect 6735 5165 6750 5185
rect 6700 5135 6750 5165
rect 6700 5115 6715 5135
rect 6735 5115 6750 5135
rect 6700 5085 6750 5115
rect 6700 5065 6715 5085
rect 6735 5065 6750 5085
rect 6700 5035 6750 5065
rect 6700 5015 6715 5035
rect 6735 5015 6750 5035
rect 6700 5000 6750 5015
rect 6850 5485 6900 5500
rect 6850 5465 6865 5485
rect 6885 5465 6900 5485
rect 6850 5435 6900 5465
rect 6850 5415 6865 5435
rect 6885 5415 6900 5435
rect 6850 5385 6900 5415
rect 6850 5365 6865 5385
rect 6885 5365 6900 5385
rect 6850 5335 6900 5365
rect 6850 5315 6865 5335
rect 6885 5315 6900 5335
rect 6850 5285 6900 5315
rect 6850 5265 6865 5285
rect 6885 5265 6900 5285
rect 6850 5235 6900 5265
rect 6850 5215 6865 5235
rect 6885 5215 6900 5235
rect 6850 5185 6900 5215
rect 6850 5165 6865 5185
rect 6885 5165 6900 5185
rect 6850 5135 6900 5165
rect 6850 5115 6865 5135
rect 6885 5115 6900 5135
rect 6850 5085 6900 5115
rect 6850 5065 6865 5085
rect 6885 5065 6900 5085
rect 6850 5035 6900 5065
rect 6850 5015 6865 5035
rect 6885 5015 6900 5035
rect 6850 5000 6900 5015
rect 7000 5485 7050 5500
rect 7000 5465 7015 5485
rect 7035 5465 7050 5485
rect 7000 5435 7050 5465
rect 7000 5415 7015 5435
rect 7035 5415 7050 5435
rect 7000 5385 7050 5415
rect 7000 5365 7015 5385
rect 7035 5365 7050 5385
rect 7000 5335 7050 5365
rect 7000 5315 7015 5335
rect 7035 5315 7050 5335
rect 7000 5285 7050 5315
rect 7000 5265 7015 5285
rect 7035 5265 7050 5285
rect 7000 5235 7050 5265
rect 7000 5215 7015 5235
rect 7035 5215 7050 5235
rect 7000 5185 7050 5215
rect 7000 5165 7015 5185
rect 7035 5165 7050 5185
rect 7000 5135 7050 5165
rect 7000 5115 7015 5135
rect 7035 5115 7050 5135
rect 7000 5085 7050 5115
rect 7000 5065 7015 5085
rect 7035 5065 7050 5085
rect 7000 5035 7050 5065
rect 7000 5015 7015 5035
rect 7035 5015 7050 5035
rect 7000 5000 7050 5015
rect 7150 5485 7200 5500
rect 7150 5465 7165 5485
rect 7185 5465 7200 5485
rect 7150 5435 7200 5465
rect 7150 5415 7165 5435
rect 7185 5415 7200 5435
rect 7150 5385 7200 5415
rect 7150 5365 7165 5385
rect 7185 5365 7200 5385
rect 7150 5335 7200 5365
rect 7150 5315 7165 5335
rect 7185 5315 7200 5335
rect 7150 5285 7200 5315
rect 7150 5265 7165 5285
rect 7185 5265 7200 5285
rect 7150 5235 7200 5265
rect 7150 5215 7165 5235
rect 7185 5215 7200 5235
rect 7150 5185 7200 5215
rect 7150 5165 7165 5185
rect 7185 5165 7200 5185
rect 7150 5135 7200 5165
rect 7150 5115 7165 5135
rect 7185 5115 7200 5135
rect 7150 5085 7200 5115
rect 7150 5065 7165 5085
rect 7185 5065 7200 5085
rect 7150 5035 7200 5065
rect 7150 5015 7165 5035
rect 7185 5015 7200 5035
rect 7150 5000 7200 5015
rect 7300 5485 7350 5500
rect 7300 5465 7315 5485
rect 7335 5465 7350 5485
rect 7300 5435 7350 5465
rect 7300 5415 7315 5435
rect 7335 5415 7350 5435
rect 7300 5385 7350 5415
rect 7300 5365 7315 5385
rect 7335 5365 7350 5385
rect 7300 5335 7350 5365
rect 7300 5315 7315 5335
rect 7335 5315 7350 5335
rect 7300 5285 7350 5315
rect 7300 5265 7315 5285
rect 7335 5265 7350 5285
rect 7300 5235 7350 5265
rect 7300 5215 7315 5235
rect 7335 5215 7350 5235
rect 7300 5185 7350 5215
rect 7300 5165 7315 5185
rect 7335 5165 7350 5185
rect 7300 5135 7350 5165
rect 7300 5115 7315 5135
rect 7335 5115 7350 5135
rect 7300 5085 7350 5115
rect 7300 5065 7315 5085
rect 7335 5065 7350 5085
rect 7300 5035 7350 5065
rect 7300 5015 7315 5035
rect 7335 5015 7350 5035
rect 7300 5000 7350 5015
rect 7450 5485 7500 5500
rect 7450 5465 7465 5485
rect 7485 5465 7500 5485
rect 7450 5435 7500 5465
rect 7450 5415 7465 5435
rect 7485 5415 7500 5435
rect 7450 5385 7500 5415
rect 7450 5365 7465 5385
rect 7485 5365 7500 5385
rect 7450 5335 7500 5365
rect 7450 5315 7465 5335
rect 7485 5315 7500 5335
rect 7450 5285 7500 5315
rect 7450 5265 7465 5285
rect 7485 5265 7500 5285
rect 7450 5235 7500 5265
rect 7450 5215 7465 5235
rect 7485 5215 7500 5235
rect 7450 5185 7500 5215
rect 7450 5165 7465 5185
rect 7485 5165 7500 5185
rect 7450 5135 7500 5165
rect 7450 5115 7465 5135
rect 7485 5115 7500 5135
rect 7450 5085 7500 5115
rect 7450 5065 7465 5085
rect 7485 5065 7500 5085
rect 7450 5035 7500 5065
rect 7450 5015 7465 5035
rect 7485 5015 7500 5035
rect 7450 5000 7500 5015
rect 7600 5485 7650 5500
rect 7600 5465 7615 5485
rect 7635 5465 7650 5485
rect 7600 5435 7650 5465
rect 7600 5415 7615 5435
rect 7635 5415 7650 5435
rect 7600 5385 7650 5415
rect 7600 5365 7615 5385
rect 7635 5365 7650 5385
rect 7600 5335 7650 5365
rect 7600 5315 7615 5335
rect 7635 5315 7650 5335
rect 7600 5285 7650 5315
rect 7600 5265 7615 5285
rect 7635 5265 7650 5285
rect 7600 5235 7650 5265
rect 7600 5215 7615 5235
rect 7635 5215 7650 5235
rect 7600 5185 7650 5215
rect 7600 5165 7615 5185
rect 7635 5165 7650 5185
rect 7600 5135 7650 5165
rect 7600 5115 7615 5135
rect 7635 5115 7650 5135
rect 7600 5085 7650 5115
rect 7600 5065 7615 5085
rect 7635 5065 7650 5085
rect 7600 5035 7650 5065
rect 7600 5015 7615 5035
rect 7635 5015 7650 5035
rect 7600 5000 7650 5015
rect 7750 5485 7800 5500
rect 7750 5465 7765 5485
rect 7785 5465 7800 5485
rect 7750 5435 7800 5465
rect 7750 5415 7765 5435
rect 7785 5415 7800 5435
rect 7750 5385 7800 5415
rect 7750 5365 7765 5385
rect 7785 5365 7800 5385
rect 7750 5335 7800 5365
rect 7750 5315 7765 5335
rect 7785 5315 7800 5335
rect 7750 5285 7800 5315
rect 7750 5265 7765 5285
rect 7785 5265 7800 5285
rect 7750 5235 7800 5265
rect 7750 5215 7765 5235
rect 7785 5215 7800 5235
rect 7750 5185 7800 5215
rect 7750 5165 7765 5185
rect 7785 5165 7800 5185
rect 7750 5135 7800 5165
rect 7750 5115 7765 5135
rect 7785 5115 7800 5135
rect 7750 5085 7800 5115
rect 7750 5065 7765 5085
rect 7785 5065 7800 5085
rect 7750 5035 7800 5065
rect 7750 5015 7765 5035
rect 7785 5015 7800 5035
rect 7750 5000 7800 5015
rect 8350 5485 8400 5500
rect 8350 5465 8365 5485
rect 8385 5465 8400 5485
rect 8350 5435 8400 5465
rect 8350 5415 8365 5435
rect 8385 5415 8400 5435
rect 8350 5385 8400 5415
rect 8350 5365 8365 5385
rect 8385 5365 8400 5385
rect 8350 5335 8400 5365
rect 8350 5315 8365 5335
rect 8385 5315 8400 5335
rect 8350 5285 8400 5315
rect 8350 5265 8365 5285
rect 8385 5265 8400 5285
rect 8350 5235 8400 5265
rect 8350 5215 8365 5235
rect 8385 5215 8400 5235
rect 8350 5185 8400 5215
rect 8350 5165 8365 5185
rect 8385 5165 8400 5185
rect 8350 5135 8400 5165
rect 8350 5115 8365 5135
rect 8385 5115 8400 5135
rect 8350 5085 8400 5115
rect 8350 5065 8365 5085
rect 8385 5065 8400 5085
rect 8350 5035 8400 5065
rect 8350 5015 8365 5035
rect 8385 5015 8400 5035
rect 8350 5000 8400 5015
rect 8500 5485 8550 5500
rect 8500 5465 8515 5485
rect 8535 5465 8550 5485
rect 8500 5435 8550 5465
rect 8500 5415 8515 5435
rect 8535 5415 8550 5435
rect 8500 5385 8550 5415
rect 8500 5365 8515 5385
rect 8535 5365 8550 5385
rect 8500 5335 8550 5365
rect 8500 5315 8515 5335
rect 8535 5315 8550 5335
rect 8500 5285 8550 5315
rect 8500 5265 8515 5285
rect 8535 5265 8550 5285
rect 8500 5235 8550 5265
rect 8500 5215 8515 5235
rect 8535 5215 8550 5235
rect 8500 5185 8550 5215
rect 8500 5165 8515 5185
rect 8535 5165 8550 5185
rect 8500 5135 8550 5165
rect 8500 5115 8515 5135
rect 8535 5115 8550 5135
rect 8500 5085 8550 5115
rect 8500 5065 8515 5085
rect 8535 5065 8550 5085
rect 8500 5035 8550 5065
rect 8500 5015 8515 5035
rect 8535 5015 8550 5035
rect 8500 4950 8550 5015
rect 8650 5485 8700 5500
rect 8650 5465 8665 5485
rect 8685 5465 8700 5485
rect 8650 5435 8700 5465
rect 8650 5415 8665 5435
rect 8685 5415 8700 5435
rect 8650 5385 8700 5415
rect 8650 5365 8665 5385
rect 8685 5365 8700 5385
rect 8650 5335 8700 5365
rect 8650 5315 8665 5335
rect 8685 5315 8700 5335
rect 8650 5285 8700 5315
rect 8650 5265 8665 5285
rect 8685 5265 8700 5285
rect 8650 5235 8700 5265
rect 8650 5215 8665 5235
rect 8685 5215 8700 5235
rect 8650 5185 8700 5215
rect 8650 5165 8665 5185
rect 8685 5165 8700 5185
rect 8650 5135 8700 5165
rect 8650 5115 8665 5135
rect 8685 5115 8700 5135
rect 8650 5085 8700 5115
rect 8650 5065 8665 5085
rect 8685 5065 8700 5085
rect 8650 5035 8700 5065
rect 8650 5015 8665 5035
rect 8685 5015 8700 5035
rect 8650 5000 8700 5015
rect 8800 5485 8850 5500
rect 8800 5465 8815 5485
rect 8835 5465 8850 5485
rect 8800 5435 8850 5465
rect 8800 5415 8815 5435
rect 8835 5415 8850 5435
rect 8800 5385 8850 5415
rect 8800 5365 8815 5385
rect 8835 5365 8850 5385
rect 8800 5335 8850 5365
rect 8800 5315 8815 5335
rect 8835 5315 8850 5335
rect 8800 5285 8850 5315
rect 8800 5265 8815 5285
rect 8835 5265 8850 5285
rect 8800 5235 8850 5265
rect 8800 5215 8815 5235
rect 8835 5215 8850 5235
rect 8800 5185 8850 5215
rect 8800 5165 8815 5185
rect 8835 5165 8850 5185
rect 8800 5135 8850 5165
rect 8800 5115 8815 5135
rect 8835 5115 8850 5135
rect 8800 5085 8850 5115
rect 8800 5065 8815 5085
rect 8835 5065 8850 5085
rect 8800 5035 8850 5065
rect 8800 5015 8815 5035
rect 8835 5015 8850 5035
rect 8800 4950 8850 5015
rect 8950 5485 9000 5500
rect 8950 5465 8965 5485
rect 8985 5465 9000 5485
rect 8950 5435 9000 5465
rect 8950 5415 8965 5435
rect 8985 5415 9000 5435
rect 8950 5385 9000 5415
rect 8950 5365 8965 5385
rect 8985 5365 9000 5385
rect 8950 5335 9000 5365
rect 8950 5315 8965 5335
rect 8985 5315 9000 5335
rect 8950 5285 9000 5315
rect 8950 5265 8965 5285
rect 8985 5265 9000 5285
rect 8950 5235 9000 5265
rect 8950 5215 8965 5235
rect 8985 5215 9000 5235
rect 8950 5185 9000 5215
rect 8950 5165 8965 5185
rect 8985 5165 9000 5185
rect 8950 5135 9000 5165
rect 8950 5115 8965 5135
rect 8985 5115 9000 5135
rect 8950 5085 9000 5115
rect 8950 5065 8965 5085
rect 8985 5065 9000 5085
rect 8950 5035 9000 5065
rect 8950 5015 8965 5035
rect 8985 5015 9000 5035
rect 8950 5000 9000 5015
rect 9100 5485 9150 5500
rect 9100 5465 9115 5485
rect 9135 5465 9150 5485
rect 9100 5435 9150 5465
rect 9100 5415 9115 5435
rect 9135 5415 9150 5435
rect 9100 5385 9150 5415
rect 9100 5365 9115 5385
rect 9135 5365 9150 5385
rect 9100 5335 9150 5365
rect 9100 5315 9115 5335
rect 9135 5315 9150 5335
rect 9100 5285 9150 5315
rect 9100 5265 9115 5285
rect 9135 5265 9150 5285
rect 9100 5235 9150 5265
rect 9100 5215 9115 5235
rect 9135 5215 9150 5235
rect 9100 5185 9150 5215
rect 9100 5165 9115 5185
rect 9135 5165 9150 5185
rect 9100 5135 9150 5165
rect 9100 5115 9115 5135
rect 9135 5115 9150 5135
rect 9100 5085 9150 5115
rect 9100 5065 9115 5085
rect 9135 5065 9150 5085
rect 9100 5035 9150 5065
rect 9100 5015 9115 5035
rect 9135 5015 9150 5035
rect 9100 4950 9150 5015
rect 9250 5485 9300 5500
rect 9250 5465 9265 5485
rect 9285 5465 9300 5485
rect 9250 5435 9300 5465
rect 9250 5415 9265 5435
rect 9285 5415 9300 5435
rect 9250 5385 9300 5415
rect 9250 5365 9265 5385
rect 9285 5365 9300 5385
rect 9250 5335 9300 5365
rect 9250 5315 9265 5335
rect 9285 5315 9300 5335
rect 9250 5285 9300 5315
rect 9250 5265 9265 5285
rect 9285 5265 9300 5285
rect 9250 5235 9300 5265
rect 9250 5215 9265 5235
rect 9285 5215 9300 5235
rect 9250 5185 9300 5215
rect 9250 5165 9265 5185
rect 9285 5165 9300 5185
rect 9250 5135 9300 5165
rect 9250 5115 9265 5135
rect 9285 5115 9300 5135
rect 9250 5085 9300 5115
rect 9250 5065 9265 5085
rect 9285 5065 9300 5085
rect 9250 5035 9300 5065
rect 9250 5015 9265 5035
rect 9285 5015 9300 5035
rect 9250 5000 9300 5015
rect 9400 5485 9450 5500
rect 9400 5465 9415 5485
rect 9435 5465 9450 5485
rect 9400 5435 9450 5465
rect 9400 5415 9415 5435
rect 9435 5415 9450 5435
rect 9400 5385 9450 5415
rect 9400 5365 9415 5385
rect 9435 5365 9450 5385
rect 9400 5335 9450 5365
rect 9400 5315 9415 5335
rect 9435 5315 9450 5335
rect 9400 5285 9450 5315
rect 9400 5265 9415 5285
rect 9435 5265 9450 5285
rect 9400 5235 9450 5265
rect 9400 5215 9415 5235
rect 9435 5215 9450 5235
rect 9400 5185 9450 5215
rect 9400 5165 9415 5185
rect 9435 5165 9450 5185
rect 9400 5135 9450 5165
rect 9400 5115 9415 5135
rect 9435 5115 9450 5135
rect 9400 5085 9450 5115
rect 9400 5065 9415 5085
rect 9435 5065 9450 5085
rect 9400 5035 9450 5065
rect 9400 5015 9415 5035
rect 9435 5015 9450 5035
rect 9400 4950 9450 5015
rect 9550 5485 9600 5500
rect 9550 5465 9565 5485
rect 9585 5465 9600 5485
rect 9550 5435 9600 5465
rect 9550 5415 9565 5435
rect 9585 5415 9600 5435
rect 9550 5385 9600 5415
rect 9550 5365 9565 5385
rect 9585 5365 9600 5385
rect 9550 5335 9600 5365
rect 9550 5315 9565 5335
rect 9585 5315 9600 5335
rect 9550 5285 9600 5315
rect 9550 5265 9565 5285
rect 9585 5265 9600 5285
rect 9550 5235 9600 5265
rect 9550 5215 9565 5235
rect 9585 5215 9600 5235
rect 9550 5185 9600 5215
rect 9550 5165 9565 5185
rect 9585 5165 9600 5185
rect 9550 5135 9600 5165
rect 9550 5115 9565 5135
rect 9585 5115 9600 5135
rect 9550 5085 9600 5115
rect 9550 5065 9565 5085
rect 9585 5065 9600 5085
rect 9550 5035 9600 5065
rect 9550 5015 9565 5035
rect 9585 5015 9600 5035
rect 9550 5000 9600 5015
rect 9700 5485 9750 5500
rect 9700 5465 9715 5485
rect 9735 5465 9750 5485
rect 9700 5435 9750 5465
rect 9700 5415 9715 5435
rect 9735 5415 9750 5435
rect 9700 5385 9750 5415
rect 9700 5365 9715 5385
rect 9735 5365 9750 5385
rect 9700 5335 9750 5365
rect 9700 5315 9715 5335
rect 9735 5315 9750 5335
rect 9700 5285 9750 5315
rect 9700 5265 9715 5285
rect 9735 5265 9750 5285
rect 9700 5235 9750 5265
rect 9700 5215 9715 5235
rect 9735 5215 9750 5235
rect 9700 5185 9750 5215
rect 9700 5165 9715 5185
rect 9735 5165 9750 5185
rect 9700 5135 9750 5165
rect 9700 5115 9715 5135
rect 9735 5115 9750 5135
rect 9700 5085 9750 5115
rect 9700 5065 9715 5085
rect 9735 5065 9750 5085
rect 9700 5035 9750 5065
rect 9700 5015 9715 5035
rect 9735 5015 9750 5035
rect 9700 4950 9750 5015
rect 9850 5485 9900 5500
rect 9850 5465 9865 5485
rect 9885 5465 9900 5485
rect 9850 5435 9900 5465
rect 9850 5415 9865 5435
rect 9885 5415 9900 5435
rect 9850 5385 9900 5415
rect 9850 5365 9865 5385
rect 9885 5365 9900 5385
rect 9850 5335 9900 5365
rect 9850 5315 9865 5335
rect 9885 5315 9900 5335
rect 9850 5285 9900 5315
rect 9850 5265 9865 5285
rect 9885 5265 9900 5285
rect 9850 5235 9900 5265
rect 9850 5215 9865 5235
rect 9885 5215 9900 5235
rect 9850 5185 9900 5215
rect 9850 5165 9865 5185
rect 9885 5165 9900 5185
rect 9850 5135 9900 5165
rect 9850 5115 9865 5135
rect 9885 5115 9900 5135
rect 9850 5085 9900 5115
rect 9850 5065 9865 5085
rect 9885 5065 9900 5085
rect 9850 5035 9900 5065
rect 9850 5015 9865 5035
rect 9885 5015 9900 5035
rect 9850 5000 9900 5015
rect 10000 5485 10050 5500
rect 10000 5465 10015 5485
rect 10035 5465 10050 5485
rect 10000 5435 10050 5465
rect 10000 5415 10015 5435
rect 10035 5415 10050 5435
rect 10000 5385 10050 5415
rect 10000 5365 10015 5385
rect 10035 5365 10050 5385
rect 10000 5335 10050 5365
rect 10000 5315 10015 5335
rect 10035 5315 10050 5335
rect 10000 5285 10050 5315
rect 10000 5265 10015 5285
rect 10035 5265 10050 5285
rect 10000 5235 10050 5265
rect 10000 5215 10015 5235
rect 10035 5215 10050 5235
rect 10000 5185 10050 5215
rect 10000 5165 10015 5185
rect 10035 5165 10050 5185
rect 10000 5135 10050 5165
rect 10000 5115 10015 5135
rect 10035 5115 10050 5135
rect 10000 5085 10050 5115
rect 10000 5065 10015 5085
rect 10035 5065 10050 5085
rect 10000 5035 10050 5065
rect 10000 5015 10015 5035
rect 10035 5015 10050 5035
rect 10000 4950 10050 5015
rect 10150 5485 10200 5500
rect 10150 5465 10165 5485
rect 10185 5465 10200 5485
rect 10150 5435 10200 5465
rect 10150 5415 10165 5435
rect 10185 5415 10200 5435
rect 10150 5385 10200 5415
rect 10150 5365 10165 5385
rect 10185 5365 10200 5385
rect 10150 5335 10200 5365
rect 10150 5315 10165 5335
rect 10185 5315 10200 5335
rect 10150 5285 10200 5315
rect 10150 5265 10165 5285
rect 10185 5265 10200 5285
rect 10150 5235 10200 5265
rect 10150 5215 10165 5235
rect 10185 5215 10200 5235
rect 10150 5185 10200 5215
rect 10150 5165 10165 5185
rect 10185 5165 10200 5185
rect 10150 5135 10200 5165
rect 10150 5115 10165 5135
rect 10185 5115 10200 5135
rect 10150 5085 10200 5115
rect 10150 5065 10165 5085
rect 10185 5065 10200 5085
rect 10150 5035 10200 5065
rect 10150 5015 10165 5035
rect 10185 5015 10200 5035
rect 10150 5000 10200 5015
rect 10300 5485 10350 5500
rect 10300 5465 10315 5485
rect 10335 5465 10350 5485
rect 10300 5435 10350 5465
rect 10300 5415 10315 5435
rect 10335 5415 10350 5435
rect 10300 5385 10350 5415
rect 10300 5365 10315 5385
rect 10335 5365 10350 5385
rect 10300 5335 10350 5365
rect 10300 5315 10315 5335
rect 10335 5315 10350 5335
rect 10300 5285 10350 5315
rect 10300 5265 10315 5285
rect 10335 5265 10350 5285
rect 10300 5235 10350 5265
rect 10300 5215 10315 5235
rect 10335 5215 10350 5235
rect 10300 5185 10350 5215
rect 10300 5165 10315 5185
rect 10335 5165 10350 5185
rect 10300 5135 10350 5165
rect 10300 5115 10315 5135
rect 10335 5115 10350 5135
rect 10300 5085 10350 5115
rect 10300 5065 10315 5085
rect 10335 5065 10350 5085
rect 10300 5035 10350 5065
rect 10300 5015 10315 5035
rect 10335 5015 10350 5035
rect 10300 4950 10350 5015
rect 10450 5485 10500 5500
rect 10450 5465 10465 5485
rect 10485 5465 10500 5485
rect 10450 5435 10500 5465
rect 10450 5415 10465 5435
rect 10485 5415 10500 5435
rect 10450 5385 10500 5415
rect 10450 5365 10465 5385
rect 10485 5365 10500 5385
rect 10450 5335 10500 5365
rect 10450 5315 10465 5335
rect 10485 5315 10500 5335
rect 10450 5285 10500 5315
rect 10450 5265 10465 5285
rect 10485 5265 10500 5285
rect 10450 5235 10500 5265
rect 10450 5215 10465 5235
rect 10485 5215 10500 5235
rect 10450 5185 10500 5215
rect 10450 5165 10465 5185
rect 10485 5165 10500 5185
rect 10450 5135 10500 5165
rect 10450 5115 10465 5135
rect 10485 5115 10500 5135
rect 10450 5085 10500 5115
rect 10450 5065 10465 5085
rect 10485 5065 10500 5085
rect 10450 5035 10500 5065
rect 10450 5015 10465 5035
rect 10485 5015 10500 5035
rect 10450 5000 10500 5015
rect 10600 5485 10650 5500
rect 10600 5465 10615 5485
rect 10635 5465 10650 5485
rect 10600 5435 10650 5465
rect 10600 5415 10615 5435
rect 10635 5415 10650 5435
rect 10600 5385 10650 5415
rect 10600 5365 10615 5385
rect 10635 5365 10650 5385
rect 10600 5335 10650 5365
rect 10600 5315 10615 5335
rect 10635 5315 10650 5335
rect 10600 5285 10650 5315
rect 10600 5265 10615 5285
rect 10635 5265 10650 5285
rect 10600 5235 10650 5265
rect 10600 5215 10615 5235
rect 10635 5215 10650 5235
rect 10600 5185 10650 5215
rect 10600 5165 10615 5185
rect 10635 5165 10650 5185
rect 10600 5135 10650 5165
rect 10600 5115 10615 5135
rect 10635 5115 10650 5135
rect 10600 5085 10650 5115
rect 10600 5065 10615 5085
rect 10635 5065 10650 5085
rect 10600 5035 10650 5065
rect 10600 5015 10615 5035
rect 10635 5015 10650 5035
rect 10600 4950 10650 5015
rect 10750 5485 10800 5500
rect 10750 5465 10765 5485
rect 10785 5465 10800 5485
rect 10750 5435 10800 5465
rect 10750 5415 10765 5435
rect 10785 5415 10800 5435
rect 10750 5385 10800 5415
rect 10750 5365 10765 5385
rect 10785 5365 10800 5385
rect 10750 5335 10800 5365
rect 10750 5315 10765 5335
rect 10785 5315 10800 5335
rect 10750 5285 10800 5315
rect 10750 5265 10765 5285
rect 10785 5265 10800 5285
rect 10750 5235 10800 5265
rect 10750 5215 10765 5235
rect 10785 5215 10800 5235
rect 10750 5185 10800 5215
rect 10750 5165 10765 5185
rect 10785 5165 10800 5185
rect 10750 5135 10800 5165
rect 10750 5115 10765 5135
rect 10785 5115 10800 5135
rect 10750 5085 10800 5115
rect 10750 5065 10765 5085
rect 10785 5065 10800 5085
rect 10750 5035 10800 5065
rect 10750 5015 10765 5035
rect 10785 5015 10800 5035
rect 10750 5000 10800 5015
rect 11350 5485 11400 5500
rect 11350 5465 11365 5485
rect 11385 5465 11400 5485
rect 11350 5435 11400 5465
rect 11350 5415 11365 5435
rect 11385 5415 11400 5435
rect 11350 5385 11400 5415
rect 11350 5365 11365 5385
rect 11385 5365 11400 5385
rect 11350 5335 11400 5365
rect 11350 5315 11365 5335
rect 11385 5315 11400 5335
rect 11350 5285 11400 5315
rect 11350 5265 11365 5285
rect 11385 5265 11400 5285
rect 11350 5235 11400 5265
rect 11350 5215 11365 5235
rect 11385 5215 11400 5235
rect 11350 5185 11400 5215
rect 11350 5165 11365 5185
rect 11385 5165 11400 5185
rect 11350 5135 11400 5165
rect 11350 5115 11365 5135
rect 11385 5115 11400 5135
rect 11350 5085 11400 5115
rect 11350 5065 11365 5085
rect 11385 5065 11400 5085
rect 11350 5035 11400 5065
rect 11350 5015 11365 5035
rect 11385 5015 11400 5035
rect 11350 5000 11400 5015
rect 11950 5485 12000 5500
rect 11950 5465 11965 5485
rect 11985 5465 12000 5485
rect 11950 5435 12000 5465
rect 11950 5415 11965 5435
rect 11985 5415 12000 5435
rect 11950 5385 12000 5415
rect 11950 5365 11965 5385
rect 11985 5365 12000 5385
rect 11950 5335 12000 5365
rect 11950 5315 11965 5335
rect 11985 5315 12000 5335
rect 11950 5285 12000 5315
rect 11950 5265 11965 5285
rect 11985 5265 12000 5285
rect 11950 5235 12000 5265
rect 11950 5215 11965 5235
rect 11985 5215 12000 5235
rect 11950 5185 12000 5215
rect 11950 5165 11965 5185
rect 11985 5165 12000 5185
rect 11950 5135 12000 5165
rect 11950 5115 11965 5135
rect 11985 5115 12000 5135
rect 11950 5085 12000 5115
rect 11950 5065 11965 5085
rect 11985 5065 12000 5085
rect 11950 5035 12000 5065
rect 11950 5015 11965 5035
rect 11985 5015 12000 5035
rect 11950 5000 12000 5015
rect 12550 5485 12600 5500
rect 12550 5465 12565 5485
rect 12585 5465 12600 5485
rect 12550 5435 12600 5465
rect 12550 5415 12565 5435
rect 12585 5415 12600 5435
rect 12550 5385 12600 5415
rect 12550 5365 12565 5385
rect 12585 5365 12600 5385
rect 12550 5335 12600 5365
rect 12550 5315 12565 5335
rect 12585 5315 12600 5335
rect 12550 5285 12600 5315
rect 12550 5265 12565 5285
rect 12585 5265 12600 5285
rect 12550 5235 12600 5265
rect 12550 5215 12565 5235
rect 12585 5215 12600 5235
rect 12550 5185 12600 5215
rect 12550 5165 12565 5185
rect 12585 5165 12600 5185
rect 12550 5135 12600 5165
rect 12550 5115 12565 5135
rect 12585 5115 12600 5135
rect 12550 5085 12600 5115
rect 12550 5065 12565 5085
rect 12585 5065 12600 5085
rect 12550 5035 12600 5065
rect 12550 5015 12565 5035
rect 12585 5015 12600 5035
rect 12550 5000 12600 5015
rect 13150 5485 13200 5500
rect 13150 5465 13165 5485
rect 13185 5465 13200 5485
rect 13150 5435 13200 5465
rect 13150 5415 13165 5435
rect 13185 5415 13200 5435
rect 13150 5385 13200 5415
rect 13150 5365 13165 5385
rect 13185 5365 13200 5385
rect 13150 5335 13200 5365
rect 13150 5315 13165 5335
rect 13185 5315 13200 5335
rect 13150 5285 13200 5315
rect 13150 5265 13165 5285
rect 13185 5265 13200 5285
rect 13150 5235 13200 5265
rect 13150 5215 13165 5235
rect 13185 5215 13200 5235
rect 13150 5185 13200 5215
rect 13150 5165 13165 5185
rect 13185 5165 13200 5185
rect 13150 5135 13200 5165
rect 13150 5115 13165 5135
rect 13185 5115 13200 5135
rect 13150 5085 13200 5115
rect 13150 5065 13165 5085
rect 13185 5065 13200 5085
rect 13150 5035 13200 5065
rect 13150 5015 13165 5035
rect 13185 5015 13200 5035
rect 13150 5000 13200 5015
rect 13750 5485 13800 5500
rect 13750 5465 13765 5485
rect 13785 5465 13800 5485
rect 13750 5435 13800 5465
rect 13750 5415 13765 5435
rect 13785 5415 13800 5435
rect 13750 5385 13800 5415
rect 13750 5365 13765 5385
rect 13785 5365 13800 5385
rect 13750 5335 13800 5365
rect 13750 5315 13765 5335
rect 13785 5315 13800 5335
rect 13750 5285 13800 5315
rect 13750 5265 13765 5285
rect 13785 5265 13800 5285
rect 13750 5235 13800 5265
rect 13750 5215 13765 5235
rect 13785 5215 13800 5235
rect 13750 5185 13800 5215
rect 13750 5165 13765 5185
rect 13785 5165 13800 5185
rect 13750 5135 13800 5165
rect 13750 5115 13765 5135
rect 13785 5115 13800 5135
rect 13750 5085 13800 5115
rect 13750 5065 13765 5085
rect 13785 5065 13800 5085
rect 13750 5035 13800 5065
rect 13750 5015 13765 5035
rect 13785 5015 13800 5035
rect 13750 5000 13800 5015
rect 14350 5485 14400 5500
rect 14350 5465 14365 5485
rect 14385 5465 14400 5485
rect 14350 5435 14400 5465
rect 14350 5415 14365 5435
rect 14385 5415 14400 5435
rect 14350 5385 14400 5415
rect 14350 5365 14365 5385
rect 14385 5365 14400 5385
rect 14350 5335 14400 5365
rect 14350 5315 14365 5335
rect 14385 5315 14400 5335
rect 14350 5285 14400 5315
rect 14350 5265 14365 5285
rect 14385 5265 14400 5285
rect 14350 5235 14400 5265
rect 14350 5215 14365 5235
rect 14385 5215 14400 5235
rect 14350 5185 14400 5215
rect 14350 5165 14365 5185
rect 14385 5165 14400 5185
rect 14350 5135 14400 5165
rect 14350 5115 14365 5135
rect 14385 5115 14400 5135
rect 14350 5085 14400 5115
rect 14350 5065 14365 5085
rect 14385 5065 14400 5085
rect 14350 5035 14400 5065
rect 14350 5015 14365 5035
rect 14385 5015 14400 5035
rect 14350 5000 14400 5015
rect 14950 5485 15000 5500
rect 14950 5465 14965 5485
rect 14985 5465 15000 5485
rect 14950 5435 15000 5465
rect 14950 5415 14965 5435
rect 14985 5415 15000 5435
rect 14950 5385 15000 5415
rect 14950 5365 14965 5385
rect 14985 5365 15000 5385
rect 14950 5335 15000 5365
rect 14950 5315 14965 5335
rect 14985 5315 15000 5335
rect 14950 5285 15000 5315
rect 14950 5265 14965 5285
rect 14985 5265 15000 5285
rect 14950 5235 15000 5265
rect 14950 5215 14965 5235
rect 14985 5215 15000 5235
rect 14950 5185 15000 5215
rect 14950 5165 14965 5185
rect 14985 5165 15000 5185
rect 14950 5135 15000 5165
rect 14950 5115 14965 5135
rect 14985 5115 15000 5135
rect 14950 5085 15000 5115
rect 14950 5065 14965 5085
rect 14985 5065 15000 5085
rect 14950 5035 15000 5065
rect 14950 5015 14965 5035
rect 14985 5015 15000 5035
rect 14950 5000 15000 5015
rect 15550 5485 15600 5500
rect 15550 5465 15565 5485
rect 15585 5465 15600 5485
rect 15550 5435 15600 5465
rect 15550 5415 15565 5435
rect 15585 5415 15600 5435
rect 15550 5385 15600 5415
rect 15550 5365 15565 5385
rect 15585 5365 15600 5385
rect 15550 5335 15600 5365
rect 15550 5315 15565 5335
rect 15585 5315 15600 5335
rect 15550 5285 15600 5315
rect 15550 5265 15565 5285
rect 15585 5265 15600 5285
rect 15550 5235 15600 5265
rect 15550 5215 15565 5235
rect 15585 5215 15600 5235
rect 15550 5185 15600 5215
rect 15550 5165 15565 5185
rect 15585 5165 15600 5185
rect 15550 5135 15600 5165
rect 15550 5115 15565 5135
rect 15585 5115 15600 5135
rect 15550 5085 15600 5115
rect 15550 5065 15565 5085
rect 15585 5065 15600 5085
rect 15550 5035 15600 5065
rect 15550 5015 15565 5035
rect 15585 5015 15600 5035
rect 15550 5000 15600 5015
rect 16150 5485 16200 5500
rect 16150 5465 16165 5485
rect 16185 5465 16200 5485
rect 16150 5435 16200 5465
rect 16150 5415 16165 5435
rect 16185 5415 16200 5435
rect 16150 5385 16200 5415
rect 16150 5365 16165 5385
rect 16185 5365 16200 5385
rect 16150 5335 16200 5365
rect 16150 5315 16165 5335
rect 16185 5315 16200 5335
rect 16150 5285 16200 5315
rect 16150 5265 16165 5285
rect 16185 5265 16200 5285
rect 16150 5235 16200 5265
rect 16150 5215 16165 5235
rect 16185 5215 16200 5235
rect 16150 5185 16200 5215
rect 16150 5165 16165 5185
rect 16185 5165 16200 5185
rect 16150 5135 16200 5165
rect 16150 5115 16165 5135
rect 16185 5115 16200 5135
rect 16150 5085 16200 5115
rect 16150 5065 16165 5085
rect 16185 5065 16200 5085
rect 16150 5035 16200 5065
rect 16150 5015 16165 5035
rect 16185 5015 16200 5035
rect 16150 5000 16200 5015
rect 16300 5485 16350 5500
rect 16300 5465 16315 5485
rect 16335 5465 16350 5485
rect 16300 5435 16350 5465
rect 16300 5415 16315 5435
rect 16335 5415 16350 5435
rect 16300 5385 16350 5415
rect 16300 5365 16315 5385
rect 16335 5365 16350 5385
rect 16300 5335 16350 5365
rect 16300 5315 16315 5335
rect 16335 5315 16350 5335
rect 16300 5285 16350 5315
rect 16300 5265 16315 5285
rect 16335 5265 16350 5285
rect 16300 5235 16350 5265
rect 16300 5215 16315 5235
rect 16335 5215 16350 5235
rect 16300 5185 16350 5215
rect 16300 5165 16315 5185
rect 16335 5165 16350 5185
rect 16300 5135 16350 5165
rect 16300 5115 16315 5135
rect 16335 5115 16350 5135
rect 16300 5085 16350 5115
rect 16300 5065 16315 5085
rect 16335 5065 16350 5085
rect 16300 5035 16350 5065
rect 16300 5015 16315 5035
rect 16335 5015 16350 5035
rect 16300 5000 16350 5015
rect 16450 5485 16500 5500
rect 16450 5465 16465 5485
rect 16485 5465 16500 5485
rect 16450 5435 16500 5465
rect 16450 5415 16465 5435
rect 16485 5415 16500 5435
rect 16450 5385 16500 5415
rect 16450 5365 16465 5385
rect 16485 5365 16500 5385
rect 16450 5335 16500 5365
rect 16450 5315 16465 5335
rect 16485 5315 16500 5335
rect 16450 5285 16500 5315
rect 16450 5265 16465 5285
rect 16485 5265 16500 5285
rect 16450 5235 16500 5265
rect 16450 5215 16465 5235
rect 16485 5215 16500 5235
rect 16450 5185 16500 5215
rect 16450 5165 16465 5185
rect 16485 5165 16500 5185
rect 16450 5135 16500 5165
rect 16450 5115 16465 5135
rect 16485 5115 16500 5135
rect 16450 5085 16500 5115
rect 16450 5065 16465 5085
rect 16485 5065 16500 5085
rect 16450 5035 16500 5065
rect 16450 5015 16465 5035
rect 16485 5015 16500 5035
rect 16450 5000 16500 5015
rect 16600 5485 16650 5500
rect 16600 5465 16615 5485
rect 16635 5465 16650 5485
rect 16600 5435 16650 5465
rect 16600 5415 16615 5435
rect 16635 5415 16650 5435
rect 16600 5385 16650 5415
rect 16600 5365 16615 5385
rect 16635 5365 16650 5385
rect 16600 5335 16650 5365
rect 16600 5315 16615 5335
rect 16635 5315 16650 5335
rect 16600 5285 16650 5315
rect 16600 5265 16615 5285
rect 16635 5265 16650 5285
rect 16600 5235 16650 5265
rect 16600 5215 16615 5235
rect 16635 5215 16650 5235
rect 16600 5185 16650 5215
rect 16600 5165 16615 5185
rect 16635 5165 16650 5185
rect 16600 5135 16650 5165
rect 16600 5115 16615 5135
rect 16635 5115 16650 5135
rect 16600 5085 16650 5115
rect 16600 5065 16615 5085
rect 16635 5065 16650 5085
rect 16600 5035 16650 5065
rect 16600 5015 16615 5035
rect 16635 5015 16650 5035
rect 16600 5000 16650 5015
rect 16750 5485 16800 5500
rect 16750 5465 16765 5485
rect 16785 5465 16800 5485
rect 16750 5435 16800 5465
rect 16750 5415 16765 5435
rect 16785 5415 16800 5435
rect 16750 5385 16800 5415
rect 16750 5365 16765 5385
rect 16785 5365 16800 5385
rect 16750 5335 16800 5365
rect 16750 5315 16765 5335
rect 16785 5315 16800 5335
rect 16750 5285 16800 5315
rect 16750 5265 16765 5285
rect 16785 5265 16800 5285
rect 16750 5235 16800 5265
rect 16750 5215 16765 5235
rect 16785 5215 16800 5235
rect 16750 5185 16800 5215
rect 16750 5165 16765 5185
rect 16785 5165 16800 5185
rect 16750 5135 16800 5165
rect 16750 5115 16765 5135
rect 16785 5115 16800 5135
rect 16750 5085 16800 5115
rect 16750 5065 16765 5085
rect 16785 5065 16800 5085
rect 16750 5035 16800 5065
rect 16750 5015 16765 5035
rect 16785 5015 16800 5035
rect 16750 5000 16800 5015
rect 16900 5485 16950 5500
rect 16900 5465 16915 5485
rect 16935 5465 16950 5485
rect 16900 5435 16950 5465
rect 16900 5415 16915 5435
rect 16935 5415 16950 5435
rect 16900 5385 16950 5415
rect 16900 5365 16915 5385
rect 16935 5365 16950 5385
rect 16900 5335 16950 5365
rect 16900 5315 16915 5335
rect 16935 5315 16950 5335
rect 16900 5285 16950 5315
rect 16900 5265 16915 5285
rect 16935 5265 16950 5285
rect 16900 5235 16950 5265
rect 16900 5215 16915 5235
rect 16935 5215 16950 5235
rect 16900 5185 16950 5215
rect 16900 5165 16915 5185
rect 16935 5165 16950 5185
rect 16900 5135 16950 5165
rect 16900 5115 16915 5135
rect 16935 5115 16950 5135
rect 16900 5085 16950 5115
rect 16900 5065 16915 5085
rect 16935 5065 16950 5085
rect 16900 5035 16950 5065
rect 16900 5015 16915 5035
rect 16935 5015 16950 5035
rect 16900 5000 16950 5015
rect 17050 5485 17100 5500
rect 17050 5465 17065 5485
rect 17085 5465 17100 5485
rect 17050 5435 17100 5465
rect 17050 5415 17065 5435
rect 17085 5415 17100 5435
rect 17050 5385 17100 5415
rect 17050 5365 17065 5385
rect 17085 5365 17100 5385
rect 17050 5335 17100 5365
rect 17050 5315 17065 5335
rect 17085 5315 17100 5335
rect 17050 5285 17100 5315
rect 17050 5265 17065 5285
rect 17085 5265 17100 5285
rect 17050 5235 17100 5265
rect 17050 5215 17065 5235
rect 17085 5215 17100 5235
rect 17050 5185 17100 5215
rect 17050 5165 17065 5185
rect 17085 5165 17100 5185
rect 17050 5135 17100 5165
rect 17050 5115 17065 5135
rect 17085 5115 17100 5135
rect 17050 5085 17100 5115
rect 17050 5065 17065 5085
rect 17085 5065 17100 5085
rect 17050 5035 17100 5065
rect 17050 5015 17065 5035
rect 17085 5015 17100 5035
rect 17050 5000 17100 5015
rect 17200 5485 17250 5500
rect 17200 5465 17215 5485
rect 17235 5465 17250 5485
rect 17200 5435 17250 5465
rect 17200 5415 17215 5435
rect 17235 5415 17250 5435
rect 17200 5385 17250 5415
rect 17200 5365 17215 5385
rect 17235 5365 17250 5385
rect 17200 5335 17250 5365
rect 17200 5315 17215 5335
rect 17235 5315 17250 5335
rect 17200 5285 17250 5315
rect 17200 5265 17215 5285
rect 17235 5265 17250 5285
rect 17200 5235 17250 5265
rect 17200 5215 17215 5235
rect 17235 5215 17250 5235
rect 17200 5185 17250 5215
rect 17200 5165 17215 5185
rect 17235 5165 17250 5185
rect 17200 5135 17250 5165
rect 17200 5115 17215 5135
rect 17235 5115 17250 5135
rect 17200 5085 17250 5115
rect 17200 5065 17215 5085
rect 17235 5065 17250 5085
rect 17200 5035 17250 5065
rect 17200 5015 17215 5035
rect 17235 5015 17250 5035
rect 17200 5000 17250 5015
rect 17350 5485 17400 5500
rect 17350 5465 17365 5485
rect 17385 5465 17400 5485
rect 17350 5435 17400 5465
rect 17350 5415 17365 5435
rect 17385 5415 17400 5435
rect 17350 5385 17400 5415
rect 17350 5365 17365 5385
rect 17385 5365 17400 5385
rect 17350 5335 17400 5365
rect 17350 5315 17365 5335
rect 17385 5315 17400 5335
rect 17350 5285 17400 5315
rect 17350 5265 17365 5285
rect 17385 5265 17400 5285
rect 17350 5235 17400 5265
rect 17350 5215 17365 5235
rect 17385 5215 17400 5235
rect 17350 5185 17400 5215
rect 17350 5165 17365 5185
rect 17385 5165 17400 5185
rect 17350 5135 17400 5165
rect 17350 5115 17365 5135
rect 17385 5115 17400 5135
rect 17350 5085 17400 5115
rect 17350 5065 17365 5085
rect 17385 5065 17400 5085
rect 17350 5035 17400 5065
rect 17350 5015 17365 5035
rect 17385 5015 17400 5035
rect 17350 5000 17400 5015
rect 17950 5485 18000 5500
rect 17950 5465 17965 5485
rect 17985 5465 18000 5485
rect 17950 5435 18000 5465
rect 17950 5415 17965 5435
rect 17985 5415 18000 5435
rect 17950 5385 18000 5415
rect 17950 5365 17965 5385
rect 17985 5365 18000 5385
rect 17950 5335 18000 5365
rect 17950 5315 17965 5335
rect 17985 5315 18000 5335
rect 17950 5285 18000 5315
rect 17950 5265 17965 5285
rect 17985 5265 18000 5285
rect 17950 5235 18000 5265
rect 17950 5215 17965 5235
rect 17985 5215 18000 5235
rect 17950 5185 18000 5215
rect 17950 5165 17965 5185
rect 17985 5165 18000 5185
rect 17950 5135 18000 5165
rect 17950 5115 17965 5135
rect 17985 5115 18000 5135
rect 17950 5085 18000 5115
rect 17950 5065 17965 5085
rect 17985 5065 18000 5085
rect 17950 5035 18000 5065
rect 17950 5015 17965 5035
rect 17985 5015 18000 5035
rect 17950 5000 18000 5015
rect 18550 5485 18600 5500
rect 18550 5465 18565 5485
rect 18585 5465 18600 5485
rect 18550 5435 18600 5465
rect 18550 5415 18565 5435
rect 18585 5415 18600 5435
rect 18550 5385 18600 5415
rect 18550 5365 18565 5385
rect 18585 5365 18600 5385
rect 18550 5335 18600 5365
rect 18550 5315 18565 5335
rect 18585 5315 18600 5335
rect 18550 5285 18600 5315
rect 18550 5265 18565 5285
rect 18585 5265 18600 5285
rect 18550 5235 18600 5265
rect 18550 5215 18565 5235
rect 18585 5215 18600 5235
rect 18550 5185 18600 5215
rect 18550 5165 18565 5185
rect 18585 5165 18600 5185
rect 18550 5135 18600 5165
rect 18550 5115 18565 5135
rect 18585 5115 18600 5135
rect 18550 5085 18600 5115
rect 18550 5065 18565 5085
rect 18585 5065 18600 5085
rect 18550 5035 18600 5065
rect 18550 5015 18565 5035
rect 18585 5015 18600 5035
rect 18550 5000 18600 5015
rect 18700 5485 18750 5500
rect 18700 5465 18715 5485
rect 18735 5465 18750 5485
rect 18700 5435 18750 5465
rect 18700 5415 18715 5435
rect 18735 5415 18750 5435
rect 18700 5385 18750 5415
rect 18700 5365 18715 5385
rect 18735 5365 18750 5385
rect 18700 5335 18750 5365
rect 18700 5315 18715 5335
rect 18735 5315 18750 5335
rect 18700 5285 18750 5315
rect 18700 5265 18715 5285
rect 18735 5265 18750 5285
rect 18700 5235 18750 5265
rect 18700 5215 18715 5235
rect 18735 5215 18750 5235
rect 18700 5185 18750 5215
rect 18700 5165 18715 5185
rect 18735 5165 18750 5185
rect 18700 5135 18750 5165
rect 18700 5115 18715 5135
rect 18735 5115 18750 5135
rect 18700 5085 18750 5115
rect 18700 5065 18715 5085
rect 18735 5065 18750 5085
rect 18700 5035 18750 5065
rect 18700 5015 18715 5035
rect 18735 5015 18750 5035
rect 18700 5000 18750 5015
rect 18850 5485 18900 5500
rect 18850 5465 18865 5485
rect 18885 5465 18900 5485
rect 18850 5435 18900 5465
rect 18850 5415 18865 5435
rect 18885 5415 18900 5435
rect 18850 5385 18900 5415
rect 18850 5365 18865 5385
rect 18885 5365 18900 5385
rect 18850 5335 18900 5365
rect 18850 5315 18865 5335
rect 18885 5315 18900 5335
rect 18850 5285 18900 5315
rect 18850 5265 18865 5285
rect 18885 5265 18900 5285
rect 18850 5235 18900 5265
rect 18850 5215 18865 5235
rect 18885 5215 18900 5235
rect 18850 5185 18900 5215
rect 18850 5165 18865 5185
rect 18885 5165 18900 5185
rect 18850 5135 18900 5165
rect 18850 5115 18865 5135
rect 18885 5115 18900 5135
rect 18850 5085 18900 5115
rect 18850 5065 18865 5085
rect 18885 5065 18900 5085
rect 18850 5035 18900 5065
rect 18850 5015 18865 5035
rect 18885 5015 18900 5035
rect 18850 5000 18900 5015
rect 19000 5485 19050 5500
rect 19000 5465 19015 5485
rect 19035 5465 19050 5485
rect 19000 5435 19050 5465
rect 19000 5415 19015 5435
rect 19035 5415 19050 5435
rect 19000 5385 19050 5415
rect 19000 5365 19015 5385
rect 19035 5365 19050 5385
rect 19000 5335 19050 5365
rect 19000 5315 19015 5335
rect 19035 5315 19050 5335
rect 19000 5285 19050 5315
rect 19000 5265 19015 5285
rect 19035 5265 19050 5285
rect 19000 5235 19050 5265
rect 19000 5215 19015 5235
rect 19035 5215 19050 5235
rect 19000 5185 19050 5215
rect 19000 5165 19015 5185
rect 19035 5165 19050 5185
rect 19000 5135 19050 5165
rect 19000 5115 19015 5135
rect 19035 5115 19050 5135
rect 19000 5085 19050 5115
rect 19000 5065 19015 5085
rect 19035 5065 19050 5085
rect 19000 5035 19050 5065
rect 19000 5015 19015 5035
rect 19035 5015 19050 5035
rect 19000 5000 19050 5015
rect 19150 5485 19200 5500
rect 19150 5465 19165 5485
rect 19185 5465 19200 5485
rect 19150 5435 19200 5465
rect 19150 5415 19165 5435
rect 19185 5415 19200 5435
rect 19150 5385 19200 5415
rect 19150 5365 19165 5385
rect 19185 5365 19200 5385
rect 19150 5335 19200 5365
rect 19150 5315 19165 5335
rect 19185 5315 19200 5335
rect 19150 5285 19200 5315
rect 19150 5265 19165 5285
rect 19185 5265 19200 5285
rect 19150 5235 19200 5265
rect 19150 5215 19165 5235
rect 19185 5215 19200 5235
rect 19150 5185 19200 5215
rect 19150 5165 19165 5185
rect 19185 5165 19200 5185
rect 19150 5135 19200 5165
rect 19150 5115 19165 5135
rect 19185 5115 19200 5135
rect 19150 5085 19200 5115
rect 19150 5065 19165 5085
rect 19185 5065 19200 5085
rect 19150 5035 19200 5065
rect 19150 5015 19165 5035
rect 19185 5015 19200 5035
rect 19150 5000 19200 5015
rect 19300 5485 19350 5500
rect 19300 5465 19315 5485
rect 19335 5465 19350 5485
rect 19300 5435 19350 5465
rect 19300 5415 19315 5435
rect 19335 5415 19350 5435
rect 19300 5385 19350 5415
rect 19300 5365 19315 5385
rect 19335 5365 19350 5385
rect 19300 5335 19350 5365
rect 19300 5315 19315 5335
rect 19335 5315 19350 5335
rect 19300 5285 19350 5315
rect 19300 5265 19315 5285
rect 19335 5265 19350 5285
rect 19300 5235 19350 5265
rect 19300 5215 19315 5235
rect 19335 5215 19350 5235
rect 19300 5185 19350 5215
rect 19300 5165 19315 5185
rect 19335 5165 19350 5185
rect 19300 5135 19350 5165
rect 19300 5115 19315 5135
rect 19335 5115 19350 5135
rect 19300 5085 19350 5115
rect 19300 5065 19315 5085
rect 19335 5065 19350 5085
rect 19300 5035 19350 5065
rect 19300 5015 19315 5035
rect 19335 5015 19350 5035
rect 19300 5000 19350 5015
rect 19450 5485 19500 5500
rect 19450 5465 19465 5485
rect 19485 5465 19500 5485
rect 19450 5435 19500 5465
rect 19450 5415 19465 5435
rect 19485 5415 19500 5435
rect 19450 5385 19500 5415
rect 19450 5365 19465 5385
rect 19485 5365 19500 5385
rect 19450 5335 19500 5365
rect 19450 5315 19465 5335
rect 19485 5315 19500 5335
rect 19450 5285 19500 5315
rect 19450 5265 19465 5285
rect 19485 5265 19500 5285
rect 19450 5235 19500 5265
rect 19450 5215 19465 5235
rect 19485 5215 19500 5235
rect 19450 5185 19500 5215
rect 19450 5165 19465 5185
rect 19485 5165 19500 5185
rect 19450 5135 19500 5165
rect 19450 5115 19465 5135
rect 19485 5115 19500 5135
rect 19450 5085 19500 5115
rect 19450 5065 19465 5085
rect 19485 5065 19500 5085
rect 19450 5035 19500 5065
rect 19450 5015 19465 5035
rect 19485 5015 19500 5035
rect 19450 5000 19500 5015
rect 19600 5485 19650 5500
rect 19600 5465 19615 5485
rect 19635 5465 19650 5485
rect 19600 5435 19650 5465
rect 19600 5415 19615 5435
rect 19635 5415 19650 5435
rect 19600 5385 19650 5415
rect 19600 5365 19615 5385
rect 19635 5365 19650 5385
rect 19600 5335 19650 5365
rect 19600 5315 19615 5335
rect 19635 5315 19650 5335
rect 19600 5285 19650 5315
rect 19600 5265 19615 5285
rect 19635 5265 19650 5285
rect 19600 5235 19650 5265
rect 19600 5215 19615 5235
rect 19635 5215 19650 5235
rect 19600 5185 19650 5215
rect 19600 5165 19615 5185
rect 19635 5165 19650 5185
rect 19600 5135 19650 5165
rect 19600 5115 19615 5135
rect 19635 5115 19650 5135
rect 19600 5085 19650 5115
rect 19600 5065 19615 5085
rect 19635 5065 19650 5085
rect 19600 5035 19650 5065
rect 19600 5015 19615 5035
rect 19635 5015 19650 5035
rect 19600 5000 19650 5015
rect 19750 5485 19800 5500
rect 19750 5465 19765 5485
rect 19785 5465 19800 5485
rect 19750 5435 19800 5465
rect 19750 5415 19765 5435
rect 19785 5415 19800 5435
rect 19750 5385 19800 5415
rect 19750 5365 19765 5385
rect 19785 5365 19800 5385
rect 19750 5335 19800 5365
rect 19750 5315 19765 5335
rect 19785 5315 19800 5335
rect 19750 5285 19800 5315
rect 19750 5265 19765 5285
rect 19785 5265 19800 5285
rect 19750 5235 19800 5265
rect 19750 5215 19765 5235
rect 19785 5215 19800 5235
rect 19750 5185 19800 5215
rect 19750 5165 19765 5185
rect 19785 5165 19800 5185
rect 19750 5135 19800 5165
rect 19750 5115 19765 5135
rect 19785 5115 19800 5135
rect 19750 5085 19800 5115
rect 19750 5065 19765 5085
rect 19785 5065 19800 5085
rect 19750 5035 19800 5065
rect 19750 5015 19765 5035
rect 19785 5015 19800 5035
rect 19750 5000 19800 5015
rect 20350 5485 20400 5500
rect 20350 5465 20365 5485
rect 20385 5465 20400 5485
rect 20350 5435 20400 5465
rect 20350 5415 20365 5435
rect 20385 5415 20400 5435
rect 20350 5385 20400 5415
rect 20350 5365 20365 5385
rect 20385 5365 20400 5385
rect 20350 5335 20400 5365
rect 20350 5315 20365 5335
rect 20385 5315 20400 5335
rect 20350 5285 20400 5315
rect 20350 5265 20365 5285
rect 20385 5265 20400 5285
rect 20350 5235 20400 5265
rect 20350 5215 20365 5235
rect 20385 5215 20400 5235
rect 20350 5185 20400 5215
rect 20350 5165 20365 5185
rect 20385 5165 20400 5185
rect 20350 5135 20400 5165
rect 20350 5115 20365 5135
rect 20385 5115 20400 5135
rect 20350 5085 20400 5115
rect 20350 5065 20365 5085
rect 20385 5065 20400 5085
rect 20350 5035 20400 5065
rect 20350 5015 20365 5035
rect 20385 5015 20400 5035
rect 20350 5000 20400 5015
rect 20950 5485 21000 5500
rect 20950 5465 20965 5485
rect 20985 5465 21000 5485
rect 20950 5435 21000 5465
rect 20950 5415 20965 5435
rect 20985 5415 21000 5435
rect 20950 5385 21000 5415
rect 20950 5365 20965 5385
rect 20985 5365 21000 5385
rect 20950 5335 21000 5365
rect 20950 5315 20965 5335
rect 20985 5315 21000 5335
rect 20950 5285 21000 5315
rect 20950 5265 20965 5285
rect 20985 5265 21000 5285
rect 20950 5235 21000 5265
rect 20950 5215 20965 5235
rect 20985 5215 21000 5235
rect 20950 5185 21000 5215
rect 20950 5165 20965 5185
rect 20985 5165 21000 5185
rect 20950 5135 21000 5165
rect 20950 5115 20965 5135
rect 20985 5115 21000 5135
rect 20950 5085 21000 5115
rect 20950 5065 20965 5085
rect 20985 5065 21000 5085
rect 20950 5035 21000 5065
rect 20950 5015 20965 5035
rect 20985 5015 21000 5035
rect 20950 5000 21000 5015
rect 21400 5485 21450 5500
rect 21400 5465 21415 5485
rect 21435 5465 21450 5485
rect 21400 5435 21450 5465
rect 21400 5415 21415 5435
rect 21435 5415 21450 5435
rect 21400 5385 21450 5415
rect 21400 5365 21415 5385
rect 21435 5365 21450 5385
rect 21400 5335 21450 5365
rect 21400 5315 21415 5335
rect 21435 5315 21450 5335
rect 21400 5285 21450 5315
rect 21400 5265 21415 5285
rect 21435 5265 21450 5285
rect 21400 5235 21450 5265
rect 21400 5215 21415 5235
rect 21435 5215 21450 5235
rect 21400 5185 21450 5215
rect 21400 5165 21415 5185
rect 21435 5165 21450 5185
rect 21400 5135 21450 5165
rect 21400 5115 21415 5135
rect 21435 5115 21450 5135
rect 21400 5085 21450 5115
rect 21400 5065 21415 5085
rect 21435 5065 21450 5085
rect 21400 5035 21450 5065
rect 21400 5015 21415 5035
rect 21435 5015 21450 5035
rect 21400 5000 21450 5015
rect 21850 5485 21900 5500
rect 21850 5465 21865 5485
rect 21885 5465 21900 5485
rect 21850 5435 21900 5465
rect 21850 5415 21865 5435
rect 21885 5415 21900 5435
rect 21850 5385 21900 5415
rect 21850 5365 21865 5385
rect 21885 5365 21900 5385
rect 21850 5335 21900 5365
rect 21850 5315 21865 5335
rect 21885 5315 21900 5335
rect 21850 5285 21900 5315
rect 21850 5265 21865 5285
rect 21885 5265 21900 5285
rect 21850 5235 21900 5265
rect 21850 5215 21865 5235
rect 21885 5215 21900 5235
rect 21850 5185 21900 5215
rect 21850 5165 21865 5185
rect 21885 5165 21900 5185
rect 21850 5135 21900 5165
rect 21850 5115 21865 5135
rect 21885 5115 21900 5135
rect 21850 5085 21900 5115
rect 21850 5065 21865 5085
rect 21885 5065 21900 5085
rect 21850 5035 21900 5065
rect 21850 5015 21865 5035
rect 21885 5015 21900 5035
rect 21850 5000 21900 5015
rect 22450 5485 22500 5500
rect 22450 5465 22465 5485
rect 22485 5465 22500 5485
rect 22450 5435 22500 5465
rect 22450 5415 22465 5435
rect 22485 5415 22500 5435
rect 22450 5385 22500 5415
rect 22450 5365 22465 5385
rect 22485 5365 22500 5385
rect 22450 5335 22500 5365
rect 22450 5315 22465 5335
rect 22485 5315 22500 5335
rect 22450 5285 22500 5315
rect 22450 5265 22465 5285
rect 22485 5265 22500 5285
rect 22450 5235 22500 5265
rect 22450 5215 22465 5235
rect 22485 5215 22500 5235
rect 22450 5185 22500 5215
rect 22450 5165 22465 5185
rect 22485 5165 22500 5185
rect 22450 5135 22500 5165
rect 22450 5115 22465 5135
rect 22485 5115 22500 5135
rect 22450 5085 22500 5115
rect 22450 5065 22465 5085
rect 22485 5065 22500 5085
rect 22450 5035 22500 5065
rect 22450 5015 22465 5035
rect 22485 5015 22500 5035
rect 22450 5000 22500 5015
rect 23050 5485 23100 5500
rect 23050 5465 23065 5485
rect 23085 5465 23100 5485
rect 23050 5435 23100 5465
rect 23050 5415 23065 5435
rect 23085 5415 23100 5435
rect 23050 5385 23100 5415
rect 23050 5365 23065 5385
rect 23085 5365 23100 5385
rect 23050 5335 23100 5365
rect 23050 5315 23065 5335
rect 23085 5315 23100 5335
rect 23050 5285 23100 5315
rect 23050 5265 23065 5285
rect 23085 5265 23100 5285
rect 23050 5235 23100 5265
rect 23050 5215 23065 5235
rect 23085 5215 23100 5235
rect 23050 5185 23100 5215
rect 23050 5165 23065 5185
rect 23085 5165 23100 5185
rect 23050 5135 23100 5165
rect 23050 5115 23065 5135
rect 23085 5115 23100 5135
rect 23050 5085 23100 5115
rect 23050 5065 23065 5085
rect 23085 5065 23100 5085
rect 23050 5035 23100 5065
rect 23050 5015 23065 5035
rect 23085 5015 23100 5035
rect 23050 5000 23100 5015
rect 23500 5485 23550 5500
rect 23500 5465 23515 5485
rect 23535 5465 23550 5485
rect 23500 5435 23550 5465
rect 23500 5415 23515 5435
rect 23535 5415 23550 5435
rect 23500 5385 23550 5415
rect 23500 5365 23515 5385
rect 23535 5365 23550 5385
rect 23500 5335 23550 5365
rect 23500 5315 23515 5335
rect 23535 5315 23550 5335
rect 23500 5285 23550 5315
rect 23500 5265 23515 5285
rect 23535 5265 23550 5285
rect 23500 5235 23550 5265
rect 23500 5215 23515 5235
rect 23535 5215 23550 5235
rect 23500 5185 23550 5215
rect 23500 5165 23515 5185
rect 23535 5165 23550 5185
rect 23500 5135 23550 5165
rect 23500 5115 23515 5135
rect 23535 5115 23550 5135
rect 23500 5085 23550 5115
rect 23500 5065 23515 5085
rect 23535 5065 23550 5085
rect 23500 5035 23550 5065
rect 23500 5015 23515 5035
rect 23535 5015 23550 5035
rect 23500 5000 23550 5015
rect 23950 5485 24000 5500
rect 23950 5465 23965 5485
rect 23985 5465 24000 5485
rect 23950 5435 24000 5465
rect 23950 5415 23965 5435
rect 23985 5415 24000 5435
rect 23950 5385 24000 5415
rect 23950 5365 23965 5385
rect 23985 5365 24000 5385
rect 23950 5335 24000 5365
rect 23950 5315 23965 5335
rect 23985 5315 24000 5335
rect 23950 5285 24000 5315
rect 23950 5265 23965 5285
rect 23985 5265 24000 5285
rect 23950 5235 24000 5265
rect 23950 5215 23965 5235
rect 23985 5215 24000 5235
rect 23950 5185 24000 5215
rect 23950 5165 23965 5185
rect 23985 5165 24000 5185
rect 23950 5135 24000 5165
rect 23950 5115 23965 5135
rect 23985 5115 24000 5135
rect 23950 5085 24000 5115
rect 23950 5065 23965 5085
rect 23985 5065 24000 5085
rect 23950 5035 24000 5065
rect 23950 5015 23965 5035
rect 23985 5015 24000 5035
rect 23950 5000 24000 5015
rect 24550 5485 24600 5500
rect 24550 5465 24565 5485
rect 24585 5465 24600 5485
rect 24550 5435 24600 5465
rect 24550 5415 24565 5435
rect 24585 5415 24600 5435
rect 24550 5385 24600 5415
rect 24550 5365 24565 5385
rect 24585 5365 24600 5385
rect 24550 5335 24600 5365
rect 24550 5315 24565 5335
rect 24585 5315 24600 5335
rect 24550 5285 24600 5315
rect 24550 5265 24565 5285
rect 24585 5265 24600 5285
rect 24550 5235 24600 5265
rect 24550 5215 24565 5235
rect 24585 5215 24600 5235
rect 24550 5185 24600 5215
rect 24550 5165 24565 5185
rect 24585 5165 24600 5185
rect 24550 5135 24600 5165
rect 24550 5115 24565 5135
rect 24585 5115 24600 5135
rect 24550 5085 24600 5115
rect 24550 5065 24565 5085
rect 24585 5065 24600 5085
rect 24550 5035 24600 5065
rect 24550 5015 24565 5035
rect 24585 5015 24600 5035
rect 24550 5000 24600 5015
rect 25150 5485 25200 5500
rect 25150 5465 25165 5485
rect 25185 5465 25200 5485
rect 25150 5435 25200 5465
rect 25150 5415 25165 5435
rect 25185 5415 25200 5435
rect 25150 5385 25200 5415
rect 25150 5365 25165 5385
rect 25185 5365 25200 5385
rect 25150 5335 25200 5365
rect 25150 5315 25165 5335
rect 25185 5315 25200 5335
rect 25150 5285 25200 5315
rect 25150 5265 25165 5285
rect 25185 5265 25200 5285
rect 25150 5235 25200 5265
rect 25150 5215 25165 5235
rect 25185 5215 25200 5235
rect 25150 5185 25200 5215
rect 25150 5165 25165 5185
rect 25185 5165 25200 5185
rect 25150 5135 25200 5165
rect 25150 5115 25165 5135
rect 25185 5115 25200 5135
rect 25150 5085 25200 5115
rect 25150 5065 25165 5085
rect 25185 5065 25200 5085
rect 25150 5035 25200 5065
rect 25150 5015 25165 5035
rect 25185 5015 25200 5035
rect 25150 5000 25200 5015
rect 25600 5485 25650 5500
rect 25600 5465 25615 5485
rect 25635 5465 25650 5485
rect 25600 5435 25650 5465
rect 25600 5415 25615 5435
rect 25635 5415 25650 5435
rect 25600 5385 25650 5415
rect 25600 5365 25615 5385
rect 25635 5365 25650 5385
rect 25600 5335 25650 5365
rect 25600 5315 25615 5335
rect 25635 5315 25650 5335
rect 25600 5285 25650 5315
rect 25600 5265 25615 5285
rect 25635 5265 25650 5285
rect 25600 5235 25650 5265
rect 25600 5215 25615 5235
rect 25635 5215 25650 5235
rect 25600 5185 25650 5215
rect 25600 5165 25615 5185
rect 25635 5165 25650 5185
rect 25600 5135 25650 5165
rect 25600 5115 25615 5135
rect 25635 5115 25650 5135
rect 25600 5085 25650 5115
rect 25600 5065 25615 5085
rect 25635 5065 25650 5085
rect 25600 5035 25650 5065
rect 25600 5015 25615 5035
rect 25635 5015 25650 5035
rect 25600 5000 25650 5015
rect 26050 5485 26100 5500
rect 26050 5465 26065 5485
rect 26085 5465 26100 5485
rect 26050 5435 26100 5465
rect 26050 5415 26065 5435
rect 26085 5415 26100 5435
rect 26050 5385 26100 5415
rect 26050 5365 26065 5385
rect 26085 5365 26100 5385
rect 26050 5335 26100 5365
rect 26050 5315 26065 5335
rect 26085 5315 26100 5335
rect 26050 5285 26100 5315
rect 26050 5265 26065 5285
rect 26085 5265 26100 5285
rect 26050 5235 26100 5265
rect 26050 5215 26065 5235
rect 26085 5215 26100 5235
rect 26050 5185 26100 5215
rect 26050 5165 26065 5185
rect 26085 5165 26100 5185
rect 26050 5135 26100 5165
rect 26050 5115 26065 5135
rect 26085 5115 26100 5135
rect 26050 5085 26100 5115
rect 26050 5065 26065 5085
rect 26085 5065 26100 5085
rect 26050 5035 26100 5065
rect 26050 5015 26065 5035
rect 26085 5015 26100 5035
rect 26050 5000 26100 5015
rect 26650 5485 26700 5500
rect 26650 5465 26665 5485
rect 26685 5465 26700 5485
rect 26650 5435 26700 5465
rect 26650 5415 26665 5435
rect 26685 5415 26700 5435
rect 26650 5385 26700 5415
rect 26650 5365 26665 5385
rect 26685 5365 26700 5385
rect 26650 5335 26700 5365
rect 26650 5315 26665 5335
rect 26685 5315 26700 5335
rect 26650 5285 26700 5315
rect 26650 5265 26665 5285
rect 26685 5265 26700 5285
rect 26650 5235 26700 5265
rect 26650 5215 26665 5235
rect 26685 5215 26700 5235
rect 26650 5185 26700 5215
rect 26650 5165 26665 5185
rect 26685 5165 26700 5185
rect 26650 5135 26700 5165
rect 26650 5115 26665 5135
rect 26685 5115 26700 5135
rect 26650 5085 26700 5115
rect 26650 5065 26665 5085
rect 26685 5065 26700 5085
rect 26650 5035 26700 5065
rect 26650 5015 26665 5035
rect 26685 5015 26700 5035
rect 26650 5000 26700 5015
rect 27250 5485 27300 5500
rect 27250 5465 27265 5485
rect 27285 5465 27300 5485
rect 27250 5435 27300 5465
rect 27250 5415 27265 5435
rect 27285 5415 27300 5435
rect 27250 5385 27300 5415
rect 27250 5365 27265 5385
rect 27285 5365 27300 5385
rect 27250 5335 27300 5365
rect 27250 5315 27265 5335
rect 27285 5315 27300 5335
rect 27250 5285 27300 5315
rect 27250 5265 27265 5285
rect 27285 5265 27300 5285
rect 27250 5235 27300 5265
rect 27250 5215 27265 5235
rect 27285 5215 27300 5235
rect 27250 5185 27300 5215
rect 27250 5165 27265 5185
rect 27285 5165 27300 5185
rect 27250 5135 27300 5165
rect 27250 5115 27265 5135
rect 27285 5115 27300 5135
rect 27250 5085 27300 5115
rect 27250 5065 27265 5085
rect 27285 5065 27300 5085
rect 27250 5035 27300 5065
rect 27250 5015 27265 5035
rect 27285 5015 27300 5035
rect 27250 5000 27300 5015
rect 27700 5485 27750 5500
rect 27700 5465 27715 5485
rect 27735 5465 27750 5485
rect 27700 5435 27750 5465
rect 27700 5415 27715 5435
rect 27735 5415 27750 5435
rect 27700 5385 27750 5415
rect 27700 5365 27715 5385
rect 27735 5365 27750 5385
rect 27700 5335 27750 5365
rect 27700 5315 27715 5335
rect 27735 5315 27750 5335
rect 27700 5285 27750 5315
rect 27700 5265 27715 5285
rect 27735 5265 27750 5285
rect 27700 5235 27750 5265
rect 27700 5215 27715 5235
rect 27735 5215 27750 5235
rect 27700 5185 27750 5215
rect 27700 5165 27715 5185
rect 27735 5165 27750 5185
rect 27700 5135 27750 5165
rect 27700 5115 27715 5135
rect 27735 5115 27750 5135
rect 27700 5085 27750 5115
rect 27700 5065 27715 5085
rect 27735 5065 27750 5085
rect 27700 5035 27750 5065
rect 27700 5015 27715 5035
rect 27735 5015 27750 5035
rect 27700 5000 27750 5015
rect 28150 5485 28200 5500
rect 28150 5465 28165 5485
rect 28185 5465 28200 5485
rect 28150 5435 28200 5465
rect 28150 5415 28165 5435
rect 28185 5415 28200 5435
rect 28150 5385 28200 5415
rect 28150 5365 28165 5385
rect 28185 5365 28200 5385
rect 28150 5335 28200 5365
rect 28150 5315 28165 5335
rect 28185 5315 28200 5335
rect 28150 5285 28200 5315
rect 28150 5265 28165 5285
rect 28185 5265 28200 5285
rect 28150 5235 28200 5265
rect 28150 5215 28165 5235
rect 28185 5215 28200 5235
rect 28150 5185 28200 5215
rect 28150 5165 28165 5185
rect 28185 5165 28200 5185
rect 28150 5135 28200 5165
rect 28150 5115 28165 5135
rect 28185 5115 28200 5135
rect 28150 5085 28200 5115
rect 28150 5065 28165 5085
rect 28185 5065 28200 5085
rect 28150 5035 28200 5065
rect 28150 5015 28165 5035
rect 28185 5015 28200 5035
rect 28150 5000 28200 5015
rect 28750 5485 28800 5500
rect 28750 5465 28765 5485
rect 28785 5465 28800 5485
rect 28750 5435 28800 5465
rect 28750 5415 28765 5435
rect 28785 5415 28800 5435
rect 28750 5385 28800 5415
rect 28750 5365 28765 5385
rect 28785 5365 28800 5385
rect 28750 5335 28800 5365
rect 28750 5315 28765 5335
rect 28785 5315 28800 5335
rect 28750 5285 28800 5315
rect 28750 5265 28765 5285
rect 28785 5265 28800 5285
rect 28750 5235 28800 5265
rect 28750 5215 28765 5235
rect 28785 5215 28800 5235
rect 28750 5185 28800 5215
rect 28750 5165 28765 5185
rect 28785 5165 28800 5185
rect 28750 5135 28800 5165
rect 28750 5115 28765 5135
rect 28785 5115 28800 5135
rect 28750 5085 28800 5115
rect 28750 5065 28765 5085
rect 28785 5065 28800 5085
rect 28750 5035 28800 5065
rect 28750 5015 28765 5035
rect 28785 5015 28800 5035
rect 28750 5000 28800 5015
rect 29350 5485 29400 5500
rect 29350 5465 29365 5485
rect 29385 5465 29400 5485
rect 29350 5435 29400 5465
rect 29350 5415 29365 5435
rect 29385 5415 29400 5435
rect 29350 5385 29400 5415
rect 29350 5365 29365 5385
rect 29385 5365 29400 5385
rect 29350 5335 29400 5365
rect 29350 5315 29365 5335
rect 29385 5315 29400 5335
rect 29350 5285 29400 5315
rect 29350 5265 29365 5285
rect 29385 5265 29400 5285
rect 29350 5235 29400 5265
rect 29350 5215 29365 5235
rect 29385 5215 29400 5235
rect 29350 5185 29400 5215
rect 29350 5165 29365 5185
rect 29385 5165 29400 5185
rect 29350 5135 29400 5165
rect 29350 5115 29365 5135
rect 29385 5115 29400 5135
rect 29350 5085 29400 5115
rect 29350 5065 29365 5085
rect 29385 5065 29400 5085
rect 29350 5035 29400 5065
rect 29350 5015 29365 5035
rect 29385 5015 29400 5035
rect 29350 5000 29400 5015
rect 29500 5485 29550 5500
rect 29500 5465 29515 5485
rect 29535 5465 29550 5485
rect 29500 5435 29550 5465
rect 29500 5415 29515 5435
rect 29535 5415 29550 5435
rect 29500 5385 29550 5415
rect 29500 5365 29515 5385
rect 29535 5365 29550 5385
rect 29500 5335 29550 5365
rect 29500 5315 29515 5335
rect 29535 5315 29550 5335
rect 29500 5285 29550 5315
rect 29500 5265 29515 5285
rect 29535 5265 29550 5285
rect 29500 5235 29550 5265
rect 29500 5215 29515 5235
rect 29535 5215 29550 5235
rect 29500 5185 29550 5215
rect 29500 5165 29515 5185
rect 29535 5165 29550 5185
rect 29500 5135 29550 5165
rect 29500 5115 29515 5135
rect 29535 5115 29550 5135
rect 29500 5085 29550 5115
rect 29500 5065 29515 5085
rect 29535 5065 29550 5085
rect 29500 5035 29550 5065
rect 29500 5015 29515 5035
rect 29535 5015 29550 5035
rect 29500 5000 29550 5015
rect 29650 5485 29700 5500
rect 29650 5465 29665 5485
rect 29685 5465 29700 5485
rect 29650 5435 29700 5465
rect 29650 5415 29665 5435
rect 29685 5415 29700 5435
rect 29650 5385 29700 5415
rect 29650 5365 29665 5385
rect 29685 5365 29700 5385
rect 29650 5335 29700 5365
rect 29650 5315 29665 5335
rect 29685 5315 29700 5335
rect 29650 5285 29700 5315
rect 29650 5265 29665 5285
rect 29685 5265 29700 5285
rect 29650 5235 29700 5265
rect 29650 5215 29665 5235
rect 29685 5215 29700 5235
rect 29650 5185 29700 5215
rect 29650 5165 29665 5185
rect 29685 5165 29700 5185
rect 29650 5135 29700 5165
rect 29650 5115 29665 5135
rect 29685 5115 29700 5135
rect 29650 5085 29700 5115
rect 29650 5065 29665 5085
rect 29685 5065 29700 5085
rect 29650 5035 29700 5065
rect 29650 5015 29665 5035
rect 29685 5015 29700 5035
rect 29650 5000 29700 5015
rect 29800 5485 29850 5500
rect 29800 5465 29815 5485
rect 29835 5465 29850 5485
rect 29800 5435 29850 5465
rect 29800 5415 29815 5435
rect 29835 5415 29850 5435
rect 29800 5385 29850 5415
rect 29800 5365 29815 5385
rect 29835 5365 29850 5385
rect 29800 5335 29850 5365
rect 29800 5315 29815 5335
rect 29835 5315 29850 5335
rect 29800 5285 29850 5315
rect 29800 5265 29815 5285
rect 29835 5265 29850 5285
rect 29800 5235 29850 5265
rect 29800 5215 29815 5235
rect 29835 5215 29850 5235
rect 29800 5185 29850 5215
rect 29800 5165 29815 5185
rect 29835 5165 29850 5185
rect 29800 5135 29850 5165
rect 29800 5115 29815 5135
rect 29835 5115 29850 5135
rect 29800 5085 29850 5115
rect 29800 5065 29815 5085
rect 29835 5065 29850 5085
rect 29800 5035 29850 5065
rect 29800 5015 29815 5035
rect 29835 5015 29850 5035
rect 29800 5000 29850 5015
rect 29950 5485 30000 5500
rect 29950 5465 29965 5485
rect 29985 5465 30000 5485
rect 29950 5435 30000 5465
rect 29950 5415 29965 5435
rect 29985 5415 30000 5435
rect 29950 5385 30000 5415
rect 29950 5365 29965 5385
rect 29985 5365 30000 5385
rect 29950 5335 30000 5365
rect 29950 5315 29965 5335
rect 29985 5315 30000 5335
rect 29950 5285 30000 5315
rect 29950 5265 29965 5285
rect 29985 5265 30000 5285
rect 29950 5235 30000 5265
rect 29950 5215 29965 5235
rect 29985 5215 30000 5235
rect 29950 5185 30000 5215
rect 29950 5165 29965 5185
rect 29985 5165 30000 5185
rect 29950 5135 30000 5165
rect 29950 5115 29965 5135
rect 29985 5115 30000 5135
rect 29950 5085 30000 5115
rect 29950 5065 29965 5085
rect 29985 5065 30000 5085
rect 29950 5035 30000 5065
rect 29950 5015 29965 5035
rect 29985 5015 30000 5035
rect 29950 5000 30000 5015
rect 30100 5485 30150 5500
rect 30100 5465 30115 5485
rect 30135 5465 30150 5485
rect 30100 5435 30150 5465
rect 30100 5415 30115 5435
rect 30135 5415 30150 5435
rect 30100 5385 30150 5415
rect 30100 5365 30115 5385
rect 30135 5365 30150 5385
rect 30100 5335 30150 5365
rect 30100 5315 30115 5335
rect 30135 5315 30150 5335
rect 30100 5285 30150 5315
rect 30100 5265 30115 5285
rect 30135 5265 30150 5285
rect 30100 5235 30150 5265
rect 30100 5215 30115 5235
rect 30135 5215 30150 5235
rect 30100 5185 30150 5215
rect 30100 5165 30115 5185
rect 30135 5165 30150 5185
rect 30100 5135 30150 5165
rect 30100 5115 30115 5135
rect 30135 5115 30150 5135
rect 30100 5085 30150 5115
rect 30100 5065 30115 5085
rect 30135 5065 30150 5085
rect 30100 5035 30150 5065
rect 30100 5015 30115 5035
rect 30135 5015 30150 5035
rect 30100 5000 30150 5015
rect 30250 5485 30300 5500
rect 30250 5465 30265 5485
rect 30285 5465 30300 5485
rect 30250 5435 30300 5465
rect 30250 5415 30265 5435
rect 30285 5415 30300 5435
rect 30250 5385 30300 5415
rect 30250 5365 30265 5385
rect 30285 5365 30300 5385
rect 30250 5335 30300 5365
rect 30250 5315 30265 5335
rect 30285 5315 30300 5335
rect 30250 5285 30300 5315
rect 30250 5265 30265 5285
rect 30285 5265 30300 5285
rect 30250 5235 30300 5265
rect 30250 5215 30265 5235
rect 30285 5215 30300 5235
rect 30250 5185 30300 5215
rect 30250 5165 30265 5185
rect 30285 5165 30300 5185
rect 30250 5135 30300 5165
rect 30250 5115 30265 5135
rect 30285 5115 30300 5135
rect 30250 5085 30300 5115
rect 30250 5065 30265 5085
rect 30285 5065 30300 5085
rect 30250 5035 30300 5065
rect 30250 5015 30265 5035
rect 30285 5015 30300 5035
rect 30250 5000 30300 5015
rect 30400 5485 30450 5500
rect 30400 5465 30415 5485
rect 30435 5465 30450 5485
rect 30400 5435 30450 5465
rect 30400 5415 30415 5435
rect 30435 5415 30450 5435
rect 30400 5385 30450 5415
rect 30400 5365 30415 5385
rect 30435 5365 30450 5385
rect 30400 5335 30450 5365
rect 30400 5315 30415 5335
rect 30435 5315 30450 5335
rect 30400 5285 30450 5315
rect 30400 5265 30415 5285
rect 30435 5265 30450 5285
rect 30400 5235 30450 5265
rect 30400 5215 30415 5235
rect 30435 5215 30450 5235
rect 30400 5185 30450 5215
rect 30400 5165 30415 5185
rect 30435 5165 30450 5185
rect 30400 5135 30450 5165
rect 30400 5115 30415 5135
rect 30435 5115 30450 5135
rect 30400 5085 30450 5115
rect 30400 5065 30415 5085
rect 30435 5065 30450 5085
rect 30400 5035 30450 5065
rect 30400 5015 30415 5035
rect 30435 5015 30450 5035
rect 30400 5000 30450 5015
rect 30550 5485 30600 5500
rect 30550 5465 30565 5485
rect 30585 5465 30600 5485
rect 30550 5435 30600 5465
rect 30550 5415 30565 5435
rect 30585 5415 30600 5435
rect 30550 5385 30600 5415
rect 30550 5365 30565 5385
rect 30585 5365 30600 5385
rect 30550 5335 30600 5365
rect 30550 5315 30565 5335
rect 30585 5315 30600 5335
rect 30550 5285 30600 5315
rect 30550 5265 30565 5285
rect 30585 5265 30600 5285
rect 30550 5235 30600 5265
rect 30550 5215 30565 5235
rect 30585 5215 30600 5235
rect 30550 5185 30600 5215
rect 30550 5165 30565 5185
rect 30585 5165 30600 5185
rect 30550 5135 30600 5165
rect 30550 5115 30565 5135
rect 30585 5115 30600 5135
rect 30550 5085 30600 5115
rect 30550 5065 30565 5085
rect 30585 5065 30600 5085
rect 30550 5035 30600 5065
rect 30550 5015 30565 5035
rect 30585 5015 30600 5035
rect 30550 5000 30600 5015
rect 30700 5485 30750 5500
rect 30700 5465 30715 5485
rect 30735 5465 30750 5485
rect 30700 5435 30750 5465
rect 30700 5415 30715 5435
rect 30735 5415 30750 5435
rect 30700 5385 30750 5415
rect 30700 5365 30715 5385
rect 30735 5365 30750 5385
rect 30700 5335 30750 5365
rect 30700 5315 30715 5335
rect 30735 5315 30750 5335
rect 30700 5285 30750 5315
rect 30700 5265 30715 5285
rect 30735 5265 30750 5285
rect 30700 5235 30750 5265
rect 30700 5215 30715 5235
rect 30735 5215 30750 5235
rect 30700 5185 30750 5215
rect 30700 5165 30715 5185
rect 30735 5165 30750 5185
rect 30700 5135 30750 5165
rect 30700 5115 30715 5135
rect 30735 5115 30750 5135
rect 30700 5085 30750 5115
rect 30700 5065 30715 5085
rect 30735 5065 30750 5085
rect 30700 5035 30750 5065
rect 30700 5015 30715 5035
rect 30735 5015 30750 5035
rect 30700 5000 30750 5015
rect 30850 5485 30900 5500
rect 30850 5465 30865 5485
rect 30885 5465 30900 5485
rect 30850 5435 30900 5465
rect 30850 5415 30865 5435
rect 30885 5415 30900 5435
rect 30850 5385 30900 5415
rect 30850 5365 30865 5385
rect 30885 5365 30900 5385
rect 30850 5335 30900 5365
rect 30850 5315 30865 5335
rect 30885 5315 30900 5335
rect 30850 5285 30900 5315
rect 30850 5265 30865 5285
rect 30885 5265 30900 5285
rect 30850 5235 30900 5265
rect 30850 5215 30865 5235
rect 30885 5215 30900 5235
rect 30850 5185 30900 5215
rect 30850 5165 30865 5185
rect 30885 5165 30900 5185
rect 30850 5135 30900 5165
rect 30850 5115 30865 5135
rect 30885 5115 30900 5135
rect 30850 5085 30900 5115
rect 30850 5065 30865 5085
rect 30885 5065 30900 5085
rect 30850 5035 30900 5065
rect 30850 5015 30865 5035
rect 30885 5015 30900 5035
rect 30850 5000 30900 5015
rect 31000 5485 31050 5500
rect 31000 5465 31015 5485
rect 31035 5465 31050 5485
rect 31000 5435 31050 5465
rect 31000 5415 31015 5435
rect 31035 5415 31050 5435
rect 31000 5385 31050 5415
rect 31000 5365 31015 5385
rect 31035 5365 31050 5385
rect 31000 5335 31050 5365
rect 31000 5315 31015 5335
rect 31035 5315 31050 5335
rect 31000 5285 31050 5315
rect 31000 5265 31015 5285
rect 31035 5265 31050 5285
rect 31000 5235 31050 5265
rect 31000 5215 31015 5235
rect 31035 5215 31050 5235
rect 31000 5185 31050 5215
rect 31000 5165 31015 5185
rect 31035 5165 31050 5185
rect 31000 5135 31050 5165
rect 31000 5115 31015 5135
rect 31035 5115 31050 5135
rect 31000 5085 31050 5115
rect 31000 5065 31015 5085
rect 31035 5065 31050 5085
rect 31000 5035 31050 5065
rect 31000 5015 31015 5035
rect 31035 5015 31050 5035
rect 31000 5000 31050 5015
rect 31150 5485 31200 5500
rect 31150 5465 31165 5485
rect 31185 5465 31200 5485
rect 31150 5435 31200 5465
rect 31150 5415 31165 5435
rect 31185 5415 31200 5435
rect 31150 5385 31200 5415
rect 31150 5365 31165 5385
rect 31185 5365 31200 5385
rect 31150 5335 31200 5365
rect 31150 5315 31165 5335
rect 31185 5315 31200 5335
rect 31150 5285 31200 5315
rect 31150 5265 31165 5285
rect 31185 5265 31200 5285
rect 31150 5235 31200 5265
rect 31150 5215 31165 5235
rect 31185 5215 31200 5235
rect 31150 5185 31200 5215
rect 31150 5165 31165 5185
rect 31185 5165 31200 5185
rect 31150 5135 31200 5165
rect 31150 5115 31165 5135
rect 31185 5115 31200 5135
rect 31150 5085 31200 5115
rect 31150 5065 31165 5085
rect 31185 5065 31200 5085
rect 31150 5035 31200 5065
rect 31150 5015 31165 5035
rect 31185 5015 31200 5035
rect 31150 5000 31200 5015
rect 31300 5485 31350 5500
rect 31300 5465 31315 5485
rect 31335 5465 31350 5485
rect 31300 5435 31350 5465
rect 31300 5415 31315 5435
rect 31335 5415 31350 5435
rect 31300 5385 31350 5415
rect 31300 5365 31315 5385
rect 31335 5365 31350 5385
rect 31300 5335 31350 5365
rect 31300 5315 31315 5335
rect 31335 5315 31350 5335
rect 31300 5285 31350 5315
rect 31300 5265 31315 5285
rect 31335 5265 31350 5285
rect 31300 5235 31350 5265
rect 31300 5215 31315 5235
rect 31335 5215 31350 5235
rect 31300 5185 31350 5215
rect 31300 5165 31315 5185
rect 31335 5165 31350 5185
rect 31300 5135 31350 5165
rect 31300 5115 31315 5135
rect 31335 5115 31350 5135
rect 31300 5085 31350 5115
rect 31300 5065 31315 5085
rect 31335 5065 31350 5085
rect 31300 5035 31350 5065
rect 31300 5015 31315 5035
rect 31335 5015 31350 5035
rect 31300 5000 31350 5015
rect 31450 5485 31500 5500
rect 31450 5465 31465 5485
rect 31485 5465 31500 5485
rect 31450 5435 31500 5465
rect 31450 5415 31465 5435
rect 31485 5415 31500 5435
rect 31450 5385 31500 5415
rect 31450 5365 31465 5385
rect 31485 5365 31500 5385
rect 31450 5335 31500 5365
rect 31450 5315 31465 5335
rect 31485 5315 31500 5335
rect 31450 5285 31500 5315
rect 31450 5265 31465 5285
rect 31485 5265 31500 5285
rect 31450 5235 31500 5265
rect 31450 5215 31465 5235
rect 31485 5215 31500 5235
rect 31450 5185 31500 5215
rect 31450 5165 31465 5185
rect 31485 5165 31500 5185
rect 31450 5135 31500 5165
rect 31450 5115 31465 5135
rect 31485 5115 31500 5135
rect 31450 5085 31500 5115
rect 31450 5065 31465 5085
rect 31485 5065 31500 5085
rect 31450 5035 31500 5065
rect 31450 5015 31465 5035
rect 31485 5015 31500 5035
rect 31450 5000 31500 5015
rect 32050 5485 32100 5500
rect 32050 5465 32065 5485
rect 32085 5465 32100 5485
rect 32050 5435 32100 5465
rect 32050 5415 32065 5435
rect 32085 5415 32100 5435
rect 32050 5385 32100 5415
rect 32050 5365 32065 5385
rect 32085 5365 32100 5385
rect 32050 5335 32100 5365
rect 32050 5315 32065 5335
rect 32085 5315 32100 5335
rect 32050 5285 32100 5315
rect 32050 5265 32065 5285
rect 32085 5265 32100 5285
rect 32050 5235 32100 5265
rect 32050 5215 32065 5235
rect 32085 5215 32100 5235
rect 32050 5185 32100 5215
rect 32050 5165 32065 5185
rect 32085 5165 32100 5185
rect 32050 5135 32100 5165
rect 32050 5115 32065 5135
rect 32085 5115 32100 5135
rect 32050 5085 32100 5115
rect 32050 5065 32065 5085
rect 32085 5065 32100 5085
rect 32050 5035 32100 5065
rect 32050 5015 32065 5035
rect 32085 5015 32100 5035
rect 32050 5000 32100 5015
rect -600 4935 -350 4950
rect -600 4915 -585 4935
rect -565 4915 -535 4935
rect -515 4915 -485 4935
rect -465 4915 -435 4935
rect -415 4915 -385 4935
rect -365 4915 -350 4935
rect -600 4900 -350 4915
rect -300 4935 -50 4950
rect -300 4915 -285 4935
rect -265 4915 -235 4935
rect -215 4915 -185 4935
rect -165 4915 -135 4935
rect -115 4915 -85 4935
rect -65 4915 -50 4935
rect -300 4900 -50 4915
rect 0 4935 250 4950
rect 0 4915 15 4935
rect 35 4915 65 4935
rect 85 4915 115 4935
rect 135 4915 165 4935
rect 185 4915 215 4935
rect 235 4915 250 4935
rect 0 4900 250 4915
rect 300 4935 550 4950
rect 300 4915 315 4935
rect 335 4915 365 4935
rect 385 4915 415 4935
rect 435 4915 465 4935
rect 485 4915 515 4935
rect 535 4915 550 4935
rect 300 4900 550 4915
rect 600 4935 850 4950
rect 600 4915 615 4935
rect 635 4915 665 4935
rect 685 4915 715 4935
rect 735 4915 765 4935
rect 785 4915 815 4935
rect 835 4915 850 4935
rect 600 4900 850 4915
rect 900 4935 1150 4950
rect 900 4915 915 4935
rect 935 4915 965 4935
rect 985 4915 1015 4935
rect 1035 4915 1065 4935
rect 1085 4915 1115 4935
rect 1135 4915 1150 4935
rect 900 4900 1150 4915
rect 1200 4935 1450 4950
rect 1200 4915 1215 4935
rect 1235 4915 1265 4935
rect 1285 4915 1315 4935
rect 1335 4915 1365 4935
rect 1385 4915 1415 4935
rect 1435 4915 1450 4935
rect 1200 4900 1450 4915
rect 1500 4935 1750 4950
rect 1500 4915 1515 4935
rect 1535 4915 1565 4935
rect 1585 4915 1615 4935
rect 1635 4915 1665 4935
rect 1685 4915 1715 4935
rect 1735 4915 1750 4935
rect 1500 4900 1750 4915
rect 1800 4935 2050 4950
rect 1800 4915 1815 4935
rect 1835 4915 1865 4935
rect 1885 4915 1915 4935
rect 1935 4915 1965 4935
rect 1985 4915 2015 4935
rect 2035 4915 2050 4935
rect 1800 4900 2050 4915
rect 2100 4935 2350 4950
rect 2100 4915 2115 4935
rect 2135 4915 2165 4935
rect 2185 4915 2215 4935
rect 2235 4915 2265 4935
rect 2285 4915 2315 4935
rect 2335 4915 2350 4935
rect 2100 4900 2350 4915
rect 2400 4935 2650 4950
rect 2400 4915 2415 4935
rect 2435 4915 2465 4935
rect 2485 4915 2515 4935
rect 2535 4915 2565 4935
rect 2585 4915 2615 4935
rect 2635 4915 2650 4935
rect 2400 4900 2650 4915
rect 2700 4935 2950 4950
rect 2700 4915 2715 4935
rect 2735 4915 2765 4935
rect 2785 4915 2815 4935
rect 2835 4915 2865 4935
rect 2885 4915 2915 4935
rect 2935 4915 2950 4935
rect 2700 4900 2950 4915
rect 3000 4935 3250 4950
rect 3000 4915 3015 4935
rect 3035 4915 3065 4935
rect 3085 4915 3115 4935
rect 3135 4915 3165 4935
rect 3185 4915 3215 4935
rect 3235 4915 3250 4935
rect 3000 4900 3250 4915
rect 3300 4935 3550 4950
rect 3300 4915 3315 4935
rect 3335 4915 3365 4935
rect 3385 4915 3415 4935
rect 3435 4915 3465 4935
rect 3485 4915 3515 4935
rect 3535 4915 3550 4935
rect 3300 4900 3550 4915
rect 3600 4935 3850 4950
rect 3600 4915 3615 4935
rect 3635 4915 3665 4935
rect 3685 4915 3715 4935
rect 3735 4915 3765 4935
rect 3785 4915 3815 4935
rect 3835 4915 3850 4935
rect 3600 4900 3850 4915
rect 3900 4935 4150 4950
rect 3900 4915 3915 4935
rect 3935 4915 3965 4935
rect 3985 4915 4015 4935
rect 4035 4915 4065 4935
rect 4085 4915 4115 4935
rect 4135 4915 4150 4935
rect 3900 4900 4150 4915
rect 4200 4935 4450 4950
rect 4200 4915 4215 4935
rect 4235 4915 4265 4935
rect 4285 4915 4315 4935
rect 4335 4915 4365 4935
rect 4385 4915 4415 4935
rect 4435 4915 4450 4935
rect 4200 4900 4450 4915
rect 4500 4935 4750 4950
rect 4500 4915 4515 4935
rect 4535 4915 4565 4935
rect 4585 4915 4615 4935
rect 4635 4915 4665 4935
rect 4685 4915 4715 4935
rect 4735 4915 4750 4935
rect 4500 4900 4750 4915
rect 4800 4935 5050 4950
rect 4800 4915 4815 4935
rect 4835 4915 4865 4935
rect 4885 4915 4915 4935
rect 4935 4915 4965 4935
rect 4985 4915 5015 4935
rect 5035 4915 5050 4935
rect 4800 4900 5050 4915
rect 5100 4935 5350 4950
rect 5100 4915 5115 4935
rect 5135 4915 5165 4935
rect 5185 4915 5215 4935
rect 5235 4915 5265 4935
rect 5285 4915 5315 4935
rect 5335 4915 5350 4935
rect 5100 4900 5350 4915
rect 5400 4935 5650 4950
rect 5400 4915 5415 4935
rect 5435 4915 5465 4935
rect 5485 4915 5515 4935
rect 5535 4915 5565 4935
rect 5585 4915 5615 4935
rect 5635 4915 5650 4935
rect 5400 4900 5650 4915
rect 5700 4935 5950 4950
rect 5700 4915 5715 4935
rect 5735 4915 5765 4935
rect 5785 4915 5815 4935
rect 5835 4915 5865 4935
rect 5885 4915 5915 4935
rect 5935 4915 5950 4935
rect 5700 4900 5950 4915
rect 6000 4935 6250 4950
rect 6000 4915 6015 4935
rect 6035 4915 6065 4935
rect 6085 4915 6115 4935
rect 6135 4915 6165 4935
rect 6185 4915 6215 4935
rect 6235 4915 6250 4935
rect 6000 4900 6250 4915
rect 6300 4935 6550 4950
rect 6300 4915 6315 4935
rect 6335 4915 6365 4935
rect 6385 4915 6415 4935
rect 6435 4915 6465 4935
rect 6485 4915 6515 4935
rect 6535 4915 6550 4935
rect 6300 4900 6550 4915
rect 6600 4935 6850 4950
rect 6600 4915 6615 4935
rect 6635 4915 6665 4935
rect 6685 4915 6715 4935
rect 6735 4915 6765 4935
rect 6785 4915 6815 4935
rect 6835 4915 6850 4935
rect 6600 4900 6850 4915
rect 6900 4935 7150 4950
rect 6900 4915 6915 4935
rect 6935 4915 6965 4935
rect 6985 4915 7015 4935
rect 7035 4915 7065 4935
rect 7085 4915 7115 4935
rect 7135 4915 7150 4935
rect 6900 4900 7150 4915
rect 7200 4935 7450 4950
rect 7200 4915 7215 4935
rect 7235 4915 7265 4935
rect 7285 4915 7315 4935
rect 7335 4915 7365 4935
rect 7385 4915 7415 4935
rect 7435 4915 7450 4935
rect 7200 4900 7450 4915
rect 7500 4935 7750 4950
rect 7500 4915 7515 4935
rect 7535 4915 7565 4935
rect 7585 4915 7615 4935
rect 7635 4915 7665 4935
rect 7685 4915 7715 4935
rect 7735 4915 7750 4935
rect 7500 4900 7750 4915
rect 7800 4935 8050 4950
rect 7800 4915 7815 4935
rect 7835 4915 7865 4935
rect 7885 4915 7915 4935
rect 7935 4915 7965 4935
rect 7985 4915 8015 4935
rect 8035 4915 8050 4935
rect 7800 4900 8050 4915
rect 8100 4935 8350 4950
rect 8100 4915 8115 4935
rect 8135 4915 8165 4935
rect 8185 4915 8215 4935
rect 8235 4915 8265 4935
rect 8285 4915 8315 4935
rect 8335 4915 8350 4935
rect 8100 4900 8350 4915
rect 8400 4935 10750 4950
rect 8400 4915 8415 4935
rect 8435 4915 8465 4935
rect 8485 4915 8515 4935
rect 8535 4915 8565 4935
rect 8585 4915 8615 4935
rect 8635 4915 8715 4935
rect 8735 4915 8765 4935
rect 8785 4915 8815 4935
rect 8835 4915 8865 4935
rect 8885 4915 8915 4935
rect 8935 4915 9015 4935
rect 9035 4915 9065 4935
rect 9085 4915 9115 4935
rect 9135 4915 9165 4935
rect 9185 4915 9215 4935
rect 9235 4915 9315 4935
rect 9335 4915 9365 4935
rect 9385 4915 9415 4935
rect 9435 4915 9465 4935
rect 9485 4915 9515 4935
rect 9535 4915 9615 4935
rect 9635 4915 9665 4935
rect 9685 4915 9715 4935
rect 9735 4915 9765 4935
rect 9785 4915 9815 4935
rect 9835 4915 9915 4935
rect 9935 4915 9965 4935
rect 9985 4915 10015 4935
rect 10035 4915 10065 4935
rect 10085 4915 10115 4935
rect 10135 4915 10215 4935
rect 10235 4915 10265 4935
rect 10285 4915 10315 4935
rect 10335 4915 10365 4935
rect 10385 4915 10415 4935
rect 10435 4915 10515 4935
rect 10535 4915 10565 4935
rect 10585 4915 10615 4935
rect 10635 4915 10665 4935
rect 10685 4915 10715 4935
rect 10735 4915 10750 4935
rect 8400 4900 10750 4915
rect 10800 4935 11050 4950
rect 10800 4915 10815 4935
rect 10835 4915 10865 4935
rect 10885 4915 10915 4935
rect 10935 4915 10965 4935
rect 10985 4915 11015 4935
rect 11035 4915 11050 4935
rect 10800 4900 11050 4915
rect 11100 4935 11350 4950
rect 11100 4915 11115 4935
rect 11135 4915 11165 4935
rect 11185 4915 11215 4935
rect 11235 4915 11265 4935
rect 11285 4915 11315 4935
rect 11335 4915 11350 4935
rect 11100 4900 11350 4915
rect 11400 4935 11650 4950
rect 11400 4915 11415 4935
rect 11435 4915 11465 4935
rect 11485 4915 11515 4935
rect 11535 4915 11565 4935
rect 11585 4915 11615 4935
rect 11635 4915 11650 4935
rect 11400 4900 11650 4915
rect 11700 4935 11950 4950
rect 11700 4915 11715 4935
rect 11735 4915 11765 4935
rect 11785 4915 11815 4935
rect 11835 4915 11865 4935
rect 11885 4915 11915 4935
rect 11935 4915 11950 4935
rect 11700 4900 11950 4915
rect 12000 4935 12250 4950
rect 12000 4915 12015 4935
rect 12035 4915 12065 4935
rect 12085 4915 12115 4935
rect 12135 4915 12165 4935
rect 12185 4915 12215 4935
rect 12235 4915 12250 4935
rect 12000 4900 12250 4915
rect 12300 4935 12550 4950
rect 12300 4915 12315 4935
rect 12335 4915 12365 4935
rect 12385 4915 12415 4935
rect 12435 4915 12465 4935
rect 12485 4915 12515 4935
rect 12535 4915 12550 4935
rect 12300 4900 12550 4915
rect 12600 4935 12850 4950
rect 12600 4915 12615 4935
rect 12635 4915 12665 4935
rect 12685 4915 12715 4935
rect 12735 4915 12765 4935
rect 12785 4915 12815 4935
rect 12835 4915 12850 4935
rect 12600 4900 12850 4915
rect 12900 4935 13150 4950
rect 12900 4915 12915 4935
rect 12935 4915 12965 4935
rect 12985 4915 13015 4935
rect 13035 4915 13065 4935
rect 13085 4915 13115 4935
rect 13135 4915 13150 4935
rect 12900 4900 13150 4915
rect 13200 4935 13450 4950
rect 13200 4915 13215 4935
rect 13235 4915 13265 4935
rect 13285 4915 13315 4935
rect 13335 4915 13365 4935
rect 13385 4915 13415 4935
rect 13435 4915 13450 4935
rect 13200 4900 13450 4915
rect 13500 4935 13750 4950
rect 13500 4915 13515 4935
rect 13535 4915 13565 4935
rect 13585 4915 13615 4935
rect 13635 4915 13665 4935
rect 13685 4915 13715 4935
rect 13735 4915 13750 4935
rect 13500 4900 13750 4915
rect 13800 4935 14050 4950
rect 13800 4915 13815 4935
rect 13835 4915 13865 4935
rect 13885 4915 13915 4935
rect 13935 4915 13965 4935
rect 13985 4915 14015 4935
rect 14035 4915 14050 4935
rect 13800 4900 14050 4915
rect 14100 4935 14350 4950
rect 14100 4915 14115 4935
rect 14135 4915 14165 4935
rect 14185 4915 14215 4935
rect 14235 4915 14265 4935
rect 14285 4915 14315 4935
rect 14335 4915 14350 4935
rect 14100 4900 14350 4915
rect 14400 4935 14650 4950
rect 14400 4915 14415 4935
rect 14435 4915 14465 4935
rect 14485 4915 14515 4935
rect 14535 4915 14565 4935
rect 14585 4915 14615 4935
rect 14635 4915 14650 4935
rect 14400 4900 14650 4915
rect 14700 4935 14950 4950
rect 14700 4915 14715 4935
rect 14735 4915 14765 4935
rect 14785 4915 14815 4935
rect 14835 4915 14865 4935
rect 14885 4915 14915 4935
rect 14935 4915 14950 4935
rect 14700 4900 14950 4915
rect 15000 4935 15250 4950
rect 15000 4915 15015 4935
rect 15035 4915 15065 4935
rect 15085 4915 15115 4935
rect 15135 4915 15165 4935
rect 15185 4915 15215 4935
rect 15235 4915 15250 4935
rect 15000 4900 15250 4915
rect 15300 4935 15550 4950
rect 15300 4915 15315 4935
rect 15335 4915 15365 4935
rect 15385 4915 15415 4935
rect 15435 4915 15465 4935
rect 15485 4915 15515 4935
rect 15535 4915 15550 4935
rect 15300 4900 15550 4915
rect 15600 4935 15850 4950
rect 15600 4915 15615 4935
rect 15635 4915 15665 4935
rect 15685 4915 15715 4935
rect 15735 4915 15765 4935
rect 15785 4915 15815 4935
rect 15835 4915 15850 4935
rect 15600 4900 15850 4915
rect 15900 4935 16150 4950
rect 15900 4915 15915 4935
rect 15935 4915 15965 4935
rect 15985 4915 16015 4935
rect 16035 4915 16065 4935
rect 16085 4915 16115 4935
rect 16135 4915 16150 4935
rect 15900 4900 16150 4915
rect 16200 4935 16450 4950
rect 16200 4915 16215 4935
rect 16235 4915 16265 4935
rect 16285 4915 16315 4935
rect 16335 4915 16365 4935
rect 16385 4915 16415 4935
rect 16435 4915 16450 4935
rect 16200 4900 16450 4915
rect 16500 4935 16750 4950
rect 16500 4915 16515 4935
rect 16535 4915 16565 4935
rect 16585 4915 16615 4935
rect 16635 4915 16665 4935
rect 16685 4915 16715 4935
rect 16735 4915 16750 4935
rect 16500 4900 16750 4915
rect 16800 4935 17050 4950
rect 16800 4915 16815 4935
rect 16835 4915 16865 4935
rect 16885 4915 16915 4935
rect 16935 4915 16965 4935
rect 16985 4915 17015 4935
rect 17035 4915 17050 4935
rect 16800 4900 17050 4915
rect 17100 4935 17350 4950
rect 17100 4915 17115 4935
rect 17135 4915 17165 4935
rect 17185 4915 17215 4935
rect 17235 4915 17265 4935
rect 17285 4915 17315 4935
rect 17335 4915 17350 4935
rect 17100 4900 17350 4915
rect 17400 4935 17650 4950
rect 17400 4915 17415 4935
rect 17435 4915 17465 4935
rect 17485 4915 17515 4935
rect 17535 4915 17565 4935
rect 17585 4915 17615 4935
rect 17635 4915 17650 4935
rect 17400 4900 17650 4915
rect 17700 4935 17950 4950
rect 17700 4915 17715 4935
rect 17735 4915 17765 4935
rect 17785 4915 17815 4935
rect 17835 4915 17865 4935
rect 17885 4915 17915 4935
rect 17935 4915 17950 4935
rect 17700 4900 17950 4915
rect 18000 4935 18250 4950
rect 18000 4915 18015 4935
rect 18035 4915 18065 4935
rect 18085 4915 18115 4935
rect 18135 4915 18165 4935
rect 18185 4915 18215 4935
rect 18235 4915 18250 4935
rect 18000 4900 18250 4915
rect 18300 4935 18550 4950
rect 18300 4915 18315 4935
rect 18335 4915 18365 4935
rect 18385 4915 18415 4935
rect 18435 4915 18465 4935
rect 18485 4915 18515 4935
rect 18535 4915 18550 4935
rect 18300 4900 18550 4915
rect 18600 4935 18850 4950
rect 18600 4915 18615 4935
rect 18635 4915 18665 4935
rect 18685 4915 18715 4935
rect 18735 4915 18765 4935
rect 18785 4915 18815 4935
rect 18835 4915 18850 4935
rect 18600 4900 18850 4915
rect 18900 4935 19150 4950
rect 18900 4915 18915 4935
rect 18935 4915 18965 4935
rect 18985 4915 19015 4935
rect 19035 4915 19065 4935
rect 19085 4915 19115 4935
rect 19135 4915 19150 4935
rect 18900 4900 19150 4915
rect 19200 4935 19450 4950
rect 19200 4915 19215 4935
rect 19235 4915 19265 4935
rect 19285 4915 19315 4935
rect 19335 4915 19365 4935
rect 19385 4915 19415 4935
rect 19435 4915 19450 4935
rect 19200 4900 19450 4915
rect 19500 4935 19750 4950
rect 19500 4915 19515 4935
rect 19535 4915 19565 4935
rect 19585 4915 19615 4935
rect 19635 4915 19665 4935
rect 19685 4915 19715 4935
rect 19735 4915 19750 4935
rect 19500 4900 19750 4915
rect 19800 4935 20050 4950
rect 19800 4915 19815 4935
rect 19835 4915 19865 4935
rect 19885 4915 19915 4935
rect 19935 4915 19965 4935
rect 19985 4915 20015 4935
rect 20035 4915 20050 4935
rect 19800 4900 20050 4915
rect 20100 4935 20350 4950
rect 20100 4915 20115 4935
rect 20135 4915 20165 4935
rect 20185 4915 20215 4935
rect 20235 4915 20265 4935
rect 20285 4915 20315 4935
rect 20335 4915 20350 4935
rect 20100 4900 20350 4915
rect 20400 4935 20650 4950
rect 20400 4915 20415 4935
rect 20435 4915 20465 4935
rect 20485 4915 20515 4935
rect 20535 4915 20565 4935
rect 20585 4915 20615 4935
rect 20635 4915 20650 4935
rect 20400 4900 20650 4915
rect 20700 4935 20950 4950
rect 20700 4915 20715 4935
rect 20735 4915 20765 4935
rect 20785 4915 20815 4935
rect 20835 4915 20865 4935
rect 20885 4915 20915 4935
rect 20935 4915 20950 4935
rect 20700 4900 20950 4915
rect 21000 4935 21400 4950
rect 21000 4915 21015 4935
rect 21035 4915 21065 4935
rect 21085 4915 21115 4935
rect 21135 4915 21165 4935
rect 21185 4915 21215 4935
rect 21235 4915 21265 4935
rect 21285 4915 21315 4935
rect 21335 4915 21365 4935
rect 21385 4915 21400 4935
rect 21000 4900 21400 4915
rect 21450 4935 21850 4950
rect 21450 4915 21465 4935
rect 21485 4915 21515 4935
rect 21535 4915 21565 4935
rect 21585 4915 21615 4935
rect 21635 4915 21665 4935
rect 21685 4915 21715 4935
rect 21735 4915 21765 4935
rect 21785 4915 21815 4935
rect 21835 4915 21850 4935
rect 21450 4900 21850 4915
rect 21900 4935 22150 4950
rect 21900 4915 21915 4935
rect 21935 4915 21965 4935
rect 21985 4915 22015 4935
rect 22035 4915 22065 4935
rect 22085 4915 22115 4935
rect 22135 4915 22150 4935
rect 21900 4900 22150 4915
rect 22200 4935 22450 4950
rect 22200 4915 22215 4935
rect 22235 4915 22265 4935
rect 22285 4915 22315 4935
rect 22335 4915 22365 4935
rect 22385 4915 22415 4935
rect 22435 4915 22450 4935
rect 22200 4900 22450 4915
rect 22500 4935 22750 4950
rect 22500 4915 22515 4935
rect 22535 4915 22565 4935
rect 22585 4915 22615 4935
rect 22635 4915 22665 4935
rect 22685 4915 22715 4935
rect 22735 4915 22750 4935
rect 22500 4900 22750 4915
rect 22800 4935 23050 4950
rect 22800 4915 22815 4935
rect 22835 4915 22865 4935
rect 22885 4915 22915 4935
rect 22935 4915 22965 4935
rect 22985 4915 23015 4935
rect 23035 4915 23050 4935
rect 22800 4900 23050 4915
rect 23100 4935 23500 4950
rect 23100 4915 23115 4935
rect 23135 4915 23165 4935
rect 23185 4915 23215 4935
rect 23235 4915 23265 4935
rect 23285 4915 23315 4935
rect 23335 4915 23365 4935
rect 23385 4915 23415 4935
rect 23435 4915 23465 4935
rect 23485 4915 23500 4935
rect 23100 4900 23500 4915
rect 23550 4935 23950 4950
rect 23550 4915 23565 4935
rect 23585 4915 23615 4935
rect 23635 4915 23665 4935
rect 23685 4915 23715 4935
rect 23735 4915 23765 4935
rect 23785 4915 23815 4935
rect 23835 4915 23865 4935
rect 23885 4915 23915 4935
rect 23935 4915 23950 4935
rect 23550 4900 23950 4915
rect 24000 4935 24250 4950
rect 24000 4915 24015 4935
rect 24035 4915 24065 4935
rect 24085 4915 24115 4935
rect 24135 4915 24165 4935
rect 24185 4915 24215 4935
rect 24235 4915 24250 4935
rect 24000 4900 24250 4915
rect 24300 4935 24550 4950
rect 24300 4915 24315 4935
rect 24335 4915 24365 4935
rect 24385 4915 24415 4935
rect 24435 4915 24465 4935
rect 24485 4915 24515 4935
rect 24535 4915 24550 4935
rect 24300 4900 24550 4915
rect 24600 4935 24850 4950
rect 24600 4915 24615 4935
rect 24635 4915 24665 4935
rect 24685 4915 24715 4935
rect 24735 4915 24765 4935
rect 24785 4915 24815 4935
rect 24835 4915 24850 4935
rect 24600 4900 24850 4915
rect 24900 4935 25150 4950
rect 24900 4915 24915 4935
rect 24935 4915 24965 4935
rect 24985 4915 25015 4935
rect 25035 4915 25065 4935
rect 25085 4915 25115 4935
rect 25135 4915 25150 4935
rect 24900 4900 25150 4915
rect 25200 4935 25600 4950
rect 25200 4915 25215 4935
rect 25235 4915 25265 4935
rect 25285 4915 25315 4935
rect 25335 4915 25365 4935
rect 25385 4915 25415 4935
rect 25435 4915 25465 4935
rect 25485 4915 25515 4935
rect 25535 4915 25565 4935
rect 25585 4915 25600 4935
rect 25200 4900 25600 4915
rect 25650 4935 26050 4950
rect 25650 4915 25665 4935
rect 25685 4915 25715 4935
rect 25735 4915 25765 4935
rect 25785 4915 25815 4935
rect 25835 4915 25865 4935
rect 25885 4915 25915 4935
rect 25935 4915 25965 4935
rect 25985 4915 26015 4935
rect 26035 4915 26050 4935
rect 25650 4900 26050 4915
rect 26100 4935 26350 4950
rect 26100 4915 26115 4935
rect 26135 4915 26165 4935
rect 26185 4915 26215 4935
rect 26235 4915 26265 4935
rect 26285 4915 26315 4935
rect 26335 4915 26350 4935
rect 26100 4900 26350 4915
rect 26400 4935 26650 4950
rect 26400 4915 26415 4935
rect 26435 4915 26465 4935
rect 26485 4915 26515 4935
rect 26535 4915 26565 4935
rect 26585 4915 26615 4935
rect 26635 4915 26650 4935
rect 26400 4900 26650 4915
rect 26700 4935 26950 4950
rect 26700 4915 26715 4935
rect 26735 4915 26765 4935
rect 26785 4915 26815 4935
rect 26835 4915 26865 4935
rect 26885 4915 26915 4935
rect 26935 4915 26950 4935
rect 26700 4900 26950 4915
rect 27000 4935 27250 4950
rect 27000 4915 27015 4935
rect 27035 4915 27065 4935
rect 27085 4915 27115 4935
rect 27135 4915 27165 4935
rect 27185 4915 27215 4935
rect 27235 4915 27250 4935
rect 27000 4900 27250 4915
rect 27300 4935 27700 4950
rect 27300 4915 27315 4935
rect 27335 4915 27365 4935
rect 27385 4915 27415 4935
rect 27435 4915 27465 4935
rect 27485 4915 27515 4935
rect 27535 4915 27565 4935
rect 27585 4915 27615 4935
rect 27635 4915 27665 4935
rect 27685 4915 27700 4935
rect 27300 4900 27700 4915
rect 27750 4935 28150 4950
rect 27750 4915 27765 4935
rect 27785 4915 27815 4935
rect 27835 4915 27865 4935
rect 27885 4915 27915 4935
rect 27935 4915 27965 4935
rect 27985 4915 28015 4935
rect 28035 4915 28065 4935
rect 28085 4915 28115 4935
rect 28135 4915 28150 4935
rect 27750 4900 28150 4915
rect 28200 4935 28450 4950
rect 28200 4915 28215 4935
rect 28235 4915 28265 4935
rect 28285 4915 28315 4935
rect 28335 4915 28365 4935
rect 28385 4915 28415 4935
rect 28435 4915 28450 4935
rect 28200 4900 28450 4915
rect 28500 4935 28750 4950
rect 28500 4915 28515 4935
rect 28535 4915 28565 4935
rect 28585 4915 28615 4935
rect 28635 4915 28665 4935
rect 28685 4915 28715 4935
rect 28735 4915 28750 4935
rect 28500 4900 28750 4915
rect 28800 4935 29050 4950
rect 28800 4915 28815 4935
rect 28835 4915 28865 4935
rect 28885 4915 28915 4935
rect 28935 4915 28965 4935
rect 28985 4915 29015 4935
rect 29035 4915 29050 4935
rect 28800 4900 29050 4915
rect 29100 4935 29350 4950
rect 29100 4915 29115 4935
rect 29135 4915 29165 4935
rect 29185 4915 29215 4935
rect 29235 4915 29265 4935
rect 29285 4915 29315 4935
rect 29335 4915 29350 4935
rect 29100 4900 29350 4915
rect 29400 4935 29800 4950
rect 29400 4915 29415 4935
rect 29435 4915 29465 4935
rect 29485 4915 29515 4935
rect 29535 4915 29565 4935
rect 29585 4915 29615 4935
rect 29635 4915 29665 4935
rect 29685 4915 29715 4935
rect 29735 4915 29765 4935
rect 29785 4915 29800 4935
rect 29400 4900 29800 4915
rect 29850 4935 30100 4950
rect 29850 4915 29865 4935
rect 29885 4915 29915 4935
rect 29935 4915 29965 4935
rect 29985 4915 30015 4935
rect 30035 4915 30065 4935
rect 30085 4915 30100 4935
rect 29850 4900 30100 4915
rect 30150 4935 30400 4950
rect 30150 4915 30165 4935
rect 30185 4915 30215 4935
rect 30235 4915 30265 4935
rect 30285 4915 30315 4935
rect 30335 4915 30365 4935
rect 30385 4915 30400 4935
rect 30150 4900 30400 4915
rect 30450 4935 30700 4950
rect 30450 4915 30465 4935
rect 30485 4915 30515 4935
rect 30535 4915 30565 4935
rect 30585 4915 30615 4935
rect 30635 4915 30665 4935
rect 30685 4915 30700 4935
rect 30450 4900 30700 4915
rect 30750 4935 31000 4950
rect 30750 4915 30765 4935
rect 30785 4915 30815 4935
rect 30835 4915 30865 4935
rect 30885 4915 30915 4935
rect 30935 4915 30965 4935
rect 30985 4915 31000 4935
rect 30750 4900 31000 4915
rect 31050 4935 31450 4950
rect 31050 4915 31065 4935
rect 31085 4915 31115 4935
rect 31135 4915 31165 4935
rect 31185 4915 31215 4935
rect 31235 4915 31265 4935
rect 31285 4915 31315 4935
rect 31335 4915 31365 4935
rect 31385 4915 31415 4935
rect 31435 4915 31450 4935
rect 31050 4900 31450 4915
rect 31500 4935 31750 4950
rect 31500 4915 31515 4935
rect 31535 4915 31565 4935
rect 31585 4915 31615 4935
rect 31635 4915 31665 4935
rect 31685 4915 31715 4935
rect 31735 4915 31750 4935
rect 31500 4900 31750 4915
rect 31800 4935 32050 4950
rect 31800 4915 31815 4935
rect 31835 4915 31865 4935
rect 31885 4915 31915 4935
rect 31935 4915 31965 4935
rect 31985 4915 32015 4935
rect 32035 4915 32050 4935
rect 31800 4900 32050 4915
rect -650 4835 -600 4850
rect -650 4815 -635 4835
rect -615 4815 -600 4835
rect -650 4785 -600 4815
rect -650 4765 -635 4785
rect -615 4765 -600 4785
rect -650 4735 -600 4765
rect -650 4715 -635 4735
rect -615 4715 -600 4735
rect -650 4685 -600 4715
rect -650 4665 -635 4685
rect -615 4665 -600 4685
rect -650 4635 -600 4665
rect -650 4615 -635 4635
rect -615 4615 -600 4635
rect -650 4585 -600 4615
rect -650 4565 -635 4585
rect -615 4565 -600 4585
rect -650 4535 -600 4565
rect -650 4515 -635 4535
rect -615 4515 -600 4535
rect -650 4485 -600 4515
rect -650 4465 -635 4485
rect -615 4465 -600 4485
rect -650 4435 -600 4465
rect -650 4415 -635 4435
rect -615 4415 -600 4435
rect -650 4385 -600 4415
rect -650 4365 -635 4385
rect -615 4365 -600 4385
rect -650 4350 -600 4365
rect -500 4835 -450 4850
rect -500 4815 -485 4835
rect -465 4815 -450 4835
rect -500 4785 -450 4815
rect -500 4765 -485 4785
rect -465 4765 -450 4785
rect -500 4735 -450 4765
rect -500 4715 -485 4735
rect -465 4715 -450 4735
rect -500 4685 -450 4715
rect -500 4665 -485 4685
rect -465 4665 -450 4685
rect -500 4635 -450 4665
rect -500 4615 -485 4635
rect -465 4615 -450 4635
rect -500 4585 -450 4615
rect -500 4565 -485 4585
rect -465 4565 -450 4585
rect -500 4535 -450 4565
rect -500 4515 -485 4535
rect -465 4515 -450 4535
rect -500 4485 -450 4515
rect -500 4465 -485 4485
rect -465 4465 -450 4485
rect -500 4435 -450 4465
rect -500 4415 -485 4435
rect -465 4415 -450 4435
rect -500 4385 -450 4415
rect -500 4365 -485 4385
rect -465 4365 -450 4385
rect -500 4350 -450 4365
rect -350 4835 -300 4850
rect -350 4815 -335 4835
rect -315 4815 -300 4835
rect -350 4785 -300 4815
rect -350 4765 -335 4785
rect -315 4765 -300 4785
rect -350 4735 -300 4765
rect -350 4715 -335 4735
rect -315 4715 -300 4735
rect -350 4685 -300 4715
rect -350 4665 -335 4685
rect -315 4665 -300 4685
rect -350 4635 -300 4665
rect -350 4615 -335 4635
rect -315 4615 -300 4635
rect -350 4585 -300 4615
rect -350 4565 -335 4585
rect -315 4565 -300 4585
rect -350 4535 -300 4565
rect -350 4515 -335 4535
rect -315 4515 -300 4535
rect -350 4485 -300 4515
rect -350 4465 -335 4485
rect -315 4465 -300 4485
rect -350 4435 -300 4465
rect -350 4415 -335 4435
rect -315 4415 -300 4435
rect -350 4385 -300 4415
rect -350 4365 -335 4385
rect -315 4365 -300 4385
rect -350 4350 -300 4365
rect -200 4835 -150 4850
rect -200 4815 -185 4835
rect -165 4815 -150 4835
rect -200 4785 -150 4815
rect -200 4765 -185 4785
rect -165 4765 -150 4785
rect -200 4735 -150 4765
rect -200 4715 -185 4735
rect -165 4715 -150 4735
rect -200 4685 -150 4715
rect -200 4665 -185 4685
rect -165 4665 -150 4685
rect -200 4635 -150 4665
rect -200 4615 -185 4635
rect -165 4615 -150 4635
rect -200 4585 -150 4615
rect -200 4565 -185 4585
rect -165 4565 -150 4585
rect -200 4535 -150 4565
rect -200 4515 -185 4535
rect -165 4515 -150 4535
rect -200 4485 -150 4515
rect -200 4465 -185 4485
rect -165 4465 -150 4485
rect -200 4435 -150 4465
rect -200 4415 -185 4435
rect -165 4415 -150 4435
rect -200 4385 -150 4415
rect -200 4365 -185 4385
rect -165 4365 -150 4385
rect -200 4350 -150 4365
rect -50 4835 0 4850
rect -50 4815 -35 4835
rect -15 4815 0 4835
rect -50 4785 0 4815
rect -50 4765 -35 4785
rect -15 4765 0 4785
rect -50 4735 0 4765
rect -50 4715 -35 4735
rect -15 4715 0 4735
rect -50 4685 0 4715
rect -50 4665 -35 4685
rect -15 4665 0 4685
rect -50 4635 0 4665
rect -50 4615 -35 4635
rect -15 4615 0 4635
rect -50 4585 0 4615
rect -50 4565 -35 4585
rect -15 4565 0 4585
rect -50 4535 0 4565
rect -50 4515 -35 4535
rect -15 4515 0 4535
rect -50 4485 0 4515
rect -50 4465 -35 4485
rect -15 4465 0 4485
rect -50 4435 0 4465
rect -50 4415 -35 4435
rect -15 4415 0 4435
rect -50 4385 0 4415
rect -50 4365 -35 4385
rect -15 4365 0 4385
rect -50 4350 0 4365
rect 550 4835 600 4850
rect 550 4815 565 4835
rect 585 4815 600 4835
rect 550 4785 600 4815
rect 550 4765 565 4785
rect 585 4765 600 4785
rect 550 4735 600 4765
rect 550 4715 565 4735
rect 585 4715 600 4735
rect 550 4685 600 4715
rect 550 4665 565 4685
rect 585 4665 600 4685
rect 550 4635 600 4665
rect 550 4615 565 4635
rect 585 4615 600 4635
rect 550 4585 600 4615
rect 550 4565 565 4585
rect 585 4565 600 4585
rect 550 4535 600 4565
rect 550 4515 565 4535
rect 585 4515 600 4535
rect 550 4485 600 4515
rect 550 4465 565 4485
rect 585 4465 600 4485
rect 550 4435 600 4465
rect 550 4415 565 4435
rect 585 4415 600 4435
rect 550 4385 600 4415
rect 550 4365 565 4385
rect 585 4365 600 4385
rect 550 4350 600 4365
rect 700 4835 750 4850
rect 700 4815 715 4835
rect 735 4815 750 4835
rect 700 4785 750 4815
rect 700 4765 715 4785
rect 735 4765 750 4785
rect 700 4735 750 4765
rect 700 4715 715 4735
rect 735 4715 750 4735
rect 700 4685 750 4715
rect 700 4665 715 4685
rect 735 4665 750 4685
rect 700 4635 750 4665
rect 700 4615 715 4635
rect 735 4615 750 4635
rect 700 4585 750 4615
rect 700 4565 715 4585
rect 735 4565 750 4585
rect 700 4535 750 4565
rect 700 4515 715 4535
rect 735 4515 750 4535
rect 700 4485 750 4515
rect 700 4465 715 4485
rect 735 4465 750 4485
rect 700 4435 750 4465
rect 700 4415 715 4435
rect 735 4415 750 4435
rect 700 4385 750 4415
rect 700 4365 715 4385
rect 735 4365 750 4385
rect 700 4350 750 4365
rect 850 4835 900 4850
rect 850 4815 865 4835
rect 885 4815 900 4835
rect 850 4785 900 4815
rect 850 4765 865 4785
rect 885 4765 900 4785
rect 850 4735 900 4765
rect 850 4715 865 4735
rect 885 4715 900 4735
rect 850 4685 900 4715
rect 850 4665 865 4685
rect 885 4665 900 4685
rect 850 4635 900 4665
rect 850 4615 865 4635
rect 885 4615 900 4635
rect 850 4585 900 4615
rect 850 4565 865 4585
rect 885 4565 900 4585
rect 850 4535 900 4565
rect 850 4515 865 4535
rect 885 4515 900 4535
rect 850 4485 900 4515
rect 850 4465 865 4485
rect 885 4465 900 4485
rect 850 4435 900 4465
rect 850 4415 865 4435
rect 885 4415 900 4435
rect 850 4385 900 4415
rect 850 4365 865 4385
rect 885 4365 900 4385
rect 850 4350 900 4365
rect 1000 4835 1050 4850
rect 1000 4815 1015 4835
rect 1035 4815 1050 4835
rect 1000 4785 1050 4815
rect 1000 4765 1015 4785
rect 1035 4765 1050 4785
rect 1000 4735 1050 4765
rect 1000 4715 1015 4735
rect 1035 4715 1050 4735
rect 1000 4685 1050 4715
rect 1000 4665 1015 4685
rect 1035 4665 1050 4685
rect 1000 4635 1050 4665
rect 1000 4615 1015 4635
rect 1035 4615 1050 4635
rect 1000 4585 1050 4615
rect 1000 4565 1015 4585
rect 1035 4565 1050 4585
rect 1000 4535 1050 4565
rect 1000 4515 1015 4535
rect 1035 4515 1050 4535
rect 1000 4485 1050 4515
rect 1000 4465 1015 4485
rect 1035 4465 1050 4485
rect 1000 4435 1050 4465
rect 1000 4415 1015 4435
rect 1035 4415 1050 4435
rect 1000 4385 1050 4415
rect 1000 4365 1015 4385
rect 1035 4365 1050 4385
rect 1000 4350 1050 4365
rect 1150 4835 1200 4850
rect 1150 4815 1165 4835
rect 1185 4815 1200 4835
rect 1150 4785 1200 4815
rect 1150 4765 1165 4785
rect 1185 4765 1200 4785
rect 1150 4735 1200 4765
rect 1150 4715 1165 4735
rect 1185 4715 1200 4735
rect 1150 4685 1200 4715
rect 1150 4665 1165 4685
rect 1185 4665 1200 4685
rect 1150 4635 1200 4665
rect 1150 4615 1165 4635
rect 1185 4615 1200 4635
rect 1150 4585 1200 4615
rect 1150 4565 1165 4585
rect 1185 4565 1200 4585
rect 1150 4535 1200 4565
rect 1150 4515 1165 4535
rect 1185 4515 1200 4535
rect 1150 4485 1200 4515
rect 1150 4465 1165 4485
rect 1185 4465 1200 4485
rect 1150 4435 1200 4465
rect 1150 4415 1165 4435
rect 1185 4415 1200 4435
rect 1150 4385 1200 4415
rect 1150 4365 1165 4385
rect 1185 4365 1200 4385
rect 1150 4350 1200 4365
rect 1300 4835 1350 4850
rect 1300 4815 1315 4835
rect 1335 4815 1350 4835
rect 1300 4785 1350 4815
rect 1300 4765 1315 4785
rect 1335 4765 1350 4785
rect 1300 4735 1350 4765
rect 1300 4715 1315 4735
rect 1335 4715 1350 4735
rect 1300 4685 1350 4715
rect 1300 4665 1315 4685
rect 1335 4665 1350 4685
rect 1300 4635 1350 4665
rect 1300 4615 1315 4635
rect 1335 4615 1350 4635
rect 1300 4585 1350 4615
rect 1300 4565 1315 4585
rect 1335 4565 1350 4585
rect 1300 4535 1350 4565
rect 1300 4515 1315 4535
rect 1335 4515 1350 4535
rect 1300 4485 1350 4515
rect 1300 4465 1315 4485
rect 1335 4465 1350 4485
rect 1300 4435 1350 4465
rect 1300 4415 1315 4435
rect 1335 4415 1350 4435
rect 1300 4385 1350 4415
rect 1300 4365 1315 4385
rect 1335 4365 1350 4385
rect 1300 4350 1350 4365
rect 1450 4835 1500 4850
rect 1450 4815 1465 4835
rect 1485 4815 1500 4835
rect 1450 4785 1500 4815
rect 1450 4765 1465 4785
rect 1485 4765 1500 4785
rect 1450 4735 1500 4765
rect 1450 4715 1465 4735
rect 1485 4715 1500 4735
rect 1450 4685 1500 4715
rect 1450 4665 1465 4685
rect 1485 4665 1500 4685
rect 1450 4635 1500 4665
rect 1450 4615 1465 4635
rect 1485 4615 1500 4635
rect 1450 4585 1500 4615
rect 1450 4565 1465 4585
rect 1485 4565 1500 4585
rect 1450 4535 1500 4565
rect 1450 4515 1465 4535
rect 1485 4515 1500 4535
rect 1450 4485 1500 4515
rect 1450 4465 1465 4485
rect 1485 4465 1500 4485
rect 1450 4435 1500 4465
rect 1450 4415 1465 4435
rect 1485 4415 1500 4435
rect 1450 4385 1500 4415
rect 1450 4365 1465 4385
rect 1485 4365 1500 4385
rect 1450 4350 1500 4365
rect 1600 4835 1650 4850
rect 1600 4815 1615 4835
rect 1635 4815 1650 4835
rect 1600 4785 1650 4815
rect 1600 4765 1615 4785
rect 1635 4765 1650 4785
rect 1600 4735 1650 4765
rect 1600 4715 1615 4735
rect 1635 4715 1650 4735
rect 1600 4685 1650 4715
rect 1600 4665 1615 4685
rect 1635 4665 1650 4685
rect 1600 4635 1650 4665
rect 1600 4615 1615 4635
rect 1635 4615 1650 4635
rect 1600 4585 1650 4615
rect 1600 4565 1615 4585
rect 1635 4565 1650 4585
rect 1600 4535 1650 4565
rect 1600 4515 1615 4535
rect 1635 4515 1650 4535
rect 1600 4485 1650 4515
rect 1600 4465 1615 4485
rect 1635 4465 1650 4485
rect 1600 4435 1650 4465
rect 1600 4415 1615 4435
rect 1635 4415 1650 4435
rect 1600 4385 1650 4415
rect 1600 4365 1615 4385
rect 1635 4365 1650 4385
rect 1600 4350 1650 4365
rect 1750 4835 1800 4850
rect 1750 4815 1765 4835
rect 1785 4815 1800 4835
rect 1750 4785 1800 4815
rect 1750 4765 1765 4785
rect 1785 4765 1800 4785
rect 1750 4735 1800 4765
rect 1750 4715 1765 4735
rect 1785 4715 1800 4735
rect 1750 4685 1800 4715
rect 1750 4665 1765 4685
rect 1785 4665 1800 4685
rect 1750 4635 1800 4665
rect 1750 4615 1765 4635
rect 1785 4615 1800 4635
rect 1750 4585 1800 4615
rect 1750 4565 1765 4585
rect 1785 4565 1800 4585
rect 1750 4535 1800 4565
rect 1750 4515 1765 4535
rect 1785 4515 1800 4535
rect 1750 4485 1800 4515
rect 1750 4465 1765 4485
rect 1785 4465 1800 4485
rect 1750 4435 1800 4465
rect 1750 4415 1765 4435
rect 1785 4415 1800 4435
rect 1750 4385 1800 4415
rect 1750 4365 1765 4385
rect 1785 4365 1800 4385
rect 1750 4350 1800 4365
rect 1900 4835 1950 4850
rect 1900 4815 1915 4835
rect 1935 4815 1950 4835
rect 1900 4785 1950 4815
rect 1900 4765 1915 4785
rect 1935 4765 1950 4785
rect 1900 4735 1950 4765
rect 1900 4715 1915 4735
rect 1935 4715 1950 4735
rect 1900 4685 1950 4715
rect 1900 4665 1915 4685
rect 1935 4665 1950 4685
rect 1900 4635 1950 4665
rect 1900 4615 1915 4635
rect 1935 4615 1950 4635
rect 1900 4585 1950 4615
rect 1900 4565 1915 4585
rect 1935 4565 1950 4585
rect 1900 4535 1950 4565
rect 1900 4515 1915 4535
rect 1935 4515 1950 4535
rect 1900 4485 1950 4515
rect 1900 4465 1915 4485
rect 1935 4465 1950 4485
rect 1900 4435 1950 4465
rect 1900 4415 1915 4435
rect 1935 4415 1950 4435
rect 1900 4385 1950 4415
rect 1900 4365 1915 4385
rect 1935 4365 1950 4385
rect 1900 4350 1950 4365
rect 2050 4835 2100 4850
rect 2050 4815 2065 4835
rect 2085 4815 2100 4835
rect 2050 4785 2100 4815
rect 2050 4765 2065 4785
rect 2085 4765 2100 4785
rect 2050 4735 2100 4765
rect 2050 4715 2065 4735
rect 2085 4715 2100 4735
rect 2050 4685 2100 4715
rect 2050 4665 2065 4685
rect 2085 4665 2100 4685
rect 2050 4635 2100 4665
rect 2050 4615 2065 4635
rect 2085 4615 2100 4635
rect 2050 4585 2100 4615
rect 2050 4565 2065 4585
rect 2085 4565 2100 4585
rect 2050 4535 2100 4565
rect 2050 4515 2065 4535
rect 2085 4515 2100 4535
rect 2050 4485 2100 4515
rect 2050 4465 2065 4485
rect 2085 4465 2100 4485
rect 2050 4435 2100 4465
rect 2050 4415 2065 4435
rect 2085 4415 2100 4435
rect 2050 4385 2100 4415
rect 2050 4365 2065 4385
rect 2085 4365 2100 4385
rect 2050 4350 2100 4365
rect 2200 4835 2250 4850
rect 2200 4815 2215 4835
rect 2235 4815 2250 4835
rect 2200 4785 2250 4815
rect 2200 4765 2215 4785
rect 2235 4765 2250 4785
rect 2200 4735 2250 4765
rect 2200 4715 2215 4735
rect 2235 4715 2250 4735
rect 2200 4685 2250 4715
rect 2200 4665 2215 4685
rect 2235 4665 2250 4685
rect 2200 4635 2250 4665
rect 2200 4615 2215 4635
rect 2235 4615 2250 4635
rect 2200 4585 2250 4615
rect 2200 4565 2215 4585
rect 2235 4565 2250 4585
rect 2200 4535 2250 4565
rect 2200 4515 2215 4535
rect 2235 4515 2250 4535
rect 2200 4485 2250 4515
rect 2200 4465 2215 4485
rect 2235 4465 2250 4485
rect 2200 4435 2250 4465
rect 2200 4415 2215 4435
rect 2235 4415 2250 4435
rect 2200 4385 2250 4415
rect 2200 4365 2215 4385
rect 2235 4365 2250 4385
rect 2200 4350 2250 4365
rect 2350 4835 2400 4850
rect 2350 4815 2365 4835
rect 2385 4815 2400 4835
rect 2350 4785 2400 4815
rect 2350 4765 2365 4785
rect 2385 4765 2400 4785
rect 2350 4735 2400 4765
rect 2350 4715 2365 4735
rect 2385 4715 2400 4735
rect 2350 4685 2400 4715
rect 2350 4665 2365 4685
rect 2385 4665 2400 4685
rect 2350 4635 2400 4665
rect 2350 4615 2365 4635
rect 2385 4615 2400 4635
rect 2350 4585 2400 4615
rect 2350 4565 2365 4585
rect 2385 4565 2400 4585
rect 2350 4535 2400 4565
rect 2350 4515 2365 4535
rect 2385 4515 2400 4535
rect 2350 4485 2400 4515
rect 2350 4465 2365 4485
rect 2385 4465 2400 4485
rect 2350 4435 2400 4465
rect 2350 4415 2365 4435
rect 2385 4415 2400 4435
rect 2350 4385 2400 4415
rect 2350 4365 2365 4385
rect 2385 4365 2400 4385
rect 2350 4350 2400 4365
rect 2500 4835 2550 4850
rect 2500 4815 2515 4835
rect 2535 4815 2550 4835
rect 2500 4785 2550 4815
rect 2500 4765 2515 4785
rect 2535 4765 2550 4785
rect 2500 4735 2550 4765
rect 2500 4715 2515 4735
rect 2535 4715 2550 4735
rect 2500 4685 2550 4715
rect 2500 4665 2515 4685
rect 2535 4665 2550 4685
rect 2500 4635 2550 4665
rect 2500 4615 2515 4635
rect 2535 4615 2550 4635
rect 2500 4585 2550 4615
rect 2500 4565 2515 4585
rect 2535 4565 2550 4585
rect 2500 4535 2550 4565
rect 2500 4515 2515 4535
rect 2535 4515 2550 4535
rect 2500 4485 2550 4515
rect 2500 4465 2515 4485
rect 2535 4465 2550 4485
rect 2500 4435 2550 4465
rect 2500 4415 2515 4435
rect 2535 4415 2550 4435
rect 2500 4385 2550 4415
rect 2500 4365 2515 4385
rect 2535 4365 2550 4385
rect 2500 4350 2550 4365
rect 2650 4835 2700 4850
rect 2650 4815 2665 4835
rect 2685 4815 2700 4835
rect 2650 4785 2700 4815
rect 2650 4765 2665 4785
rect 2685 4765 2700 4785
rect 2650 4735 2700 4765
rect 2650 4715 2665 4735
rect 2685 4715 2700 4735
rect 2650 4685 2700 4715
rect 2650 4665 2665 4685
rect 2685 4665 2700 4685
rect 2650 4635 2700 4665
rect 2650 4615 2665 4635
rect 2685 4615 2700 4635
rect 2650 4585 2700 4615
rect 2650 4565 2665 4585
rect 2685 4565 2700 4585
rect 2650 4535 2700 4565
rect 2650 4515 2665 4535
rect 2685 4515 2700 4535
rect 2650 4485 2700 4515
rect 2650 4465 2665 4485
rect 2685 4465 2700 4485
rect 2650 4435 2700 4465
rect 2650 4415 2665 4435
rect 2685 4415 2700 4435
rect 2650 4385 2700 4415
rect 2650 4365 2665 4385
rect 2685 4365 2700 4385
rect 2650 4350 2700 4365
rect 2800 4835 2850 4850
rect 2800 4815 2815 4835
rect 2835 4815 2850 4835
rect 2800 4785 2850 4815
rect 2800 4765 2815 4785
rect 2835 4765 2850 4785
rect 2800 4735 2850 4765
rect 2800 4715 2815 4735
rect 2835 4715 2850 4735
rect 2800 4685 2850 4715
rect 2800 4665 2815 4685
rect 2835 4665 2850 4685
rect 2800 4635 2850 4665
rect 2800 4615 2815 4635
rect 2835 4615 2850 4635
rect 2800 4585 2850 4615
rect 2800 4565 2815 4585
rect 2835 4565 2850 4585
rect 2800 4535 2850 4565
rect 2800 4515 2815 4535
rect 2835 4515 2850 4535
rect 2800 4485 2850 4515
rect 2800 4465 2815 4485
rect 2835 4465 2850 4485
rect 2800 4435 2850 4465
rect 2800 4415 2815 4435
rect 2835 4415 2850 4435
rect 2800 4385 2850 4415
rect 2800 4365 2815 4385
rect 2835 4365 2850 4385
rect 2800 4350 2850 4365
rect 2950 4835 3000 4850
rect 2950 4815 2965 4835
rect 2985 4815 3000 4835
rect 2950 4785 3000 4815
rect 2950 4765 2965 4785
rect 2985 4765 3000 4785
rect 2950 4735 3000 4765
rect 2950 4715 2965 4735
rect 2985 4715 3000 4735
rect 2950 4685 3000 4715
rect 2950 4665 2965 4685
rect 2985 4665 3000 4685
rect 2950 4635 3000 4665
rect 2950 4615 2965 4635
rect 2985 4615 3000 4635
rect 2950 4585 3000 4615
rect 2950 4565 2965 4585
rect 2985 4565 3000 4585
rect 2950 4535 3000 4565
rect 2950 4515 2965 4535
rect 2985 4515 3000 4535
rect 2950 4485 3000 4515
rect 2950 4465 2965 4485
rect 2985 4465 3000 4485
rect 2950 4435 3000 4465
rect 2950 4415 2965 4435
rect 2985 4415 3000 4435
rect 2950 4385 3000 4415
rect 2950 4365 2965 4385
rect 2985 4365 3000 4385
rect 2950 4350 3000 4365
rect 3100 4835 3150 4850
rect 3100 4815 3115 4835
rect 3135 4815 3150 4835
rect 3100 4785 3150 4815
rect 3100 4765 3115 4785
rect 3135 4765 3150 4785
rect 3100 4735 3150 4765
rect 3100 4715 3115 4735
rect 3135 4715 3150 4735
rect 3100 4685 3150 4715
rect 3100 4665 3115 4685
rect 3135 4665 3150 4685
rect 3100 4635 3150 4665
rect 3100 4615 3115 4635
rect 3135 4615 3150 4635
rect 3100 4585 3150 4615
rect 3100 4565 3115 4585
rect 3135 4565 3150 4585
rect 3100 4535 3150 4565
rect 3100 4515 3115 4535
rect 3135 4515 3150 4535
rect 3100 4485 3150 4515
rect 3100 4465 3115 4485
rect 3135 4465 3150 4485
rect 3100 4435 3150 4465
rect 3100 4415 3115 4435
rect 3135 4415 3150 4435
rect 3100 4385 3150 4415
rect 3100 4365 3115 4385
rect 3135 4365 3150 4385
rect 3100 4350 3150 4365
rect 3250 4835 3300 4850
rect 3250 4815 3265 4835
rect 3285 4815 3300 4835
rect 3250 4785 3300 4815
rect 3250 4765 3265 4785
rect 3285 4765 3300 4785
rect 3250 4735 3300 4765
rect 3250 4715 3265 4735
rect 3285 4715 3300 4735
rect 3250 4685 3300 4715
rect 3250 4665 3265 4685
rect 3285 4665 3300 4685
rect 3250 4635 3300 4665
rect 3250 4615 3265 4635
rect 3285 4615 3300 4635
rect 3250 4585 3300 4615
rect 3250 4565 3265 4585
rect 3285 4565 3300 4585
rect 3250 4535 3300 4565
rect 3250 4515 3265 4535
rect 3285 4515 3300 4535
rect 3250 4485 3300 4515
rect 3250 4465 3265 4485
rect 3285 4465 3300 4485
rect 3250 4435 3300 4465
rect 3250 4415 3265 4435
rect 3285 4415 3300 4435
rect 3250 4385 3300 4415
rect 3250 4365 3265 4385
rect 3285 4365 3300 4385
rect 3250 4350 3300 4365
rect 3400 4835 3450 4850
rect 3400 4815 3415 4835
rect 3435 4815 3450 4835
rect 3400 4785 3450 4815
rect 3400 4765 3415 4785
rect 3435 4765 3450 4785
rect 3400 4735 3450 4765
rect 3400 4715 3415 4735
rect 3435 4715 3450 4735
rect 3400 4685 3450 4715
rect 3400 4665 3415 4685
rect 3435 4665 3450 4685
rect 3400 4635 3450 4665
rect 3400 4615 3415 4635
rect 3435 4615 3450 4635
rect 3400 4585 3450 4615
rect 3400 4565 3415 4585
rect 3435 4565 3450 4585
rect 3400 4535 3450 4565
rect 3400 4515 3415 4535
rect 3435 4515 3450 4535
rect 3400 4485 3450 4515
rect 3400 4465 3415 4485
rect 3435 4465 3450 4485
rect 3400 4435 3450 4465
rect 3400 4415 3415 4435
rect 3435 4415 3450 4435
rect 3400 4385 3450 4415
rect 3400 4365 3415 4385
rect 3435 4365 3450 4385
rect 3400 4350 3450 4365
rect 3550 4835 3600 4850
rect 3550 4815 3565 4835
rect 3585 4815 3600 4835
rect 3550 4785 3600 4815
rect 3550 4765 3565 4785
rect 3585 4765 3600 4785
rect 3550 4735 3600 4765
rect 3550 4715 3565 4735
rect 3585 4715 3600 4735
rect 3550 4685 3600 4715
rect 3550 4665 3565 4685
rect 3585 4665 3600 4685
rect 3550 4635 3600 4665
rect 3550 4615 3565 4635
rect 3585 4615 3600 4635
rect 3550 4585 3600 4615
rect 3550 4565 3565 4585
rect 3585 4565 3600 4585
rect 3550 4535 3600 4565
rect 3550 4515 3565 4535
rect 3585 4515 3600 4535
rect 3550 4485 3600 4515
rect 3550 4465 3565 4485
rect 3585 4465 3600 4485
rect 3550 4435 3600 4465
rect 3550 4415 3565 4435
rect 3585 4415 3600 4435
rect 3550 4385 3600 4415
rect 3550 4365 3565 4385
rect 3585 4365 3600 4385
rect 3550 4350 3600 4365
rect 4150 4835 4200 4850
rect 4150 4815 4165 4835
rect 4185 4815 4200 4835
rect 4150 4785 4200 4815
rect 4150 4765 4165 4785
rect 4185 4765 4200 4785
rect 4150 4735 4200 4765
rect 4150 4715 4165 4735
rect 4185 4715 4200 4735
rect 4150 4685 4200 4715
rect 4150 4665 4165 4685
rect 4185 4665 4200 4685
rect 4150 4635 4200 4665
rect 4150 4615 4165 4635
rect 4185 4615 4200 4635
rect 4150 4585 4200 4615
rect 4150 4565 4165 4585
rect 4185 4565 4200 4585
rect 4150 4535 4200 4565
rect 4150 4515 4165 4535
rect 4185 4515 4200 4535
rect 4150 4485 4200 4515
rect 4150 4465 4165 4485
rect 4185 4465 4200 4485
rect 4150 4435 4200 4465
rect 4150 4415 4165 4435
rect 4185 4415 4200 4435
rect 4150 4385 4200 4415
rect 4150 4365 4165 4385
rect 4185 4365 4200 4385
rect 4150 4350 4200 4365
rect 4750 4835 4800 4850
rect 4750 4815 4765 4835
rect 4785 4815 4800 4835
rect 4750 4785 4800 4815
rect 4750 4765 4765 4785
rect 4785 4765 4800 4785
rect 4750 4735 4800 4765
rect 4750 4715 4765 4735
rect 4785 4715 4800 4735
rect 4750 4685 4800 4715
rect 4750 4665 4765 4685
rect 4785 4665 4800 4685
rect 4750 4635 4800 4665
rect 4750 4615 4765 4635
rect 4785 4615 4800 4635
rect 4750 4585 4800 4615
rect 4750 4565 4765 4585
rect 4785 4565 4800 4585
rect 4750 4535 4800 4565
rect 4750 4515 4765 4535
rect 4785 4515 4800 4535
rect 4750 4485 4800 4515
rect 4750 4465 4765 4485
rect 4785 4465 4800 4485
rect 4750 4435 4800 4465
rect 4750 4415 4765 4435
rect 4785 4415 4800 4435
rect 4750 4385 4800 4415
rect 4750 4365 4765 4385
rect 4785 4365 4800 4385
rect 4750 4350 4800 4365
rect 4900 4835 4950 4850
rect 4900 4815 4915 4835
rect 4935 4815 4950 4835
rect 4900 4785 4950 4815
rect 4900 4765 4915 4785
rect 4935 4765 4950 4785
rect 4900 4735 4950 4765
rect 4900 4715 4915 4735
rect 4935 4715 4950 4735
rect 4900 4685 4950 4715
rect 4900 4665 4915 4685
rect 4935 4665 4950 4685
rect 4900 4635 4950 4665
rect 4900 4615 4915 4635
rect 4935 4615 4950 4635
rect 4900 4585 4950 4615
rect 4900 4565 4915 4585
rect 4935 4565 4950 4585
rect 4900 4535 4950 4565
rect 4900 4515 4915 4535
rect 4935 4515 4950 4535
rect 4900 4485 4950 4515
rect 4900 4465 4915 4485
rect 4935 4465 4950 4485
rect 4900 4435 4950 4465
rect 4900 4415 4915 4435
rect 4935 4415 4950 4435
rect 4900 4385 4950 4415
rect 4900 4365 4915 4385
rect 4935 4365 4950 4385
rect 4900 4350 4950 4365
rect 5050 4835 5100 4850
rect 5050 4815 5065 4835
rect 5085 4815 5100 4835
rect 5050 4785 5100 4815
rect 5050 4765 5065 4785
rect 5085 4765 5100 4785
rect 5050 4735 5100 4765
rect 5050 4715 5065 4735
rect 5085 4715 5100 4735
rect 5050 4685 5100 4715
rect 5050 4665 5065 4685
rect 5085 4665 5100 4685
rect 5050 4635 5100 4665
rect 5050 4615 5065 4635
rect 5085 4615 5100 4635
rect 5050 4585 5100 4615
rect 5050 4565 5065 4585
rect 5085 4565 5100 4585
rect 5050 4535 5100 4565
rect 5050 4515 5065 4535
rect 5085 4515 5100 4535
rect 5050 4485 5100 4515
rect 5050 4465 5065 4485
rect 5085 4465 5100 4485
rect 5050 4435 5100 4465
rect 5050 4415 5065 4435
rect 5085 4415 5100 4435
rect 5050 4385 5100 4415
rect 5050 4365 5065 4385
rect 5085 4365 5100 4385
rect 5050 4350 5100 4365
rect 5200 4835 5250 4850
rect 5200 4815 5215 4835
rect 5235 4815 5250 4835
rect 5200 4785 5250 4815
rect 5200 4765 5215 4785
rect 5235 4765 5250 4785
rect 5200 4735 5250 4765
rect 5200 4715 5215 4735
rect 5235 4715 5250 4735
rect 5200 4685 5250 4715
rect 5200 4665 5215 4685
rect 5235 4665 5250 4685
rect 5200 4635 5250 4665
rect 5200 4615 5215 4635
rect 5235 4615 5250 4635
rect 5200 4585 5250 4615
rect 5200 4565 5215 4585
rect 5235 4565 5250 4585
rect 5200 4535 5250 4565
rect 5200 4515 5215 4535
rect 5235 4515 5250 4535
rect 5200 4485 5250 4515
rect 5200 4465 5215 4485
rect 5235 4465 5250 4485
rect 5200 4435 5250 4465
rect 5200 4415 5215 4435
rect 5235 4415 5250 4435
rect 5200 4385 5250 4415
rect 5200 4365 5215 4385
rect 5235 4365 5250 4385
rect 5200 4350 5250 4365
rect 5350 4835 5400 4850
rect 5350 4815 5365 4835
rect 5385 4815 5400 4835
rect 5350 4785 5400 4815
rect 5350 4765 5365 4785
rect 5385 4765 5400 4785
rect 5350 4735 5400 4765
rect 5350 4715 5365 4735
rect 5385 4715 5400 4735
rect 5350 4685 5400 4715
rect 5350 4665 5365 4685
rect 5385 4665 5400 4685
rect 5350 4635 5400 4665
rect 5350 4615 5365 4635
rect 5385 4615 5400 4635
rect 5350 4585 5400 4615
rect 5350 4565 5365 4585
rect 5385 4565 5400 4585
rect 5350 4535 5400 4565
rect 5350 4515 5365 4535
rect 5385 4515 5400 4535
rect 5350 4485 5400 4515
rect 5350 4465 5365 4485
rect 5385 4465 5400 4485
rect 5350 4435 5400 4465
rect 5350 4415 5365 4435
rect 5385 4415 5400 4435
rect 5350 4385 5400 4415
rect 5350 4365 5365 4385
rect 5385 4365 5400 4385
rect 5350 4350 5400 4365
rect 5500 4835 5550 4850
rect 5500 4815 5515 4835
rect 5535 4815 5550 4835
rect 5500 4785 5550 4815
rect 5500 4765 5515 4785
rect 5535 4765 5550 4785
rect 5500 4735 5550 4765
rect 5500 4715 5515 4735
rect 5535 4715 5550 4735
rect 5500 4685 5550 4715
rect 5500 4665 5515 4685
rect 5535 4665 5550 4685
rect 5500 4635 5550 4665
rect 5500 4615 5515 4635
rect 5535 4615 5550 4635
rect 5500 4585 5550 4615
rect 5500 4565 5515 4585
rect 5535 4565 5550 4585
rect 5500 4535 5550 4565
rect 5500 4515 5515 4535
rect 5535 4515 5550 4535
rect 5500 4485 5550 4515
rect 5500 4465 5515 4485
rect 5535 4465 5550 4485
rect 5500 4435 5550 4465
rect 5500 4415 5515 4435
rect 5535 4415 5550 4435
rect 5500 4385 5550 4415
rect 5500 4365 5515 4385
rect 5535 4365 5550 4385
rect 5500 4350 5550 4365
rect 5650 4835 5700 4850
rect 5650 4815 5665 4835
rect 5685 4815 5700 4835
rect 5650 4785 5700 4815
rect 5650 4765 5665 4785
rect 5685 4765 5700 4785
rect 5650 4735 5700 4765
rect 5650 4715 5665 4735
rect 5685 4715 5700 4735
rect 5650 4685 5700 4715
rect 5650 4665 5665 4685
rect 5685 4665 5700 4685
rect 5650 4635 5700 4665
rect 5650 4615 5665 4635
rect 5685 4615 5700 4635
rect 5650 4585 5700 4615
rect 5650 4565 5665 4585
rect 5685 4565 5700 4585
rect 5650 4535 5700 4565
rect 5650 4515 5665 4535
rect 5685 4515 5700 4535
rect 5650 4485 5700 4515
rect 5650 4465 5665 4485
rect 5685 4465 5700 4485
rect 5650 4435 5700 4465
rect 5650 4415 5665 4435
rect 5685 4415 5700 4435
rect 5650 4385 5700 4415
rect 5650 4365 5665 4385
rect 5685 4365 5700 4385
rect 5650 4350 5700 4365
rect 5800 4835 5850 4850
rect 5800 4815 5815 4835
rect 5835 4815 5850 4835
rect 5800 4785 5850 4815
rect 5800 4765 5815 4785
rect 5835 4765 5850 4785
rect 5800 4735 5850 4765
rect 5800 4715 5815 4735
rect 5835 4715 5850 4735
rect 5800 4685 5850 4715
rect 5800 4665 5815 4685
rect 5835 4665 5850 4685
rect 5800 4635 5850 4665
rect 5800 4615 5815 4635
rect 5835 4615 5850 4635
rect 5800 4585 5850 4615
rect 5800 4565 5815 4585
rect 5835 4565 5850 4585
rect 5800 4535 5850 4565
rect 5800 4515 5815 4535
rect 5835 4515 5850 4535
rect 5800 4485 5850 4515
rect 5800 4465 5815 4485
rect 5835 4465 5850 4485
rect 5800 4435 5850 4465
rect 5800 4415 5815 4435
rect 5835 4415 5850 4435
rect 5800 4385 5850 4415
rect 5800 4365 5815 4385
rect 5835 4365 5850 4385
rect 5800 4350 5850 4365
rect 5950 4835 6000 4850
rect 5950 4815 5965 4835
rect 5985 4815 6000 4835
rect 5950 4785 6000 4815
rect 5950 4765 5965 4785
rect 5985 4765 6000 4785
rect 5950 4735 6000 4765
rect 5950 4715 5965 4735
rect 5985 4715 6000 4735
rect 5950 4685 6000 4715
rect 5950 4665 5965 4685
rect 5985 4665 6000 4685
rect 5950 4635 6000 4665
rect 5950 4615 5965 4635
rect 5985 4615 6000 4635
rect 5950 4585 6000 4615
rect 5950 4565 5965 4585
rect 5985 4565 6000 4585
rect 5950 4535 6000 4565
rect 5950 4515 5965 4535
rect 5985 4515 6000 4535
rect 5950 4485 6000 4515
rect 5950 4465 5965 4485
rect 5985 4465 6000 4485
rect 5950 4435 6000 4465
rect 5950 4415 5965 4435
rect 5985 4415 6000 4435
rect 5950 4385 6000 4415
rect 5950 4365 5965 4385
rect 5985 4365 6000 4385
rect 5950 4350 6000 4365
rect 6100 4835 6150 4850
rect 6100 4815 6115 4835
rect 6135 4815 6150 4835
rect 6100 4785 6150 4815
rect 6100 4765 6115 4785
rect 6135 4765 6150 4785
rect 6100 4735 6150 4765
rect 6100 4715 6115 4735
rect 6135 4715 6150 4735
rect 6100 4685 6150 4715
rect 6100 4665 6115 4685
rect 6135 4665 6150 4685
rect 6100 4635 6150 4665
rect 6100 4615 6115 4635
rect 6135 4615 6150 4635
rect 6100 4585 6150 4615
rect 6100 4565 6115 4585
rect 6135 4565 6150 4585
rect 6100 4535 6150 4565
rect 6100 4515 6115 4535
rect 6135 4515 6150 4535
rect 6100 4485 6150 4515
rect 6100 4465 6115 4485
rect 6135 4465 6150 4485
rect 6100 4435 6150 4465
rect 6100 4415 6115 4435
rect 6135 4415 6150 4435
rect 6100 4385 6150 4415
rect 6100 4365 6115 4385
rect 6135 4365 6150 4385
rect 6100 4350 6150 4365
rect 6250 4835 6300 4850
rect 6250 4815 6265 4835
rect 6285 4815 6300 4835
rect 6250 4785 6300 4815
rect 6250 4765 6265 4785
rect 6285 4765 6300 4785
rect 6250 4735 6300 4765
rect 6250 4715 6265 4735
rect 6285 4715 6300 4735
rect 6250 4685 6300 4715
rect 6250 4665 6265 4685
rect 6285 4665 6300 4685
rect 6250 4635 6300 4665
rect 6250 4615 6265 4635
rect 6285 4615 6300 4635
rect 6250 4585 6300 4615
rect 6250 4565 6265 4585
rect 6285 4565 6300 4585
rect 6250 4535 6300 4565
rect 6250 4515 6265 4535
rect 6285 4515 6300 4535
rect 6250 4485 6300 4515
rect 6250 4465 6265 4485
rect 6285 4465 6300 4485
rect 6250 4435 6300 4465
rect 6250 4415 6265 4435
rect 6285 4415 6300 4435
rect 6250 4385 6300 4415
rect 6250 4365 6265 4385
rect 6285 4365 6300 4385
rect 6250 4350 6300 4365
rect 6400 4835 6450 4850
rect 6400 4815 6415 4835
rect 6435 4815 6450 4835
rect 6400 4785 6450 4815
rect 6400 4765 6415 4785
rect 6435 4765 6450 4785
rect 6400 4735 6450 4765
rect 6400 4715 6415 4735
rect 6435 4715 6450 4735
rect 6400 4685 6450 4715
rect 6400 4665 6415 4685
rect 6435 4665 6450 4685
rect 6400 4635 6450 4665
rect 6400 4615 6415 4635
rect 6435 4615 6450 4635
rect 6400 4585 6450 4615
rect 6400 4565 6415 4585
rect 6435 4565 6450 4585
rect 6400 4535 6450 4565
rect 6400 4515 6415 4535
rect 6435 4515 6450 4535
rect 6400 4485 6450 4515
rect 6400 4465 6415 4485
rect 6435 4465 6450 4485
rect 6400 4435 6450 4465
rect 6400 4415 6415 4435
rect 6435 4415 6450 4435
rect 6400 4385 6450 4415
rect 6400 4365 6415 4385
rect 6435 4365 6450 4385
rect 6400 4350 6450 4365
rect 6550 4835 6600 4850
rect 6550 4815 6565 4835
rect 6585 4815 6600 4835
rect 6550 4785 6600 4815
rect 6550 4765 6565 4785
rect 6585 4765 6600 4785
rect 6550 4735 6600 4765
rect 6550 4715 6565 4735
rect 6585 4715 6600 4735
rect 6550 4685 6600 4715
rect 6550 4665 6565 4685
rect 6585 4665 6600 4685
rect 6550 4635 6600 4665
rect 6550 4615 6565 4635
rect 6585 4615 6600 4635
rect 6550 4585 6600 4615
rect 6550 4565 6565 4585
rect 6585 4565 6600 4585
rect 6550 4535 6600 4565
rect 6550 4515 6565 4535
rect 6585 4515 6600 4535
rect 6550 4485 6600 4515
rect 6550 4465 6565 4485
rect 6585 4465 6600 4485
rect 6550 4435 6600 4465
rect 6550 4415 6565 4435
rect 6585 4415 6600 4435
rect 6550 4385 6600 4415
rect 6550 4365 6565 4385
rect 6585 4365 6600 4385
rect 6550 4350 6600 4365
rect 6700 4835 6750 4850
rect 6700 4815 6715 4835
rect 6735 4815 6750 4835
rect 6700 4785 6750 4815
rect 6700 4765 6715 4785
rect 6735 4765 6750 4785
rect 6700 4735 6750 4765
rect 6700 4715 6715 4735
rect 6735 4715 6750 4735
rect 6700 4685 6750 4715
rect 6700 4665 6715 4685
rect 6735 4665 6750 4685
rect 6700 4635 6750 4665
rect 6700 4615 6715 4635
rect 6735 4615 6750 4635
rect 6700 4585 6750 4615
rect 6700 4565 6715 4585
rect 6735 4565 6750 4585
rect 6700 4535 6750 4565
rect 6700 4515 6715 4535
rect 6735 4515 6750 4535
rect 6700 4485 6750 4515
rect 6700 4465 6715 4485
rect 6735 4465 6750 4485
rect 6700 4435 6750 4465
rect 6700 4415 6715 4435
rect 6735 4415 6750 4435
rect 6700 4385 6750 4415
rect 6700 4365 6715 4385
rect 6735 4365 6750 4385
rect 6700 4350 6750 4365
rect 6850 4835 6900 4850
rect 6850 4815 6865 4835
rect 6885 4815 6900 4835
rect 6850 4785 6900 4815
rect 6850 4765 6865 4785
rect 6885 4765 6900 4785
rect 6850 4735 6900 4765
rect 6850 4715 6865 4735
rect 6885 4715 6900 4735
rect 6850 4685 6900 4715
rect 6850 4665 6865 4685
rect 6885 4665 6900 4685
rect 6850 4635 6900 4665
rect 6850 4615 6865 4635
rect 6885 4615 6900 4635
rect 6850 4585 6900 4615
rect 6850 4565 6865 4585
rect 6885 4565 6900 4585
rect 6850 4535 6900 4565
rect 6850 4515 6865 4535
rect 6885 4515 6900 4535
rect 6850 4485 6900 4515
rect 6850 4465 6865 4485
rect 6885 4465 6900 4485
rect 6850 4435 6900 4465
rect 6850 4415 6865 4435
rect 6885 4415 6900 4435
rect 6850 4385 6900 4415
rect 6850 4365 6865 4385
rect 6885 4365 6900 4385
rect 6850 4350 6900 4365
rect 7000 4835 7050 4850
rect 7000 4815 7015 4835
rect 7035 4815 7050 4835
rect 7000 4785 7050 4815
rect 7000 4765 7015 4785
rect 7035 4765 7050 4785
rect 7000 4735 7050 4765
rect 7000 4715 7015 4735
rect 7035 4715 7050 4735
rect 7000 4685 7050 4715
rect 7000 4665 7015 4685
rect 7035 4665 7050 4685
rect 7000 4635 7050 4665
rect 7000 4615 7015 4635
rect 7035 4615 7050 4635
rect 7000 4585 7050 4615
rect 7000 4565 7015 4585
rect 7035 4565 7050 4585
rect 7000 4535 7050 4565
rect 7000 4515 7015 4535
rect 7035 4515 7050 4535
rect 7000 4485 7050 4515
rect 7000 4465 7015 4485
rect 7035 4465 7050 4485
rect 7000 4435 7050 4465
rect 7000 4415 7015 4435
rect 7035 4415 7050 4435
rect 7000 4385 7050 4415
rect 7000 4365 7015 4385
rect 7035 4365 7050 4385
rect 7000 4350 7050 4365
rect 7150 4835 7200 4850
rect 7150 4815 7165 4835
rect 7185 4815 7200 4835
rect 7150 4785 7200 4815
rect 7150 4765 7165 4785
rect 7185 4765 7200 4785
rect 7150 4735 7200 4765
rect 7150 4715 7165 4735
rect 7185 4715 7200 4735
rect 7150 4685 7200 4715
rect 7150 4665 7165 4685
rect 7185 4665 7200 4685
rect 7150 4635 7200 4665
rect 7150 4615 7165 4635
rect 7185 4615 7200 4635
rect 7150 4585 7200 4615
rect 7150 4565 7165 4585
rect 7185 4565 7200 4585
rect 7150 4535 7200 4565
rect 7150 4515 7165 4535
rect 7185 4515 7200 4535
rect 7150 4485 7200 4515
rect 7150 4465 7165 4485
rect 7185 4465 7200 4485
rect 7150 4435 7200 4465
rect 7150 4415 7165 4435
rect 7185 4415 7200 4435
rect 7150 4385 7200 4415
rect 7150 4365 7165 4385
rect 7185 4365 7200 4385
rect 7150 4350 7200 4365
rect 7300 4835 7350 4850
rect 7300 4815 7315 4835
rect 7335 4815 7350 4835
rect 7300 4785 7350 4815
rect 7300 4765 7315 4785
rect 7335 4765 7350 4785
rect 7300 4735 7350 4765
rect 7300 4715 7315 4735
rect 7335 4715 7350 4735
rect 7300 4685 7350 4715
rect 7300 4665 7315 4685
rect 7335 4665 7350 4685
rect 7300 4635 7350 4665
rect 7300 4615 7315 4635
rect 7335 4615 7350 4635
rect 7300 4585 7350 4615
rect 7300 4565 7315 4585
rect 7335 4565 7350 4585
rect 7300 4535 7350 4565
rect 7300 4515 7315 4535
rect 7335 4515 7350 4535
rect 7300 4485 7350 4515
rect 7300 4465 7315 4485
rect 7335 4465 7350 4485
rect 7300 4435 7350 4465
rect 7300 4415 7315 4435
rect 7335 4415 7350 4435
rect 7300 4385 7350 4415
rect 7300 4365 7315 4385
rect 7335 4365 7350 4385
rect 7300 4350 7350 4365
rect 7450 4835 7500 4850
rect 7450 4815 7465 4835
rect 7485 4815 7500 4835
rect 7450 4785 7500 4815
rect 7450 4765 7465 4785
rect 7485 4765 7500 4785
rect 7450 4735 7500 4765
rect 7450 4715 7465 4735
rect 7485 4715 7500 4735
rect 7450 4685 7500 4715
rect 7450 4665 7465 4685
rect 7485 4665 7500 4685
rect 7450 4635 7500 4665
rect 7450 4615 7465 4635
rect 7485 4615 7500 4635
rect 7450 4585 7500 4615
rect 7450 4565 7465 4585
rect 7485 4565 7500 4585
rect 7450 4535 7500 4565
rect 7450 4515 7465 4535
rect 7485 4515 7500 4535
rect 7450 4485 7500 4515
rect 7450 4465 7465 4485
rect 7485 4465 7500 4485
rect 7450 4435 7500 4465
rect 7450 4415 7465 4435
rect 7485 4415 7500 4435
rect 7450 4385 7500 4415
rect 7450 4365 7465 4385
rect 7485 4365 7500 4385
rect 7450 4350 7500 4365
rect 7600 4835 7650 4850
rect 7600 4815 7615 4835
rect 7635 4815 7650 4835
rect 7600 4785 7650 4815
rect 7600 4765 7615 4785
rect 7635 4765 7650 4785
rect 7600 4735 7650 4765
rect 7600 4715 7615 4735
rect 7635 4715 7650 4735
rect 7600 4685 7650 4715
rect 7600 4665 7615 4685
rect 7635 4665 7650 4685
rect 7600 4635 7650 4665
rect 7600 4615 7615 4635
rect 7635 4615 7650 4635
rect 7600 4585 7650 4615
rect 7600 4565 7615 4585
rect 7635 4565 7650 4585
rect 7600 4535 7650 4565
rect 7600 4515 7615 4535
rect 7635 4515 7650 4535
rect 7600 4485 7650 4515
rect 7600 4465 7615 4485
rect 7635 4465 7650 4485
rect 7600 4435 7650 4465
rect 7600 4415 7615 4435
rect 7635 4415 7650 4435
rect 7600 4385 7650 4415
rect 7600 4365 7615 4385
rect 7635 4365 7650 4385
rect 7600 4350 7650 4365
rect 7750 4835 7800 4850
rect 7750 4815 7765 4835
rect 7785 4815 7800 4835
rect 7750 4785 7800 4815
rect 7750 4765 7765 4785
rect 7785 4765 7800 4785
rect 7750 4735 7800 4765
rect 7750 4715 7765 4735
rect 7785 4715 7800 4735
rect 7750 4685 7800 4715
rect 7750 4665 7765 4685
rect 7785 4665 7800 4685
rect 7750 4635 7800 4665
rect 7750 4615 7765 4635
rect 7785 4615 7800 4635
rect 7750 4585 7800 4615
rect 7750 4565 7765 4585
rect 7785 4565 7800 4585
rect 7750 4535 7800 4565
rect 7750 4515 7765 4535
rect 7785 4515 7800 4535
rect 7750 4485 7800 4515
rect 7750 4465 7765 4485
rect 7785 4465 7800 4485
rect 7750 4435 7800 4465
rect 7750 4415 7765 4435
rect 7785 4415 7800 4435
rect 7750 4385 7800 4415
rect 7750 4365 7765 4385
rect 7785 4365 7800 4385
rect 7750 4350 7800 4365
rect 8350 4835 8400 4850
rect 8350 4815 8365 4835
rect 8385 4815 8400 4835
rect 8350 4785 8400 4815
rect 8350 4765 8365 4785
rect 8385 4765 8400 4785
rect 8350 4735 8400 4765
rect 8350 4715 8365 4735
rect 8385 4715 8400 4735
rect 8350 4685 8400 4715
rect 8350 4665 8365 4685
rect 8385 4665 8400 4685
rect 8350 4635 8400 4665
rect 8350 4615 8365 4635
rect 8385 4615 8400 4635
rect 8350 4585 8400 4615
rect 8350 4565 8365 4585
rect 8385 4565 8400 4585
rect 8350 4535 8400 4565
rect 8350 4515 8365 4535
rect 8385 4515 8400 4535
rect 8350 4485 8400 4515
rect 8350 4465 8365 4485
rect 8385 4465 8400 4485
rect 8350 4435 8400 4465
rect 8350 4415 8365 4435
rect 8385 4415 8400 4435
rect 8350 4385 8400 4415
rect 8350 4365 8365 4385
rect 8385 4365 8400 4385
rect 8350 4350 8400 4365
rect 8500 4835 8550 4900
rect 8500 4815 8515 4835
rect 8535 4815 8550 4835
rect 8500 4785 8550 4815
rect 8500 4765 8515 4785
rect 8535 4765 8550 4785
rect 8500 4735 8550 4765
rect 8500 4715 8515 4735
rect 8535 4715 8550 4735
rect 8500 4685 8550 4715
rect 8500 4665 8515 4685
rect 8535 4665 8550 4685
rect 8500 4635 8550 4665
rect 8500 4615 8515 4635
rect 8535 4615 8550 4635
rect 8500 4585 8550 4615
rect 8500 4565 8515 4585
rect 8535 4565 8550 4585
rect 8500 4535 8550 4565
rect 8500 4515 8515 4535
rect 8535 4515 8550 4535
rect 8500 4485 8550 4515
rect 8500 4465 8515 4485
rect 8535 4465 8550 4485
rect 8500 4435 8550 4465
rect 8500 4415 8515 4435
rect 8535 4415 8550 4435
rect 8500 4385 8550 4415
rect 8500 4365 8515 4385
rect 8535 4365 8550 4385
rect 8500 4350 8550 4365
rect 8650 4835 8700 4850
rect 8650 4815 8665 4835
rect 8685 4815 8700 4835
rect 8650 4785 8700 4815
rect 8650 4765 8665 4785
rect 8685 4765 8700 4785
rect 8650 4735 8700 4765
rect 8650 4715 8665 4735
rect 8685 4715 8700 4735
rect 8650 4685 8700 4715
rect 8650 4665 8665 4685
rect 8685 4665 8700 4685
rect 8650 4635 8700 4665
rect 8650 4615 8665 4635
rect 8685 4615 8700 4635
rect 8650 4585 8700 4615
rect 8650 4565 8665 4585
rect 8685 4565 8700 4585
rect 8650 4535 8700 4565
rect 8650 4515 8665 4535
rect 8685 4515 8700 4535
rect 8650 4485 8700 4515
rect 8650 4465 8665 4485
rect 8685 4465 8700 4485
rect 8650 4435 8700 4465
rect 8650 4415 8665 4435
rect 8685 4415 8700 4435
rect 8650 4385 8700 4415
rect 8650 4365 8665 4385
rect 8685 4365 8700 4385
rect 8650 4350 8700 4365
rect 8800 4835 8850 4900
rect 8800 4815 8815 4835
rect 8835 4815 8850 4835
rect 8800 4785 8850 4815
rect 8800 4765 8815 4785
rect 8835 4765 8850 4785
rect 8800 4735 8850 4765
rect 8800 4715 8815 4735
rect 8835 4715 8850 4735
rect 8800 4685 8850 4715
rect 8800 4665 8815 4685
rect 8835 4665 8850 4685
rect 8800 4635 8850 4665
rect 8800 4615 8815 4635
rect 8835 4615 8850 4635
rect 8800 4585 8850 4615
rect 8800 4565 8815 4585
rect 8835 4565 8850 4585
rect 8800 4535 8850 4565
rect 8800 4515 8815 4535
rect 8835 4515 8850 4535
rect 8800 4485 8850 4515
rect 8800 4465 8815 4485
rect 8835 4465 8850 4485
rect 8800 4435 8850 4465
rect 8800 4415 8815 4435
rect 8835 4415 8850 4435
rect 8800 4385 8850 4415
rect 8800 4365 8815 4385
rect 8835 4365 8850 4385
rect 8800 4350 8850 4365
rect 8950 4835 9000 4850
rect 8950 4815 8965 4835
rect 8985 4815 9000 4835
rect 8950 4785 9000 4815
rect 8950 4765 8965 4785
rect 8985 4765 9000 4785
rect 8950 4735 9000 4765
rect 8950 4715 8965 4735
rect 8985 4715 9000 4735
rect 8950 4685 9000 4715
rect 8950 4665 8965 4685
rect 8985 4665 9000 4685
rect 8950 4635 9000 4665
rect 8950 4615 8965 4635
rect 8985 4615 9000 4635
rect 8950 4585 9000 4615
rect 8950 4565 8965 4585
rect 8985 4565 9000 4585
rect 8950 4535 9000 4565
rect 8950 4515 8965 4535
rect 8985 4515 9000 4535
rect 8950 4485 9000 4515
rect 8950 4465 8965 4485
rect 8985 4465 9000 4485
rect 8950 4435 9000 4465
rect 8950 4415 8965 4435
rect 8985 4415 9000 4435
rect 8950 4385 9000 4415
rect 8950 4365 8965 4385
rect 8985 4365 9000 4385
rect 8950 4350 9000 4365
rect 9100 4835 9150 4900
rect 9100 4815 9115 4835
rect 9135 4815 9150 4835
rect 9100 4785 9150 4815
rect 9100 4765 9115 4785
rect 9135 4765 9150 4785
rect 9100 4735 9150 4765
rect 9100 4715 9115 4735
rect 9135 4715 9150 4735
rect 9100 4685 9150 4715
rect 9100 4665 9115 4685
rect 9135 4665 9150 4685
rect 9100 4635 9150 4665
rect 9100 4615 9115 4635
rect 9135 4615 9150 4635
rect 9100 4585 9150 4615
rect 9100 4565 9115 4585
rect 9135 4565 9150 4585
rect 9100 4535 9150 4565
rect 9100 4515 9115 4535
rect 9135 4515 9150 4535
rect 9100 4485 9150 4515
rect 9100 4465 9115 4485
rect 9135 4465 9150 4485
rect 9100 4435 9150 4465
rect 9100 4415 9115 4435
rect 9135 4415 9150 4435
rect 9100 4385 9150 4415
rect 9100 4365 9115 4385
rect 9135 4365 9150 4385
rect 9100 4350 9150 4365
rect 9250 4835 9300 4850
rect 9250 4815 9265 4835
rect 9285 4815 9300 4835
rect 9250 4785 9300 4815
rect 9250 4765 9265 4785
rect 9285 4765 9300 4785
rect 9250 4735 9300 4765
rect 9250 4715 9265 4735
rect 9285 4715 9300 4735
rect 9250 4685 9300 4715
rect 9250 4665 9265 4685
rect 9285 4665 9300 4685
rect 9250 4635 9300 4665
rect 9250 4615 9265 4635
rect 9285 4615 9300 4635
rect 9250 4585 9300 4615
rect 9250 4565 9265 4585
rect 9285 4565 9300 4585
rect 9250 4535 9300 4565
rect 9250 4515 9265 4535
rect 9285 4515 9300 4535
rect 9250 4485 9300 4515
rect 9250 4465 9265 4485
rect 9285 4465 9300 4485
rect 9250 4435 9300 4465
rect 9250 4415 9265 4435
rect 9285 4415 9300 4435
rect 9250 4385 9300 4415
rect 9250 4365 9265 4385
rect 9285 4365 9300 4385
rect 9250 4350 9300 4365
rect 9400 4835 9450 4900
rect 9400 4815 9415 4835
rect 9435 4815 9450 4835
rect 9400 4785 9450 4815
rect 9400 4765 9415 4785
rect 9435 4765 9450 4785
rect 9400 4735 9450 4765
rect 9400 4715 9415 4735
rect 9435 4715 9450 4735
rect 9400 4685 9450 4715
rect 9400 4665 9415 4685
rect 9435 4665 9450 4685
rect 9400 4635 9450 4665
rect 9400 4615 9415 4635
rect 9435 4615 9450 4635
rect 9400 4585 9450 4615
rect 9400 4565 9415 4585
rect 9435 4565 9450 4585
rect 9400 4535 9450 4565
rect 9400 4515 9415 4535
rect 9435 4515 9450 4535
rect 9400 4485 9450 4515
rect 9400 4465 9415 4485
rect 9435 4465 9450 4485
rect 9400 4435 9450 4465
rect 9400 4415 9415 4435
rect 9435 4415 9450 4435
rect 9400 4385 9450 4415
rect 9400 4365 9415 4385
rect 9435 4365 9450 4385
rect 9400 4350 9450 4365
rect 9550 4835 9600 4850
rect 9550 4815 9565 4835
rect 9585 4815 9600 4835
rect 9550 4785 9600 4815
rect 9550 4765 9565 4785
rect 9585 4765 9600 4785
rect 9550 4735 9600 4765
rect 9550 4715 9565 4735
rect 9585 4715 9600 4735
rect 9550 4685 9600 4715
rect 9550 4665 9565 4685
rect 9585 4665 9600 4685
rect 9550 4635 9600 4665
rect 9550 4615 9565 4635
rect 9585 4615 9600 4635
rect 9550 4585 9600 4615
rect 9550 4565 9565 4585
rect 9585 4565 9600 4585
rect 9550 4535 9600 4565
rect 9550 4515 9565 4535
rect 9585 4515 9600 4535
rect 9550 4485 9600 4515
rect 9550 4465 9565 4485
rect 9585 4465 9600 4485
rect 9550 4435 9600 4465
rect 9550 4415 9565 4435
rect 9585 4415 9600 4435
rect 9550 4385 9600 4415
rect 9550 4365 9565 4385
rect 9585 4365 9600 4385
rect 9550 4350 9600 4365
rect 9700 4835 9750 4900
rect 9700 4815 9715 4835
rect 9735 4815 9750 4835
rect 9700 4785 9750 4815
rect 9700 4765 9715 4785
rect 9735 4765 9750 4785
rect 9700 4735 9750 4765
rect 9700 4715 9715 4735
rect 9735 4715 9750 4735
rect 9700 4685 9750 4715
rect 9700 4665 9715 4685
rect 9735 4665 9750 4685
rect 9700 4635 9750 4665
rect 9700 4615 9715 4635
rect 9735 4615 9750 4635
rect 9700 4585 9750 4615
rect 9700 4565 9715 4585
rect 9735 4565 9750 4585
rect 9700 4535 9750 4565
rect 9700 4515 9715 4535
rect 9735 4515 9750 4535
rect 9700 4485 9750 4515
rect 9700 4465 9715 4485
rect 9735 4465 9750 4485
rect 9700 4435 9750 4465
rect 9700 4415 9715 4435
rect 9735 4415 9750 4435
rect 9700 4385 9750 4415
rect 9700 4365 9715 4385
rect 9735 4365 9750 4385
rect 9700 4350 9750 4365
rect 9850 4835 9900 4850
rect 9850 4815 9865 4835
rect 9885 4815 9900 4835
rect 9850 4785 9900 4815
rect 9850 4765 9865 4785
rect 9885 4765 9900 4785
rect 9850 4735 9900 4765
rect 9850 4715 9865 4735
rect 9885 4715 9900 4735
rect 9850 4685 9900 4715
rect 9850 4665 9865 4685
rect 9885 4665 9900 4685
rect 9850 4635 9900 4665
rect 9850 4615 9865 4635
rect 9885 4615 9900 4635
rect 9850 4585 9900 4615
rect 9850 4565 9865 4585
rect 9885 4565 9900 4585
rect 9850 4535 9900 4565
rect 9850 4515 9865 4535
rect 9885 4515 9900 4535
rect 9850 4485 9900 4515
rect 9850 4465 9865 4485
rect 9885 4465 9900 4485
rect 9850 4435 9900 4465
rect 9850 4415 9865 4435
rect 9885 4415 9900 4435
rect 9850 4385 9900 4415
rect 9850 4365 9865 4385
rect 9885 4365 9900 4385
rect 9850 4350 9900 4365
rect 10000 4835 10050 4900
rect 10000 4815 10015 4835
rect 10035 4815 10050 4835
rect 10000 4785 10050 4815
rect 10000 4765 10015 4785
rect 10035 4765 10050 4785
rect 10000 4735 10050 4765
rect 10000 4715 10015 4735
rect 10035 4715 10050 4735
rect 10000 4685 10050 4715
rect 10000 4665 10015 4685
rect 10035 4665 10050 4685
rect 10000 4635 10050 4665
rect 10000 4615 10015 4635
rect 10035 4615 10050 4635
rect 10000 4585 10050 4615
rect 10000 4565 10015 4585
rect 10035 4565 10050 4585
rect 10000 4535 10050 4565
rect 10000 4515 10015 4535
rect 10035 4515 10050 4535
rect 10000 4485 10050 4515
rect 10000 4465 10015 4485
rect 10035 4465 10050 4485
rect 10000 4435 10050 4465
rect 10000 4415 10015 4435
rect 10035 4415 10050 4435
rect 10000 4385 10050 4415
rect 10000 4365 10015 4385
rect 10035 4365 10050 4385
rect 10000 4350 10050 4365
rect 10150 4835 10200 4850
rect 10150 4815 10165 4835
rect 10185 4815 10200 4835
rect 10150 4785 10200 4815
rect 10150 4765 10165 4785
rect 10185 4765 10200 4785
rect 10150 4735 10200 4765
rect 10150 4715 10165 4735
rect 10185 4715 10200 4735
rect 10150 4685 10200 4715
rect 10150 4665 10165 4685
rect 10185 4665 10200 4685
rect 10150 4635 10200 4665
rect 10150 4615 10165 4635
rect 10185 4615 10200 4635
rect 10150 4585 10200 4615
rect 10150 4565 10165 4585
rect 10185 4565 10200 4585
rect 10150 4535 10200 4565
rect 10150 4515 10165 4535
rect 10185 4515 10200 4535
rect 10150 4485 10200 4515
rect 10150 4465 10165 4485
rect 10185 4465 10200 4485
rect 10150 4435 10200 4465
rect 10150 4415 10165 4435
rect 10185 4415 10200 4435
rect 10150 4385 10200 4415
rect 10150 4365 10165 4385
rect 10185 4365 10200 4385
rect 10150 4350 10200 4365
rect 10300 4835 10350 4900
rect 10300 4815 10315 4835
rect 10335 4815 10350 4835
rect 10300 4785 10350 4815
rect 10300 4765 10315 4785
rect 10335 4765 10350 4785
rect 10300 4735 10350 4765
rect 10300 4715 10315 4735
rect 10335 4715 10350 4735
rect 10300 4685 10350 4715
rect 10300 4665 10315 4685
rect 10335 4665 10350 4685
rect 10300 4635 10350 4665
rect 10300 4615 10315 4635
rect 10335 4615 10350 4635
rect 10300 4585 10350 4615
rect 10300 4565 10315 4585
rect 10335 4565 10350 4585
rect 10300 4535 10350 4565
rect 10300 4515 10315 4535
rect 10335 4515 10350 4535
rect 10300 4485 10350 4515
rect 10300 4465 10315 4485
rect 10335 4465 10350 4485
rect 10300 4435 10350 4465
rect 10300 4415 10315 4435
rect 10335 4415 10350 4435
rect 10300 4385 10350 4415
rect 10300 4365 10315 4385
rect 10335 4365 10350 4385
rect 10300 4350 10350 4365
rect 10450 4835 10500 4850
rect 10450 4815 10465 4835
rect 10485 4815 10500 4835
rect 10450 4785 10500 4815
rect 10450 4765 10465 4785
rect 10485 4765 10500 4785
rect 10450 4735 10500 4765
rect 10450 4715 10465 4735
rect 10485 4715 10500 4735
rect 10450 4685 10500 4715
rect 10450 4665 10465 4685
rect 10485 4665 10500 4685
rect 10450 4635 10500 4665
rect 10450 4615 10465 4635
rect 10485 4615 10500 4635
rect 10450 4585 10500 4615
rect 10450 4565 10465 4585
rect 10485 4565 10500 4585
rect 10450 4535 10500 4565
rect 10450 4515 10465 4535
rect 10485 4515 10500 4535
rect 10450 4485 10500 4515
rect 10450 4465 10465 4485
rect 10485 4465 10500 4485
rect 10450 4435 10500 4465
rect 10450 4415 10465 4435
rect 10485 4415 10500 4435
rect 10450 4385 10500 4415
rect 10450 4365 10465 4385
rect 10485 4365 10500 4385
rect 10450 4350 10500 4365
rect 10600 4835 10650 4900
rect 10600 4815 10615 4835
rect 10635 4815 10650 4835
rect 10600 4785 10650 4815
rect 10600 4765 10615 4785
rect 10635 4765 10650 4785
rect 10600 4735 10650 4765
rect 10600 4715 10615 4735
rect 10635 4715 10650 4735
rect 10600 4685 10650 4715
rect 10600 4665 10615 4685
rect 10635 4665 10650 4685
rect 10600 4635 10650 4665
rect 10600 4615 10615 4635
rect 10635 4615 10650 4635
rect 10600 4585 10650 4615
rect 10600 4565 10615 4585
rect 10635 4565 10650 4585
rect 10600 4535 10650 4565
rect 10600 4515 10615 4535
rect 10635 4515 10650 4535
rect 10600 4485 10650 4515
rect 10600 4465 10615 4485
rect 10635 4465 10650 4485
rect 10600 4435 10650 4465
rect 10600 4415 10615 4435
rect 10635 4415 10650 4435
rect 10600 4385 10650 4415
rect 10600 4365 10615 4385
rect 10635 4365 10650 4385
rect 10600 4350 10650 4365
rect 10750 4835 10800 4850
rect 10750 4815 10765 4835
rect 10785 4815 10800 4835
rect 10750 4785 10800 4815
rect 10750 4765 10765 4785
rect 10785 4765 10800 4785
rect 10750 4735 10800 4765
rect 10750 4715 10765 4735
rect 10785 4715 10800 4735
rect 10750 4685 10800 4715
rect 10750 4665 10765 4685
rect 10785 4665 10800 4685
rect 10750 4635 10800 4665
rect 10750 4615 10765 4635
rect 10785 4615 10800 4635
rect 10750 4585 10800 4615
rect 10750 4565 10765 4585
rect 10785 4565 10800 4585
rect 10750 4535 10800 4565
rect 10750 4515 10765 4535
rect 10785 4515 10800 4535
rect 10750 4485 10800 4515
rect 10750 4465 10765 4485
rect 10785 4465 10800 4485
rect 10750 4435 10800 4465
rect 10750 4415 10765 4435
rect 10785 4415 10800 4435
rect 10750 4385 10800 4415
rect 10750 4365 10765 4385
rect 10785 4365 10800 4385
rect 10750 4350 10800 4365
rect 11350 4835 11400 4850
rect 11350 4815 11365 4835
rect 11385 4815 11400 4835
rect 11350 4785 11400 4815
rect 11350 4765 11365 4785
rect 11385 4765 11400 4785
rect 11350 4735 11400 4765
rect 11350 4715 11365 4735
rect 11385 4715 11400 4735
rect 11350 4685 11400 4715
rect 11350 4665 11365 4685
rect 11385 4665 11400 4685
rect 11350 4635 11400 4665
rect 11350 4615 11365 4635
rect 11385 4615 11400 4635
rect 11350 4585 11400 4615
rect 11350 4565 11365 4585
rect 11385 4565 11400 4585
rect 11350 4535 11400 4565
rect 11350 4515 11365 4535
rect 11385 4515 11400 4535
rect 11350 4485 11400 4515
rect 11350 4465 11365 4485
rect 11385 4465 11400 4485
rect 11350 4435 11400 4465
rect 11350 4415 11365 4435
rect 11385 4415 11400 4435
rect 11350 4385 11400 4415
rect 11350 4365 11365 4385
rect 11385 4365 11400 4385
rect 11350 4350 11400 4365
rect 11950 4835 12000 4850
rect 11950 4815 11965 4835
rect 11985 4815 12000 4835
rect 11950 4785 12000 4815
rect 11950 4765 11965 4785
rect 11985 4765 12000 4785
rect 11950 4735 12000 4765
rect 11950 4715 11965 4735
rect 11985 4715 12000 4735
rect 11950 4685 12000 4715
rect 11950 4665 11965 4685
rect 11985 4665 12000 4685
rect 11950 4635 12000 4665
rect 11950 4615 11965 4635
rect 11985 4615 12000 4635
rect 11950 4585 12000 4615
rect 11950 4565 11965 4585
rect 11985 4565 12000 4585
rect 11950 4535 12000 4565
rect 11950 4515 11965 4535
rect 11985 4515 12000 4535
rect 11950 4485 12000 4515
rect 11950 4465 11965 4485
rect 11985 4465 12000 4485
rect 11950 4435 12000 4465
rect 11950 4415 11965 4435
rect 11985 4415 12000 4435
rect 11950 4385 12000 4415
rect 11950 4365 11965 4385
rect 11985 4365 12000 4385
rect 11950 4350 12000 4365
rect 12550 4835 12600 4850
rect 12550 4815 12565 4835
rect 12585 4815 12600 4835
rect 12550 4785 12600 4815
rect 12550 4765 12565 4785
rect 12585 4765 12600 4785
rect 12550 4735 12600 4765
rect 12550 4715 12565 4735
rect 12585 4715 12600 4735
rect 12550 4685 12600 4715
rect 12550 4665 12565 4685
rect 12585 4665 12600 4685
rect 12550 4635 12600 4665
rect 12550 4615 12565 4635
rect 12585 4615 12600 4635
rect 12550 4585 12600 4615
rect 12550 4565 12565 4585
rect 12585 4565 12600 4585
rect 12550 4535 12600 4565
rect 12550 4515 12565 4535
rect 12585 4515 12600 4535
rect 12550 4485 12600 4515
rect 12550 4465 12565 4485
rect 12585 4465 12600 4485
rect 12550 4435 12600 4465
rect 12550 4415 12565 4435
rect 12585 4415 12600 4435
rect 12550 4385 12600 4415
rect 12550 4365 12565 4385
rect 12585 4365 12600 4385
rect 12550 4350 12600 4365
rect 13150 4835 13200 4850
rect 13150 4815 13165 4835
rect 13185 4815 13200 4835
rect 13150 4785 13200 4815
rect 13150 4765 13165 4785
rect 13185 4765 13200 4785
rect 13150 4735 13200 4765
rect 13150 4715 13165 4735
rect 13185 4715 13200 4735
rect 13150 4685 13200 4715
rect 13150 4665 13165 4685
rect 13185 4665 13200 4685
rect 13150 4635 13200 4665
rect 13150 4615 13165 4635
rect 13185 4615 13200 4635
rect 13150 4585 13200 4615
rect 13150 4565 13165 4585
rect 13185 4565 13200 4585
rect 13150 4535 13200 4565
rect 13150 4515 13165 4535
rect 13185 4515 13200 4535
rect 13150 4485 13200 4515
rect 13150 4465 13165 4485
rect 13185 4465 13200 4485
rect 13150 4435 13200 4465
rect 13150 4415 13165 4435
rect 13185 4415 13200 4435
rect 13150 4385 13200 4415
rect 13150 4365 13165 4385
rect 13185 4365 13200 4385
rect 13150 4350 13200 4365
rect 13750 4835 13800 4850
rect 13750 4815 13765 4835
rect 13785 4815 13800 4835
rect 13750 4785 13800 4815
rect 13750 4765 13765 4785
rect 13785 4765 13800 4785
rect 13750 4735 13800 4765
rect 13750 4715 13765 4735
rect 13785 4715 13800 4735
rect 13750 4685 13800 4715
rect 13750 4665 13765 4685
rect 13785 4665 13800 4685
rect 13750 4635 13800 4665
rect 13750 4615 13765 4635
rect 13785 4615 13800 4635
rect 13750 4585 13800 4615
rect 13750 4565 13765 4585
rect 13785 4565 13800 4585
rect 13750 4535 13800 4565
rect 13750 4515 13765 4535
rect 13785 4515 13800 4535
rect 13750 4485 13800 4515
rect 13750 4465 13765 4485
rect 13785 4465 13800 4485
rect 13750 4435 13800 4465
rect 13750 4415 13765 4435
rect 13785 4415 13800 4435
rect 13750 4385 13800 4415
rect 13750 4365 13765 4385
rect 13785 4365 13800 4385
rect 13750 4350 13800 4365
rect 14350 4835 14400 4850
rect 14350 4815 14365 4835
rect 14385 4815 14400 4835
rect 14350 4785 14400 4815
rect 14350 4765 14365 4785
rect 14385 4765 14400 4785
rect 14350 4735 14400 4765
rect 14350 4715 14365 4735
rect 14385 4715 14400 4735
rect 14350 4685 14400 4715
rect 14350 4665 14365 4685
rect 14385 4665 14400 4685
rect 14350 4635 14400 4665
rect 14350 4615 14365 4635
rect 14385 4615 14400 4635
rect 14350 4585 14400 4615
rect 14350 4565 14365 4585
rect 14385 4565 14400 4585
rect 14350 4535 14400 4565
rect 14350 4515 14365 4535
rect 14385 4515 14400 4535
rect 14350 4485 14400 4515
rect 14350 4465 14365 4485
rect 14385 4465 14400 4485
rect 14350 4435 14400 4465
rect 14350 4415 14365 4435
rect 14385 4415 14400 4435
rect 14350 4385 14400 4415
rect 14350 4365 14365 4385
rect 14385 4365 14400 4385
rect 14350 4350 14400 4365
rect 14950 4835 15000 4850
rect 14950 4815 14965 4835
rect 14985 4815 15000 4835
rect 14950 4785 15000 4815
rect 14950 4765 14965 4785
rect 14985 4765 15000 4785
rect 14950 4735 15000 4765
rect 14950 4715 14965 4735
rect 14985 4715 15000 4735
rect 14950 4685 15000 4715
rect 14950 4665 14965 4685
rect 14985 4665 15000 4685
rect 14950 4635 15000 4665
rect 14950 4615 14965 4635
rect 14985 4615 15000 4635
rect 14950 4585 15000 4615
rect 14950 4565 14965 4585
rect 14985 4565 15000 4585
rect 14950 4535 15000 4565
rect 14950 4515 14965 4535
rect 14985 4515 15000 4535
rect 14950 4485 15000 4515
rect 14950 4465 14965 4485
rect 14985 4465 15000 4485
rect 14950 4435 15000 4465
rect 14950 4415 14965 4435
rect 14985 4415 15000 4435
rect 14950 4385 15000 4415
rect 14950 4365 14965 4385
rect 14985 4365 15000 4385
rect 14950 4350 15000 4365
rect 15550 4835 15600 4850
rect 15550 4815 15565 4835
rect 15585 4815 15600 4835
rect 15550 4785 15600 4815
rect 15550 4765 15565 4785
rect 15585 4765 15600 4785
rect 15550 4735 15600 4765
rect 15550 4715 15565 4735
rect 15585 4715 15600 4735
rect 15550 4685 15600 4715
rect 15550 4665 15565 4685
rect 15585 4665 15600 4685
rect 15550 4635 15600 4665
rect 15550 4615 15565 4635
rect 15585 4615 15600 4635
rect 15550 4585 15600 4615
rect 15550 4565 15565 4585
rect 15585 4565 15600 4585
rect 15550 4535 15600 4565
rect 15550 4515 15565 4535
rect 15585 4515 15600 4535
rect 15550 4485 15600 4515
rect 15550 4465 15565 4485
rect 15585 4465 15600 4485
rect 15550 4435 15600 4465
rect 15550 4415 15565 4435
rect 15585 4415 15600 4435
rect 15550 4385 15600 4415
rect 15550 4365 15565 4385
rect 15585 4365 15600 4385
rect 15550 4350 15600 4365
rect 16150 4835 16200 4850
rect 16150 4815 16165 4835
rect 16185 4815 16200 4835
rect 16150 4785 16200 4815
rect 16150 4765 16165 4785
rect 16185 4765 16200 4785
rect 16150 4735 16200 4765
rect 16150 4715 16165 4735
rect 16185 4715 16200 4735
rect 16150 4685 16200 4715
rect 16150 4665 16165 4685
rect 16185 4665 16200 4685
rect 16150 4635 16200 4665
rect 16150 4615 16165 4635
rect 16185 4615 16200 4635
rect 16150 4585 16200 4615
rect 16150 4565 16165 4585
rect 16185 4565 16200 4585
rect 16150 4535 16200 4565
rect 16150 4515 16165 4535
rect 16185 4515 16200 4535
rect 16150 4485 16200 4515
rect 16150 4465 16165 4485
rect 16185 4465 16200 4485
rect 16150 4435 16200 4465
rect 16150 4415 16165 4435
rect 16185 4415 16200 4435
rect 16150 4385 16200 4415
rect 16150 4365 16165 4385
rect 16185 4365 16200 4385
rect 16150 4350 16200 4365
rect 16300 4835 16350 4850
rect 16300 4815 16315 4835
rect 16335 4815 16350 4835
rect 16300 4785 16350 4815
rect 16300 4765 16315 4785
rect 16335 4765 16350 4785
rect 16300 4735 16350 4765
rect 16300 4715 16315 4735
rect 16335 4715 16350 4735
rect 16300 4685 16350 4715
rect 16300 4665 16315 4685
rect 16335 4665 16350 4685
rect 16300 4635 16350 4665
rect 16300 4615 16315 4635
rect 16335 4615 16350 4635
rect 16300 4585 16350 4615
rect 16300 4565 16315 4585
rect 16335 4565 16350 4585
rect 16300 4535 16350 4565
rect 16300 4515 16315 4535
rect 16335 4515 16350 4535
rect 16300 4485 16350 4515
rect 16300 4465 16315 4485
rect 16335 4465 16350 4485
rect 16300 4435 16350 4465
rect 16300 4415 16315 4435
rect 16335 4415 16350 4435
rect 16300 4385 16350 4415
rect 16300 4365 16315 4385
rect 16335 4365 16350 4385
rect 16300 4350 16350 4365
rect 16450 4835 16500 4850
rect 16450 4815 16465 4835
rect 16485 4815 16500 4835
rect 16450 4785 16500 4815
rect 16450 4765 16465 4785
rect 16485 4765 16500 4785
rect 16450 4735 16500 4765
rect 16450 4715 16465 4735
rect 16485 4715 16500 4735
rect 16450 4685 16500 4715
rect 16450 4665 16465 4685
rect 16485 4665 16500 4685
rect 16450 4635 16500 4665
rect 16450 4615 16465 4635
rect 16485 4615 16500 4635
rect 16450 4585 16500 4615
rect 16450 4565 16465 4585
rect 16485 4565 16500 4585
rect 16450 4535 16500 4565
rect 16450 4515 16465 4535
rect 16485 4515 16500 4535
rect 16450 4485 16500 4515
rect 16450 4465 16465 4485
rect 16485 4465 16500 4485
rect 16450 4435 16500 4465
rect 16450 4415 16465 4435
rect 16485 4415 16500 4435
rect 16450 4385 16500 4415
rect 16450 4365 16465 4385
rect 16485 4365 16500 4385
rect 16450 4350 16500 4365
rect 16600 4835 16650 4850
rect 16600 4815 16615 4835
rect 16635 4815 16650 4835
rect 16600 4785 16650 4815
rect 16600 4765 16615 4785
rect 16635 4765 16650 4785
rect 16600 4735 16650 4765
rect 16600 4715 16615 4735
rect 16635 4715 16650 4735
rect 16600 4685 16650 4715
rect 16600 4665 16615 4685
rect 16635 4665 16650 4685
rect 16600 4635 16650 4665
rect 16600 4615 16615 4635
rect 16635 4615 16650 4635
rect 16600 4585 16650 4615
rect 16600 4565 16615 4585
rect 16635 4565 16650 4585
rect 16600 4535 16650 4565
rect 16600 4515 16615 4535
rect 16635 4515 16650 4535
rect 16600 4485 16650 4515
rect 16600 4465 16615 4485
rect 16635 4465 16650 4485
rect 16600 4435 16650 4465
rect 16600 4415 16615 4435
rect 16635 4415 16650 4435
rect 16600 4385 16650 4415
rect 16600 4365 16615 4385
rect 16635 4365 16650 4385
rect 16600 4350 16650 4365
rect 16750 4835 16800 4850
rect 16750 4815 16765 4835
rect 16785 4815 16800 4835
rect 16750 4785 16800 4815
rect 16750 4765 16765 4785
rect 16785 4765 16800 4785
rect 16750 4735 16800 4765
rect 16750 4715 16765 4735
rect 16785 4715 16800 4735
rect 16750 4685 16800 4715
rect 16750 4665 16765 4685
rect 16785 4665 16800 4685
rect 16750 4635 16800 4665
rect 16750 4615 16765 4635
rect 16785 4615 16800 4635
rect 16750 4585 16800 4615
rect 16750 4565 16765 4585
rect 16785 4565 16800 4585
rect 16750 4535 16800 4565
rect 16750 4515 16765 4535
rect 16785 4515 16800 4535
rect 16750 4485 16800 4515
rect 16750 4465 16765 4485
rect 16785 4465 16800 4485
rect 16750 4435 16800 4465
rect 16750 4415 16765 4435
rect 16785 4415 16800 4435
rect 16750 4385 16800 4415
rect 16750 4365 16765 4385
rect 16785 4365 16800 4385
rect 16750 4350 16800 4365
rect 16900 4835 16950 4850
rect 16900 4815 16915 4835
rect 16935 4815 16950 4835
rect 16900 4785 16950 4815
rect 16900 4765 16915 4785
rect 16935 4765 16950 4785
rect 16900 4735 16950 4765
rect 16900 4715 16915 4735
rect 16935 4715 16950 4735
rect 16900 4685 16950 4715
rect 16900 4665 16915 4685
rect 16935 4665 16950 4685
rect 16900 4635 16950 4665
rect 16900 4615 16915 4635
rect 16935 4615 16950 4635
rect 16900 4585 16950 4615
rect 16900 4565 16915 4585
rect 16935 4565 16950 4585
rect 16900 4535 16950 4565
rect 16900 4515 16915 4535
rect 16935 4515 16950 4535
rect 16900 4485 16950 4515
rect 16900 4465 16915 4485
rect 16935 4465 16950 4485
rect 16900 4435 16950 4465
rect 16900 4415 16915 4435
rect 16935 4415 16950 4435
rect 16900 4385 16950 4415
rect 16900 4365 16915 4385
rect 16935 4365 16950 4385
rect 16900 4350 16950 4365
rect 17050 4835 17100 4850
rect 17050 4815 17065 4835
rect 17085 4815 17100 4835
rect 17050 4785 17100 4815
rect 17050 4765 17065 4785
rect 17085 4765 17100 4785
rect 17050 4735 17100 4765
rect 17050 4715 17065 4735
rect 17085 4715 17100 4735
rect 17050 4685 17100 4715
rect 17050 4665 17065 4685
rect 17085 4665 17100 4685
rect 17050 4635 17100 4665
rect 17050 4615 17065 4635
rect 17085 4615 17100 4635
rect 17050 4585 17100 4615
rect 17050 4565 17065 4585
rect 17085 4565 17100 4585
rect 17050 4535 17100 4565
rect 17050 4515 17065 4535
rect 17085 4515 17100 4535
rect 17050 4485 17100 4515
rect 17050 4465 17065 4485
rect 17085 4465 17100 4485
rect 17050 4435 17100 4465
rect 17050 4415 17065 4435
rect 17085 4415 17100 4435
rect 17050 4385 17100 4415
rect 17050 4365 17065 4385
rect 17085 4365 17100 4385
rect 17050 4350 17100 4365
rect 17200 4835 17250 4850
rect 17200 4815 17215 4835
rect 17235 4815 17250 4835
rect 17200 4785 17250 4815
rect 17200 4765 17215 4785
rect 17235 4765 17250 4785
rect 17200 4735 17250 4765
rect 17200 4715 17215 4735
rect 17235 4715 17250 4735
rect 17200 4685 17250 4715
rect 17200 4665 17215 4685
rect 17235 4665 17250 4685
rect 17200 4635 17250 4665
rect 17200 4615 17215 4635
rect 17235 4615 17250 4635
rect 17200 4585 17250 4615
rect 17200 4565 17215 4585
rect 17235 4565 17250 4585
rect 17200 4535 17250 4565
rect 17200 4515 17215 4535
rect 17235 4515 17250 4535
rect 17200 4485 17250 4515
rect 17200 4465 17215 4485
rect 17235 4465 17250 4485
rect 17200 4435 17250 4465
rect 17200 4415 17215 4435
rect 17235 4415 17250 4435
rect 17200 4385 17250 4415
rect 17200 4365 17215 4385
rect 17235 4365 17250 4385
rect 17200 4350 17250 4365
rect 17350 4835 17400 4850
rect 17350 4815 17365 4835
rect 17385 4815 17400 4835
rect 17350 4785 17400 4815
rect 17350 4765 17365 4785
rect 17385 4765 17400 4785
rect 17350 4735 17400 4765
rect 17350 4715 17365 4735
rect 17385 4715 17400 4735
rect 17350 4685 17400 4715
rect 17350 4665 17365 4685
rect 17385 4665 17400 4685
rect 17350 4635 17400 4665
rect 17350 4615 17365 4635
rect 17385 4615 17400 4635
rect 17350 4585 17400 4615
rect 17350 4565 17365 4585
rect 17385 4565 17400 4585
rect 17350 4535 17400 4565
rect 17350 4515 17365 4535
rect 17385 4515 17400 4535
rect 17350 4485 17400 4515
rect 17350 4465 17365 4485
rect 17385 4465 17400 4485
rect 17350 4435 17400 4465
rect 17350 4415 17365 4435
rect 17385 4415 17400 4435
rect 17350 4385 17400 4415
rect 17350 4365 17365 4385
rect 17385 4365 17400 4385
rect 17350 4350 17400 4365
rect 17950 4835 18000 4850
rect 17950 4815 17965 4835
rect 17985 4815 18000 4835
rect 17950 4785 18000 4815
rect 17950 4765 17965 4785
rect 17985 4765 18000 4785
rect 17950 4735 18000 4765
rect 17950 4715 17965 4735
rect 17985 4715 18000 4735
rect 17950 4685 18000 4715
rect 17950 4665 17965 4685
rect 17985 4665 18000 4685
rect 17950 4635 18000 4665
rect 17950 4615 17965 4635
rect 17985 4615 18000 4635
rect 17950 4585 18000 4615
rect 17950 4565 17965 4585
rect 17985 4565 18000 4585
rect 17950 4535 18000 4565
rect 17950 4515 17965 4535
rect 17985 4515 18000 4535
rect 17950 4485 18000 4515
rect 17950 4465 17965 4485
rect 17985 4465 18000 4485
rect 17950 4435 18000 4465
rect 17950 4415 17965 4435
rect 17985 4415 18000 4435
rect 17950 4385 18000 4415
rect 17950 4365 17965 4385
rect 17985 4365 18000 4385
rect 17950 4350 18000 4365
rect 18550 4835 18600 4850
rect 18550 4815 18565 4835
rect 18585 4815 18600 4835
rect 18550 4785 18600 4815
rect 18550 4765 18565 4785
rect 18585 4765 18600 4785
rect 18550 4735 18600 4765
rect 18550 4715 18565 4735
rect 18585 4715 18600 4735
rect 18550 4685 18600 4715
rect 18550 4665 18565 4685
rect 18585 4665 18600 4685
rect 18550 4635 18600 4665
rect 18550 4615 18565 4635
rect 18585 4615 18600 4635
rect 18550 4585 18600 4615
rect 18550 4565 18565 4585
rect 18585 4565 18600 4585
rect 18550 4535 18600 4565
rect 18550 4515 18565 4535
rect 18585 4515 18600 4535
rect 18550 4485 18600 4515
rect 18550 4465 18565 4485
rect 18585 4465 18600 4485
rect 18550 4435 18600 4465
rect 18550 4415 18565 4435
rect 18585 4415 18600 4435
rect 18550 4385 18600 4415
rect 18550 4365 18565 4385
rect 18585 4365 18600 4385
rect 18550 4350 18600 4365
rect 18700 4835 18750 4850
rect 18700 4815 18715 4835
rect 18735 4815 18750 4835
rect 18700 4785 18750 4815
rect 18700 4765 18715 4785
rect 18735 4765 18750 4785
rect 18700 4735 18750 4765
rect 18700 4715 18715 4735
rect 18735 4715 18750 4735
rect 18700 4685 18750 4715
rect 18700 4665 18715 4685
rect 18735 4665 18750 4685
rect 18700 4635 18750 4665
rect 18700 4615 18715 4635
rect 18735 4615 18750 4635
rect 18700 4585 18750 4615
rect 18700 4565 18715 4585
rect 18735 4565 18750 4585
rect 18700 4535 18750 4565
rect 18700 4515 18715 4535
rect 18735 4515 18750 4535
rect 18700 4485 18750 4515
rect 18700 4465 18715 4485
rect 18735 4465 18750 4485
rect 18700 4435 18750 4465
rect 18700 4415 18715 4435
rect 18735 4415 18750 4435
rect 18700 4385 18750 4415
rect 18700 4365 18715 4385
rect 18735 4365 18750 4385
rect 18700 4350 18750 4365
rect 18850 4835 18900 4850
rect 18850 4815 18865 4835
rect 18885 4815 18900 4835
rect 18850 4785 18900 4815
rect 18850 4765 18865 4785
rect 18885 4765 18900 4785
rect 18850 4735 18900 4765
rect 18850 4715 18865 4735
rect 18885 4715 18900 4735
rect 18850 4685 18900 4715
rect 18850 4665 18865 4685
rect 18885 4665 18900 4685
rect 18850 4635 18900 4665
rect 18850 4615 18865 4635
rect 18885 4615 18900 4635
rect 18850 4585 18900 4615
rect 18850 4565 18865 4585
rect 18885 4565 18900 4585
rect 18850 4535 18900 4565
rect 18850 4515 18865 4535
rect 18885 4515 18900 4535
rect 18850 4485 18900 4515
rect 18850 4465 18865 4485
rect 18885 4465 18900 4485
rect 18850 4435 18900 4465
rect 18850 4415 18865 4435
rect 18885 4415 18900 4435
rect 18850 4385 18900 4415
rect 18850 4365 18865 4385
rect 18885 4365 18900 4385
rect 18850 4350 18900 4365
rect 19000 4835 19050 4850
rect 19000 4815 19015 4835
rect 19035 4815 19050 4835
rect 19000 4785 19050 4815
rect 19000 4765 19015 4785
rect 19035 4765 19050 4785
rect 19000 4735 19050 4765
rect 19000 4715 19015 4735
rect 19035 4715 19050 4735
rect 19000 4685 19050 4715
rect 19000 4665 19015 4685
rect 19035 4665 19050 4685
rect 19000 4635 19050 4665
rect 19000 4615 19015 4635
rect 19035 4615 19050 4635
rect 19000 4585 19050 4615
rect 19000 4565 19015 4585
rect 19035 4565 19050 4585
rect 19000 4535 19050 4565
rect 19000 4515 19015 4535
rect 19035 4515 19050 4535
rect 19000 4485 19050 4515
rect 19000 4465 19015 4485
rect 19035 4465 19050 4485
rect 19000 4435 19050 4465
rect 19000 4415 19015 4435
rect 19035 4415 19050 4435
rect 19000 4385 19050 4415
rect 19000 4365 19015 4385
rect 19035 4365 19050 4385
rect 19000 4350 19050 4365
rect 19150 4835 19200 4850
rect 19150 4815 19165 4835
rect 19185 4815 19200 4835
rect 19150 4785 19200 4815
rect 19150 4765 19165 4785
rect 19185 4765 19200 4785
rect 19150 4735 19200 4765
rect 19150 4715 19165 4735
rect 19185 4715 19200 4735
rect 19150 4685 19200 4715
rect 19150 4665 19165 4685
rect 19185 4665 19200 4685
rect 19150 4635 19200 4665
rect 19150 4615 19165 4635
rect 19185 4615 19200 4635
rect 19150 4585 19200 4615
rect 19150 4565 19165 4585
rect 19185 4565 19200 4585
rect 19150 4535 19200 4565
rect 19150 4515 19165 4535
rect 19185 4515 19200 4535
rect 19150 4485 19200 4515
rect 19150 4465 19165 4485
rect 19185 4465 19200 4485
rect 19150 4435 19200 4465
rect 19150 4415 19165 4435
rect 19185 4415 19200 4435
rect 19150 4385 19200 4415
rect 19150 4365 19165 4385
rect 19185 4365 19200 4385
rect 19150 4350 19200 4365
rect 19300 4835 19350 4850
rect 19300 4815 19315 4835
rect 19335 4815 19350 4835
rect 19300 4785 19350 4815
rect 19300 4765 19315 4785
rect 19335 4765 19350 4785
rect 19300 4735 19350 4765
rect 19300 4715 19315 4735
rect 19335 4715 19350 4735
rect 19300 4685 19350 4715
rect 19300 4665 19315 4685
rect 19335 4665 19350 4685
rect 19300 4635 19350 4665
rect 19300 4615 19315 4635
rect 19335 4615 19350 4635
rect 19300 4585 19350 4615
rect 19300 4565 19315 4585
rect 19335 4565 19350 4585
rect 19300 4535 19350 4565
rect 19300 4515 19315 4535
rect 19335 4515 19350 4535
rect 19300 4485 19350 4515
rect 19300 4465 19315 4485
rect 19335 4465 19350 4485
rect 19300 4435 19350 4465
rect 19300 4415 19315 4435
rect 19335 4415 19350 4435
rect 19300 4385 19350 4415
rect 19300 4365 19315 4385
rect 19335 4365 19350 4385
rect 19300 4350 19350 4365
rect 19450 4835 19500 4850
rect 19450 4815 19465 4835
rect 19485 4815 19500 4835
rect 19450 4785 19500 4815
rect 19450 4765 19465 4785
rect 19485 4765 19500 4785
rect 19450 4735 19500 4765
rect 19450 4715 19465 4735
rect 19485 4715 19500 4735
rect 19450 4685 19500 4715
rect 19450 4665 19465 4685
rect 19485 4665 19500 4685
rect 19450 4635 19500 4665
rect 19450 4615 19465 4635
rect 19485 4615 19500 4635
rect 19450 4585 19500 4615
rect 19450 4565 19465 4585
rect 19485 4565 19500 4585
rect 19450 4535 19500 4565
rect 19450 4515 19465 4535
rect 19485 4515 19500 4535
rect 19450 4485 19500 4515
rect 19450 4465 19465 4485
rect 19485 4465 19500 4485
rect 19450 4435 19500 4465
rect 19450 4415 19465 4435
rect 19485 4415 19500 4435
rect 19450 4385 19500 4415
rect 19450 4365 19465 4385
rect 19485 4365 19500 4385
rect 19450 4350 19500 4365
rect 19600 4835 19650 4850
rect 19600 4815 19615 4835
rect 19635 4815 19650 4835
rect 19600 4785 19650 4815
rect 19600 4765 19615 4785
rect 19635 4765 19650 4785
rect 19600 4735 19650 4765
rect 19600 4715 19615 4735
rect 19635 4715 19650 4735
rect 19600 4685 19650 4715
rect 19600 4665 19615 4685
rect 19635 4665 19650 4685
rect 19600 4635 19650 4665
rect 19600 4615 19615 4635
rect 19635 4615 19650 4635
rect 19600 4585 19650 4615
rect 19600 4565 19615 4585
rect 19635 4565 19650 4585
rect 19600 4535 19650 4565
rect 19600 4515 19615 4535
rect 19635 4515 19650 4535
rect 19600 4485 19650 4515
rect 19600 4465 19615 4485
rect 19635 4465 19650 4485
rect 19600 4435 19650 4465
rect 19600 4415 19615 4435
rect 19635 4415 19650 4435
rect 19600 4385 19650 4415
rect 19600 4365 19615 4385
rect 19635 4365 19650 4385
rect 19600 4350 19650 4365
rect 19750 4835 19800 4850
rect 19750 4815 19765 4835
rect 19785 4815 19800 4835
rect 19750 4785 19800 4815
rect 19750 4765 19765 4785
rect 19785 4765 19800 4785
rect 19750 4735 19800 4765
rect 19750 4715 19765 4735
rect 19785 4715 19800 4735
rect 19750 4685 19800 4715
rect 19750 4665 19765 4685
rect 19785 4665 19800 4685
rect 19750 4635 19800 4665
rect 19750 4615 19765 4635
rect 19785 4615 19800 4635
rect 19750 4585 19800 4615
rect 19750 4565 19765 4585
rect 19785 4565 19800 4585
rect 19750 4535 19800 4565
rect 19750 4515 19765 4535
rect 19785 4515 19800 4535
rect 19750 4485 19800 4515
rect 19750 4465 19765 4485
rect 19785 4465 19800 4485
rect 19750 4435 19800 4465
rect 19750 4415 19765 4435
rect 19785 4415 19800 4435
rect 19750 4385 19800 4415
rect 19750 4365 19765 4385
rect 19785 4365 19800 4385
rect 19750 4350 19800 4365
rect 20350 4835 20400 4850
rect 20350 4815 20365 4835
rect 20385 4815 20400 4835
rect 20350 4785 20400 4815
rect 20350 4765 20365 4785
rect 20385 4765 20400 4785
rect 20350 4735 20400 4765
rect 20350 4715 20365 4735
rect 20385 4715 20400 4735
rect 20350 4685 20400 4715
rect 20350 4665 20365 4685
rect 20385 4665 20400 4685
rect 20350 4635 20400 4665
rect 20350 4615 20365 4635
rect 20385 4615 20400 4635
rect 20350 4585 20400 4615
rect 20350 4565 20365 4585
rect 20385 4565 20400 4585
rect 20350 4535 20400 4565
rect 20350 4515 20365 4535
rect 20385 4515 20400 4535
rect 20350 4485 20400 4515
rect 20350 4465 20365 4485
rect 20385 4465 20400 4485
rect 20350 4435 20400 4465
rect 20350 4415 20365 4435
rect 20385 4415 20400 4435
rect 20350 4385 20400 4415
rect 20350 4365 20365 4385
rect 20385 4365 20400 4385
rect 20350 4350 20400 4365
rect 20950 4835 21000 4850
rect 20950 4815 20965 4835
rect 20985 4815 21000 4835
rect 20950 4785 21000 4815
rect 20950 4765 20965 4785
rect 20985 4765 21000 4785
rect 20950 4735 21000 4765
rect 20950 4715 20965 4735
rect 20985 4715 21000 4735
rect 20950 4685 21000 4715
rect 20950 4665 20965 4685
rect 20985 4665 21000 4685
rect 20950 4635 21000 4665
rect 20950 4615 20965 4635
rect 20985 4615 21000 4635
rect 20950 4585 21000 4615
rect 20950 4565 20965 4585
rect 20985 4565 21000 4585
rect 20950 4535 21000 4565
rect 20950 4515 20965 4535
rect 20985 4515 21000 4535
rect 20950 4485 21000 4515
rect 20950 4465 20965 4485
rect 20985 4465 21000 4485
rect 20950 4435 21000 4465
rect 20950 4415 20965 4435
rect 20985 4415 21000 4435
rect 20950 4385 21000 4415
rect 20950 4365 20965 4385
rect 20985 4365 21000 4385
rect 20950 4350 21000 4365
rect 21400 4835 21450 4850
rect 21400 4815 21415 4835
rect 21435 4815 21450 4835
rect 21400 4785 21450 4815
rect 21400 4765 21415 4785
rect 21435 4765 21450 4785
rect 21400 4735 21450 4765
rect 21400 4715 21415 4735
rect 21435 4715 21450 4735
rect 21400 4685 21450 4715
rect 21400 4665 21415 4685
rect 21435 4665 21450 4685
rect 21400 4635 21450 4665
rect 21400 4615 21415 4635
rect 21435 4615 21450 4635
rect 21400 4585 21450 4615
rect 21400 4565 21415 4585
rect 21435 4565 21450 4585
rect 21400 4535 21450 4565
rect 21400 4515 21415 4535
rect 21435 4515 21450 4535
rect 21400 4485 21450 4515
rect 21400 4465 21415 4485
rect 21435 4465 21450 4485
rect 21400 4435 21450 4465
rect 21400 4415 21415 4435
rect 21435 4415 21450 4435
rect 21400 4385 21450 4415
rect 21400 4365 21415 4385
rect 21435 4365 21450 4385
rect 21400 4350 21450 4365
rect 21850 4835 21900 4850
rect 21850 4815 21865 4835
rect 21885 4815 21900 4835
rect 21850 4785 21900 4815
rect 21850 4765 21865 4785
rect 21885 4765 21900 4785
rect 21850 4735 21900 4765
rect 21850 4715 21865 4735
rect 21885 4715 21900 4735
rect 21850 4685 21900 4715
rect 21850 4665 21865 4685
rect 21885 4665 21900 4685
rect 21850 4635 21900 4665
rect 21850 4615 21865 4635
rect 21885 4615 21900 4635
rect 21850 4585 21900 4615
rect 21850 4565 21865 4585
rect 21885 4565 21900 4585
rect 21850 4535 21900 4565
rect 21850 4515 21865 4535
rect 21885 4515 21900 4535
rect 21850 4485 21900 4515
rect 21850 4465 21865 4485
rect 21885 4465 21900 4485
rect 21850 4435 21900 4465
rect 21850 4415 21865 4435
rect 21885 4415 21900 4435
rect 21850 4385 21900 4415
rect 21850 4365 21865 4385
rect 21885 4365 21900 4385
rect 21850 4350 21900 4365
rect 22450 4835 22500 4850
rect 22450 4815 22465 4835
rect 22485 4815 22500 4835
rect 22450 4785 22500 4815
rect 22450 4765 22465 4785
rect 22485 4765 22500 4785
rect 22450 4735 22500 4765
rect 22450 4715 22465 4735
rect 22485 4715 22500 4735
rect 22450 4685 22500 4715
rect 22450 4665 22465 4685
rect 22485 4665 22500 4685
rect 22450 4635 22500 4665
rect 22450 4615 22465 4635
rect 22485 4615 22500 4635
rect 22450 4585 22500 4615
rect 22450 4565 22465 4585
rect 22485 4565 22500 4585
rect 22450 4535 22500 4565
rect 22450 4515 22465 4535
rect 22485 4515 22500 4535
rect 22450 4485 22500 4515
rect 22450 4465 22465 4485
rect 22485 4465 22500 4485
rect 22450 4435 22500 4465
rect 22450 4415 22465 4435
rect 22485 4415 22500 4435
rect 22450 4385 22500 4415
rect 22450 4365 22465 4385
rect 22485 4365 22500 4385
rect 22450 4350 22500 4365
rect 23050 4835 23100 4850
rect 23050 4815 23065 4835
rect 23085 4815 23100 4835
rect 23050 4785 23100 4815
rect 23050 4765 23065 4785
rect 23085 4765 23100 4785
rect 23050 4735 23100 4765
rect 23050 4715 23065 4735
rect 23085 4715 23100 4735
rect 23050 4685 23100 4715
rect 23050 4665 23065 4685
rect 23085 4665 23100 4685
rect 23050 4635 23100 4665
rect 23050 4615 23065 4635
rect 23085 4615 23100 4635
rect 23050 4585 23100 4615
rect 23050 4565 23065 4585
rect 23085 4565 23100 4585
rect 23050 4535 23100 4565
rect 23050 4515 23065 4535
rect 23085 4515 23100 4535
rect 23050 4485 23100 4515
rect 23050 4465 23065 4485
rect 23085 4465 23100 4485
rect 23050 4435 23100 4465
rect 23050 4415 23065 4435
rect 23085 4415 23100 4435
rect 23050 4385 23100 4415
rect 23050 4365 23065 4385
rect 23085 4365 23100 4385
rect 23050 4350 23100 4365
rect 23500 4835 23550 4850
rect 23500 4815 23515 4835
rect 23535 4815 23550 4835
rect 23500 4785 23550 4815
rect 23500 4765 23515 4785
rect 23535 4765 23550 4785
rect 23500 4735 23550 4765
rect 23500 4715 23515 4735
rect 23535 4715 23550 4735
rect 23500 4685 23550 4715
rect 23500 4665 23515 4685
rect 23535 4665 23550 4685
rect 23500 4635 23550 4665
rect 23500 4615 23515 4635
rect 23535 4615 23550 4635
rect 23500 4585 23550 4615
rect 23500 4565 23515 4585
rect 23535 4565 23550 4585
rect 23500 4535 23550 4565
rect 23500 4515 23515 4535
rect 23535 4515 23550 4535
rect 23500 4485 23550 4515
rect 23500 4465 23515 4485
rect 23535 4465 23550 4485
rect 23500 4435 23550 4465
rect 23500 4415 23515 4435
rect 23535 4415 23550 4435
rect 23500 4385 23550 4415
rect 23500 4365 23515 4385
rect 23535 4365 23550 4385
rect 23500 4350 23550 4365
rect 23950 4835 24000 4850
rect 23950 4815 23965 4835
rect 23985 4815 24000 4835
rect 23950 4785 24000 4815
rect 23950 4765 23965 4785
rect 23985 4765 24000 4785
rect 23950 4735 24000 4765
rect 23950 4715 23965 4735
rect 23985 4715 24000 4735
rect 23950 4685 24000 4715
rect 23950 4665 23965 4685
rect 23985 4665 24000 4685
rect 23950 4635 24000 4665
rect 23950 4615 23965 4635
rect 23985 4615 24000 4635
rect 23950 4585 24000 4615
rect 23950 4565 23965 4585
rect 23985 4565 24000 4585
rect 23950 4535 24000 4565
rect 23950 4515 23965 4535
rect 23985 4515 24000 4535
rect 23950 4485 24000 4515
rect 23950 4465 23965 4485
rect 23985 4465 24000 4485
rect 23950 4435 24000 4465
rect 23950 4415 23965 4435
rect 23985 4415 24000 4435
rect 23950 4385 24000 4415
rect 23950 4365 23965 4385
rect 23985 4365 24000 4385
rect 23950 4350 24000 4365
rect 24550 4835 24600 4850
rect 24550 4815 24565 4835
rect 24585 4815 24600 4835
rect 24550 4785 24600 4815
rect 24550 4765 24565 4785
rect 24585 4765 24600 4785
rect 24550 4735 24600 4765
rect 24550 4715 24565 4735
rect 24585 4715 24600 4735
rect 24550 4685 24600 4715
rect 24550 4665 24565 4685
rect 24585 4665 24600 4685
rect 24550 4635 24600 4665
rect 24550 4615 24565 4635
rect 24585 4615 24600 4635
rect 24550 4585 24600 4615
rect 24550 4565 24565 4585
rect 24585 4565 24600 4585
rect 24550 4535 24600 4565
rect 24550 4515 24565 4535
rect 24585 4515 24600 4535
rect 24550 4485 24600 4515
rect 24550 4465 24565 4485
rect 24585 4465 24600 4485
rect 24550 4435 24600 4465
rect 24550 4415 24565 4435
rect 24585 4415 24600 4435
rect 24550 4385 24600 4415
rect 24550 4365 24565 4385
rect 24585 4365 24600 4385
rect 24550 4350 24600 4365
rect 25150 4835 25200 4850
rect 25150 4815 25165 4835
rect 25185 4815 25200 4835
rect 25150 4785 25200 4815
rect 25150 4765 25165 4785
rect 25185 4765 25200 4785
rect 25150 4735 25200 4765
rect 25150 4715 25165 4735
rect 25185 4715 25200 4735
rect 25150 4685 25200 4715
rect 25150 4665 25165 4685
rect 25185 4665 25200 4685
rect 25150 4635 25200 4665
rect 25150 4615 25165 4635
rect 25185 4615 25200 4635
rect 25150 4585 25200 4615
rect 25150 4565 25165 4585
rect 25185 4565 25200 4585
rect 25150 4535 25200 4565
rect 25150 4515 25165 4535
rect 25185 4515 25200 4535
rect 25150 4485 25200 4515
rect 25150 4465 25165 4485
rect 25185 4465 25200 4485
rect 25150 4435 25200 4465
rect 25150 4415 25165 4435
rect 25185 4415 25200 4435
rect 25150 4385 25200 4415
rect 25150 4365 25165 4385
rect 25185 4365 25200 4385
rect 25150 4350 25200 4365
rect 25600 4835 25650 4850
rect 25600 4815 25615 4835
rect 25635 4815 25650 4835
rect 25600 4785 25650 4815
rect 25600 4765 25615 4785
rect 25635 4765 25650 4785
rect 25600 4735 25650 4765
rect 25600 4715 25615 4735
rect 25635 4715 25650 4735
rect 25600 4685 25650 4715
rect 25600 4665 25615 4685
rect 25635 4665 25650 4685
rect 25600 4635 25650 4665
rect 25600 4615 25615 4635
rect 25635 4615 25650 4635
rect 25600 4585 25650 4615
rect 25600 4565 25615 4585
rect 25635 4565 25650 4585
rect 25600 4535 25650 4565
rect 25600 4515 25615 4535
rect 25635 4515 25650 4535
rect 25600 4485 25650 4515
rect 25600 4465 25615 4485
rect 25635 4465 25650 4485
rect 25600 4435 25650 4465
rect 25600 4415 25615 4435
rect 25635 4415 25650 4435
rect 25600 4385 25650 4415
rect 25600 4365 25615 4385
rect 25635 4365 25650 4385
rect 25600 4350 25650 4365
rect 26050 4835 26100 4850
rect 26050 4815 26065 4835
rect 26085 4815 26100 4835
rect 26050 4785 26100 4815
rect 26050 4765 26065 4785
rect 26085 4765 26100 4785
rect 26050 4735 26100 4765
rect 26050 4715 26065 4735
rect 26085 4715 26100 4735
rect 26050 4685 26100 4715
rect 26050 4665 26065 4685
rect 26085 4665 26100 4685
rect 26050 4635 26100 4665
rect 26050 4615 26065 4635
rect 26085 4615 26100 4635
rect 26050 4585 26100 4615
rect 26050 4565 26065 4585
rect 26085 4565 26100 4585
rect 26050 4535 26100 4565
rect 26050 4515 26065 4535
rect 26085 4515 26100 4535
rect 26050 4485 26100 4515
rect 26050 4465 26065 4485
rect 26085 4465 26100 4485
rect 26050 4435 26100 4465
rect 26050 4415 26065 4435
rect 26085 4415 26100 4435
rect 26050 4385 26100 4415
rect 26050 4365 26065 4385
rect 26085 4365 26100 4385
rect 26050 4350 26100 4365
rect 26650 4835 26700 4850
rect 26650 4815 26665 4835
rect 26685 4815 26700 4835
rect 26650 4785 26700 4815
rect 26650 4765 26665 4785
rect 26685 4765 26700 4785
rect 26650 4735 26700 4765
rect 26650 4715 26665 4735
rect 26685 4715 26700 4735
rect 26650 4685 26700 4715
rect 26650 4665 26665 4685
rect 26685 4665 26700 4685
rect 26650 4635 26700 4665
rect 26650 4615 26665 4635
rect 26685 4615 26700 4635
rect 26650 4585 26700 4615
rect 26650 4565 26665 4585
rect 26685 4565 26700 4585
rect 26650 4535 26700 4565
rect 26650 4515 26665 4535
rect 26685 4515 26700 4535
rect 26650 4485 26700 4515
rect 26650 4465 26665 4485
rect 26685 4465 26700 4485
rect 26650 4435 26700 4465
rect 26650 4415 26665 4435
rect 26685 4415 26700 4435
rect 26650 4385 26700 4415
rect 26650 4365 26665 4385
rect 26685 4365 26700 4385
rect 26650 4350 26700 4365
rect 27250 4835 27300 4850
rect 27250 4815 27265 4835
rect 27285 4815 27300 4835
rect 27250 4785 27300 4815
rect 27250 4765 27265 4785
rect 27285 4765 27300 4785
rect 27250 4735 27300 4765
rect 27250 4715 27265 4735
rect 27285 4715 27300 4735
rect 27250 4685 27300 4715
rect 27250 4665 27265 4685
rect 27285 4665 27300 4685
rect 27250 4635 27300 4665
rect 27250 4615 27265 4635
rect 27285 4615 27300 4635
rect 27250 4585 27300 4615
rect 27250 4565 27265 4585
rect 27285 4565 27300 4585
rect 27250 4535 27300 4565
rect 27250 4515 27265 4535
rect 27285 4515 27300 4535
rect 27250 4485 27300 4515
rect 27250 4465 27265 4485
rect 27285 4465 27300 4485
rect 27250 4435 27300 4465
rect 27250 4415 27265 4435
rect 27285 4415 27300 4435
rect 27250 4385 27300 4415
rect 27250 4365 27265 4385
rect 27285 4365 27300 4385
rect 27250 4350 27300 4365
rect 27700 4835 27750 4850
rect 27700 4815 27715 4835
rect 27735 4815 27750 4835
rect 27700 4785 27750 4815
rect 27700 4765 27715 4785
rect 27735 4765 27750 4785
rect 27700 4735 27750 4765
rect 27700 4715 27715 4735
rect 27735 4715 27750 4735
rect 27700 4685 27750 4715
rect 27700 4665 27715 4685
rect 27735 4665 27750 4685
rect 27700 4635 27750 4665
rect 27700 4615 27715 4635
rect 27735 4615 27750 4635
rect 27700 4585 27750 4615
rect 27700 4565 27715 4585
rect 27735 4565 27750 4585
rect 27700 4535 27750 4565
rect 27700 4515 27715 4535
rect 27735 4515 27750 4535
rect 27700 4485 27750 4515
rect 27700 4465 27715 4485
rect 27735 4465 27750 4485
rect 27700 4435 27750 4465
rect 27700 4415 27715 4435
rect 27735 4415 27750 4435
rect 27700 4385 27750 4415
rect 27700 4365 27715 4385
rect 27735 4365 27750 4385
rect 27700 4350 27750 4365
rect 28150 4835 28200 4850
rect 28150 4815 28165 4835
rect 28185 4815 28200 4835
rect 28150 4785 28200 4815
rect 28150 4765 28165 4785
rect 28185 4765 28200 4785
rect 28150 4735 28200 4765
rect 28150 4715 28165 4735
rect 28185 4715 28200 4735
rect 28150 4685 28200 4715
rect 28150 4665 28165 4685
rect 28185 4665 28200 4685
rect 28150 4635 28200 4665
rect 28150 4615 28165 4635
rect 28185 4615 28200 4635
rect 28150 4585 28200 4615
rect 28150 4565 28165 4585
rect 28185 4565 28200 4585
rect 28150 4535 28200 4565
rect 28150 4515 28165 4535
rect 28185 4515 28200 4535
rect 28150 4485 28200 4515
rect 28150 4465 28165 4485
rect 28185 4465 28200 4485
rect 28150 4435 28200 4465
rect 28150 4415 28165 4435
rect 28185 4415 28200 4435
rect 28150 4385 28200 4415
rect 28150 4365 28165 4385
rect 28185 4365 28200 4385
rect 28150 4350 28200 4365
rect 28750 4835 28800 4850
rect 28750 4815 28765 4835
rect 28785 4815 28800 4835
rect 28750 4785 28800 4815
rect 28750 4765 28765 4785
rect 28785 4765 28800 4785
rect 28750 4735 28800 4765
rect 28750 4715 28765 4735
rect 28785 4715 28800 4735
rect 28750 4685 28800 4715
rect 28750 4665 28765 4685
rect 28785 4665 28800 4685
rect 28750 4635 28800 4665
rect 28750 4615 28765 4635
rect 28785 4615 28800 4635
rect 28750 4585 28800 4615
rect 28750 4565 28765 4585
rect 28785 4565 28800 4585
rect 28750 4535 28800 4565
rect 28750 4515 28765 4535
rect 28785 4515 28800 4535
rect 28750 4485 28800 4515
rect 28750 4465 28765 4485
rect 28785 4465 28800 4485
rect 28750 4435 28800 4465
rect 28750 4415 28765 4435
rect 28785 4415 28800 4435
rect 28750 4385 28800 4415
rect 28750 4365 28765 4385
rect 28785 4365 28800 4385
rect 28750 4350 28800 4365
rect 29350 4835 29400 4850
rect 29350 4815 29365 4835
rect 29385 4815 29400 4835
rect 29350 4785 29400 4815
rect 29350 4765 29365 4785
rect 29385 4765 29400 4785
rect 29350 4735 29400 4765
rect 29350 4715 29365 4735
rect 29385 4715 29400 4735
rect 29350 4685 29400 4715
rect 29350 4665 29365 4685
rect 29385 4665 29400 4685
rect 29350 4635 29400 4665
rect 29350 4615 29365 4635
rect 29385 4615 29400 4635
rect 29350 4585 29400 4615
rect 29350 4565 29365 4585
rect 29385 4565 29400 4585
rect 29350 4535 29400 4565
rect 29350 4515 29365 4535
rect 29385 4515 29400 4535
rect 29350 4485 29400 4515
rect 29350 4465 29365 4485
rect 29385 4465 29400 4485
rect 29350 4435 29400 4465
rect 29350 4415 29365 4435
rect 29385 4415 29400 4435
rect 29350 4385 29400 4415
rect 29350 4365 29365 4385
rect 29385 4365 29400 4385
rect 29350 4350 29400 4365
rect 29500 4835 29550 4850
rect 29500 4815 29515 4835
rect 29535 4815 29550 4835
rect 29500 4785 29550 4815
rect 29500 4765 29515 4785
rect 29535 4765 29550 4785
rect 29500 4735 29550 4765
rect 29500 4715 29515 4735
rect 29535 4715 29550 4735
rect 29500 4685 29550 4715
rect 29500 4665 29515 4685
rect 29535 4665 29550 4685
rect 29500 4635 29550 4665
rect 29500 4615 29515 4635
rect 29535 4615 29550 4635
rect 29500 4585 29550 4615
rect 29500 4565 29515 4585
rect 29535 4565 29550 4585
rect 29500 4535 29550 4565
rect 29500 4515 29515 4535
rect 29535 4515 29550 4535
rect 29500 4485 29550 4515
rect 29500 4465 29515 4485
rect 29535 4465 29550 4485
rect 29500 4435 29550 4465
rect 29500 4415 29515 4435
rect 29535 4415 29550 4435
rect 29500 4385 29550 4415
rect 29500 4365 29515 4385
rect 29535 4365 29550 4385
rect 29500 4350 29550 4365
rect 29650 4835 29700 4850
rect 29650 4815 29665 4835
rect 29685 4815 29700 4835
rect 29650 4785 29700 4815
rect 29650 4765 29665 4785
rect 29685 4765 29700 4785
rect 29650 4735 29700 4765
rect 29650 4715 29665 4735
rect 29685 4715 29700 4735
rect 29650 4685 29700 4715
rect 29650 4665 29665 4685
rect 29685 4665 29700 4685
rect 29650 4635 29700 4665
rect 29650 4615 29665 4635
rect 29685 4615 29700 4635
rect 29650 4585 29700 4615
rect 29650 4565 29665 4585
rect 29685 4565 29700 4585
rect 29650 4535 29700 4565
rect 29650 4515 29665 4535
rect 29685 4515 29700 4535
rect 29650 4485 29700 4515
rect 29650 4465 29665 4485
rect 29685 4465 29700 4485
rect 29650 4435 29700 4465
rect 29650 4415 29665 4435
rect 29685 4415 29700 4435
rect 29650 4385 29700 4415
rect 29650 4365 29665 4385
rect 29685 4365 29700 4385
rect 29650 4350 29700 4365
rect 29800 4835 29850 4850
rect 29800 4815 29815 4835
rect 29835 4815 29850 4835
rect 29800 4785 29850 4815
rect 29800 4765 29815 4785
rect 29835 4765 29850 4785
rect 29800 4735 29850 4765
rect 29800 4715 29815 4735
rect 29835 4715 29850 4735
rect 29800 4685 29850 4715
rect 29800 4665 29815 4685
rect 29835 4665 29850 4685
rect 29800 4635 29850 4665
rect 29800 4615 29815 4635
rect 29835 4615 29850 4635
rect 29800 4585 29850 4615
rect 29800 4565 29815 4585
rect 29835 4565 29850 4585
rect 29800 4535 29850 4565
rect 29800 4515 29815 4535
rect 29835 4515 29850 4535
rect 29800 4485 29850 4515
rect 29800 4465 29815 4485
rect 29835 4465 29850 4485
rect 29800 4435 29850 4465
rect 29800 4415 29815 4435
rect 29835 4415 29850 4435
rect 29800 4385 29850 4415
rect 29800 4365 29815 4385
rect 29835 4365 29850 4385
rect 29800 4350 29850 4365
rect 29950 4835 30000 4850
rect 29950 4815 29965 4835
rect 29985 4815 30000 4835
rect 29950 4785 30000 4815
rect 29950 4765 29965 4785
rect 29985 4765 30000 4785
rect 29950 4735 30000 4765
rect 29950 4715 29965 4735
rect 29985 4715 30000 4735
rect 29950 4685 30000 4715
rect 29950 4665 29965 4685
rect 29985 4665 30000 4685
rect 29950 4635 30000 4665
rect 29950 4615 29965 4635
rect 29985 4615 30000 4635
rect 29950 4585 30000 4615
rect 29950 4565 29965 4585
rect 29985 4565 30000 4585
rect 29950 4535 30000 4565
rect 29950 4515 29965 4535
rect 29985 4515 30000 4535
rect 29950 4485 30000 4515
rect 29950 4465 29965 4485
rect 29985 4465 30000 4485
rect 29950 4435 30000 4465
rect 29950 4415 29965 4435
rect 29985 4415 30000 4435
rect 29950 4385 30000 4415
rect 29950 4365 29965 4385
rect 29985 4365 30000 4385
rect 29950 4350 30000 4365
rect 30100 4835 30150 4850
rect 30100 4815 30115 4835
rect 30135 4815 30150 4835
rect 30100 4785 30150 4815
rect 30100 4765 30115 4785
rect 30135 4765 30150 4785
rect 30100 4735 30150 4765
rect 30100 4715 30115 4735
rect 30135 4715 30150 4735
rect 30100 4685 30150 4715
rect 30100 4665 30115 4685
rect 30135 4665 30150 4685
rect 30100 4635 30150 4665
rect 30100 4615 30115 4635
rect 30135 4615 30150 4635
rect 30100 4585 30150 4615
rect 30100 4565 30115 4585
rect 30135 4565 30150 4585
rect 30100 4535 30150 4565
rect 30100 4515 30115 4535
rect 30135 4515 30150 4535
rect 30100 4485 30150 4515
rect 30100 4465 30115 4485
rect 30135 4465 30150 4485
rect 30100 4435 30150 4465
rect 30100 4415 30115 4435
rect 30135 4415 30150 4435
rect 30100 4385 30150 4415
rect 30100 4365 30115 4385
rect 30135 4365 30150 4385
rect 30100 4350 30150 4365
rect 30250 4835 30300 4850
rect 30250 4815 30265 4835
rect 30285 4815 30300 4835
rect 30250 4785 30300 4815
rect 30250 4765 30265 4785
rect 30285 4765 30300 4785
rect 30250 4735 30300 4765
rect 30250 4715 30265 4735
rect 30285 4715 30300 4735
rect 30250 4685 30300 4715
rect 30250 4665 30265 4685
rect 30285 4665 30300 4685
rect 30250 4635 30300 4665
rect 30250 4615 30265 4635
rect 30285 4615 30300 4635
rect 30250 4585 30300 4615
rect 30250 4565 30265 4585
rect 30285 4565 30300 4585
rect 30250 4535 30300 4565
rect 30250 4515 30265 4535
rect 30285 4515 30300 4535
rect 30250 4485 30300 4515
rect 30250 4465 30265 4485
rect 30285 4465 30300 4485
rect 30250 4435 30300 4465
rect 30250 4415 30265 4435
rect 30285 4415 30300 4435
rect 30250 4385 30300 4415
rect 30250 4365 30265 4385
rect 30285 4365 30300 4385
rect 30250 4350 30300 4365
rect 30400 4835 30450 4850
rect 30400 4815 30415 4835
rect 30435 4815 30450 4835
rect 30400 4785 30450 4815
rect 30400 4765 30415 4785
rect 30435 4765 30450 4785
rect 30400 4735 30450 4765
rect 30400 4715 30415 4735
rect 30435 4715 30450 4735
rect 30400 4685 30450 4715
rect 30400 4665 30415 4685
rect 30435 4665 30450 4685
rect 30400 4635 30450 4665
rect 30400 4615 30415 4635
rect 30435 4615 30450 4635
rect 30400 4585 30450 4615
rect 30400 4565 30415 4585
rect 30435 4565 30450 4585
rect 30400 4535 30450 4565
rect 30400 4515 30415 4535
rect 30435 4515 30450 4535
rect 30400 4485 30450 4515
rect 30400 4465 30415 4485
rect 30435 4465 30450 4485
rect 30400 4435 30450 4465
rect 30400 4415 30415 4435
rect 30435 4415 30450 4435
rect 30400 4385 30450 4415
rect 30400 4365 30415 4385
rect 30435 4365 30450 4385
rect 30400 4350 30450 4365
rect 30550 4835 30600 4850
rect 30550 4815 30565 4835
rect 30585 4815 30600 4835
rect 30550 4785 30600 4815
rect 30550 4765 30565 4785
rect 30585 4765 30600 4785
rect 30550 4735 30600 4765
rect 30550 4715 30565 4735
rect 30585 4715 30600 4735
rect 30550 4685 30600 4715
rect 30550 4665 30565 4685
rect 30585 4665 30600 4685
rect 30550 4635 30600 4665
rect 30550 4615 30565 4635
rect 30585 4615 30600 4635
rect 30550 4585 30600 4615
rect 30550 4565 30565 4585
rect 30585 4565 30600 4585
rect 30550 4535 30600 4565
rect 30550 4515 30565 4535
rect 30585 4515 30600 4535
rect 30550 4485 30600 4515
rect 30550 4465 30565 4485
rect 30585 4465 30600 4485
rect 30550 4435 30600 4465
rect 30550 4415 30565 4435
rect 30585 4415 30600 4435
rect 30550 4385 30600 4415
rect 30550 4365 30565 4385
rect 30585 4365 30600 4385
rect 30550 4350 30600 4365
rect 30700 4835 30750 4850
rect 30700 4815 30715 4835
rect 30735 4815 30750 4835
rect 30700 4785 30750 4815
rect 30700 4765 30715 4785
rect 30735 4765 30750 4785
rect 30700 4735 30750 4765
rect 30700 4715 30715 4735
rect 30735 4715 30750 4735
rect 30700 4685 30750 4715
rect 30700 4665 30715 4685
rect 30735 4665 30750 4685
rect 30700 4635 30750 4665
rect 30700 4615 30715 4635
rect 30735 4615 30750 4635
rect 30700 4585 30750 4615
rect 30700 4565 30715 4585
rect 30735 4565 30750 4585
rect 30700 4535 30750 4565
rect 30700 4515 30715 4535
rect 30735 4515 30750 4535
rect 30700 4485 30750 4515
rect 30700 4465 30715 4485
rect 30735 4465 30750 4485
rect 30700 4435 30750 4465
rect 30700 4415 30715 4435
rect 30735 4415 30750 4435
rect 30700 4385 30750 4415
rect 30700 4365 30715 4385
rect 30735 4365 30750 4385
rect 30700 4350 30750 4365
rect 30850 4835 30900 4850
rect 30850 4815 30865 4835
rect 30885 4815 30900 4835
rect 30850 4785 30900 4815
rect 30850 4765 30865 4785
rect 30885 4765 30900 4785
rect 30850 4735 30900 4765
rect 30850 4715 30865 4735
rect 30885 4715 30900 4735
rect 30850 4685 30900 4715
rect 30850 4665 30865 4685
rect 30885 4665 30900 4685
rect 30850 4635 30900 4665
rect 30850 4615 30865 4635
rect 30885 4615 30900 4635
rect 30850 4585 30900 4615
rect 30850 4565 30865 4585
rect 30885 4565 30900 4585
rect 30850 4535 30900 4565
rect 30850 4515 30865 4535
rect 30885 4515 30900 4535
rect 30850 4485 30900 4515
rect 30850 4465 30865 4485
rect 30885 4465 30900 4485
rect 30850 4435 30900 4465
rect 30850 4415 30865 4435
rect 30885 4415 30900 4435
rect 30850 4385 30900 4415
rect 30850 4365 30865 4385
rect 30885 4365 30900 4385
rect 30850 4350 30900 4365
rect 31000 4835 31050 4850
rect 31000 4815 31015 4835
rect 31035 4815 31050 4835
rect 31000 4785 31050 4815
rect 31000 4765 31015 4785
rect 31035 4765 31050 4785
rect 31000 4735 31050 4765
rect 31000 4715 31015 4735
rect 31035 4715 31050 4735
rect 31000 4685 31050 4715
rect 31000 4665 31015 4685
rect 31035 4665 31050 4685
rect 31000 4635 31050 4665
rect 31000 4615 31015 4635
rect 31035 4615 31050 4635
rect 31000 4585 31050 4615
rect 31000 4565 31015 4585
rect 31035 4565 31050 4585
rect 31000 4535 31050 4565
rect 31000 4515 31015 4535
rect 31035 4515 31050 4535
rect 31000 4485 31050 4515
rect 31000 4465 31015 4485
rect 31035 4465 31050 4485
rect 31000 4435 31050 4465
rect 31000 4415 31015 4435
rect 31035 4415 31050 4435
rect 31000 4385 31050 4415
rect 31000 4365 31015 4385
rect 31035 4365 31050 4385
rect 31000 4350 31050 4365
rect 31150 4835 31200 4850
rect 31150 4815 31165 4835
rect 31185 4815 31200 4835
rect 31150 4785 31200 4815
rect 31150 4765 31165 4785
rect 31185 4765 31200 4785
rect 31150 4735 31200 4765
rect 31150 4715 31165 4735
rect 31185 4715 31200 4735
rect 31150 4685 31200 4715
rect 31150 4665 31165 4685
rect 31185 4665 31200 4685
rect 31150 4635 31200 4665
rect 31150 4615 31165 4635
rect 31185 4615 31200 4635
rect 31150 4585 31200 4615
rect 31150 4565 31165 4585
rect 31185 4565 31200 4585
rect 31150 4535 31200 4565
rect 31150 4515 31165 4535
rect 31185 4515 31200 4535
rect 31150 4485 31200 4515
rect 31150 4465 31165 4485
rect 31185 4465 31200 4485
rect 31150 4435 31200 4465
rect 31150 4415 31165 4435
rect 31185 4415 31200 4435
rect 31150 4385 31200 4415
rect 31150 4365 31165 4385
rect 31185 4365 31200 4385
rect 31150 4350 31200 4365
rect 31300 4835 31350 4850
rect 31300 4815 31315 4835
rect 31335 4815 31350 4835
rect 31300 4785 31350 4815
rect 31300 4765 31315 4785
rect 31335 4765 31350 4785
rect 31300 4735 31350 4765
rect 31300 4715 31315 4735
rect 31335 4715 31350 4735
rect 31300 4685 31350 4715
rect 31300 4665 31315 4685
rect 31335 4665 31350 4685
rect 31300 4635 31350 4665
rect 31300 4615 31315 4635
rect 31335 4615 31350 4635
rect 31300 4585 31350 4615
rect 31300 4565 31315 4585
rect 31335 4565 31350 4585
rect 31300 4535 31350 4565
rect 31300 4515 31315 4535
rect 31335 4515 31350 4535
rect 31300 4485 31350 4515
rect 31300 4465 31315 4485
rect 31335 4465 31350 4485
rect 31300 4435 31350 4465
rect 31300 4415 31315 4435
rect 31335 4415 31350 4435
rect 31300 4385 31350 4415
rect 31300 4365 31315 4385
rect 31335 4365 31350 4385
rect 31300 4350 31350 4365
rect 31450 4835 31500 4850
rect 31450 4815 31465 4835
rect 31485 4815 31500 4835
rect 31450 4785 31500 4815
rect 31450 4765 31465 4785
rect 31485 4765 31500 4785
rect 31450 4735 31500 4765
rect 31450 4715 31465 4735
rect 31485 4715 31500 4735
rect 31450 4685 31500 4715
rect 31450 4665 31465 4685
rect 31485 4665 31500 4685
rect 31450 4635 31500 4665
rect 31450 4615 31465 4635
rect 31485 4615 31500 4635
rect 31450 4585 31500 4615
rect 31450 4565 31465 4585
rect 31485 4565 31500 4585
rect 31450 4535 31500 4565
rect 31450 4515 31465 4535
rect 31485 4515 31500 4535
rect 31450 4485 31500 4515
rect 31450 4465 31465 4485
rect 31485 4465 31500 4485
rect 31450 4435 31500 4465
rect 31450 4415 31465 4435
rect 31485 4415 31500 4435
rect 31450 4385 31500 4415
rect 31450 4365 31465 4385
rect 31485 4365 31500 4385
rect 31450 4350 31500 4365
rect 32050 4835 32100 4850
rect 32050 4815 32065 4835
rect 32085 4815 32100 4835
rect 32050 4785 32100 4815
rect 32050 4765 32065 4785
rect 32085 4765 32100 4785
rect 32050 4735 32100 4765
rect 32050 4715 32065 4735
rect 32085 4715 32100 4735
rect 32050 4685 32100 4715
rect 32050 4665 32065 4685
rect 32085 4665 32100 4685
rect 32050 4635 32100 4665
rect 32050 4615 32065 4635
rect 32085 4615 32100 4635
rect 32050 4585 32100 4615
rect 32050 4565 32065 4585
rect 32085 4565 32100 4585
rect 32050 4535 32100 4565
rect 32050 4515 32065 4535
rect 32085 4515 32100 4535
rect 32050 4485 32100 4515
rect 32050 4465 32065 4485
rect 32085 4465 32100 4485
rect 32050 4435 32100 4465
rect 32050 4415 32065 4435
rect 32085 4415 32100 4435
rect 32050 4385 32100 4415
rect 32050 4365 32065 4385
rect 32085 4365 32100 4385
rect 32050 4350 32100 4365
rect -650 4285 32100 4300
rect -650 4265 -635 4285
rect -615 4265 -585 4285
rect -565 4265 -535 4285
rect -515 4265 -485 4285
rect -465 4265 -435 4285
rect -415 4265 -385 4285
rect -365 4265 -335 4285
rect -315 4265 -285 4285
rect -265 4265 -235 4285
rect -215 4265 -185 4285
rect -165 4265 -135 4285
rect -115 4265 -85 4285
rect -65 4265 -35 4285
rect -15 4265 15 4285
rect 35 4265 65 4285
rect 85 4265 115 4285
rect 135 4265 165 4285
rect 185 4265 215 4285
rect 235 4265 265 4285
rect 285 4265 315 4285
rect 335 4265 365 4285
rect 385 4265 415 4285
rect 435 4265 465 4285
rect 485 4265 515 4285
rect 535 4265 565 4285
rect 585 4265 615 4285
rect 635 4265 665 4285
rect 685 4265 715 4285
rect 735 4265 765 4285
rect 785 4265 815 4285
rect 835 4265 865 4285
rect 885 4265 915 4285
rect 935 4265 965 4285
rect 985 4265 1015 4285
rect 1035 4265 1065 4285
rect 1085 4265 1115 4285
rect 1135 4265 1165 4285
rect 1185 4265 1215 4285
rect 1235 4265 1265 4285
rect 1285 4265 1315 4285
rect 1335 4265 1365 4285
rect 1385 4265 1415 4285
rect 1435 4265 1465 4285
rect 1485 4265 1515 4285
rect 1535 4265 1565 4285
rect 1585 4265 1615 4285
rect 1635 4265 1665 4285
rect 1685 4265 1715 4285
rect 1735 4265 1765 4285
rect 1785 4265 1815 4285
rect 1835 4265 1865 4285
rect 1885 4265 1915 4285
rect 1935 4265 1965 4285
rect 1985 4265 2015 4285
rect 2035 4265 2065 4285
rect 2085 4265 2115 4285
rect 2135 4265 2165 4285
rect 2185 4265 2215 4285
rect 2235 4265 2265 4285
rect 2285 4265 2315 4285
rect 2335 4265 2365 4285
rect 2385 4265 2415 4285
rect 2435 4265 2465 4285
rect 2485 4265 2515 4285
rect 2535 4265 2565 4285
rect 2585 4265 2615 4285
rect 2635 4265 2665 4285
rect 2685 4265 2715 4285
rect 2735 4265 2765 4285
rect 2785 4265 2815 4285
rect 2835 4265 2865 4285
rect 2885 4265 2915 4285
rect 2935 4265 2965 4285
rect 2985 4265 3015 4285
rect 3035 4265 3065 4285
rect 3085 4265 3115 4285
rect 3135 4265 3165 4285
rect 3185 4265 3215 4285
rect 3235 4265 3265 4285
rect 3285 4265 3315 4285
rect 3335 4265 3365 4285
rect 3385 4265 3415 4285
rect 3435 4265 3465 4285
rect 3485 4265 3515 4285
rect 3535 4265 3565 4285
rect 3585 4265 3615 4285
rect 3635 4265 3665 4285
rect 3685 4265 3715 4285
rect 3735 4265 3765 4285
rect 3785 4265 3815 4285
rect 3835 4265 3865 4285
rect 3885 4265 3915 4285
rect 3935 4265 3965 4285
rect 3985 4265 4015 4285
rect 4035 4265 4065 4285
rect 4085 4265 4115 4285
rect 4135 4265 4165 4285
rect 4185 4265 4215 4285
rect 4235 4265 4265 4285
rect 4285 4265 4315 4285
rect 4335 4265 4365 4285
rect 4385 4265 4415 4285
rect 4435 4265 4465 4285
rect 4485 4265 4515 4285
rect 4535 4265 4565 4285
rect 4585 4265 4615 4285
rect 4635 4265 4665 4285
rect 4685 4265 4715 4285
rect 4735 4265 4765 4285
rect 4785 4265 4815 4285
rect 4835 4265 4865 4285
rect 4885 4265 4915 4285
rect 4935 4265 4965 4285
rect 4985 4265 5015 4285
rect 5035 4265 5065 4285
rect 5085 4265 5115 4285
rect 5135 4265 5165 4285
rect 5185 4265 5215 4285
rect 5235 4265 5265 4285
rect 5285 4265 5315 4285
rect 5335 4265 5365 4285
rect 5385 4265 5415 4285
rect 5435 4265 5465 4285
rect 5485 4265 5515 4285
rect 5535 4265 5565 4285
rect 5585 4265 5615 4285
rect 5635 4265 5665 4285
rect 5685 4265 5715 4285
rect 5735 4265 5765 4285
rect 5785 4265 5815 4285
rect 5835 4265 5865 4285
rect 5885 4265 5915 4285
rect 5935 4265 5965 4285
rect 5985 4265 6015 4285
rect 6035 4265 6065 4285
rect 6085 4265 6115 4285
rect 6135 4265 6165 4285
rect 6185 4265 6215 4285
rect 6235 4265 6265 4285
rect 6285 4265 6315 4285
rect 6335 4265 6365 4285
rect 6385 4265 6415 4285
rect 6435 4265 6465 4285
rect 6485 4265 6515 4285
rect 6535 4265 6565 4285
rect 6585 4265 6615 4285
rect 6635 4265 6665 4285
rect 6685 4265 6715 4285
rect 6735 4265 6765 4285
rect 6785 4265 6815 4285
rect 6835 4265 6865 4285
rect 6885 4265 6915 4285
rect 6935 4265 6965 4285
rect 6985 4265 7015 4285
rect 7035 4265 7065 4285
rect 7085 4265 7115 4285
rect 7135 4265 7165 4285
rect 7185 4265 7215 4285
rect 7235 4265 7265 4285
rect 7285 4265 7315 4285
rect 7335 4265 7365 4285
rect 7385 4265 7415 4285
rect 7435 4265 7465 4285
rect 7485 4265 7515 4285
rect 7535 4265 7565 4285
rect 7585 4265 7615 4285
rect 7635 4265 7665 4285
rect 7685 4265 7715 4285
rect 7735 4265 7765 4285
rect 7785 4265 7815 4285
rect 7835 4265 7865 4285
rect 7885 4265 7915 4285
rect 7935 4265 7965 4285
rect 7985 4265 8015 4285
rect 8035 4265 8065 4285
rect 8085 4265 8115 4285
rect 8135 4265 8165 4285
rect 8185 4265 8215 4285
rect 8235 4265 8265 4285
rect 8285 4265 8315 4285
rect 8335 4265 8365 4285
rect 8385 4265 8415 4285
rect 8435 4265 8465 4285
rect 8485 4265 8515 4285
rect 8535 4265 8565 4285
rect 8585 4265 8615 4285
rect 8635 4265 8665 4285
rect 8685 4265 8715 4285
rect 8735 4265 8765 4285
rect 8785 4265 8815 4285
rect 8835 4265 8865 4285
rect 8885 4265 8915 4285
rect 8935 4265 8965 4285
rect 8985 4265 9015 4285
rect 9035 4265 9065 4285
rect 9085 4265 9115 4285
rect 9135 4265 9165 4285
rect 9185 4265 9215 4285
rect 9235 4265 9265 4285
rect 9285 4265 9315 4285
rect 9335 4265 9365 4285
rect 9385 4265 9415 4285
rect 9435 4265 9465 4285
rect 9485 4265 9515 4285
rect 9535 4265 9565 4285
rect 9585 4265 9615 4285
rect 9635 4265 9665 4285
rect 9685 4265 9715 4285
rect 9735 4265 9765 4285
rect 9785 4265 9815 4285
rect 9835 4265 9865 4285
rect 9885 4265 9915 4285
rect 9935 4265 9965 4285
rect 9985 4265 10015 4285
rect 10035 4265 10065 4285
rect 10085 4265 10115 4285
rect 10135 4265 10165 4285
rect 10185 4265 10215 4285
rect 10235 4265 10265 4285
rect 10285 4265 10315 4285
rect 10335 4265 10365 4285
rect 10385 4265 10415 4285
rect 10435 4265 10465 4285
rect 10485 4265 10515 4285
rect 10535 4265 10565 4285
rect 10585 4265 10615 4285
rect 10635 4265 10665 4285
rect 10685 4265 10715 4285
rect 10735 4265 10765 4285
rect 10785 4265 10815 4285
rect 10835 4265 10865 4285
rect 10885 4265 10915 4285
rect 10935 4265 10965 4285
rect 10985 4265 11015 4285
rect 11035 4265 11065 4285
rect 11085 4265 11115 4285
rect 11135 4265 11165 4285
rect 11185 4265 11215 4285
rect 11235 4265 11265 4285
rect 11285 4265 11315 4285
rect 11335 4265 11365 4285
rect 11385 4265 11415 4285
rect 11435 4265 11465 4285
rect 11485 4265 11515 4285
rect 11535 4265 11565 4285
rect 11585 4265 11615 4285
rect 11635 4265 11665 4285
rect 11685 4265 11715 4285
rect 11735 4265 11765 4285
rect 11785 4265 11815 4285
rect 11835 4265 11865 4285
rect 11885 4265 11915 4285
rect 11935 4265 11965 4285
rect 11985 4265 12015 4285
rect 12035 4265 12065 4285
rect 12085 4265 12115 4285
rect 12135 4265 12165 4285
rect 12185 4265 12215 4285
rect 12235 4265 12265 4285
rect 12285 4265 12315 4285
rect 12335 4265 12365 4285
rect 12385 4265 12415 4285
rect 12435 4265 12465 4285
rect 12485 4265 12515 4285
rect 12535 4265 12565 4285
rect 12585 4265 12615 4285
rect 12635 4265 12665 4285
rect 12685 4265 12715 4285
rect 12735 4265 12765 4285
rect 12785 4265 12815 4285
rect 12835 4265 12865 4285
rect 12885 4265 12915 4285
rect 12935 4265 12965 4285
rect 12985 4265 13015 4285
rect 13035 4265 13065 4285
rect 13085 4265 13115 4285
rect 13135 4265 13165 4285
rect 13185 4265 13215 4285
rect 13235 4265 13265 4285
rect 13285 4265 13315 4285
rect 13335 4265 13365 4285
rect 13385 4265 13415 4285
rect 13435 4265 13465 4285
rect 13485 4265 13515 4285
rect 13535 4265 13565 4285
rect 13585 4265 13615 4285
rect 13635 4265 13665 4285
rect 13685 4265 13715 4285
rect 13735 4265 13765 4285
rect 13785 4265 13815 4285
rect 13835 4265 13865 4285
rect 13885 4265 13915 4285
rect 13935 4265 13965 4285
rect 13985 4265 14015 4285
rect 14035 4265 14065 4285
rect 14085 4265 14115 4285
rect 14135 4265 14165 4285
rect 14185 4265 14215 4285
rect 14235 4265 14265 4285
rect 14285 4265 14315 4285
rect 14335 4265 14365 4285
rect 14385 4265 14415 4285
rect 14435 4265 14465 4285
rect 14485 4265 14515 4285
rect 14535 4265 14565 4285
rect 14585 4265 14615 4285
rect 14635 4265 14665 4285
rect 14685 4265 14715 4285
rect 14735 4265 14765 4285
rect 14785 4265 14815 4285
rect 14835 4265 14865 4285
rect 14885 4265 14915 4285
rect 14935 4265 14965 4285
rect 14985 4265 15015 4285
rect 15035 4265 15065 4285
rect 15085 4265 15115 4285
rect 15135 4265 15165 4285
rect 15185 4265 15215 4285
rect 15235 4265 15265 4285
rect 15285 4265 15315 4285
rect 15335 4265 15365 4285
rect 15385 4265 15415 4285
rect 15435 4265 15465 4285
rect 15485 4265 15515 4285
rect 15535 4265 15565 4285
rect 15585 4265 15615 4285
rect 15635 4265 15665 4285
rect 15685 4265 15715 4285
rect 15735 4265 15765 4285
rect 15785 4265 15815 4285
rect 15835 4265 15865 4285
rect 15885 4265 15915 4285
rect 15935 4265 15965 4285
rect 15985 4265 16015 4285
rect 16035 4265 16065 4285
rect 16085 4265 16115 4285
rect 16135 4265 16165 4285
rect 16185 4265 16215 4285
rect 16235 4265 16265 4285
rect 16285 4265 16315 4285
rect 16335 4265 16365 4285
rect 16385 4265 16415 4285
rect 16435 4265 16465 4285
rect 16485 4265 16515 4285
rect 16535 4265 16565 4285
rect 16585 4265 16615 4285
rect 16635 4265 16665 4285
rect 16685 4265 16715 4285
rect 16735 4265 16765 4285
rect 16785 4265 16815 4285
rect 16835 4265 16865 4285
rect 16885 4265 16915 4285
rect 16935 4265 16965 4285
rect 16985 4265 17015 4285
rect 17035 4265 17065 4285
rect 17085 4265 17115 4285
rect 17135 4265 17165 4285
rect 17185 4265 17215 4285
rect 17235 4265 17265 4285
rect 17285 4265 17315 4285
rect 17335 4265 17365 4285
rect 17385 4265 17415 4285
rect 17435 4265 17465 4285
rect 17485 4265 17515 4285
rect 17535 4265 17565 4285
rect 17585 4265 17615 4285
rect 17635 4265 17665 4285
rect 17685 4265 17715 4285
rect 17735 4265 17765 4285
rect 17785 4265 17815 4285
rect 17835 4265 17865 4285
rect 17885 4265 17915 4285
rect 17935 4265 17965 4285
rect 17985 4265 18015 4285
rect 18035 4265 18065 4285
rect 18085 4265 18115 4285
rect 18135 4265 18165 4285
rect 18185 4265 18215 4285
rect 18235 4265 18265 4285
rect 18285 4265 18315 4285
rect 18335 4265 18365 4285
rect 18385 4265 18415 4285
rect 18435 4265 18465 4285
rect 18485 4265 18515 4285
rect 18535 4265 18565 4285
rect 18585 4265 18615 4285
rect 18635 4265 18665 4285
rect 18685 4265 18715 4285
rect 18735 4265 18765 4285
rect 18785 4265 18815 4285
rect 18835 4265 18865 4285
rect 18885 4265 18915 4285
rect 18935 4265 18965 4285
rect 18985 4265 19015 4285
rect 19035 4265 19065 4285
rect 19085 4265 19115 4285
rect 19135 4265 19165 4285
rect 19185 4265 19215 4285
rect 19235 4265 19265 4285
rect 19285 4265 19315 4285
rect 19335 4265 19365 4285
rect 19385 4265 19415 4285
rect 19435 4265 19465 4285
rect 19485 4265 19515 4285
rect 19535 4265 19565 4285
rect 19585 4265 19615 4285
rect 19635 4265 19665 4285
rect 19685 4265 19715 4285
rect 19735 4265 19765 4285
rect 19785 4265 19815 4285
rect 19835 4265 19865 4285
rect 19885 4265 19915 4285
rect 19935 4265 19965 4285
rect 19985 4265 20015 4285
rect 20035 4265 20065 4285
rect 20085 4265 20115 4285
rect 20135 4265 20165 4285
rect 20185 4265 20215 4285
rect 20235 4265 20265 4285
rect 20285 4265 20315 4285
rect 20335 4265 20365 4285
rect 20385 4265 20415 4285
rect 20435 4265 20465 4285
rect 20485 4265 20515 4285
rect 20535 4265 20565 4285
rect 20585 4265 20615 4285
rect 20635 4265 20665 4285
rect 20685 4265 20715 4285
rect 20735 4265 20765 4285
rect 20785 4265 20815 4285
rect 20835 4265 20865 4285
rect 20885 4265 20915 4285
rect 20935 4265 20965 4285
rect 20985 4265 21015 4285
rect 21035 4265 21065 4285
rect 21085 4265 21115 4285
rect 21135 4265 21165 4285
rect 21185 4265 21215 4285
rect 21235 4265 21265 4285
rect 21285 4265 21315 4285
rect 21335 4265 21365 4285
rect 21385 4265 21415 4285
rect 21435 4265 21465 4285
rect 21485 4265 21515 4285
rect 21535 4265 21565 4285
rect 21585 4265 21615 4285
rect 21635 4265 21665 4285
rect 21685 4265 21715 4285
rect 21735 4265 21765 4285
rect 21785 4265 21815 4285
rect 21835 4265 21865 4285
rect 21885 4265 21915 4285
rect 21935 4265 21965 4285
rect 21985 4265 22015 4285
rect 22035 4265 22065 4285
rect 22085 4265 22115 4285
rect 22135 4265 22165 4285
rect 22185 4265 22215 4285
rect 22235 4265 22265 4285
rect 22285 4265 22315 4285
rect 22335 4265 22365 4285
rect 22385 4265 22415 4285
rect 22435 4265 22465 4285
rect 22485 4265 22515 4285
rect 22535 4265 22565 4285
rect 22585 4265 22615 4285
rect 22635 4265 22665 4285
rect 22685 4265 22715 4285
rect 22735 4265 22765 4285
rect 22785 4265 22815 4285
rect 22835 4265 22865 4285
rect 22885 4265 22915 4285
rect 22935 4265 22965 4285
rect 22985 4265 23015 4285
rect 23035 4265 23065 4285
rect 23085 4265 23115 4285
rect 23135 4265 23165 4285
rect 23185 4265 23215 4285
rect 23235 4265 23265 4285
rect 23285 4265 23315 4285
rect 23335 4265 23365 4285
rect 23385 4265 23415 4285
rect 23435 4265 23465 4285
rect 23485 4265 23515 4285
rect 23535 4265 23565 4285
rect 23585 4265 23615 4285
rect 23635 4265 23665 4285
rect 23685 4265 23715 4285
rect 23735 4265 23765 4285
rect 23785 4265 23815 4285
rect 23835 4265 23865 4285
rect 23885 4265 23915 4285
rect 23935 4265 23965 4285
rect 23985 4265 24015 4285
rect 24035 4265 24065 4285
rect 24085 4265 24115 4285
rect 24135 4265 24165 4285
rect 24185 4265 24215 4285
rect 24235 4265 24265 4285
rect 24285 4265 24315 4285
rect 24335 4265 24365 4285
rect 24385 4265 24415 4285
rect 24435 4265 24465 4285
rect 24485 4265 24515 4285
rect 24535 4265 24565 4285
rect 24585 4265 24615 4285
rect 24635 4265 24665 4285
rect 24685 4265 24715 4285
rect 24735 4265 24765 4285
rect 24785 4265 24815 4285
rect 24835 4265 24865 4285
rect 24885 4265 24915 4285
rect 24935 4265 24965 4285
rect 24985 4265 25015 4285
rect 25035 4265 25065 4285
rect 25085 4265 25115 4285
rect 25135 4265 25165 4285
rect 25185 4265 25215 4285
rect 25235 4265 25265 4285
rect 25285 4265 25315 4285
rect 25335 4265 25365 4285
rect 25385 4265 25415 4285
rect 25435 4265 25465 4285
rect 25485 4265 25515 4285
rect 25535 4265 25565 4285
rect 25585 4265 25615 4285
rect 25635 4265 25665 4285
rect 25685 4265 25715 4285
rect 25735 4265 25765 4285
rect 25785 4265 25815 4285
rect 25835 4265 25865 4285
rect 25885 4265 25915 4285
rect 25935 4265 25965 4285
rect 25985 4265 26015 4285
rect 26035 4265 26065 4285
rect 26085 4265 26115 4285
rect 26135 4265 26165 4285
rect 26185 4265 26215 4285
rect 26235 4265 26265 4285
rect 26285 4265 26315 4285
rect 26335 4265 26365 4285
rect 26385 4265 26415 4285
rect 26435 4265 26465 4285
rect 26485 4265 26515 4285
rect 26535 4265 26565 4285
rect 26585 4265 26615 4285
rect 26635 4265 26665 4285
rect 26685 4265 26715 4285
rect 26735 4265 26765 4285
rect 26785 4265 26815 4285
rect 26835 4265 26865 4285
rect 26885 4265 26915 4285
rect 26935 4265 26965 4285
rect 26985 4265 27015 4285
rect 27035 4265 27065 4285
rect 27085 4265 27115 4285
rect 27135 4265 27165 4285
rect 27185 4265 27215 4285
rect 27235 4265 27265 4285
rect 27285 4265 27315 4285
rect 27335 4265 27365 4285
rect 27385 4265 27415 4285
rect 27435 4265 27465 4285
rect 27485 4265 27515 4285
rect 27535 4265 27565 4285
rect 27585 4265 27615 4285
rect 27635 4265 27665 4285
rect 27685 4265 27715 4285
rect 27735 4265 27765 4285
rect 27785 4265 27815 4285
rect 27835 4265 27865 4285
rect 27885 4265 27915 4285
rect 27935 4265 27965 4285
rect 27985 4265 28015 4285
rect 28035 4265 28065 4285
rect 28085 4265 28115 4285
rect 28135 4265 28165 4285
rect 28185 4265 28215 4285
rect 28235 4265 28265 4285
rect 28285 4265 28315 4285
rect 28335 4265 28365 4285
rect 28385 4265 28415 4285
rect 28435 4265 28465 4285
rect 28485 4265 28515 4285
rect 28535 4265 28565 4285
rect 28585 4265 28615 4285
rect 28635 4265 28665 4285
rect 28685 4265 28715 4285
rect 28735 4265 28765 4285
rect 28785 4265 28815 4285
rect 28835 4265 28865 4285
rect 28885 4265 28915 4285
rect 28935 4265 28965 4285
rect 28985 4265 29015 4285
rect 29035 4265 29065 4285
rect 29085 4265 29115 4285
rect 29135 4265 29165 4285
rect 29185 4265 29215 4285
rect 29235 4265 29265 4285
rect 29285 4265 29315 4285
rect 29335 4265 29365 4285
rect 29385 4265 29415 4285
rect 29435 4265 29465 4285
rect 29485 4265 29515 4285
rect 29535 4265 29565 4285
rect 29585 4265 29615 4285
rect 29635 4265 29665 4285
rect 29685 4265 29715 4285
rect 29735 4265 29765 4285
rect 29785 4265 29815 4285
rect 29835 4265 29865 4285
rect 29885 4265 29915 4285
rect 29935 4265 29965 4285
rect 29985 4265 30015 4285
rect 30035 4265 30065 4285
rect 30085 4265 30115 4285
rect 30135 4265 30165 4285
rect 30185 4265 30215 4285
rect 30235 4265 30265 4285
rect 30285 4265 30315 4285
rect 30335 4265 30365 4285
rect 30385 4265 30415 4285
rect 30435 4265 30465 4285
rect 30485 4265 30515 4285
rect 30535 4265 30565 4285
rect 30585 4265 30615 4285
rect 30635 4265 30665 4285
rect 30685 4265 30715 4285
rect 30735 4265 30765 4285
rect 30785 4265 30815 4285
rect 30835 4265 30865 4285
rect 30885 4265 30915 4285
rect 30935 4265 30965 4285
rect 30985 4265 31015 4285
rect 31035 4265 31065 4285
rect 31085 4265 31115 4285
rect 31135 4265 31165 4285
rect 31185 4265 31215 4285
rect 31235 4265 31265 4285
rect 31285 4265 31315 4285
rect 31335 4265 31365 4285
rect 31385 4265 31415 4285
rect 31435 4265 31465 4285
rect 31485 4265 31515 4285
rect 31535 4265 31565 4285
rect 31585 4265 31615 4285
rect 31635 4265 31665 4285
rect 31685 4265 31715 4285
rect 31735 4265 31765 4285
rect 31785 4265 31815 4285
rect 31835 4265 31865 4285
rect 31885 4265 31915 4285
rect 31935 4265 31965 4285
rect 31985 4265 32015 4285
rect 32035 4265 32065 4285
rect 32085 4265 32100 4285
rect -650 4250 32100 4265
rect -650 4185 -600 4200
rect -650 4165 -635 4185
rect -615 4165 -600 4185
rect -650 4135 -600 4165
rect -650 4115 -635 4135
rect -615 4115 -600 4135
rect -650 4085 -600 4115
rect -650 4065 -635 4085
rect -615 4065 -600 4085
rect -650 4035 -600 4065
rect -650 4015 -635 4035
rect -615 4015 -600 4035
rect -650 3985 -600 4015
rect -650 3965 -635 3985
rect -615 3965 -600 3985
rect -650 3935 -600 3965
rect -650 3915 -635 3935
rect -615 3915 -600 3935
rect -650 3885 -600 3915
rect -650 3865 -635 3885
rect -615 3865 -600 3885
rect -650 3835 -600 3865
rect -650 3815 -635 3835
rect -615 3815 -600 3835
rect -650 3785 -600 3815
rect -650 3765 -635 3785
rect -615 3765 -600 3785
rect -650 3735 -600 3765
rect -650 3715 -635 3735
rect -615 3715 -600 3735
rect -650 3700 -600 3715
rect -500 4185 -450 4200
rect -500 4165 -485 4185
rect -465 4165 -450 4185
rect -500 4135 -450 4165
rect -500 4115 -485 4135
rect -465 4115 -450 4135
rect -500 4085 -450 4115
rect -500 4065 -485 4085
rect -465 4065 -450 4085
rect -500 4035 -450 4065
rect -500 4015 -485 4035
rect -465 4015 -450 4035
rect -500 3985 -450 4015
rect -500 3965 -485 3985
rect -465 3965 -450 3985
rect -500 3935 -450 3965
rect -500 3915 -485 3935
rect -465 3915 -450 3935
rect -500 3885 -450 3915
rect -500 3865 -485 3885
rect -465 3865 -450 3885
rect -500 3835 -450 3865
rect -500 3815 -485 3835
rect -465 3815 -450 3835
rect -500 3785 -450 3815
rect -500 3765 -485 3785
rect -465 3765 -450 3785
rect -500 3735 -450 3765
rect -500 3715 -485 3735
rect -465 3715 -450 3735
rect -500 3700 -450 3715
rect -350 4185 -300 4200
rect -350 4165 -335 4185
rect -315 4165 -300 4185
rect -350 4135 -300 4165
rect -350 4115 -335 4135
rect -315 4115 -300 4135
rect -350 4085 -300 4115
rect -350 4065 -335 4085
rect -315 4065 -300 4085
rect -350 4035 -300 4065
rect -350 4015 -335 4035
rect -315 4015 -300 4035
rect -350 3985 -300 4015
rect -350 3965 -335 3985
rect -315 3965 -300 3985
rect -350 3935 -300 3965
rect -350 3915 -335 3935
rect -315 3915 -300 3935
rect -350 3885 -300 3915
rect -350 3865 -335 3885
rect -315 3865 -300 3885
rect -350 3835 -300 3865
rect -350 3815 -335 3835
rect -315 3815 -300 3835
rect -350 3785 -300 3815
rect -350 3765 -335 3785
rect -315 3765 -300 3785
rect -350 3735 -300 3765
rect -350 3715 -335 3735
rect -315 3715 -300 3735
rect -350 3700 -300 3715
rect -200 4185 -150 4200
rect -200 4165 -185 4185
rect -165 4165 -150 4185
rect -200 4135 -150 4165
rect -200 4115 -185 4135
rect -165 4115 -150 4135
rect -200 4085 -150 4115
rect -200 4065 -185 4085
rect -165 4065 -150 4085
rect -200 4035 -150 4065
rect -200 4015 -185 4035
rect -165 4015 -150 4035
rect -200 3985 -150 4015
rect -200 3965 -185 3985
rect -165 3965 -150 3985
rect -200 3935 -150 3965
rect -200 3915 -185 3935
rect -165 3915 -150 3935
rect -200 3885 -150 3915
rect -200 3865 -185 3885
rect -165 3865 -150 3885
rect -200 3835 -150 3865
rect -200 3815 -185 3835
rect -165 3815 -150 3835
rect -200 3785 -150 3815
rect -200 3765 -185 3785
rect -165 3765 -150 3785
rect -200 3735 -150 3765
rect -200 3715 -185 3735
rect -165 3715 -150 3735
rect -200 3700 -150 3715
rect -50 4185 0 4200
rect -50 4165 -35 4185
rect -15 4165 0 4185
rect -50 4135 0 4165
rect -50 4115 -35 4135
rect -15 4115 0 4135
rect -50 4085 0 4115
rect -50 4065 -35 4085
rect -15 4065 0 4085
rect -50 4035 0 4065
rect -50 4015 -35 4035
rect -15 4015 0 4035
rect -50 3985 0 4015
rect -50 3965 -35 3985
rect -15 3965 0 3985
rect -50 3935 0 3965
rect -50 3915 -35 3935
rect -15 3915 0 3935
rect -50 3885 0 3915
rect -50 3865 -35 3885
rect -15 3865 0 3885
rect -50 3835 0 3865
rect -50 3815 -35 3835
rect -15 3815 0 3835
rect -50 3785 0 3815
rect -50 3765 -35 3785
rect -15 3765 0 3785
rect -50 3735 0 3765
rect -50 3715 -35 3735
rect -15 3715 0 3735
rect -50 3700 0 3715
rect 550 4185 600 4200
rect 550 4165 565 4185
rect 585 4165 600 4185
rect 550 4135 600 4165
rect 550 4115 565 4135
rect 585 4115 600 4135
rect 550 4085 600 4115
rect 550 4065 565 4085
rect 585 4065 600 4085
rect 550 4035 600 4065
rect 550 4015 565 4035
rect 585 4015 600 4035
rect 550 3985 600 4015
rect 550 3965 565 3985
rect 585 3965 600 3985
rect 550 3935 600 3965
rect 550 3915 565 3935
rect 585 3915 600 3935
rect 550 3885 600 3915
rect 550 3865 565 3885
rect 585 3865 600 3885
rect 550 3835 600 3865
rect 550 3815 565 3835
rect 585 3815 600 3835
rect 550 3785 600 3815
rect 550 3765 565 3785
rect 585 3765 600 3785
rect 550 3735 600 3765
rect 550 3715 565 3735
rect 585 3715 600 3735
rect 550 3700 600 3715
rect 700 4185 750 4200
rect 700 4165 715 4185
rect 735 4165 750 4185
rect 700 4135 750 4165
rect 700 4115 715 4135
rect 735 4115 750 4135
rect 700 4085 750 4115
rect 700 4065 715 4085
rect 735 4065 750 4085
rect 700 4035 750 4065
rect 700 4015 715 4035
rect 735 4015 750 4035
rect 700 3985 750 4015
rect 700 3965 715 3985
rect 735 3965 750 3985
rect 700 3935 750 3965
rect 700 3915 715 3935
rect 735 3915 750 3935
rect 700 3885 750 3915
rect 700 3865 715 3885
rect 735 3865 750 3885
rect 700 3835 750 3865
rect 700 3815 715 3835
rect 735 3815 750 3835
rect 700 3785 750 3815
rect 700 3765 715 3785
rect 735 3765 750 3785
rect 700 3735 750 3765
rect 700 3715 715 3735
rect 735 3715 750 3735
rect 700 3700 750 3715
rect 850 4185 900 4200
rect 850 4165 865 4185
rect 885 4165 900 4185
rect 850 4135 900 4165
rect 850 4115 865 4135
rect 885 4115 900 4135
rect 850 4085 900 4115
rect 850 4065 865 4085
rect 885 4065 900 4085
rect 850 4035 900 4065
rect 850 4015 865 4035
rect 885 4015 900 4035
rect 850 3985 900 4015
rect 850 3965 865 3985
rect 885 3965 900 3985
rect 850 3935 900 3965
rect 850 3915 865 3935
rect 885 3915 900 3935
rect 850 3885 900 3915
rect 850 3865 865 3885
rect 885 3865 900 3885
rect 850 3835 900 3865
rect 850 3815 865 3835
rect 885 3815 900 3835
rect 850 3785 900 3815
rect 850 3765 865 3785
rect 885 3765 900 3785
rect 850 3735 900 3765
rect 850 3715 865 3735
rect 885 3715 900 3735
rect 850 3700 900 3715
rect 1000 4185 1050 4200
rect 1000 4165 1015 4185
rect 1035 4165 1050 4185
rect 1000 4135 1050 4165
rect 1000 4115 1015 4135
rect 1035 4115 1050 4135
rect 1000 4085 1050 4115
rect 1000 4065 1015 4085
rect 1035 4065 1050 4085
rect 1000 4035 1050 4065
rect 1000 4015 1015 4035
rect 1035 4015 1050 4035
rect 1000 3985 1050 4015
rect 1000 3965 1015 3985
rect 1035 3965 1050 3985
rect 1000 3935 1050 3965
rect 1000 3915 1015 3935
rect 1035 3915 1050 3935
rect 1000 3885 1050 3915
rect 1000 3865 1015 3885
rect 1035 3865 1050 3885
rect 1000 3835 1050 3865
rect 1000 3815 1015 3835
rect 1035 3815 1050 3835
rect 1000 3785 1050 3815
rect 1000 3765 1015 3785
rect 1035 3765 1050 3785
rect 1000 3735 1050 3765
rect 1000 3715 1015 3735
rect 1035 3715 1050 3735
rect 1000 3700 1050 3715
rect 1150 4185 1200 4200
rect 1150 4165 1165 4185
rect 1185 4165 1200 4185
rect 1150 4135 1200 4165
rect 1150 4115 1165 4135
rect 1185 4115 1200 4135
rect 1150 4085 1200 4115
rect 1150 4065 1165 4085
rect 1185 4065 1200 4085
rect 1150 4035 1200 4065
rect 1150 4015 1165 4035
rect 1185 4015 1200 4035
rect 1150 3985 1200 4015
rect 1150 3965 1165 3985
rect 1185 3965 1200 3985
rect 1150 3935 1200 3965
rect 1150 3915 1165 3935
rect 1185 3915 1200 3935
rect 1150 3885 1200 3915
rect 1150 3865 1165 3885
rect 1185 3865 1200 3885
rect 1150 3835 1200 3865
rect 1150 3815 1165 3835
rect 1185 3815 1200 3835
rect 1150 3785 1200 3815
rect 1150 3765 1165 3785
rect 1185 3765 1200 3785
rect 1150 3735 1200 3765
rect 1150 3715 1165 3735
rect 1185 3715 1200 3735
rect 1150 3700 1200 3715
rect 1300 4185 1350 4200
rect 1300 4165 1315 4185
rect 1335 4165 1350 4185
rect 1300 4135 1350 4165
rect 1300 4115 1315 4135
rect 1335 4115 1350 4135
rect 1300 4085 1350 4115
rect 1300 4065 1315 4085
rect 1335 4065 1350 4085
rect 1300 4035 1350 4065
rect 1300 4015 1315 4035
rect 1335 4015 1350 4035
rect 1300 3985 1350 4015
rect 1300 3965 1315 3985
rect 1335 3965 1350 3985
rect 1300 3935 1350 3965
rect 1300 3915 1315 3935
rect 1335 3915 1350 3935
rect 1300 3885 1350 3915
rect 1300 3865 1315 3885
rect 1335 3865 1350 3885
rect 1300 3835 1350 3865
rect 1300 3815 1315 3835
rect 1335 3815 1350 3835
rect 1300 3785 1350 3815
rect 1300 3765 1315 3785
rect 1335 3765 1350 3785
rect 1300 3735 1350 3765
rect 1300 3715 1315 3735
rect 1335 3715 1350 3735
rect 1300 3700 1350 3715
rect 1450 4185 1500 4200
rect 1450 4165 1465 4185
rect 1485 4165 1500 4185
rect 1450 4135 1500 4165
rect 1450 4115 1465 4135
rect 1485 4115 1500 4135
rect 1450 4085 1500 4115
rect 1450 4065 1465 4085
rect 1485 4065 1500 4085
rect 1450 4035 1500 4065
rect 1450 4015 1465 4035
rect 1485 4015 1500 4035
rect 1450 3985 1500 4015
rect 1450 3965 1465 3985
rect 1485 3965 1500 3985
rect 1450 3935 1500 3965
rect 1450 3915 1465 3935
rect 1485 3915 1500 3935
rect 1450 3885 1500 3915
rect 1450 3865 1465 3885
rect 1485 3865 1500 3885
rect 1450 3835 1500 3865
rect 1450 3815 1465 3835
rect 1485 3815 1500 3835
rect 1450 3785 1500 3815
rect 1450 3765 1465 3785
rect 1485 3765 1500 3785
rect 1450 3735 1500 3765
rect 1450 3715 1465 3735
rect 1485 3715 1500 3735
rect 1450 3700 1500 3715
rect 1600 4185 1650 4200
rect 1600 4165 1615 4185
rect 1635 4165 1650 4185
rect 1600 4135 1650 4165
rect 1600 4115 1615 4135
rect 1635 4115 1650 4135
rect 1600 4085 1650 4115
rect 1600 4065 1615 4085
rect 1635 4065 1650 4085
rect 1600 4035 1650 4065
rect 1600 4015 1615 4035
rect 1635 4015 1650 4035
rect 1600 3985 1650 4015
rect 1600 3965 1615 3985
rect 1635 3965 1650 3985
rect 1600 3935 1650 3965
rect 1600 3915 1615 3935
rect 1635 3915 1650 3935
rect 1600 3885 1650 3915
rect 1600 3865 1615 3885
rect 1635 3865 1650 3885
rect 1600 3835 1650 3865
rect 1600 3815 1615 3835
rect 1635 3815 1650 3835
rect 1600 3785 1650 3815
rect 1600 3765 1615 3785
rect 1635 3765 1650 3785
rect 1600 3735 1650 3765
rect 1600 3715 1615 3735
rect 1635 3715 1650 3735
rect 1600 3700 1650 3715
rect 1750 4185 1800 4200
rect 1750 4165 1765 4185
rect 1785 4165 1800 4185
rect 1750 4135 1800 4165
rect 1750 4115 1765 4135
rect 1785 4115 1800 4135
rect 1750 4085 1800 4115
rect 1750 4065 1765 4085
rect 1785 4065 1800 4085
rect 1750 4035 1800 4065
rect 1750 4015 1765 4035
rect 1785 4015 1800 4035
rect 1750 3985 1800 4015
rect 1750 3965 1765 3985
rect 1785 3965 1800 3985
rect 1750 3935 1800 3965
rect 1750 3915 1765 3935
rect 1785 3915 1800 3935
rect 1750 3885 1800 3915
rect 1750 3865 1765 3885
rect 1785 3865 1800 3885
rect 1750 3835 1800 3865
rect 1750 3815 1765 3835
rect 1785 3815 1800 3835
rect 1750 3785 1800 3815
rect 1750 3765 1765 3785
rect 1785 3765 1800 3785
rect 1750 3735 1800 3765
rect 1750 3715 1765 3735
rect 1785 3715 1800 3735
rect 1750 3700 1800 3715
rect 1900 4185 1950 4200
rect 1900 4165 1915 4185
rect 1935 4165 1950 4185
rect 1900 4135 1950 4165
rect 1900 4115 1915 4135
rect 1935 4115 1950 4135
rect 1900 4085 1950 4115
rect 1900 4065 1915 4085
rect 1935 4065 1950 4085
rect 1900 4035 1950 4065
rect 1900 4015 1915 4035
rect 1935 4015 1950 4035
rect 1900 3985 1950 4015
rect 1900 3965 1915 3985
rect 1935 3965 1950 3985
rect 1900 3935 1950 3965
rect 1900 3915 1915 3935
rect 1935 3915 1950 3935
rect 1900 3885 1950 3915
rect 1900 3865 1915 3885
rect 1935 3865 1950 3885
rect 1900 3835 1950 3865
rect 1900 3815 1915 3835
rect 1935 3815 1950 3835
rect 1900 3785 1950 3815
rect 1900 3765 1915 3785
rect 1935 3765 1950 3785
rect 1900 3735 1950 3765
rect 1900 3715 1915 3735
rect 1935 3715 1950 3735
rect 1900 3700 1950 3715
rect 2050 4185 2100 4200
rect 2050 4165 2065 4185
rect 2085 4165 2100 4185
rect 2050 4135 2100 4165
rect 2050 4115 2065 4135
rect 2085 4115 2100 4135
rect 2050 4085 2100 4115
rect 2050 4065 2065 4085
rect 2085 4065 2100 4085
rect 2050 4035 2100 4065
rect 2050 4015 2065 4035
rect 2085 4015 2100 4035
rect 2050 3985 2100 4015
rect 2050 3965 2065 3985
rect 2085 3965 2100 3985
rect 2050 3935 2100 3965
rect 2050 3915 2065 3935
rect 2085 3915 2100 3935
rect 2050 3885 2100 3915
rect 2050 3865 2065 3885
rect 2085 3865 2100 3885
rect 2050 3835 2100 3865
rect 2050 3815 2065 3835
rect 2085 3815 2100 3835
rect 2050 3785 2100 3815
rect 2050 3765 2065 3785
rect 2085 3765 2100 3785
rect 2050 3735 2100 3765
rect 2050 3715 2065 3735
rect 2085 3715 2100 3735
rect 2050 3700 2100 3715
rect 2200 4185 2250 4200
rect 2200 4165 2215 4185
rect 2235 4165 2250 4185
rect 2200 4135 2250 4165
rect 2200 4115 2215 4135
rect 2235 4115 2250 4135
rect 2200 4085 2250 4115
rect 2200 4065 2215 4085
rect 2235 4065 2250 4085
rect 2200 4035 2250 4065
rect 2200 4015 2215 4035
rect 2235 4015 2250 4035
rect 2200 3985 2250 4015
rect 2200 3965 2215 3985
rect 2235 3965 2250 3985
rect 2200 3935 2250 3965
rect 2200 3915 2215 3935
rect 2235 3915 2250 3935
rect 2200 3885 2250 3915
rect 2200 3865 2215 3885
rect 2235 3865 2250 3885
rect 2200 3835 2250 3865
rect 2200 3815 2215 3835
rect 2235 3815 2250 3835
rect 2200 3785 2250 3815
rect 2200 3765 2215 3785
rect 2235 3765 2250 3785
rect 2200 3735 2250 3765
rect 2200 3715 2215 3735
rect 2235 3715 2250 3735
rect 2200 3700 2250 3715
rect 2350 4185 2400 4200
rect 2350 4165 2365 4185
rect 2385 4165 2400 4185
rect 2350 4135 2400 4165
rect 2350 4115 2365 4135
rect 2385 4115 2400 4135
rect 2350 4085 2400 4115
rect 2350 4065 2365 4085
rect 2385 4065 2400 4085
rect 2350 4035 2400 4065
rect 2350 4015 2365 4035
rect 2385 4015 2400 4035
rect 2350 3985 2400 4015
rect 2350 3965 2365 3985
rect 2385 3965 2400 3985
rect 2350 3935 2400 3965
rect 2350 3915 2365 3935
rect 2385 3915 2400 3935
rect 2350 3885 2400 3915
rect 2350 3865 2365 3885
rect 2385 3865 2400 3885
rect 2350 3835 2400 3865
rect 2350 3815 2365 3835
rect 2385 3815 2400 3835
rect 2350 3785 2400 3815
rect 2350 3765 2365 3785
rect 2385 3765 2400 3785
rect 2350 3735 2400 3765
rect 2350 3715 2365 3735
rect 2385 3715 2400 3735
rect 2350 3700 2400 3715
rect 2500 4185 2550 4200
rect 2500 4165 2515 4185
rect 2535 4165 2550 4185
rect 2500 4135 2550 4165
rect 2500 4115 2515 4135
rect 2535 4115 2550 4135
rect 2500 4085 2550 4115
rect 2500 4065 2515 4085
rect 2535 4065 2550 4085
rect 2500 4035 2550 4065
rect 2500 4015 2515 4035
rect 2535 4015 2550 4035
rect 2500 3985 2550 4015
rect 2500 3965 2515 3985
rect 2535 3965 2550 3985
rect 2500 3935 2550 3965
rect 2500 3915 2515 3935
rect 2535 3915 2550 3935
rect 2500 3885 2550 3915
rect 2500 3865 2515 3885
rect 2535 3865 2550 3885
rect 2500 3835 2550 3865
rect 2500 3815 2515 3835
rect 2535 3815 2550 3835
rect 2500 3785 2550 3815
rect 2500 3765 2515 3785
rect 2535 3765 2550 3785
rect 2500 3735 2550 3765
rect 2500 3715 2515 3735
rect 2535 3715 2550 3735
rect 2500 3700 2550 3715
rect 2650 4185 2700 4200
rect 2650 4165 2665 4185
rect 2685 4165 2700 4185
rect 2650 4135 2700 4165
rect 2650 4115 2665 4135
rect 2685 4115 2700 4135
rect 2650 4085 2700 4115
rect 2650 4065 2665 4085
rect 2685 4065 2700 4085
rect 2650 4035 2700 4065
rect 2650 4015 2665 4035
rect 2685 4015 2700 4035
rect 2650 3985 2700 4015
rect 2650 3965 2665 3985
rect 2685 3965 2700 3985
rect 2650 3935 2700 3965
rect 2650 3915 2665 3935
rect 2685 3915 2700 3935
rect 2650 3885 2700 3915
rect 2650 3865 2665 3885
rect 2685 3865 2700 3885
rect 2650 3835 2700 3865
rect 2650 3815 2665 3835
rect 2685 3815 2700 3835
rect 2650 3785 2700 3815
rect 2650 3765 2665 3785
rect 2685 3765 2700 3785
rect 2650 3735 2700 3765
rect 2650 3715 2665 3735
rect 2685 3715 2700 3735
rect 2650 3700 2700 3715
rect 2800 4185 2850 4200
rect 2800 4165 2815 4185
rect 2835 4165 2850 4185
rect 2800 4135 2850 4165
rect 2800 4115 2815 4135
rect 2835 4115 2850 4135
rect 2800 4085 2850 4115
rect 2800 4065 2815 4085
rect 2835 4065 2850 4085
rect 2800 4035 2850 4065
rect 2800 4015 2815 4035
rect 2835 4015 2850 4035
rect 2800 3985 2850 4015
rect 2800 3965 2815 3985
rect 2835 3965 2850 3985
rect 2800 3935 2850 3965
rect 2800 3915 2815 3935
rect 2835 3915 2850 3935
rect 2800 3885 2850 3915
rect 2800 3865 2815 3885
rect 2835 3865 2850 3885
rect 2800 3835 2850 3865
rect 2800 3815 2815 3835
rect 2835 3815 2850 3835
rect 2800 3785 2850 3815
rect 2800 3765 2815 3785
rect 2835 3765 2850 3785
rect 2800 3735 2850 3765
rect 2800 3715 2815 3735
rect 2835 3715 2850 3735
rect 2800 3700 2850 3715
rect 2950 4185 3000 4200
rect 2950 4165 2965 4185
rect 2985 4165 3000 4185
rect 2950 4135 3000 4165
rect 2950 4115 2965 4135
rect 2985 4115 3000 4135
rect 2950 4085 3000 4115
rect 2950 4065 2965 4085
rect 2985 4065 3000 4085
rect 2950 4035 3000 4065
rect 2950 4015 2965 4035
rect 2985 4015 3000 4035
rect 2950 3985 3000 4015
rect 2950 3965 2965 3985
rect 2985 3965 3000 3985
rect 2950 3935 3000 3965
rect 2950 3915 2965 3935
rect 2985 3915 3000 3935
rect 2950 3885 3000 3915
rect 2950 3865 2965 3885
rect 2985 3865 3000 3885
rect 2950 3835 3000 3865
rect 2950 3815 2965 3835
rect 2985 3815 3000 3835
rect 2950 3785 3000 3815
rect 2950 3765 2965 3785
rect 2985 3765 3000 3785
rect 2950 3735 3000 3765
rect 2950 3715 2965 3735
rect 2985 3715 3000 3735
rect 2950 3700 3000 3715
rect 3100 4185 3150 4200
rect 3100 4165 3115 4185
rect 3135 4165 3150 4185
rect 3100 4135 3150 4165
rect 3100 4115 3115 4135
rect 3135 4115 3150 4135
rect 3100 4085 3150 4115
rect 3100 4065 3115 4085
rect 3135 4065 3150 4085
rect 3100 4035 3150 4065
rect 3100 4015 3115 4035
rect 3135 4015 3150 4035
rect 3100 3985 3150 4015
rect 3100 3965 3115 3985
rect 3135 3965 3150 3985
rect 3100 3935 3150 3965
rect 3100 3915 3115 3935
rect 3135 3915 3150 3935
rect 3100 3885 3150 3915
rect 3100 3865 3115 3885
rect 3135 3865 3150 3885
rect 3100 3835 3150 3865
rect 3100 3815 3115 3835
rect 3135 3815 3150 3835
rect 3100 3785 3150 3815
rect 3100 3765 3115 3785
rect 3135 3765 3150 3785
rect 3100 3735 3150 3765
rect 3100 3715 3115 3735
rect 3135 3715 3150 3735
rect 3100 3700 3150 3715
rect 3250 4185 3300 4200
rect 3250 4165 3265 4185
rect 3285 4165 3300 4185
rect 3250 4135 3300 4165
rect 3250 4115 3265 4135
rect 3285 4115 3300 4135
rect 3250 4085 3300 4115
rect 3250 4065 3265 4085
rect 3285 4065 3300 4085
rect 3250 4035 3300 4065
rect 3250 4015 3265 4035
rect 3285 4015 3300 4035
rect 3250 3985 3300 4015
rect 3250 3965 3265 3985
rect 3285 3965 3300 3985
rect 3250 3935 3300 3965
rect 3250 3915 3265 3935
rect 3285 3915 3300 3935
rect 3250 3885 3300 3915
rect 3250 3865 3265 3885
rect 3285 3865 3300 3885
rect 3250 3835 3300 3865
rect 3250 3815 3265 3835
rect 3285 3815 3300 3835
rect 3250 3785 3300 3815
rect 3250 3765 3265 3785
rect 3285 3765 3300 3785
rect 3250 3735 3300 3765
rect 3250 3715 3265 3735
rect 3285 3715 3300 3735
rect 3250 3700 3300 3715
rect 3400 4185 3450 4200
rect 3400 4165 3415 4185
rect 3435 4165 3450 4185
rect 3400 4135 3450 4165
rect 3400 4115 3415 4135
rect 3435 4115 3450 4135
rect 3400 4085 3450 4115
rect 3400 4065 3415 4085
rect 3435 4065 3450 4085
rect 3400 4035 3450 4065
rect 3400 4015 3415 4035
rect 3435 4015 3450 4035
rect 3400 3985 3450 4015
rect 3400 3965 3415 3985
rect 3435 3965 3450 3985
rect 3400 3935 3450 3965
rect 3400 3915 3415 3935
rect 3435 3915 3450 3935
rect 3400 3885 3450 3915
rect 3400 3865 3415 3885
rect 3435 3865 3450 3885
rect 3400 3835 3450 3865
rect 3400 3815 3415 3835
rect 3435 3815 3450 3835
rect 3400 3785 3450 3815
rect 3400 3765 3415 3785
rect 3435 3765 3450 3785
rect 3400 3735 3450 3765
rect 3400 3715 3415 3735
rect 3435 3715 3450 3735
rect 3400 3700 3450 3715
rect 3550 4185 3600 4200
rect 3550 4165 3565 4185
rect 3585 4165 3600 4185
rect 3550 4135 3600 4165
rect 3550 4115 3565 4135
rect 3585 4115 3600 4135
rect 3550 4085 3600 4115
rect 3550 4065 3565 4085
rect 3585 4065 3600 4085
rect 3550 4035 3600 4065
rect 3550 4015 3565 4035
rect 3585 4015 3600 4035
rect 3550 3985 3600 4015
rect 3550 3965 3565 3985
rect 3585 3965 3600 3985
rect 3550 3935 3600 3965
rect 3550 3915 3565 3935
rect 3585 3915 3600 3935
rect 3550 3885 3600 3915
rect 3550 3865 3565 3885
rect 3585 3865 3600 3885
rect 3550 3835 3600 3865
rect 3550 3815 3565 3835
rect 3585 3815 3600 3835
rect 3550 3785 3600 3815
rect 3550 3765 3565 3785
rect 3585 3765 3600 3785
rect 3550 3735 3600 3765
rect 3550 3715 3565 3735
rect 3585 3715 3600 3735
rect 3550 3700 3600 3715
rect 4150 4185 4200 4200
rect 4150 4165 4165 4185
rect 4185 4165 4200 4185
rect 4150 4135 4200 4165
rect 4150 4115 4165 4135
rect 4185 4115 4200 4135
rect 4150 4085 4200 4115
rect 4150 4065 4165 4085
rect 4185 4065 4200 4085
rect 4150 4035 4200 4065
rect 4150 4015 4165 4035
rect 4185 4015 4200 4035
rect 4150 3985 4200 4015
rect 4150 3965 4165 3985
rect 4185 3965 4200 3985
rect 4150 3935 4200 3965
rect 4150 3915 4165 3935
rect 4185 3915 4200 3935
rect 4150 3885 4200 3915
rect 4150 3865 4165 3885
rect 4185 3865 4200 3885
rect 4150 3835 4200 3865
rect 4150 3815 4165 3835
rect 4185 3815 4200 3835
rect 4150 3785 4200 3815
rect 4150 3765 4165 3785
rect 4185 3765 4200 3785
rect 4150 3735 4200 3765
rect 4150 3715 4165 3735
rect 4185 3715 4200 3735
rect 4150 3700 4200 3715
rect 4750 4185 4800 4200
rect 4750 4165 4765 4185
rect 4785 4165 4800 4185
rect 4750 4135 4800 4165
rect 4750 4115 4765 4135
rect 4785 4115 4800 4135
rect 4750 4085 4800 4115
rect 4750 4065 4765 4085
rect 4785 4065 4800 4085
rect 4750 4035 4800 4065
rect 4750 4015 4765 4035
rect 4785 4015 4800 4035
rect 4750 3985 4800 4015
rect 4750 3965 4765 3985
rect 4785 3965 4800 3985
rect 4750 3935 4800 3965
rect 4750 3915 4765 3935
rect 4785 3915 4800 3935
rect 4750 3885 4800 3915
rect 4750 3865 4765 3885
rect 4785 3865 4800 3885
rect 4750 3835 4800 3865
rect 4750 3815 4765 3835
rect 4785 3815 4800 3835
rect 4750 3785 4800 3815
rect 4750 3765 4765 3785
rect 4785 3765 4800 3785
rect 4750 3735 4800 3765
rect 4750 3715 4765 3735
rect 4785 3715 4800 3735
rect 4750 3700 4800 3715
rect 4900 4185 4950 4200
rect 4900 4165 4915 4185
rect 4935 4165 4950 4185
rect 4900 4135 4950 4165
rect 4900 4115 4915 4135
rect 4935 4115 4950 4135
rect 4900 4085 4950 4115
rect 4900 4065 4915 4085
rect 4935 4065 4950 4085
rect 4900 4035 4950 4065
rect 4900 4015 4915 4035
rect 4935 4015 4950 4035
rect 4900 3985 4950 4015
rect 4900 3965 4915 3985
rect 4935 3965 4950 3985
rect 4900 3935 4950 3965
rect 4900 3915 4915 3935
rect 4935 3915 4950 3935
rect 4900 3885 4950 3915
rect 4900 3865 4915 3885
rect 4935 3865 4950 3885
rect 4900 3835 4950 3865
rect 4900 3815 4915 3835
rect 4935 3815 4950 3835
rect 4900 3785 4950 3815
rect 4900 3765 4915 3785
rect 4935 3765 4950 3785
rect 4900 3735 4950 3765
rect 4900 3715 4915 3735
rect 4935 3715 4950 3735
rect 4900 3700 4950 3715
rect 5050 4185 5100 4200
rect 5050 4165 5065 4185
rect 5085 4165 5100 4185
rect 5050 4135 5100 4165
rect 5050 4115 5065 4135
rect 5085 4115 5100 4135
rect 5050 4085 5100 4115
rect 5050 4065 5065 4085
rect 5085 4065 5100 4085
rect 5050 4035 5100 4065
rect 5050 4015 5065 4035
rect 5085 4015 5100 4035
rect 5050 3985 5100 4015
rect 5050 3965 5065 3985
rect 5085 3965 5100 3985
rect 5050 3935 5100 3965
rect 5050 3915 5065 3935
rect 5085 3915 5100 3935
rect 5050 3885 5100 3915
rect 5050 3865 5065 3885
rect 5085 3865 5100 3885
rect 5050 3835 5100 3865
rect 5050 3815 5065 3835
rect 5085 3815 5100 3835
rect 5050 3785 5100 3815
rect 5050 3765 5065 3785
rect 5085 3765 5100 3785
rect 5050 3735 5100 3765
rect 5050 3715 5065 3735
rect 5085 3715 5100 3735
rect 5050 3700 5100 3715
rect 5200 4185 5250 4200
rect 5200 4165 5215 4185
rect 5235 4165 5250 4185
rect 5200 4135 5250 4165
rect 5200 4115 5215 4135
rect 5235 4115 5250 4135
rect 5200 4085 5250 4115
rect 5200 4065 5215 4085
rect 5235 4065 5250 4085
rect 5200 4035 5250 4065
rect 5200 4015 5215 4035
rect 5235 4015 5250 4035
rect 5200 3985 5250 4015
rect 5200 3965 5215 3985
rect 5235 3965 5250 3985
rect 5200 3935 5250 3965
rect 5200 3915 5215 3935
rect 5235 3915 5250 3935
rect 5200 3885 5250 3915
rect 5200 3865 5215 3885
rect 5235 3865 5250 3885
rect 5200 3835 5250 3865
rect 5200 3815 5215 3835
rect 5235 3815 5250 3835
rect 5200 3785 5250 3815
rect 5200 3765 5215 3785
rect 5235 3765 5250 3785
rect 5200 3735 5250 3765
rect 5200 3715 5215 3735
rect 5235 3715 5250 3735
rect 5200 3700 5250 3715
rect 5350 4185 5400 4200
rect 5350 4165 5365 4185
rect 5385 4165 5400 4185
rect 5350 4135 5400 4165
rect 5350 4115 5365 4135
rect 5385 4115 5400 4135
rect 5350 4085 5400 4115
rect 5350 4065 5365 4085
rect 5385 4065 5400 4085
rect 5350 4035 5400 4065
rect 5350 4015 5365 4035
rect 5385 4015 5400 4035
rect 5350 3985 5400 4015
rect 5350 3965 5365 3985
rect 5385 3965 5400 3985
rect 5350 3935 5400 3965
rect 5350 3915 5365 3935
rect 5385 3915 5400 3935
rect 5350 3885 5400 3915
rect 5350 3865 5365 3885
rect 5385 3865 5400 3885
rect 5350 3835 5400 3865
rect 5350 3815 5365 3835
rect 5385 3815 5400 3835
rect 5350 3785 5400 3815
rect 5350 3765 5365 3785
rect 5385 3765 5400 3785
rect 5350 3735 5400 3765
rect 5350 3715 5365 3735
rect 5385 3715 5400 3735
rect 5350 3700 5400 3715
rect 5500 4185 5550 4200
rect 5500 4165 5515 4185
rect 5535 4165 5550 4185
rect 5500 4135 5550 4165
rect 5500 4115 5515 4135
rect 5535 4115 5550 4135
rect 5500 4085 5550 4115
rect 5500 4065 5515 4085
rect 5535 4065 5550 4085
rect 5500 4035 5550 4065
rect 5500 4015 5515 4035
rect 5535 4015 5550 4035
rect 5500 3985 5550 4015
rect 5500 3965 5515 3985
rect 5535 3965 5550 3985
rect 5500 3935 5550 3965
rect 5500 3915 5515 3935
rect 5535 3915 5550 3935
rect 5500 3885 5550 3915
rect 5500 3865 5515 3885
rect 5535 3865 5550 3885
rect 5500 3835 5550 3865
rect 5500 3815 5515 3835
rect 5535 3815 5550 3835
rect 5500 3785 5550 3815
rect 5500 3765 5515 3785
rect 5535 3765 5550 3785
rect 5500 3735 5550 3765
rect 5500 3715 5515 3735
rect 5535 3715 5550 3735
rect 5500 3700 5550 3715
rect 5650 4185 5700 4200
rect 5650 4165 5665 4185
rect 5685 4165 5700 4185
rect 5650 4135 5700 4165
rect 5650 4115 5665 4135
rect 5685 4115 5700 4135
rect 5650 4085 5700 4115
rect 5650 4065 5665 4085
rect 5685 4065 5700 4085
rect 5650 4035 5700 4065
rect 5650 4015 5665 4035
rect 5685 4015 5700 4035
rect 5650 3985 5700 4015
rect 5650 3965 5665 3985
rect 5685 3965 5700 3985
rect 5650 3935 5700 3965
rect 5650 3915 5665 3935
rect 5685 3915 5700 3935
rect 5650 3885 5700 3915
rect 5650 3865 5665 3885
rect 5685 3865 5700 3885
rect 5650 3835 5700 3865
rect 5650 3815 5665 3835
rect 5685 3815 5700 3835
rect 5650 3785 5700 3815
rect 5650 3765 5665 3785
rect 5685 3765 5700 3785
rect 5650 3735 5700 3765
rect 5650 3715 5665 3735
rect 5685 3715 5700 3735
rect 5650 3700 5700 3715
rect 5800 4185 5850 4200
rect 5800 4165 5815 4185
rect 5835 4165 5850 4185
rect 5800 4135 5850 4165
rect 5800 4115 5815 4135
rect 5835 4115 5850 4135
rect 5800 4085 5850 4115
rect 5800 4065 5815 4085
rect 5835 4065 5850 4085
rect 5800 4035 5850 4065
rect 5800 4015 5815 4035
rect 5835 4015 5850 4035
rect 5800 3985 5850 4015
rect 5800 3965 5815 3985
rect 5835 3965 5850 3985
rect 5800 3935 5850 3965
rect 5800 3915 5815 3935
rect 5835 3915 5850 3935
rect 5800 3885 5850 3915
rect 5800 3865 5815 3885
rect 5835 3865 5850 3885
rect 5800 3835 5850 3865
rect 5800 3815 5815 3835
rect 5835 3815 5850 3835
rect 5800 3785 5850 3815
rect 5800 3765 5815 3785
rect 5835 3765 5850 3785
rect 5800 3735 5850 3765
rect 5800 3715 5815 3735
rect 5835 3715 5850 3735
rect 5800 3700 5850 3715
rect 5950 4185 6000 4200
rect 5950 4165 5965 4185
rect 5985 4165 6000 4185
rect 5950 4135 6000 4165
rect 5950 4115 5965 4135
rect 5985 4115 6000 4135
rect 5950 4085 6000 4115
rect 5950 4065 5965 4085
rect 5985 4065 6000 4085
rect 5950 4035 6000 4065
rect 5950 4015 5965 4035
rect 5985 4015 6000 4035
rect 5950 3985 6000 4015
rect 5950 3965 5965 3985
rect 5985 3965 6000 3985
rect 5950 3935 6000 3965
rect 5950 3915 5965 3935
rect 5985 3915 6000 3935
rect 5950 3885 6000 3915
rect 5950 3865 5965 3885
rect 5985 3865 6000 3885
rect 5950 3835 6000 3865
rect 5950 3815 5965 3835
rect 5985 3815 6000 3835
rect 5950 3785 6000 3815
rect 5950 3765 5965 3785
rect 5985 3765 6000 3785
rect 5950 3735 6000 3765
rect 5950 3715 5965 3735
rect 5985 3715 6000 3735
rect 5950 3700 6000 3715
rect 6100 4185 6150 4200
rect 6100 4165 6115 4185
rect 6135 4165 6150 4185
rect 6100 4135 6150 4165
rect 6100 4115 6115 4135
rect 6135 4115 6150 4135
rect 6100 4085 6150 4115
rect 6100 4065 6115 4085
rect 6135 4065 6150 4085
rect 6100 4035 6150 4065
rect 6100 4015 6115 4035
rect 6135 4015 6150 4035
rect 6100 3985 6150 4015
rect 6100 3965 6115 3985
rect 6135 3965 6150 3985
rect 6100 3935 6150 3965
rect 6100 3915 6115 3935
rect 6135 3915 6150 3935
rect 6100 3885 6150 3915
rect 6100 3865 6115 3885
rect 6135 3865 6150 3885
rect 6100 3835 6150 3865
rect 6100 3815 6115 3835
rect 6135 3815 6150 3835
rect 6100 3785 6150 3815
rect 6100 3765 6115 3785
rect 6135 3765 6150 3785
rect 6100 3735 6150 3765
rect 6100 3715 6115 3735
rect 6135 3715 6150 3735
rect 6100 3700 6150 3715
rect 6250 4185 6300 4200
rect 6250 4165 6265 4185
rect 6285 4165 6300 4185
rect 6250 4135 6300 4165
rect 6250 4115 6265 4135
rect 6285 4115 6300 4135
rect 6250 4085 6300 4115
rect 6250 4065 6265 4085
rect 6285 4065 6300 4085
rect 6250 4035 6300 4065
rect 6250 4015 6265 4035
rect 6285 4015 6300 4035
rect 6250 3985 6300 4015
rect 6250 3965 6265 3985
rect 6285 3965 6300 3985
rect 6250 3935 6300 3965
rect 6250 3915 6265 3935
rect 6285 3915 6300 3935
rect 6250 3885 6300 3915
rect 6250 3865 6265 3885
rect 6285 3865 6300 3885
rect 6250 3835 6300 3865
rect 6250 3815 6265 3835
rect 6285 3815 6300 3835
rect 6250 3785 6300 3815
rect 6250 3765 6265 3785
rect 6285 3765 6300 3785
rect 6250 3735 6300 3765
rect 6250 3715 6265 3735
rect 6285 3715 6300 3735
rect 6250 3700 6300 3715
rect 6400 4185 6450 4200
rect 6400 4165 6415 4185
rect 6435 4165 6450 4185
rect 6400 4135 6450 4165
rect 6400 4115 6415 4135
rect 6435 4115 6450 4135
rect 6400 4085 6450 4115
rect 6400 4065 6415 4085
rect 6435 4065 6450 4085
rect 6400 4035 6450 4065
rect 6400 4015 6415 4035
rect 6435 4015 6450 4035
rect 6400 3985 6450 4015
rect 6400 3965 6415 3985
rect 6435 3965 6450 3985
rect 6400 3935 6450 3965
rect 6400 3915 6415 3935
rect 6435 3915 6450 3935
rect 6400 3885 6450 3915
rect 6400 3865 6415 3885
rect 6435 3865 6450 3885
rect 6400 3835 6450 3865
rect 6400 3815 6415 3835
rect 6435 3815 6450 3835
rect 6400 3785 6450 3815
rect 6400 3765 6415 3785
rect 6435 3765 6450 3785
rect 6400 3735 6450 3765
rect 6400 3715 6415 3735
rect 6435 3715 6450 3735
rect 6400 3700 6450 3715
rect 6550 4185 6600 4200
rect 6550 4165 6565 4185
rect 6585 4165 6600 4185
rect 6550 4135 6600 4165
rect 6550 4115 6565 4135
rect 6585 4115 6600 4135
rect 6550 4085 6600 4115
rect 6550 4065 6565 4085
rect 6585 4065 6600 4085
rect 6550 4035 6600 4065
rect 6550 4015 6565 4035
rect 6585 4015 6600 4035
rect 6550 3985 6600 4015
rect 6550 3965 6565 3985
rect 6585 3965 6600 3985
rect 6550 3935 6600 3965
rect 6550 3915 6565 3935
rect 6585 3915 6600 3935
rect 6550 3885 6600 3915
rect 6550 3865 6565 3885
rect 6585 3865 6600 3885
rect 6550 3835 6600 3865
rect 6550 3815 6565 3835
rect 6585 3815 6600 3835
rect 6550 3785 6600 3815
rect 6550 3765 6565 3785
rect 6585 3765 6600 3785
rect 6550 3735 6600 3765
rect 6550 3715 6565 3735
rect 6585 3715 6600 3735
rect 6550 3700 6600 3715
rect 6700 4185 6750 4200
rect 6700 4165 6715 4185
rect 6735 4165 6750 4185
rect 6700 4135 6750 4165
rect 6700 4115 6715 4135
rect 6735 4115 6750 4135
rect 6700 4085 6750 4115
rect 6700 4065 6715 4085
rect 6735 4065 6750 4085
rect 6700 4035 6750 4065
rect 6700 4015 6715 4035
rect 6735 4015 6750 4035
rect 6700 3985 6750 4015
rect 6700 3965 6715 3985
rect 6735 3965 6750 3985
rect 6700 3935 6750 3965
rect 6700 3915 6715 3935
rect 6735 3915 6750 3935
rect 6700 3885 6750 3915
rect 6700 3865 6715 3885
rect 6735 3865 6750 3885
rect 6700 3835 6750 3865
rect 6700 3815 6715 3835
rect 6735 3815 6750 3835
rect 6700 3785 6750 3815
rect 6700 3765 6715 3785
rect 6735 3765 6750 3785
rect 6700 3735 6750 3765
rect 6700 3715 6715 3735
rect 6735 3715 6750 3735
rect 6700 3700 6750 3715
rect 6850 4185 6900 4200
rect 6850 4165 6865 4185
rect 6885 4165 6900 4185
rect 6850 4135 6900 4165
rect 6850 4115 6865 4135
rect 6885 4115 6900 4135
rect 6850 4085 6900 4115
rect 6850 4065 6865 4085
rect 6885 4065 6900 4085
rect 6850 4035 6900 4065
rect 6850 4015 6865 4035
rect 6885 4015 6900 4035
rect 6850 3985 6900 4015
rect 6850 3965 6865 3985
rect 6885 3965 6900 3985
rect 6850 3935 6900 3965
rect 6850 3915 6865 3935
rect 6885 3915 6900 3935
rect 6850 3885 6900 3915
rect 6850 3865 6865 3885
rect 6885 3865 6900 3885
rect 6850 3835 6900 3865
rect 6850 3815 6865 3835
rect 6885 3815 6900 3835
rect 6850 3785 6900 3815
rect 6850 3765 6865 3785
rect 6885 3765 6900 3785
rect 6850 3735 6900 3765
rect 6850 3715 6865 3735
rect 6885 3715 6900 3735
rect 6850 3700 6900 3715
rect 7000 4185 7050 4200
rect 7000 4165 7015 4185
rect 7035 4165 7050 4185
rect 7000 4135 7050 4165
rect 7000 4115 7015 4135
rect 7035 4115 7050 4135
rect 7000 4085 7050 4115
rect 7000 4065 7015 4085
rect 7035 4065 7050 4085
rect 7000 4035 7050 4065
rect 7000 4015 7015 4035
rect 7035 4015 7050 4035
rect 7000 3985 7050 4015
rect 7000 3965 7015 3985
rect 7035 3965 7050 3985
rect 7000 3935 7050 3965
rect 7000 3915 7015 3935
rect 7035 3915 7050 3935
rect 7000 3885 7050 3915
rect 7000 3865 7015 3885
rect 7035 3865 7050 3885
rect 7000 3835 7050 3865
rect 7000 3815 7015 3835
rect 7035 3815 7050 3835
rect 7000 3785 7050 3815
rect 7000 3765 7015 3785
rect 7035 3765 7050 3785
rect 7000 3735 7050 3765
rect 7000 3715 7015 3735
rect 7035 3715 7050 3735
rect 7000 3700 7050 3715
rect 7150 4185 7200 4200
rect 7150 4165 7165 4185
rect 7185 4165 7200 4185
rect 7150 4135 7200 4165
rect 7150 4115 7165 4135
rect 7185 4115 7200 4135
rect 7150 4085 7200 4115
rect 7150 4065 7165 4085
rect 7185 4065 7200 4085
rect 7150 4035 7200 4065
rect 7150 4015 7165 4035
rect 7185 4015 7200 4035
rect 7150 3985 7200 4015
rect 7150 3965 7165 3985
rect 7185 3965 7200 3985
rect 7150 3935 7200 3965
rect 7150 3915 7165 3935
rect 7185 3915 7200 3935
rect 7150 3885 7200 3915
rect 7150 3865 7165 3885
rect 7185 3865 7200 3885
rect 7150 3835 7200 3865
rect 7150 3815 7165 3835
rect 7185 3815 7200 3835
rect 7150 3785 7200 3815
rect 7150 3765 7165 3785
rect 7185 3765 7200 3785
rect 7150 3735 7200 3765
rect 7150 3715 7165 3735
rect 7185 3715 7200 3735
rect 7150 3700 7200 3715
rect 7300 4185 7350 4200
rect 7300 4165 7315 4185
rect 7335 4165 7350 4185
rect 7300 4135 7350 4165
rect 7300 4115 7315 4135
rect 7335 4115 7350 4135
rect 7300 4085 7350 4115
rect 7300 4065 7315 4085
rect 7335 4065 7350 4085
rect 7300 4035 7350 4065
rect 7300 4015 7315 4035
rect 7335 4015 7350 4035
rect 7300 3985 7350 4015
rect 7300 3965 7315 3985
rect 7335 3965 7350 3985
rect 7300 3935 7350 3965
rect 7300 3915 7315 3935
rect 7335 3915 7350 3935
rect 7300 3885 7350 3915
rect 7300 3865 7315 3885
rect 7335 3865 7350 3885
rect 7300 3835 7350 3865
rect 7300 3815 7315 3835
rect 7335 3815 7350 3835
rect 7300 3785 7350 3815
rect 7300 3765 7315 3785
rect 7335 3765 7350 3785
rect 7300 3735 7350 3765
rect 7300 3715 7315 3735
rect 7335 3715 7350 3735
rect 7300 3700 7350 3715
rect 7450 4185 7500 4200
rect 7450 4165 7465 4185
rect 7485 4165 7500 4185
rect 7450 4135 7500 4165
rect 7450 4115 7465 4135
rect 7485 4115 7500 4135
rect 7450 4085 7500 4115
rect 7450 4065 7465 4085
rect 7485 4065 7500 4085
rect 7450 4035 7500 4065
rect 7450 4015 7465 4035
rect 7485 4015 7500 4035
rect 7450 3985 7500 4015
rect 7450 3965 7465 3985
rect 7485 3965 7500 3985
rect 7450 3935 7500 3965
rect 7450 3915 7465 3935
rect 7485 3915 7500 3935
rect 7450 3885 7500 3915
rect 7450 3865 7465 3885
rect 7485 3865 7500 3885
rect 7450 3835 7500 3865
rect 7450 3815 7465 3835
rect 7485 3815 7500 3835
rect 7450 3785 7500 3815
rect 7450 3765 7465 3785
rect 7485 3765 7500 3785
rect 7450 3735 7500 3765
rect 7450 3715 7465 3735
rect 7485 3715 7500 3735
rect 7450 3700 7500 3715
rect 7600 4185 7650 4200
rect 7600 4165 7615 4185
rect 7635 4165 7650 4185
rect 7600 4135 7650 4165
rect 7600 4115 7615 4135
rect 7635 4115 7650 4135
rect 7600 4085 7650 4115
rect 7600 4065 7615 4085
rect 7635 4065 7650 4085
rect 7600 4035 7650 4065
rect 7600 4015 7615 4035
rect 7635 4015 7650 4035
rect 7600 3985 7650 4015
rect 7600 3965 7615 3985
rect 7635 3965 7650 3985
rect 7600 3935 7650 3965
rect 7600 3915 7615 3935
rect 7635 3915 7650 3935
rect 7600 3885 7650 3915
rect 7600 3865 7615 3885
rect 7635 3865 7650 3885
rect 7600 3835 7650 3865
rect 7600 3815 7615 3835
rect 7635 3815 7650 3835
rect 7600 3785 7650 3815
rect 7600 3765 7615 3785
rect 7635 3765 7650 3785
rect 7600 3735 7650 3765
rect 7600 3715 7615 3735
rect 7635 3715 7650 3735
rect 7600 3700 7650 3715
rect 7750 4185 7800 4200
rect 7750 4165 7765 4185
rect 7785 4165 7800 4185
rect 7750 4135 7800 4165
rect 7750 4115 7765 4135
rect 7785 4115 7800 4135
rect 7750 4085 7800 4115
rect 7750 4065 7765 4085
rect 7785 4065 7800 4085
rect 7750 4035 7800 4065
rect 7750 4015 7765 4035
rect 7785 4015 7800 4035
rect 7750 3985 7800 4015
rect 7750 3965 7765 3985
rect 7785 3965 7800 3985
rect 7750 3935 7800 3965
rect 7750 3915 7765 3935
rect 7785 3915 7800 3935
rect 7750 3885 7800 3915
rect 7750 3865 7765 3885
rect 7785 3865 7800 3885
rect 7750 3835 7800 3865
rect 7750 3815 7765 3835
rect 7785 3815 7800 3835
rect 7750 3785 7800 3815
rect 7750 3765 7765 3785
rect 7785 3765 7800 3785
rect 7750 3735 7800 3765
rect 7750 3715 7765 3735
rect 7785 3715 7800 3735
rect 7750 3700 7800 3715
rect 8350 4185 8400 4200
rect 8350 4165 8365 4185
rect 8385 4165 8400 4185
rect 8350 4135 8400 4165
rect 8350 4115 8365 4135
rect 8385 4115 8400 4135
rect 8350 4085 8400 4115
rect 8350 4065 8365 4085
rect 8385 4065 8400 4085
rect 8350 4035 8400 4065
rect 8350 4015 8365 4035
rect 8385 4015 8400 4035
rect 8350 3985 8400 4015
rect 8350 3965 8365 3985
rect 8385 3965 8400 3985
rect 8350 3935 8400 3965
rect 8350 3915 8365 3935
rect 8385 3915 8400 3935
rect 8350 3885 8400 3915
rect 8350 3865 8365 3885
rect 8385 3865 8400 3885
rect 8350 3835 8400 3865
rect 8350 3815 8365 3835
rect 8385 3815 8400 3835
rect 8350 3785 8400 3815
rect 8350 3765 8365 3785
rect 8385 3765 8400 3785
rect 8350 3735 8400 3765
rect 8350 3715 8365 3735
rect 8385 3715 8400 3735
rect 8350 3700 8400 3715
rect 8500 4185 8550 4200
rect 8500 4165 8515 4185
rect 8535 4165 8550 4185
rect 8500 4135 8550 4165
rect 8500 4115 8515 4135
rect 8535 4115 8550 4135
rect 8500 4085 8550 4115
rect 8500 4065 8515 4085
rect 8535 4065 8550 4085
rect 8500 4035 8550 4065
rect 8500 4015 8515 4035
rect 8535 4015 8550 4035
rect 8500 3985 8550 4015
rect 8500 3965 8515 3985
rect 8535 3965 8550 3985
rect 8500 3935 8550 3965
rect 8500 3915 8515 3935
rect 8535 3915 8550 3935
rect 8500 3885 8550 3915
rect 8500 3865 8515 3885
rect 8535 3865 8550 3885
rect 8500 3835 8550 3865
rect 8500 3815 8515 3835
rect 8535 3815 8550 3835
rect 8500 3785 8550 3815
rect 8500 3765 8515 3785
rect 8535 3765 8550 3785
rect 8500 3735 8550 3765
rect 8500 3715 8515 3735
rect 8535 3715 8550 3735
rect 8500 3650 8550 3715
rect 8650 4185 8700 4200
rect 8650 4165 8665 4185
rect 8685 4165 8700 4185
rect 8650 4135 8700 4165
rect 8650 4115 8665 4135
rect 8685 4115 8700 4135
rect 8650 4085 8700 4115
rect 8650 4065 8665 4085
rect 8685 4065 8700 4085
rect 8650 4035 8700 4065
rect 8650 4015 8665 4035
rect 8685 4015 8700 4035
rect 8650 3985 8700 4015
rect 8650 3965 8665 3985
rect 8685 3965 8700 3985
rect 8650 3935 8700 3965
rect 8650 3915 8665 3935
rect 8685 3915 8700 3935
rect 8650 3885 8700 3915
rect 8650 3865 8665 3885
rect 8685 3865 8700 3885
rect 8650 3835 8700 3865
rect 8650 3815 8665 3835
rect 8685 3815 8700 3835
rect 8650 3785 8700 3815
rect 8650 3765 8665 3785
rect 8685 3765 8700 3785
rect 8650 3735 8700 3765
rect 8650 3715 8665 3735
rect 8685 3715 8700 3735
rect 8650 3700 8700 3715
rect 8800 4185 8850 4200
rect 8800 4165 8815 4185
rect 8835 4165 8850 4185
rect 8800 4135 8850 4165
rect 8800 4115 8815 4135
rect 8835 4115 8850 4135
rect 8800 4085 8850 4115
rect 8800 4065 8815 4085
rect 8835 4065 8850 4085
rect 8800 4035 8850 4065
rect 8800 4015 8815 4035
rect 8835 4015 8850 4035
rect 8800 3985 8850 4015
rect 8800 3965 8815 3985
rect 8835 3965 8850 3985
rect 8800 3935 8850 3965
rect 8800 3915 8815 3935
rect 8835 3915 8850 3935
rect 8800 3885 8850 3915
rect 8800 3865 8815 3885
rect 8835 3865 8850 3885
rect 8800 3835 8850 3865
rect 8800 3815 8815 3835
rect 8835 3815 8850 3835
rect 8800 3785 8850 3815
rect 8800 3765 8815 3785
rect 8835 3765 8850 3785
rect 8800 3735 8850 3765
rect 8800 3715 8815 3735
rect 8835 3715 8850 3735
rect 8800 3650 8850 3715
rect 8950 4185 9000 4200
rect 8950 4165 8965 4185
rect 8985 4165 9000 4185
rect 8950 4135 9000 4165
rect 8950 4115 8965 4135
rect 8985 4115 9000 4135
rect 8950 4085 9000 4115
rect 8950 4065 8965 4085
rect 8985 4065 9000 4085
rect 8950 4035 9000 4065
rect 8950 4015 8965 4035
rect 8985 4015 9000 4035
rect 8950 3985 9000 4015
rect 8950 3965 8965 3985
rect 8985 3965 9000 3985
rect 8950 3935 9000 3965
rect 8950 3915 8965 3935
rect 8985 3915 9000 3935
rect 8950 3885 9000 3915
rect 8950 3865 8965 3885
rect 8985 3865 9000 3885
rect 8950 3835 9000 3865
rect 8950 3815 8965 3835
rect 8985 3815 9000 3835
rect 8950 3785 9000 3815
rect 8950 3765 8965 3785
rect 8985 3765 9000 3785
rect 8950 3735 9000 3765
rect 8950 3715 8965 3735
rect 8985 3715 9000 3735
rect 8950 3700 9000 3715
rect 9100 4185 9150 4200
rect 9100 4165 9115 4185
rect 9135 4165 9150 4185
rect 9100 4135 9150 4165
rect 9100 4115 9115 4135
rect 9135 4115 9150 4135
rect 9100 4085 9150 4115
rect 9100 4065 9115 4085
rect 9135 4065 9150 4085
rect 9100 4035 9150 4065
rect 9100 4015 9115 4035
rect 9135 4015 9150 4035
rect 9100 3985 9150 4015
rect 9100 3965 9115 3985
rect 9135 3965 9150 3985
rect 9100 3935 9150 3965
rect 9100 3915 9115 3935
rect 9135 3915 9150 3935
rect 9100 3885 9150 3915
rect 9100 3865 9115 3885
rect 9135 3865 9150 3885
rect 9100 3835 9150 3865
rect 9100 3815 9115 3835
rect 9135 3815 9150 3835
rect 9100 3785 9150 3815
rect 9100 3765 9115 3785
rect 9135 3765 9150 3785
rect 9100 3735 9150 3765
rect 9100 3715 9115 3735
rect 9135 3715 9150 3735
rect 9100 3650 9150 3715
rect 9250 4185 9300 4200
rect 9250 4165 9265 4185
rect 9285 4165 9300 4185
rect 9250 4135 9300 4165
rect 9250 4115 9265 4135
rect 9285 4115 9300 4135
rect 9250 4085 9300 4115
rect 9250 4065 9265 4085
rect 9285 4065 9300 4085
rect 9250 4035 9300 4065
rect 9250 4015 9265 4035
rect 9285 4015 9300 4035
rect 9250 3985 9300 4015
rect 9250 3965 9265 3985
rect 9285 3965 9300 3985
rect 9250 3935 9300 3965
rect 9250 3915 9265 3935
rect 9285 3915 9300 3935
rect 9250 3885 9300 3915
rect 9250 3865 9265 3885
rect 9285 3865 9300 3885
rect 9250 3835 9300 3865
rect 9250 3815 9265 3835
rect 9285 3815 9300 3835
rect 9250 3785 9300 3815
rect 9250 3765 9265 3785
rect 9285 3765 9300 3785
rect 9250 3735 9300 3765
rect 9250 3715 9265 3735
rect 9285 3715 9300 3735
rect 9250 3700 9300 3715
rect 9400 4185 9450 4200
rect 9400 4165 9415 4185
rect 9435 4165 9450 4185
rect 9400 4135 9450 4165
rect 9400 4115 9415 4135
rect 9435 4115 9450 4135
rect 9400 4085 9450 4115
rect 9400 4065 9415 4085
rect 9435 4065 9450 4085
rect 9400 4035 9450 4065
rect 9400 4015 9415 4035
rect 9435 4015 9450 4035
rect 9400 3985 9450 4015
rect 9400 3965 9415 3985
rect 9435 3965 9450 3985
rect 9400 3935 9450 3965
rect 9400 3915 9415 3935
rect 9435 3915 9450 3935
rect 9400 3885 9450 3915
rect 9400 3865 9415 3885
rect 9435 3865 9450 3885
rect 9400 3835 9450 3865
rect 9400 3815 9415 3835
rect 9435 3815 9450 3835
rect 9400 3785 9450 3815
rect 9400 3765 9415 3785
rect 9435 3765 9450 3785
rect 9400 3735 9450 3765
rect 9400 3715 9415 3735
rect 9435 3715 9450 3735
rect 9400 3650 9450 3715
rect 9550 4185 9600 4200
rect 9550 4165 9565 4185
rect 9585 4165 9600 4185
rect 9550 4135 9600 4165
rect 9550 4115 9565 4135
rect 9585 4115 9600 4135
rect 9550 4085 9600 4115
rect 9550 4065 9565 4085
rect 9585 4065 9600 4085
rect 9550 4035 9600 4065
rect 9550 4015 9565 4035
rect 9585 4015 9600 4035
rect 9550 3985 9600 4015
rect 9550 3965 9565 3985
rect 9585 3965 9600 3985
rect 9550 3935 9600 3965
rect 9550 3915 9565 3935
rect 9585 3915 9600 3935
rect 9550 3885 9600 3915
rect 9550 3865 9565 3885
rect 9585 3865 9600 3885
rect 9550 3835 9600 3865
rect 9550 3815 9565 3835
rect 9585 3815 9600 3835
rect 9550 3785 9600 3815
rect 9550 3765 9565 3785
rect 9585 3765 9600 3785
rect 9550 3735 9600 3765
rect 9550 3715 9565 3735
rect 9585 3715 9600 3735
rect 9550 3700 9600 3715
rect 9700 4185 9750 4200
rect 9700 4165 9715 4185
rect 9735 4165 9750 4185
rect 9700 4135 9750 4165
rect 9700 4115 9715 4135
rect 9735 4115 9750 4135
rect 9700 4085 9750 4115
rect 9700 4065 9715 4085
rect 9735 4065 9750 4085
rect 9700 4035 9750 4065
rect 9700 4015 9715 4035
rect 9735 4015 9750 4035
rect 9700 3985 9750 4015
rect 9700 3965 9715 3985
rect 9735 3965 9750 3985
rect 9700 3935 9750 3965
rect 9700 3915 9715 3935
rect 9735 3915 9750 3935
rect 9700 3885 9750 3915
rect 9700 3865 9715 3885
rect 9735 3865 9750 3885
rect 9700 3835 9750 3865
rect 9700 3815 9715 3835
rect 9735 3815 9750 3835
rect 9700 3785 9750 3815
rect 9700 3765 9715 3785
rect 9735 3765 9750 3785
rect 9700 3735 9750 3765
rect 9700 3715 9715 3735
rect 9735 3715 9750 3735
rect 9700 3650 9750 3715
rect 9850 4185 9900 4200
rect 9850 4165 9865 4185
rect 9885 4165 9900 4185
rect 9850 4135 9900 4165
rect 9850 4115 9865 4135
rect 9885 4115 9900 4135
rect 9850 4085 9900 4115
rect 9850 4065 9865 4085
rect 9885 4065 9900 4085
rect 9850 4035 9900 4065
rect 9850 4015 9865 4035
rect 9885 4015 9900 4035
rect 9850 3985 9900 4015
rect 9850 3965 9865 3985
rect 9885 3965 9900 3985
rect 9850 3935 9900 3965
rect 9850 3915 9865 3935
rect 9885 3915 9900 3935
rect 9850 3885 9900 3915
rect 9850 3865 9865 3885
rect 9885 3865 9900 3885
rect 9850 3835 9900 3865
rect 9850 3815 9865 3835
rect 9885 3815 9900 3835
rect 9850 3785 9900 3815
rect 9850 3765 9865 3785
rect 9885 3765 9900 3785
rect 9850 3735 9900 3765
rect 9850 3715 9865 3735
rect 9885 3715 9900 3735
rect 9850 3700 9900 3715
rect 10000 4185 10050 4200
rect 10000 4165 10015 4185
rect 10035 4165 10050 4185
rect 10000 4135 10050 4165
rect 10000 4115 10015 4135
rect 10035 4115 10050 4135
rect 10000 4085 10050 4115
rect 10000 4065 10015 4085
rect 10035 4065 10050 4085
rect 10000 4035 10050 4065
rect 10000 4015 10015 4035
rect 10035 4015 10050 4035
rect 10000 3985 10050 4015
rect 10000 3965 10015 3985
rect 10035 3965 10050 3985
rect 10000 3935 10050 3965
rect 10000 3915 10015 3935
rect 10035 3915 10050 3935
rect 10000 3885 10050 3915
rect 10000 3865 10015 3885
rect 10035 3865 10050 3885
rect 10000 3835 10050 3865
rect 10000 3815 10015 3835
rect 10035 3815 10050 3835
rect 10000 3785 10050 3815
rect 10000 3765 10015 3785
rect 10035 3765 10050 3785
rect 10000 3735 10050 3765
rect 10000 3715 10015 3735
rect 10035 3715 10050 3735
rect 10000 3650 10050 3715
rect 10150 4185 10200 4200
rect 10150 4165 10165 4185
rect 10185 4165 10200 4185
rect 10150 4135 10200 4165
rect 10150 4115 10165 4135
rect 10185 4115 10200 4135
rect 10150 4085 10200 4115
rect 10150 4065 10165 4085
rect 10185 4065 10200 4085
rect 10150 4035 10200 4065
rect 10150 4015 10165 4035
rect 10185 4015 10200 4035
rect 10150 3985 10200 4015
rect 10150 3965 10165 3985
rect 10185 3965 10200 3985
rect 10150 3935 10200 3965
rect 10150 3915 10165 3935
rect 10185 3915 10200 3935
rect 10150 3885 10200 3915
rect 10150 3865 10165 3885
rect 10185 3865 10200 3885
rect 10150 3835 10200 3865
rect 10150 3815 10165 3835
rect 10185 3815 10200 3835
rect 10150 3785 10200 3815
rect 10150 3765 10165 3785
rect 10185 3765 10200 3785
rect 10150 3735 10200 3765
rect 10150 3715 10165 3735
rect 10185 3715 10200 3735
rect 10150 3700 10200 3715
rect 10300 4185 10350 4200
rect 10300 4165 10315 4185
rect 10335 4165 10350 4185
rect 10300 4135 10350 4165
rect 10300 4115 10315 4135
rect 10335 4115 10350 4135
rect 10300 4085 10350 4115
rect 10300 4065 10315 4085
rect 10335 4065 10350 4085
rect 10300 4035 10350 4065
rect 10300 4015 10315 4035
rect 10335 4015 10350 4035
rect 10300 3985 10350 4015
rect 10300 3965 10315 3985
rect 10335 3965 10350 3985
rect 10300 3935 10350 3965
rect 10300 3915 10315 3935
rect 10335 3915 10350 3935
rect 10300 3885 10350 3915
rect 10300 3865 10315 3885
rect 10335 3865 10350 3885
rect 10300 3835 10350 3865
rect 10300 3815 10315 3835
rect 10335 3815 10350 3835
rect 10300 3785 10350 3815
rect 10300 3765 10315 3785
rect 10335 3765 10350 3785
rect 10300 3735 10350 3765
rect 10300 3715 10315 3735
rect 10335 3715 10350 3735
rect 10300 3650 10350 3715
rect 10450 4185 10500 4200
rect 10450 4165 10465 4185
rect 10485 4165 10500 4185
rect 10450 4135 10500 4165
rect 10450 4115 10465 4135
rect 10485 4115 10500 4135
rect 10450 4085 10500 4115
rect 10450 4065 10465 4085
rect 10485 4065 10500 4085
rect 10450 4035 10500 4065
rect 10450 4015 10465 4035
rect 10485 4015 10500 4035
rect 10450 3985 10500 4015
rect 10450 3965 10465 3985
rect 10485 3965 10500 3985
rect 10450 3935 10500 3965
rect 10450 3915 10465 3935
rect 10485 3915 10500 3935
rect 10450 3885 10500 3915
rect 10450 3865 10465 3885
rect 10485 3865 10500 3885
rect 10450 3835 10500 3865
rect 10450 3815 10465 3835
rect 10485 3815 10500 3835
rect 10450 3785 10500 3815
rect 10450 3765 10465 3785
rect 10485 3765 10500 3785
rect 10450 3735 10500 3765
rect 10450 3715 10465 3735
rect 10485 3715 10500 3735
rect 10450 3700 10500 3715
rect 10600 4185 10650 4200
rect 10600 4165 10615 4185
rect 10635 4165 10650 4185
rect 10600 4135 10650 4165
rect 10600 4115 10615 4135
rect 10635 4115 10650 4135
rect 10600 4085 10650 4115
rect 10600 4065 10615 4085
rect 10635 4065 10650 4085
rect 10600 4035 10650 4065
rect 10600 4015 10615 4035
rect 10635 4015 10650 4035
rect 10600 3985 10650 4015
rect 10600 3965 10615 3985
rect 10635 3965 10650 3985
rect 10600 3935 10650 3965
rect 10600 3915 10615 3935
rect 10635 3915 10650 3935
rect 10600 3885 10650 3915
rect 10600 3865 10615 3885
rect 10635 3865 10650 3885
rect 10600 3835 10650 3865
rect 10600 3815 10615 3835
rect 10635 3815 10650 3835
rect 10600 3785 10650 3815
rect 10600 3765 10615 3785
rect 10635 3765 10650 3785
rect 10600 3735 10650 3765
rect 10600 3715 10615 3735
rect 10635 3715 10650 3735
rect 10600 3650 10650 3715
rect 10750 4185 10800 4200
rect 10750 4165 10765 4185
rect 10785 4165 10800 4185
rect 10750 4135 10800 4165
rect 10750 4115 10765 4135
rect 10785 4115 10800 4135
rect 10750 4085 10800 4115
rect 10750 4065 10765 4085
rect 10785 4065 10800 4085
rect 10750 4035 10800 4065
rect 10750 4015 10765 4035
rect 10785 4015 10800 4035
rect 10750 3985 10800 4015
rect 10750 3965 10765 3985
rect 10785 3965 10800 3985
rect 10750 3935 10800 3965
rect 10750 3915 10765 3935
rect 10785 3915 10800 3935
rect 10750 3885 10800 3915
rect 10750 3865 10765 3885
rect 10785 3865 10800 3885
rect 10750 3835 10800 3865
rect 10750 3815 10765 3835
rect 10785 3815 10800 3835
rect 10750 3785 10800 3815
rect 10750 3765 10765 3785
rect 10785 3765 10800 3785
rect 10750 3735 10800 3765
rect 10750 3715 10765 3735
rect 10785 3715 10800 3735
rect 10750 3700 10800 3715
rect 11350 4185 11400 4200
rect 11350 4165 11365 4185
rect 11385 4165 11400 4185
rect 11350 4135 11400 4165
rect 11350 4115 11365 4135
rect 11385 4115 11400 4135
rect 11350 4085 11400 4115
rect 11350 4065 11365 4085
rect 11385 4065 11400 4085
rect 11350 4035 11400 4065
rect 11350 4015 11365 4035
rect 11385 4015 11400 4035
rect 11350 3985 11400 4015
rect 11350 3965 11365 3985
rect 11385 3965 11400 3985
rect 11350 3935 11400 3965
rect 11350 3915 11365 3935
rect 11385 3915 11400 3935
rect 11350 3885 11400 3915
rect 11350 3865 11365 3885
rect 11385 3865 11400 3885
rect 11350 3835 11400 3865
rect 11350 3815 11365 3835
rect 11385 3815 11400 3835
rect 11350 3785 11400 3815
rect 11350 3765 11365 3785
rect 11385 3765 11400 3785
rect 11350 3735 11400 3765
rect 11350 3715 11365 3735
rect 11385 3715 11400 3735
rect 11350 3700 11400 3715
rect 11950 4185 12000 4200
rect 11950 4165 11965 4185
rect 11985 4165 12000 4185
rect 11950 4135 12000 4165
rect 11950 4115 11965 4135
rect 11985 4115 12000 4135
rect 11950 4085 12000 4115
rect 11950 4065 11965 4085
rect 11985 4065 12000 4085
rect 11950 4035 12000 4065
rect 11950 4015 11965 4035
rect 11985 4015 12000 4035
rect 11950 3985 12000 4015
rect 11950 3965 11965 3985
rect 11985 3965 12000 3985
rect 11950 3935 12000 3965
rect 11950 3915 11965 3935
rect 11985 3915 12000 3935
rect 11950 3885 12000 3915
rect 11950 3865 11965 3885
rect 11985 3865 12000 3885
rect 11950 3835 12000 3865
rect 11950 3815 11965 3835
rect 11985 3815 12000 3835
rect 11950 3785 12000 3815
rect 11950 3765 11965 3785
rect 11985 3765 12000 3785
rect 11950 3735 12000 3765
rect 11950 3715 11965 3735
rect 11985 3715 12000 3735
rect 11950 3700 12000 3715
rect 12550 4185 12600 4200
rect 12550 4165 12565 4185
rect 12585 4165 12600 4185
rect 12550 4135 12600 4165
rect 12550 4115 12565 4135
rect 12585 4115 12600 4135
rect 12550 4085 12600 4115
rect 12550 4065 12565 4085
rect 12585 4065 12600 4085
rect 12550 4035 12600 4065
rect 12550 4015 12565 4035
rect 12585 4015 12600 4035
rect 12550 3985 12600 4015
rect 12550 3965 12565 3985
rect 12585 3965 12600 3985
rect 12550 3935 12600 3965
rect 12550 3915 12565 3935
rect 12585 3915 12600 3935
rect 12550 3885 12600 3915
rect 12550 3865 12565 3885
rect 12585 3865 12600 3885
rect 12550 3835 12600 3865
rect 12550 3815 12565 3835
rect 12585 3815 12600 3835
rect 12550 3785 12600 3815
rect 12550 3765 12565 3785
rect 12585 3765 12600 3785
rect 12550 3735 12600 3765
rect 12550 3715 12565 3735
rect 12585 3715 12600 3735
rect 12550 3700 12600 3715
rect 13150 4185 13200 4200
rect 13150 4165 13165 4185
rect 13185 4165 13200 4185
rect 13150 4135 13200 4165
rect 13150 4115 13165 4135
rect 13185 4115 13200 4135
rect 13150 4085 13200 4115
rect 13150 4065 13165 4085
rect 13185 4065 13200 4085
rect 13150 4035 13200 4065
rect 13150 4015 13165 4035
rect 13185 4015 13200 4035
rect 13150 3985 13200 4015
rect 13150 3965 13165 3985
rect 13185 3965 13200 3985
rect 13150 3935 13200 3965
rect 13150 3915 13165 3935
rect 13185 3915 13200 3935
rect 13150 3885 13200 3915
rect 13150 3865 13165 3885
rect 13185 3865 13200 3885
rect 13150 3835 13200 3865
rect 13150 3815 13165 3835
rect 13185 3815 13200 3835
rect 13150 3785 13200 3815
rect 13150 3765 13165 3785
rect 13185 3765 13200 3785
rect 13150 3735 13200 3765
rect 13150 3715 13165 3735
rect 13185 3715 13200 3735
rect 13150 3700 13200 3715
rect 13750 4185 13800 4200
rect 13750 4165 13765 4185
rect 13785 4165 13800 4185
rect 13750 4135 13800 4165
rect 13750 4115 13765 4135
rect 13785 4115 13800 4135
rect 13750 4085 13800 4115
rect 13750 4065 13765 4085
rect 13785 4065 13800 4085
rect 13750 4035 13800 4065
rect 13750 4015 13765 4035
rect 13785 4015 13800 4035
rect 13750 3985 13800 4015
rect 13750 3965 13765 3985
rect 13785 3965 13800 3985
rect 13750 3935 13800 3965
rect 13750 3915 13765 3935
rect 13785 3915 13800 3935
rect 13750 3885 13800 3915
rect 13750 3865 13765 3885
rect 13785 3865 13800 3885
rect 13750 3835 13800 3865
rect 13750 3815 13765 3835
rect 13785 3815 13800 3835
rect 13750 3785 13800 3815
rect 13750 3765 13765 3785
rect 13785 3765 13800 3785
rect 13750 3735 13800 3765
rect 13750 3715 13765 3735
rect 13785 3715 13800 3735
rect 13750 3700 13800 3715
rect 14350 4185 14400 4200
rect 14350 4165 14365 4185
rect 14385 4165 14400 4185
rect 14350 4135 14400 4165
rect 14350 4115 14365 4135
rect 14385 4115 14400 4135
rect 14350 4085 14400 4115
rect 14350 4065 14365 4085
rect 14385 4065 14400 4085
rect 14350 4035 14400 4065
rect 14350 4015 14365 4035
rect 14385 4015 14400 4035
rect 14350 3985 14400 4015
rect 14350 3965 14365 3985
rect 14385 3965 14400 3985
rect 14350 3935 14400 3965
rect 14350 3915 14365 3935
rect 14385 3915 14400 3935
rect 14350 3885 14400 3915
rect 14350 3865 14365 3885
rect 14385 3865 14400 3885
rect 14350 3835 14400 3865
rect 14350 3815 14365 3835
rect 14385 3815 14400 3835
rect 14350 3785 14400 3815
rect 14350 3765 14365 3785
rect 14385 3765 14400 3785
rect 14350 3735 14400 3765
rect 14350 3715 14365 3735
rect 14385 3715 14400 3735
rect 14350 3700 14400 3715
rect 14950 4185 15000 4200
rect 14950 4165 14965 4185
rect 14985 4165 15000 4185
rect 14950 4135 15000 4165
rect 14950 4115 14965 4135
rect 14985 4115 15000 4135
rect 14950 4085 15000 4115
rect 14950 4065 14965 4085
rect 14985 4065 15000 4085
rect 14950 4035 15000 4065
rect 14950 4015 14965 4035
rect 14985 4015 15000 4035
rect 14950 3985 15000 4015
rect 14950 3965 14965 3985
rect 14985 3965 15000 3985
rect 14950 3935 15000 3965
rect 14950 3915 14965 3935
rect 14985 3915 15000 3935
rect 14950 3885 15000 3915
rect 14950 3865 14965 3885
rect 14985 3865 15000 3885
rect 14950 3835 15000 3865
rect 14950 3815 14965 3835
rect 14985 3815 15000 3835
rect 14950 3785 15000 3815
rect 14950 3765 14965 3785
rect 14985 3765 15000 3785
rect 14950 3735 15000 3765
rect 14950 3715 14965 3735
rect 14985 3715 15000 3735
rect 14950 3700 15000 3715
rect 15550 4185 15600 4200
rect 15550 4165 15565 4185
rect 15585 4165 15600 4185
rect 15550 4135 15600 4165
rect 15550 4115 15565 4135
rect 15585 4115 15600 4135
rect 15550 4085 15600 4115
rect 15550 4065 15565 4085
rect 15585 4065 15600 4085
rect 15550 4035 15600 4065
rect 15550 4015 15565 4035
rect 15585 4015 15600 4035
rect 15550 3985 15600 4015
rect 15550 3965 15565 3985
rect 15585 3965 15600 3985
rect 15550 3935 15600 3965
rect 15550 3915 15565 3935
rect 15585 3915 15600 3935
rect 15550 3885 15600 3915
rect 15550 3865 15565 3885
rect 15585 3865 15600 3885
rect 15550 3835 15600 3865
rect 15550 3815 15565 3835
rect 15585 3815 15600 3835
rect 15550 3785 15600 3815
rect 15550 3765 15565 3785
rect 15585 3765 15600 3785
rect 15550 3735 15600 3765
rect 15550 3715 15565 3735
rect 15585 3715 15600 3735
rect 15550 3700 15600 3715
rect 16150 4185 16200 4200
rect 16150 4165 16165 4185
rect 16185 4165 16200 4185
rect 16150 4135 16200 4165
rect 16150 4115 16165 4135
rect 16185 4115 16200 4135
rect 16150 4085 16200 4115
rect 16150 4065 16165 4085
rect 16185 4065 16200 4085
rect 16150 4035 16200 4065
rect 16150 4015 16165 4035
rect 16185 4015 16200 4035
rect 16150 3985 16200 4015
rect 16150 3965 16165 3985
rect 16185 3965 16200 3985
rect 16150 3935 16200 3965
rect 16150 3915 16165 3935
rect 16185 3915 16200 3935
rect 16150 3885 16200 3915
rect 16150 3865 16165 3885
rect 16185 3865 16200 3885
rect 16150 3835 16200 3865
rect 16150 3815 16165 3835
rect 16185 3815 16200 3835
rect 16150 3785 16200 3815
rect 16150 3765 16165 3785
rect 16185 3765 16200 3785
rect 16150 3735 16200 3765
rect 16150 3715 16165 3735
rect 16185 3715 16200 3735
rect 16150 3700 16200 3715
rect 16300 4185 16350 4200
rect 16300 4165 16315 4185
rect 16335 4165 16350 4185
rect 16300 4135 16350 4165
rect 16300 4115 16315 4135
rect 16335 4115 16350 4135
rect 16300 4085 16350 4115
rect 16300 4065 16315 4085
rect 16335 4065 16350 4085
rect 16300 4035 16350 4065
rect 16300 4015 16315 4035
rect 16335 4015 16350 4035
rect 16300 3985 16350 4015
rect 16300 3965 16315 3985
rect 16335 3965 16350 3985
rect 16300 3935 16350 3965
rect 16300 3915 16315 3935
rect 16335 3915 16350 3935
rect 16300 3885 16350 3915
rect 16300 3865 16315 3885
rect 16335 3865 16350 3885
rect 16300 3835 16350 3865
rect 16300 3815 16315 3835
rect 16335 3815 16350 3835
rect 16300 3785 16350 3815
rect 16300 3765 16315 3785
rect 16335 3765 16350 3785
rect 16300 3735 16350 3765
rect 16300 3715 16315 3735
rect 16335 3715 16350 3735
rect 16300 3700 16350 3715
rect 16450 4185 16500 4200
rect 16450 4165 16465 4185
rect 16485 4165 16500 4185
rect 16450 4135 16500 4165
rect 16450 4115 16465 4135
rect 16485 4115 16500 4135
rect 16450 4085 16500 4115
rect 16450 4065 16465 4085
rect 16485 4065 16500 4085
rect 16450 4035 16500 4065
rect 16450 4015 16465 4035
rect 16485 4015 16500 4035
rect 16450 3985 16500 4015
rect 16450 3965 16465 3985
rect 16485 3965 16500 3985
rect 16450 3935 16500 3965
rect 16450 3915 16465 3935
rect 16485 3915 16500 3935
rect 16450 3885 16500 3915
rect 16450 3865 16465 3885
rect 16485 3865 16500 3885
rect 16450 3835 16500 3865
rect 16450 3815 16465 3835
rect 16485 3815 16500 3835
rect 16450 3785 16500 3815
rect 16450 3765 16465 3785
rect 16485 3765 16500 3785
rect 16450 3735 16500 3765
rect 16450 3715 16465 3735
rect 16485 3715 16500 3735
rect 16450 3700 16500 3715
rect 16600 4185 16650 4200
rect 16600 4165 16615 4185
rect 16635 4165 16650 4185
rect 16600 4135 16650 4165
rect 16600 4115 16615 4135
rect 16635 4115 16650 4135
rect 16600 4085 16650 4115
rect 16600 4065 16615 4085
rect 16635 4065 16650 4085
rect 16600 4035 16650 4065
rect 16600 4015 16615 4035
rect 16635 4015 16650 4035
rect 16600 3985 16650 4015
rect 16600 3965 16615 3985
rect 16635 3965 16650 3985
rect 16600 3935 16650 3965
rect 16600 3915 16615 3935
rect 16635 3915 16650 3935
rect 16600 3885 16650 3915
rect 16600 3865 16615 3885
rect 16635 3865 16650 3885
rect 16600 3835 16650 3865
rect 16600 3815 16615 3835
rect 16635 3815 16650 3835
rect 16600 3785 16650 3815
rect 16600 3765 16615 3785
rect 16635 3765 16650 3785
rect 16600 3735 16650 3765
rect 16600 3715 16615 3735
rect 16635 3715 16650 3735
rect 16600 3700 16650 3715
rect 16750 4185 16800 4200
rect 16750 4165 16765 4185
rect 16785 4165 16800 4185
rect 16750 4135 16800 4165
rect 16750 4115 16765 4135
rect 16785 4115 16800 4135
rect 16750 4085 16800 4115
rect 16750 4065 16765 4085
rect 16785 4065 16800 4085
rect 16750 4035 16800 4065
rect 16750 4015 16765 4035
rect 16785 4015 16800 4035
rect 16750 3985 16800 4015
rect 16750 3965 16765 3985
rect 16785 3965 16800 3985
rect 16750 3935 16800 3965
rect 16750 3915 16765 3935
rect 16785 3915 16800 3935
rect 16750 3885 16800 3915
rect 16750 3865 16765 3885
rect 16785 3865 16800 3885
rect 16750 3835 16800 3865
rect 16750 3815 16765 3835
rect 16785 3815 16800 3835
rect 16750 3785 16800 3815
rect 16750 3765 16765 3785
rect 16785 3765 16800 3785
rect 16750 3735 16800 3765
rect 16750 3715 16765 3735
rect 16785 3715 16800 3735
rect 16750 3700 16800 3715
rect 16900 4185 16950 4200
rect 16900 4165 16915 4185
rect 16935 4165 16950 4185
rect 16900 4135 16950 4165
rect 16900 4115 16915 4135
rect 16935 4115 16950 4135
rect 16900 4085 16950 4115
rect 16900 4065 16915 4085
rect 16935 4065 16950 4085
rect 16900 4035 16950 4065
rect 16900 4015 16915 4035
rect 16935 4015 16950 4035
rect 16900 3985 16950 4015
rect 16900 3965 16915 3985
rect 16935 3965 16950 3985
rect 16900 3935 16950 3965
rect 16900 3915 16915 3935
rect 16935 3915 16950 3935
rect 16900 3885 16950 3915
rect 16900 3865 16915 3885
rect 16935 3865 16950 3885
rect 16900 3835 16950 3865
rect 16900 3815 16915 3835
rect 16935 3815 16950 3835
rect 16900 3785 16950 3815
rect 16900 3765 16915 3785
rect 16935 3765 16950 3785
rect 16900 3735 16950 3765
rect 16900 3715 16915 3735
rect 16935 3715 16950 3735
rect 16900 3700 16950 3715
rect 17050 4185 17100 4200
rect 17050 4165 17065 4185
rect 17085 4165 17100 4185
rect 17050 4135 17100 4165
rect 17050 4115 17065 4135
rect 17085 4115 17100 4135
rect 17050 4085 17100 4115
rect 17050 4065 17065 4085
rect 17085 4065 17100 4085
rect 17050 4035 17100 4065
rect 17050 4015 17065 4035
rect 17085 4015 17100 4035
rect 17050 3985 17100 4015
rect 17050 3965 17065 3985
rect 17085 3965 17100 3985
rect 17050 3935 17100 3965
rect 17050 3915 17065 3935
rect 17085 3915 17100 3935
rect 17050 3885 17100 3915
rect 17050 3865 17065 3885
rect 17085 3865 17100 3885
rect 17050 3835 17100 3865
rect 17050 3815 17065 3835
rect 17085 3815 17100 3835
rect 17050 3785 17100 3815
rect 17050 3765 17065 3785
rect 17085 3765 17100 3785
rect 17050 3735 17100 3765
rect 17050 3715 17065 3735
rect 17085 3715 17100 3735
rect 17050 3700 17100 3715
rect 17200 4185 17250 4200
rect 17200 4165 17215 4185
rect 17235 4165 17250 4185
rect 17200 4135 17250 4165
rect 17200 4115 17215 4135
rect 17235 4115 17250 4135
rect 17200 4085 17250 4115
rect 17200 4065 17215 4085
rect 17235 4065 17250 4085
rect 17200 4035 17250 4065
rect 17200 4015 17215 4035
rect 17235 4015 17250 4035
rect 17200 3985 17250 4015
rect 17200 3965 17215 3985
rect 17235 3965 17250 3985
rect 17200 3935 17250 3965
rect 17200 3915 17215 3935
rect 17235 3915 17250 3935
rect 17200 3885 17250 3915
rect 17200 3865 17215 3885
rect 17235 3865 17250 3885
rect 17200 3835 17250 3865
rect 17200 3815 17215 3835
rect 17235 3815 17250 3835
rect 17200 3785 17250 3815
rect 17200 3765 17215 3785
rect 17235 3765 17250 3785
rect 17200 3735 17250 3765
rect 17200 3715 17215 3735
rect 17235 3715 17250 3735
rect 17200 3700 17250 3715
rect 17350 4185 17400 4200
rect 17350 4165 17365 4185
rect 17385 4165 17400 4185
rect 17350 4135 17400 4165
rect 17350 4115 17365 4135
rect 17385 4115 17400 4135
rect 17350 4085 17400 4115
rect 17350 4065 17365 4085
rect 17385 4065 17400 4085
rect 17350 4035 17400 4065
rect 17350 4015 17365 4035
rect 17385 4015 17400 4035
rect 17350 3985 17400 4015
rect 17350 3965 17365 3985
rect 17385 3965 17400 3985
rect 17350 3935 17400 3965
rect 17350 3915 17365 3935
rect 17385 3915 17400 3935
rect 17350 3885 17400 3915
rect 17350 3865 17365 3885
rect 17385 3865 17400 3885
rect 17350 3835 17400 3865
rect 17350 3815 17365 3835
rect 17385 3815 17400 3835
rect 17350 3785 17400 3815
rect 17350 3765 17365 3785
rect 17385 3765 17400 3785
rect 17350 3735 17400 3765
rect 17350 3715 17365 3735
rect 17385 3715 17400 3735
rect 17350 3700 17400 3715
rect 17950 4185 18000 4200
rect 17950 4165 17965 4185
rect 17985 4165 18000 4185
rect 17950 4135 18000 4165
rect 17950 4115 17965 4135
rect 17985 4115 18000 4135
rect 17950 4085 18000 4115
rect 17950 4065 17965 4085
rect 17985 4065 18000 4085
rect 17950 4035 18000 4065
rect 17950 4015 17965 4035
rect 17985 4015 18000 4035
rect 17950 3985 18000 4015
rect 17950 3965 17965 3985
rect 17985 3965 18000 3985
rect 17950 3935 18000 3965
rect 17950 3915 17965 3935
rect 17985 3915 18000 3935
rect 17950 3885 18000 3915
rect 17950 3865 17965 3885
rect 17985 3865 18000 3885
rect 17950 3835 18000 3865
rect 17950 3815 17965 3835
rect 17985 3815 18000 3835
rect 17950 3785 18000 3815
rect 17950 3765 17965 3785
rect 17985 3765 18000 3785
rect 17950 3735 18000 3765
rect 17950 3715 17965 3735
rect 17985 3715 18000 3735
rect 17950 3700 18000 3715
rect 18550 4185 18600 4200
rect 18550 4165 18565 4185
rect 18585 4165 18600 4185
rect 18550 4135 18600 4165
rect 18550 4115 18565 4135
rect 18585 4115 18600 4135
rect 18550 4085 18600 4115
rect 18550 4065 18565 4085
rect 18585 4065 18600 4085
rect 18550 4035 18600 4065
rect 18550 4015 18565 4035
rect 18585 4015 18600 4035
rect 18550 3985 18600 4015
rect 18550 3965 18565 3985
rect 18585 3965 18600 3985
rect 18550 3935 18600 3965
rect 18550 3915 18565 3935
rect 18585 3915 18600 3935
rect 18550 3885 18600 3915
rect 18550 3865 18565 3885
rect 18585 3865 18600 3885
rect 18550 3835 18600 3865
rect 18550 3815 18565 3835
rect 18585 3815 18600 3835
rect 18550 3785 18600 3815
rect 18550 3765 18565 3785
rect 18585 3765 18600 3785
rect 18550 3735 18600 3765
rect 18550 3715 18565 3735
rect 18585 3715 18600 3735
rect 18550 3700 18600 3715
rect 18700 4185 18750 4200
rect 18700 4165 18715 4185
rect 18735 4165 18750 4185
rect 18700 4135 18750 4165
rect 18700 4115 18715 4135
rect 18735 4115 18750 4135
rect 18700 4085 18750 4115
rect 18700 4065 18715 4085
rect 18735 4065 18750 4085
rect 18700 4035 18750 4065
rect 18700 4015 18715 4035
rect 18735 4015 18750 4035
rect 18700 3985 18750 4015
rect 18700 3965 18715 3985
rect 18735 3965 18750 3985
rect 18700 3935 18750 3965
rect 18700 3915 18715 3935
rect 18735 3915 18750 3935
rect 18700 3885 18750 3915
rect 18700 3865 18715 3885
rect 18735 3865 18750 3885
rect 18700 3835 18750 3865
rect 18700 3815 18715 3835
rect 18735 3815 18750 3835
rect 18700 3785 18750 3815
rect 18700 3765 18715 3785
rect 18735 3765 18750 3785
rect 18700 3735 18750 3765
rect 18700 3715 18715 3735
rect 18735 3715 18750 3735
rect 18700 3700 18750 3715
rect 18850 4185 18900 4200
rect 18850 4165 18865 4185
rect 18885 4165 18900 4185
rect 18850 4135 18900 4165
rect 18850 4115 18865 4135
rect 18885 4115 18900 4135
rect 18850 4085 18900 4115
rect 18850 4065 18865 4085
rect 18885 4065 18900 4085
rect 18850 4035 18900 4065
rect 18850 4015 18865 4035
rect 18885 4015 18900 4035
rect 18850 3985 18900 4015
rect 18850 3965 18865 3985
rect 18885 3965 18900 3985
rect 18850 3935 18900 3965
rect 18850 3915 18865 3935
rect 18885 3915 18900 3935
rect 18850 3885 18900 3915
rect 18850 3865 18865 3885
rect 18885 3865 18900 3885
rect 18850 3835 18900 3865
rect 18850 3815 18865 3835
rect 18885 3815 18900 3835
rect 18850 3785 18900 3815
rect 18850 3765 18865 3785
rect 18885 3765 18900 3785
rect 18850 3735 18900 3765
rect 18850 3715 18865 3735
rect 18885 3715 18900 3735
rect 18850 3700 18900 3715
rect 19000 4185 19050 4200
rect 19000 4165 19015 4185
rect 19035 4165 19050 4185
rect 19000 4135 19050 4165
rect 19000 4115 19015 4135
rect 19035 4115 19050 4135
rect 19000 4085 19050 4115
rect 19000 4065 19015 4085
rect 19035 4065 19050 4085
rect 19000 4035 19050 4065
rect 19000 4015 19015 4035
rect 19035 4015 19050 4035
rect 19000 3985 19050 4015
rect 19000 3965 19015 3985
rect 19035 3965 19050 3985
rect 19000 3935 19050 3965
rect 19000 3915 19015 3935
rect 19035 3915 19050 3935
rect 19000 3885 19050 3915
rect 19000 3865 19015 3885
rect 19035 3865 19050 3885
rect 19000 3835 19050 3865
rect 19000 3815 19015 3835
rect 19035 3815 19050 3835
rect 19000 3785 19050 3815
rect 19000 3765 19015 3785
rect 19035 3765 19050 3785
rect 19000 3735 19050 3765
rect 19000 3715 19015 3735
rect 19035 3715 19050 3735
rect 19000 3700 19050 3715
rect 19150 4185 19200 4200
rect 19150 4165 19165 4185
rect 19185 4165 19200 4185
rect 19150 4135 19200 4165
rect 19150 4115 19165 4135
rect 19185 4115 19200 4135
rect 19150 4085 19200 4115
rect 19150 4065 19165 4085
rect 19185 4065 19200 4085
rect 19150 4035 19200 4065
rect 19150 4015 19165 4035
rect 19185 4015 19200 4035
rect 19150 3985 19200 4015
rect 19150 3965 19165 3985
rect 19185 3965 19200 3985
rect 19150 3935 19200 3965
rect 19150 3915 19165 3935
rect 19185 3915 19200 3935
rect 19150 3885 19200 3915
rect 19150 3865 19165 3885
rect 19185 3865 19200 3885
rect 19150 3835 19200 3865
rect 19150 3815 19165 3835
rect 19185 3815 19200 3835
rect 19150 3785 19200 3815
rect 19150 3765 19165 3785
rect 19185 3765 19200 3785
rect 19150 3735 19200 3765
rect 19150 3715 19165 3735
rect 19185 3715 19200 3735
rect 19150 3700 19200 3715
rect 19300 4185 19350 4200
rect 19300 4165 19315 4185
rect 19335 4165 19350 4185
rect 19300 4135 19350 4165
rect 19300 4115 19315 4135
rect 19335 4115 19350 4135
rect 19300 4085 19350 4115
rect 19300 4065 19315 4085
rect 19335 4065 19350 4085
rect 19300 4035 19350 4065
rect 19300 4015 19315 4035
rect 19335 4015 19350 4035
rect 19300 3985 19350 4015
rect 19300 3965 19315 3985
rect 19335 3965 19350 3985
rect 19300 3935 19350 3965
rect 19300 3915 19315 3935
rect 19335 3915 19350 3935
rect 19300 3885 19350 3915
rect 19300 3865 19315 3885
rect 19335 3865 19350 3885
rect 19300 3835 19350 3865
rect 19300 3815 19315 3835
rect 19335 3815 19350 3835
rect 19300 3785 19350 3815
rect 19300 3765 19315 3785
rect 19335 3765 19350 3785
rect 19300 3735 19350 3765
rect 19300 3715 19315 3735
rect 19335 3715 19350 3735
rect 19300 3700 19350 3715
rect 19450 4185 19500 4200
rect 19450 4165 19465 4185
rect 19485 4165 19500 4185
rect 19450 4135 19500 4165
rect 19450 4115 19465 4135
rect 19485 4115 19500 4135
rect 19450 4085 19500 4115
rect 19450 4065 19465 4085
rect 19485 4065 19500 4085
rect 19450 4035 19500 4065
rect 19450 4015 19465 4035
rect 19485 4015 19500 4035
rect 19450 3985 19500 4015
rect 19450 3965 19465 3985
rect 19485 3965 19500 3985
rect 19450 3935 19500 3965
rect 19450 3915 19465 3935
rect 19485 3915 19500 3935
rect 19450 3885 19500 3915
rect 19450 3865 19465 3885
rect 19485 3865 19500 3885
rect 19450 3835 19500 3865
rect 19450 3815 19465 3835
rect 19485 3815 19500 3835
rect 19450 3785 19500 3815
rect 19450 3765 19465 3785
rect 19485 3765 19500 3785
rect 19450 3735 19500 3765
rect 19450 3715 19465 3735
rect 19485 3715 19500 3735
rect 19450 3700 19500 3715
rect 19600 4185 19650 4200
rect 19600 4165 19615 4185
rect 19635 4165 19650 4185
rect 19600 4135 19650 4165
rect 19600 4115 19615 4135
rect 19635 4115 19650 4135
rect 19600 4085 19650 4115
rect 19600 4065 19615 4085
rect 19635 4065 19650 4085
rect 19600 4035 19650 4065
rect 19600 4015 19615 4035
rect 19635 4015 19650 4035
rect 19600 3985 19650 4015
rect 19600 3965 19615 3985
rect 19635 3965 19650 3985
rect 19600 3935 19650 3965
rect 19600 3915 19615 3935
rect 19635 3915 19650 3935
rect 19600 3885 19650 3915
rect 19600 3865 19615 3885
rect 19635 3865 19650 3885
rect 19600 3835 19650 3865
rect 19600 3815 19615 3835
rect 19635 3815 19650 3835
rect 19600 3785 19650 3815
rect 19600 3765 19615 3785
rect 19635 3765 19650 3785
rect 19600 3735 19650 3765
rect 19600 3715 19615 3735
rect 19635 3715 19650 3735
rect 19600 3700 19650 3715
rect 19750 4185 19800 4200
rect 19750 4165 19765 4185
rect 19785 4165 19800 4185
rect 19750 4135 19800 4165
rect 19750 4115 19765 4135
rect 19785 4115 19800 4135
rect 19750 4085 19800 4115
rect 19750 4065 19765 4085
rect 19785 4065 19800 4085
rect 19750 4035 19800 4065
rect 19750 4015 19765 4035
rect 19785 4015 19800 4035
rect 19750 3985 19800 4015
rect 19750 3965 19765 3985
rect 19785 3965 19800 3985
rect 19750 3935 19800 3965
rect 19750 3915 19765 3935
rect 19785 3915 19800 3935
rect 19750 3885 19800 3915
rect 19750 3865 19765 3885
rect 19785 3865 19800 3885
rect 19750 3835 19800 3865
rect 19750 3815 19765 3835
rect 19785 3815 19800 3835
rect 19750 3785 19800 3815
rect 19750 3765 19765 3785
rect 19785 3765 19800 3785
rect 19750 3735 19800 3765
rect 19750 3715 19765 3735
rect 19785 3715 19800 3735
rect 19750 3700 19800 3715
rect 20350 4185 20400 4200
rect 20350 4165 20365 4185
rect 20385 4165 20400 4185
rect 20350 4135 20400 4165
rect 20350 4115 20365 4135
rect 20385 4115 20400 4135
rect 20350 4085 20400 4115
rect 20350 4065 20365 4085
rect 20385 4065 20400 4085
rect 20350 4035 20400 4065
rect 20350 4015 20365 4035
rect 20385 4015 20400 4035
rect 20350 3985 20400 4015
rect 20350 3965 20365 3985
rect 20385 3965 20400 3985
rect 20350 3935 20400 3965
rect 20350 3915 20365 3935
rect 20385 3915 20400 3935
rect 20350 3885 20400 3915
rect 20350 3865 20365 3885
rect 20385 3865 20400 3885
rect 20350 3835 20400 3865
rect 20350 3815 20365 3835
rect 20385 3815 20400 3835
rect 20350 3785 20400 3815
rect 20350 3765 20365 3785
rect 20385 3765 20400 3785
rect 20350 3735 20400 3765
rect 20350 3715 20365 3735
rect 20385 3715 20400 3735
rect 20350 3700 20400 3715
rect 20950 4185 21000 4200
rect 20950 4165 20965 4185
rect 20985 4165 21000 4185
rect 20950 4135 21000 4165
rect 20950 4115 20965 4135
rect 20985 4115 21000 4135
rect 20950 4085 21000 4115
rect 20950 4065 20965 4085
rect 20985 4065 21000 4085
rect 20950 4035 21000 4065
rect 20950 4015 20965 4035
rect 20985 4015 21000 4035
rect 20950 3985 21000 4015
rect 20950 3965 20965 3985
rect 20985 3965 21000 3985
rect 20950 3935 21000 3965
rect 20950 3915 20965 3935
rect 20985 3915 21000 3935
rect 20950 3885 21000 3915
rect 20950 3865 20965 3885
rect 20985 3865 21000 3885
rect 20950 3835 21000 3865
rect 20950 3815 20965 3835
rect 20985 3815 21000 3835
rect 20950 3785 21000 3815
rect 20950 3765 20965 3785
rect 20985 3765 21000 3785
rect 20950 3735 21000 3765
rect 20950 3715 20965 3735
rect 20985 3715 21000 3735
rect 20950 3700 21000 3715
rect 21400 4185 21450 4200
rect 21400 4165 21415 4185
rect 21435 4165 21450 4185
rect 21400 4135 21450 4165
rect 21400 4115 21415 4135
rect 21435 4115 21450 4135
rect 21400 4085 21450 4115
rect 21400 4065 21415 4085
rect 21435 4065 21450 4085
rect 21400 4035 21450 4065
rect 21400 4015 21415 4035
rect 21435 4015 21450 4035
rect 21400 3985 21450 4015
rect 21400 3965 21415 3985
rect 21435 3965 21450 3985
rect 21400 3935 21450 3965
rect 21400 3915 21415 3935
rect 21435 3915 21450 3935
rect 21400 3885 21450 3915
rect 21400 3865 21415 3885
rect 21435 3865 21450 3885
rect 21400 3835 21450 3865
rect 21400 3815 21415 3835
rect 21435 3815 21450 3835
rect 21400 3785 21450 3815
rect 21400 3765 21415 3785
rect 21435 3765 21450 3785
rect 21400 3735 21450 3765
rect 21400 3715 21415 3735
rect 21435 3715 21450 3735
rect 21400 3700 21450 3715
rect 21850 4185 21900 4200
rect 21850 4165 21865 4185
rect 21885 4165 21900 4185
rect 21850 4135 21900 4165
rect 21850 4115 21865 4135
rect 21885 4115 21900 4135
rect 21850 4085 21900 4115
rect 21850 4065 21865 4085
rect 21885 4065 21900 4085
rect 21850 4035 21900 4065
rect 21850 4015 21865 4035
rect 21885 4015 21900 4035
rect 21850 3985 21900 4015
rect 21850 3965 21865 3985
rect 21885 3965 21900 3985
rect 21850 3935 21900 3965
rect 21850 3915 21865 3935
rect 21885 3915 21900 3935
rect 21850 3885 21900 3915
rect 21850 3865 21865 3885
rect 21885 3865 21900 3885
rect 21850 3835 21900 3865
rect 21850 3815 21865 3835
rect 21885 3815 21900 3835
rect 21850 3785 21900 3815
rect 21850 3765 21865 3785
rect 21885 3765 21900 3785
rect 21850 3735 21900 3765
rect 21850 3715 21865 3735
rect 21885 3715 21900 3735
rect 21850 3700 21900 3715
rect 22450 4185 22500 4200
rect 22450 4165 22465 4185
rect 22485 4165 22500 4185
rect 22450 4135 22500 4165
rect 22450 4115 22465 4135
rect 22485 4115 22500 4135
rect 22450 4085 22500 4115
rect 22450 4065 22465 4085
rect 22485 4065 22500 4085
rect 22450 4035 22500 4065
rect 22450 4015 22465 4035
rect 22485 4015 22500 4035
rect 22450 3985 22500 4015
rect 22450 3965 22465 3985
rect 22485 3965 22500 3985
rect 22450 3935 22500 3965
rect 22450 3915 22465 3935
rect 22485 3915 22500 3935
rect 22450 3885 22500 3915
rect 22450 3865 22465 3885
rect 22485 3865 22500 3885
rect 22450 3835 22500 3865
rect 22450 3815 22465 3835
rect 22485 3815 22500 3835
rect 22450 3785 22500 3815
rect 22450 3765 22465 3785
rect 22485 3765 22500 3785
rect 22450 3735 22500 3765
rect 22450 3715 22465 3735
rect 22485 3715 22500 3735
rect 22450 3700 22500 3715
rect 23050 4185 23100 4200
rect 23050 4165 23065 4185
rect 23085 4165 23100 4185
rect 23050 4135 23100 4165
rect 23050 4115 23065 4135
rect 23085 4115 23100 4135
rect 23050 4085 23100 4115
rect 23050 4065 23065 4085
rect 23085 4065 23100 4085
rect 23050 4035 23100 4065
rect 23050 4015 23065 4035
rect 23085 4015 23100 4035
rect 23050 3985 23100 4015
rect 23050 3965 23065 3985
rect 23085 3965 23100 3985
rect 23050 3935 23100 3965
rect 23050 3915 23065 3935
rect 23085 3915 23100 3935
rect 23050 3885 23100 3915
rect 23050 3865 23065 3885
rect 23085 3865 23100 3885
rect 23050 3835 23100 3865
rect 23050 3815 23065 3835
rect 23085 3815 23100 3835
rect 23050 3785 23100 3815
rect 23050 3765 23065 3785
rect 23085 3765 23100 3785
rect 23050 3735 23100 3765
rect 23050 3715 23065 3735
rect 23085 3715 23100 3735
rect 23050 3700 23100 3715
rect 23500 4185 23550 4200
rect 23500 4165 23515 4185
rect 23535 4165 23550 4185
rect 23500 4135 23550 4165
rect 23500 4115 23515 4135
rect 23535 4115 23550 4135
rect 23500 4085 23550 4115
rect 23500 4065 23515 4085
rect 23535 4065 23550 4085
rect 23500 4035 23550 4065
rect 23500 4015 23515 4035
rect 23535 4015 23550 4035
rect 23500 3985 23550 4015
rect 23500 3965 23515 3985
rect 23535 3965 23550 3985
rect 23500 3935 23550 3965
rect 23500 3915 23515 3935
rect 23535 3915 23550 3935
rect 23500 3885 23550 3915
rect 23500 3865 23515 3885
rect 23535 3865 23550 3885
rect 23500 3835 23550 3865
rect 23500 3815 23515 3835
rect 23535 3815 23550 3835
rect 23500 3785 23550 3815
rect 23500 3765 23515 3785
rect 23535 3765 23550 3785
rect 23500 3735 23550 3765
rect 23500 3715 23515 3735
rect 23535 3715 23550 3735
rect 23500 3700 23550 3715
rect 23950 4185 24000 4200
rect 23950 4165 23965 4185
rect 23985 4165 24000 4185
rect 23950 4135 24000 4165
rect 23950 4115 23965 4135
rect 23985 4115 24000 4135
rect 23950 4085 24000 4115
rect 23950 4065 23965 4085
rect 23985 4065 24000 4085
rect 23950 4035 24000 4065
rect 23950 4015 23965 4035
rect 23985 4015 24000 4035
rect 23950 3985 24000 4015
rect 23950 3965 23965 3985
rect 23985 3965 24000 3985
rect 23950 3935 24000 3965
rect 23950 3915 23965 3935
rect 23985 3915 24000 3935
rect 23950 3885 24000 3915
rect 23950 3865 23965 3885
rect 23985 3865 24000 3885
rect 23950 3835 24000 3865
rect 23950 3815 23965 3835
rect 23985 3815 24000 3835
rect 23950 3785 24000 3815
rect 23950 3765 23965 3785
rect 23985 3765 24000 3785
rect 23950 3735 24000 3765
rect 23950 3715 23965 3735
rect 23985 3715 24000 3735
rect 23950 3700 24000 3715
rect 24550 4185 24600 4200
rect 24550 4165 24565 4185
rect 24585 4165 24600 4185
rect 24550 4135 24600 4165
rect 24550 4115 24565 4135
rect 24585 4115 24600 4135
rect 24550 4085 24600 4115
rect 24550 4065 24565 4085
rect 24585 4065 24600 4085
rect 24550 4035 24600 4065
rect 24550 4015 24565 4035
rect 24585 4015 24600 4035
rect 24550 3985 24600 4015
rect 24550 3965 24565 3985
rect 24585 3965 24600 3985
rect 24550 3935 24600 3965
rect 24550 3915 24565 3935
rect 24585 3915 24600 3935
rect 24550 3885 24600 3915
rect 24550 3865 24565 3885
rect 24585 3865 24600 3885
rect 24550 3835 24600 3865
rect 24550 3815 24565 3835
rect 24585 3815 24600 3835
rect 24550 3785 24600 3815
rect 24550 3765 24565 3785
rect 24585 3765 24600 3785
rect 24550 3735 24600 3765
rect 24550 3715 24565 3735
rect 24585 3715 24600 3735
rect 24550 3700 24600 3715
rect 25150 4185 25200 4200
rect 25150 4165 25165 4185
rect 25185 4165 25200 4185
rect 25150 4135 25200 4165
rect 25150 4115 25165 4135
rect 25185 4115 25200 4135
rect 25150 4085 25200 4115
rect 25150 4065 25165 4085
rect 25185 4065 25200 4085
rect 25150 4035 25200 4065
rect 25150 4015 25165 4035
rect 25185 4015 25200 4035
rect 25150 3985 25200 4015
rect 25150 3965 25165 3985
rect 25185 3965 25200 3985
rect 25150 3935 25200 3965
rect 25150 3915 25165 3935
rect 25185 3915 25200 3935
rect 25150 3885 25200 3915
rect 25150 3865 25165 3885
rect 25185 3865 25200 3885
rect 25150 3835 25200 3865
rect 25150 3815 25165 3835
rect 25185 3815 25200 3835
rect 25150 3785 25200 3815
rect 25150 3765 25165 3785
rect 25185 3765 25200 3785
rect 25150 3735 25200 3765
rect 25150 3715 25165 3735
rect 25185 3715 25200 3735
rect 25150 3700 25200 3715
rect 25600 4185 25650 4200
rect 25600 4165 25615 4185
rect 25635 4165 25650 4185
rect 25600 4135 25650 4165
rect 25600 4115 25615 4135
rect 25635 4115 25650 4135
rect 25600 4085 25650 4115
rect 25600 4065 25615 4085
rect 25635 4065 25650 4085
rect 25600 4035 25650 4065
rect 25600 4015 25615 4035
rect 25635 4015 25650 4035
rect 25600 3985 25650 4015
rect 25600 3965 25615 3985
rect 25635 3965 25650 3985
rect 25600 3935 25650 3965
rect 25600 3915 25615 3935
rect 25635 3915 25650 3935
rect 25600 3885 25650 3915
rect 25600 3865 25615 3885
rect 25635 3865 25650 3885
rect 25600 3835 25650 3865
rect 25600 3815 25615 3835
rect 25635 3815 25650 3835
rect 25600 3785 25650 3815
rect 25600 3765 25615 3785
rect 25635 3765 25650 3785
rect 25600 3735 25650 3765
rect 25600 3715 25615 3735
rect 25635 3715 25650 3735
rect 25600 3700 25650 3715
rect 26050 4185 26100 4200
rect 26050 4165 26065 4185
rect 26085 4165 26100 4185
rect 26050 4135 26100 4165
rect 26050 4115 26065 4135
rect 26085 4115 26100 4135
rect 26050 4085 26100 4115
rect 26050 4065 26065 4085
rect 26085 4065 26100 4085
rect 26050 4035 26100 4065
rect 26050 4015 26065 4035
rect 26085 4015 26100 4035
rect 26050 3985 26100 4015
rect 26050 3965 26065 3985
rect 26085 3965 26100 3985
rect 26050 3935 26100 3965
rect 26050 3915 26065 3935
rect 26085 3915 26100 3935
rect 26050 3885 26100 3915
rect 26050 3865 26065 3885
rect 26085 3865 26100 3885
rect 26050 3835 26100 3865
rect 26050 3815 26065 3835
rect 26085 3815 26100 3835
rect 26050 3785 26100 3815
rect 26050 3765 26065 3785
rect 26085 3765 26100 3785
rect 26050 3735 26100 3765
rect 26050 3715 26065 3735
rect 26085 3715 26100 3735
rect 26050 3700 26100 3715
rect 26650 4185 26700 4200
rect 26650 4165 26665 4185
rect 26685 4165 26700 4185
rect 26650 4135 26700 4165
rect 26650 4115 26665 4135
rect 26685 4115 26700 4135
rect 26650 4085 26700 4115
rect 26650 4065 26665 4085
rect 26685 4065 26700 4085
rect 26650 4035 26700 4065
rect 26650 4015 26665 4035
rect 26685 4015 26700 4035
rect 26650 3985 26700 4015
rect 26650 3965 26665 3985
rect 26685 3965 26700 3985
rect 26650 3935 26700 3965
rect 26650 3915 26665 3935
rect 26685 3915 26700 3935
rect 26650 3885 26700 3915
rect 26650 3865 26665 3885
rect 26685 3865 26700 3885
rect 26650 3835 26700 3865
rect 26650 3815 26665 3835
rect 26685 3815 26700 3835
rect 26650 3785 26700 3815
rect 26650 3765 26665 3785
rect 26685 3765 26700 3785
rect 26650 3735 26700 3765
rect 26650 3715 26665 3735
rect 26685 3715 26700 3735
rect 26650 3700 26700 3715
rect 27250 4185 27300 4200
rect 27250 4165 27265 4185
rect 27285 4165 27300 4185
rect 27250 4135 27300 4165
rect 27250 4115 27265 4135
rect 27285 4115 27300 4135
rect 27250 4085 27300 4115
rect 27250 4065 27265 4085
rect 27285 4065 27300 4085
rect 27250 4035 27300 4065
rect 27250 4015 27265 4035
rect 27285 4015 27300 4035
rect 27250 3985 27300 4015
rect 27250 3965 27265 3985
rect 27285 3965 27300 3985
rect 27250 3935 27300 3965
rect 27250 3915 27265 3935
rect 27285 3915 27300 3935
rect 27250 3885 27300 3915
rect 27250 3865 27265 3885
rect 27285 3865 27300 3885
rect 27250 3835 27300 3865
rect 27250 3815 27265 3835
rect 27285 3815 27300 3835
rect 27250 3785 27300 3815
rect 27250 3765 27265 3785
rect 27285 3765 27300 3785
rect 27250 3735 27300 3765
rect 27250 3715 27265 3735
rect 27285 3715 27300 3735
rect 27250 3700 27300 3715
rect 27700 4185 27750 4200
rect 27700 4165 27715 4185
rect 27735 4165 27750 4185
rect 27700 4135 27750 4165
rect 27700 4115 27715 4135
rect 27735 4115 27750 4135
rect 27700 4085 27750 4115
rect 27700 4065 27715 4085
rect 27735 4065 27750 4085
rect 27700 4035 27750 4065
rect 27700 4015 27715 4035
rect 27735 4015 27750 4035
rect 27700 3985 27750 4015
rect 27700 3965 27715 3985
rect 27735 3965 27750 3985
rect 27700 3935 27750 3965
rect 27700 3915 27715 3935
rect 27735 3915 27750 3935
rect 27700 3885 27750 3915
rect 27700 3865 27715 3885
rect 27735 3865 27750 3885
rect 27700 3835 27750 3865
rect 27700 3815 27715 3835
rect 27735 3815 27750 3835
rect 27700 3785 27750 3815
rect 27700 3765 27715 3785
rect 27735 3765 27750 3785
rect 27700 3735 27750 3765
rect 27700 3715 27715 3735
rect 27735 3715 27750 3735
rect 27700 3700 27750 3715
rect 28150 4185 28200 4200
rect 28150 4165 28165 4185
rect 28185 4165 28200 4185
rect 28150 4135 28200 4165
rect 28150 4115 28165 4135
rect 28185 4115 28200 4135
rect 28150 4085 28200 4115
rect 28150 4065 28165 4085
rect 28185 4065 28200 4085
rect 28150 4035 28200 4065
rect 28150 4015 28165 4035
rect 28185 4015 28200 4035
rect 28150 3985 28200 4015
rect 28150 3965 28165 3985
rect 28185 3965 28200 3985
rect 28150 3935 28200 3965
rect 28150 3915 28165 3935
rect 28185 3915 28200 3935
rect 28150 3885 28200 3915
rect 28150 3865 28165 3885
rect 28185 3865 28200 3885
rect 28150 3835 28200 3865
rect 28150 3815 28165 3835
rect 28185 3815 28200 3835
rect 28150 3785 28200 3815
rect 28150 3765 28165 3785
rect 28185 3765 28200 3785
rect 28150 3735 28200 3765
rect 28150 3715 28165 3735
rect 28185 3715 28200 3735
rect 28150 3700 28200 3715
rect 28750 4185 28800 4200
rect 28750 4165 28765 4185
rect 28785 4165 28800 4185
rect 28750 4135 28800 4165
rect 28750 4115 28765 4135
rect 28785 4115 28800 4135
rect 28750 4085 28800 4115
rect 28750 4065 28765 4085
rect 28785 4065 28800 4085
rect 28750 4035 28800 4065
rect 28750 4015 28765 4035
rect 28785 4015 28800 4035
rect 28750 3985 28800 4015
rect 28750 3965 28765 3985
rect 28785 3965 28800 3985
rect 28750 3935 28800 3965
rect 28750 3915 28765 3935
rect 28785 3915 28800 3935
rect 28750 3885 28800 3915
rect 28750 3865 28765 3885
rect 28785 3865 28800 3885
rect 28750 3835 28800 3865
rect 28750 3815 28765 3835
rect 28785 3815 28800 3835
rect 28750 3785 28800 3815
rect 28750 3765 28765 3785
rect 28785 3765 28800 3785
rect 28750 3735 28800 3765
rect 28750 3715 28765 3735
rect 28785 3715 28800 3735
rect 28750 3700 28800 3715
rect 29350 4185 29400 4200
rect 29350 4165 29365 4185
rect 29385 4165 29400 4185
rect 29350 4135 29400 4165
rect 29350 4115 29365 4135
rect 29385 4115 29400 4135
rect 29350 4085 29400 4115
rect 29350 4065 29365 4085
rect 29385 4065 29400 4085
rect 29350 4035 29400 4065
rect 29350 4015 29365 4035
rect 29385 4015 29400 4035
rect 29350 3985 29400 4015
rect 29350 3965 29365 3985
rect 29385 3965 29400 3985
rect 29350 3935 29400 3965
rect 29350 3915 29365 3935
rect 29385 3915 29400 3935
rect 29350 3885 29400 3915
rect 29350 3865 29365 3885
rect 29385 3865 29400 3885
rect 29350 3835 29400 3865
rect 29350 3815 29365 3835
rect 29385 3815 29400 3835
rect 29350 3785 29400 3815
rect 29350 3765 29365 3785
rect 29385 3765 29400 3785
rect 29350 3735 29400 3765
rect 29350 3715 29365 3735
rect 29385 3715 29400 3735
rect 29350 3700 29400 3715
rect 29500 4185 29550 4200
rect 29500 4165 29515 4185
rect 29535 4165 29550 4185
rect 29500 4135 29550 4165
rect 29500 4115 29515 4135
rect 29535 4115 29550 4135
rect 29500 4085 29550 4115
rect 29500 4065 29515 4085
rect 29535 4065 29550 4085
rect 29500 4035 29550 4065
rect 29500 4015 29515 4035
rect 29535 4015 29550 4035
rect 29500 3985 29550 4015
rect 29500 3965 29515 3985
rect 29535 3965 29550 3985
rect 29500 3935 29550 3965
rect 29500 3915 29515 3935
rect 29535 3915 29550 3935
rect 29500 3885 29550 3915
rect 29500 3865 29515 3885
rect 29535 3865 29550 3885
rect 29500 3835 29550 3865
rect 29500 3815 29515 3835
rect 29535 3815 29550 3835
rect 29500 3785 29550 3815
rect 29500 3765 29515 3785
rect 29535 3765 29550 3785
rect 29500 3735 29550 3765
rect 29500 3715 29515 3735
rect 29535 3715 29550 3735
rect 29500 3700 29550 3715
rect 29650 4185 29700 4200
rect 29650 4165 29665 4185
rect 29685 4165 29700 4185
rect 29650 4135 29700 4165
rect 29650 4115 29665 4135
rect 29685 4115 29700 4135
rect 29650 4085 29700 4115
rect 29650 4065 29665 4085
rect 29685 4065 29700 4085
rect 29650 4035 29700 4065
rect 29650 4015 29665 4035
rect 29685 4015 29700 4035
rect 29650 3985 29700 4015
rect 29650 3965 29665 3985
rect 29685 3965 29700 3985
rect 29650 3935 29700 3965
rect 29650 3915 29665 3935
rect 29685 3915 29700 3935
rect 29650 3885 29700 3915
rect 29650 3865 29665 3885
rect 29685 3865 29700 3885
rect 29650 3835 29700 3865
rect 29650 3815 29665 3835
rect 29685 3815 29700 3835
rect 29650 3785 29700 3815
rect 29650 3765 29665 3785
rect 29685 3765 29700 3785
rect 29650 3735 29700 3765
rect 29650 3715 29665 3735
rect 29685 3715 29700 3735
rect 29650 3700 29700 3715
rect 29800 4185 29850 4200
rect 29800 4165 29815 4185
rect 29835 4165 29850 4185
rect 29800 4135 29850 4165
rect 29800 4115 29815 4135
rect 29835 4115 29850 4135
rect 29800 4085 29850 4115
rect 29800 4065 29815 4085
rect 29835 4065 29850 4085
rect 29800 4035 29850 4065
rect 29800 4015 29815 4035
rect 29835 4015 29850 4035
rect 29800 3985 29850 4015
rect 29800 3965 29815 3985
rect 29835 3965 29850 3985
rect 29800 3935 29850 3965
rect 29800 3915 29815 3935
rect 29835 3915 29850 3935
rect 29800 3885 29850 3915
rect 29800 3865 29815 3885
rect 29835 3865 29850 3885
rect 29800 3835 29850 3865
rect 29800 3815 29815 3835
rect 29835 3815 29850 3835
rect 29800 3785 29850 3815
rect 29800 3765 29815 3785
rect 29835 3765 29850 3785
rect 29800 3735 29850 3765
rect 29800 3715 29815 3735
rect 29835 3715 29850 3735
rect 29800 3700 29850 3715
rect 29950 4185 30000 4200
rect 29950 4165 29965 4185
rect 29985 4165 30000 4185
rect 29950 4135 30000 4165
rect 29950 4115 29965 4135
rect 29985 4115 30000 4135
rect 29950 4085 30000 4115
rect 29950 4065 29965 4085
rect 29985 4065 30000 4085
rect 29950 4035 30000 4065
rect 29950 4015 29965 4035
rect 29985 4015 30000 4035
rect 29950 3985 30000 4015
rect 29950 3965 29965 3985
rect 29985 3965 30000 3985
rect 29950 3935 30000 3965
rect 29950 3915 29965 3935
rect 29985 3915 30000 3935
rect 29950 3885 30000 3915
rect 29950 3865 29965 3885
rect 29985 3865 30000 3885
rect 29950 3835 30000 3865
rect 29950 3815 29965 3835
rect 29985 3815 30000 3835
rect 29950 3785 30000 3815
rect 29950 3765 29965 3785
rect 29985 3765 30000 3785
rect 29950 3735 30000 3765
rect 29950 3715 29965 3735
rect 29985 3715 30000 3735
rect 29950 3700 30000 3715
rect 30100 4185 30150 4200
rect 30100 4165 30115 4185
rect 30135 4165 30150 4185
rect 30100 4135 30150 4165
rect 30100 4115 30115 4135
rect 30135 4115 30150 4135
rect 30100 4085 30150 4115
rect 30100 4065 30115 4085
rect 30135 4065 30150 4085
rect 30100 4035 30150 4065
rect 30100 4015 30115 4035
rect 30135 4015 30150 4035
rect 30100 3985 30150 4015
rect 30100 3965 30115 3985
rect 30135 3965 30150 3985
rect 30100 3935 30150 3965
rect 30100 3915 30115 3935
rect 30135 3915 30150 3935
rect 30100 3885 30150 3915
rect 30100 3865 30115 3885
rect 30135 3865 30150 3885
rect 30100 3835 30150 3865
rect 30100 3815 30115 3835
rect 30135 3815 30150 3835
rect 30100 3785 30150 3815
rect 30100 3765 30115 3785
rect 30135 3765 30150 3785
rect 30100 3735 30150 3765
rect 30100 3715 30115 3735
rect 30135 3715 30150 3735
rect 30100 3700 30150 3715
rect 30250 4185 30300 4200
rect 30250 4165 30265 4185
rect 30285 4165 30300 4185
rect 30250 4135 30300 4165
rect 30250 4115 30265 4135
rect 30285 4115 30300 4135
rect 30250 4085 30300 4115
rect 30250 4065 30265 4085
rect 30285 4065 30300 4085
rect 30250 4035 30300 4065
rect 30250 4015 30265 4035
rect 30285 4015 30300 4035
rect 30250 3985 30300 4015
rect 30250 3965 30265 3985
rect 30285 3965 30300 3985
rect 30250 3935 30300 3965
rect 30250 3915 30265 3935
rect 30285 3915 30300 3935
rect 30250 3885 30300 3915
rect 30250 3865 30265 3885
rect 30285 3865 30300 3885
rect 30250 3835 30300 3865
rect 30250 3815 30265 3835
rect 30285 3815 30300 3835
rect 30250 3785 30300 3815
rect 30250 3765 30265 3785
rect 30285 3765 30300 3785
rect 30250 3735 30300 3765
rect 30250 3715 30265 3735
rect 30285 3715 30300 3735
rect 30250 3700 30300 3715
rect 30400 4185 30450 4200
rect 30400 4165 30415 4185
rect 30435 4165 30450 4185
rect 30400 4135 30450 4165
rect 30400 4115 30415 4135
rect 30435 4115 30450 4135
rect 30400 4085 30450 4115
rect 30400 4065 30415 4085
rect 30435 4065 30450 4085
rect 30400 4035 30450 4065
rect 30400 4015 30415 4035
rect 30435 4015 30450 4035
rect 30400 3985 30450 4015
rect 30400 3965 30415 3985
rect 30435 3965 30450 3985
rect 30400 3935 30450 3965
rect 30400 3915 30415 3935
rect 30435 3915 30450 3935
rect 30400 3885 30450 3915
rect 30400 3865 30415 3885
rect 30435 3865 30450 3885
rect 30400 3835 30450 3865
rect 30400 3815 30415 3835
rect 30435 3815 30450 3835
rect 30400 3785 30450 3815
rect 30400 3765 30415 3785
rect 30435 3765 30450 3785
rect 30400 3735 30450 3765
rect 30400 3715 30415 3735
rect 30435 3715 30450 3735
rect 30400 3700 30450 3715
rect 30550 4185 30600 4200
rect 30550 4165 30565 4185
rect 30585 4165 30600 4185
rect 30550 4135 30600 4165
rect 30550 4115 30565 4135
rect 30585 4115 30600 4135
rect 30550 4085 30600 4115
rect 30550 4065 30565 4085
rect 30585 4065 30600 4085
rect 30550 4035 30600 4065
rect 30550 4015 30565 4035
rect 30585 4015 30600 4035
rect 30550 3985 30600 4015
rect 30550 3965 30565 3985
rect 30585 3965 30600 3985
rect 30550 3935 30600 3965
rect 30550 3915 30565 3935
rect 30585 3915 30600 3935
rect 30550 3885 30600 3915
rect 30550 3865 30565 3885
rect 30585 3865 30600 3885
rect 30550 3835 30600 3865
rect 30550 3815 30565 3835
rect 30585 3815 30600 3835
rect 30550 3785 30600 3815
rect 30550 3765 30565 3785
rect 30585 3765 30600 3785
rect 30550 3735 30600 3765
rect 30550 3715 30565 3735
rect 30585 3715 30600 3735
rect 30550 3700 30600 3715
rect 30700 4185 30750 4200
rect 30700 4165 30715 4185
rect 30735 4165 30750 4185
rect 30700 4135 30750 4165
rect 30700 4115 30715 4135
rect 30735 4115 30750 4135
rect 30700 4085 30750 4115
rect 30700 4065 30715 4085
rect 30735 4065 30750 4085
rect 30700 4035 30750 4065
rect 30700 4015 30715 4035
rect 30735 4015 30750 4035
rect 30700 3985 30750 4015
rect 30700 3965 30715 3985
rect 30735 3965 30750 3985
rect 30700 3935 30750 3965
rect 30700 3915 30715 3935
rect 30735 3915 30750 3935
rect 30700 3885 30750 3915
rect 30700 3865 30715 3885
rect 30735 3865 30750 3885
rect 30700 3835 30750 3865
rect 30700 3815 30715 3835
rect 30735 3815 30750 3835
rect 30700 3785 30750 3815
rect 30700 3765 30715 3785
rect 30735 3765 30750 3785
rect 30700 3735 30750 3765
rect 30700 3715 30715 3735
rect 30735 3715 30750 3735
rect 30700 3700 30750 3715
rect 30850 4185 30900 4200
rect 30850 4165 30865 4185
rect 30885 4165 30900 4185
rect 30850 4135 30900 4165
rect 30850 4115 30865 4135
rect 30885 4115 30900 4135
rect 30850 4085 30900 4115
rect 30850 4065 30865 4085
rect 30885 4065 30900 4085
rect 30850 4035 30900 4065
rect 30850 4015 30865 4035
rect 30885 4015 30900 4035
rect 30850 3985 30900 4015
rect 30850 3965 30865 3985
rect 30885 3965 30900 3985
rect 30850 3935 30900 3965
rect 30850 3915 30865 3935
rect 30885 3915 30900 3935
rect 30850 3885 30900 3915
rect 30850 3865 30865 3885
rect 30885 3865 30900 3885
rect 30850 3835 30900 3865
rect 30850 3815 30865 3835
rect 30885 3815 30900 3835
rect 30850 3785 30900 3815
rect 30850 3765 30865 3785
rect 30885 3765 30900 3785
rect 30850 3735 30900 3765
rect 30850 3715 30865 3735
rect 30885 3715 30900 3735
rect 30850 3700 30900 3715
rect 31000 4185 31050 4200
rect 31000 4165 31015 4185
rect 31035 4165 31050 4185
rect 31000 4135 31050 4165
rect 31000 4115 31015 4135
rect 31035 4115 31050 4135
rect 31000 4085 31050 4115
rect 31000 4065 31015 4085
rect 31035 4065 31050 4085
rect 31000 4035 31050 4065
rect 31000 4015 31015 4035
rect 31035 4015 31050 4035
rect 31000 3985 31050 4015
rect 31000 3965 31015 3985
rect 31035 3965 31050 3985
rect 31000 3935 31050 3965
rect 31000 3915 31015 3935
rect 31035 3915 31050 3935
rect 31000 3885 31050 3915
rect 31000 3865 31015 3885
rect 31035 3865 31050 3885
rect 31000 3835 31050 3865
rect 31000 3815 31015 3835
rect 31035 3815 31050 3835
rect 31000 3785 31050 3815
rect 31000 3765 31015 3785
rect 31035 3765 31050 3785
rect 31000 3735 31050 3765
rect 31000 3715 31015 3735
rect 31035 3715 31050 3735
rect 31000 3700 31050 3715
rect 31150 4185 31200 4200
rect 31150 4165 31165 4185
rect 31185 4165 31200 4185
rect 31150 4135 31200 4165
rect 31150 4115 31165 4135
rect 31185 4115 31200 4135
rect 31150 4085 31200 4115
rect 31150 4065 31165 4085
rect 31185 4065 31200 4085
rect 31150 4035 31200 4065
rect 31150 4015 31165 4035
rect 31185 4015 31200 4035
rect 31150 3985 31200 4015
rect 31150 3965 31165 3985
rect 31185 3965 31200 3985
rect 31150 3935 31200 3965
rect 31150 3915 31165 3935
rect 31185 3915 31200 3935
rect 31150 3885 31200 3915
rect 31150 3865 31165 3885
rect 31185 3865 31200 3885
rect 31150 3835 31200 3865
rect 31150 3815 31165 3835
rect 31185 3815 31200 3835
rect 31150 3785 31200 3815
rect 31150 3765 31165 3785
rect 31185 3765 31200 3785
rect 31150 3735 31200 3765
rect 31150 3715 31165 3735
rect 31185 3715 31200 3735
rect 31150 3700 31200 3715
rect 31300 4185 31350 4200
rect 31300 4165 31315 4185
rect 31335 4165 31350 4185
rect 31300 4135 31350 4165
rect 31300 4115 31315 4135
rect 31335 4115 31350 4135
rect 31300 4085 31350 4115
rect 31300 4065 31315 4085
rect 31335 4065 31350 4085
rect 31300 4035 31350 4065
rect 31300 4015 31315 4035
rect 31335 4015 31350 4035
rect 31300 3985 31350 4015
rect 31300 3965 31315 3985
rect 31335 3965 31350 3985
rect 31300 3935 31350 3965
rect 31300 3915 31315 3935
rect 31335 3915 31350 3935
rect 31300 3885 31350 3915
rect 31300 3865 31315 3885
rect 31335 3865 31350 3885
rect 31300 3835 31350 3865
rect 31300 3815 31315 3835
rect 31335 3815 31350 3835
rect 31300 3785 31350 3815
rect 31300 3765 31315 3785
rect 31335 3765 31350 3785
rect 31300 3735 31350 3765
rect 31300 3715 31315 3735
rect 31335 3715 31350 3735
rect 31300 3700 31350 3715
rect 31450 4185 31500 4200
rect 31450 4165 31465 4185
rect 31485 4165 31500 4185
rect 31450 4135 31500 4165
rect 31450 4115 31465 4135
rect 31485 4115 31500 4135
rect 31450 4085 31500 4115
rect 31450 4065 31465 4085
rect 31485 4065 31500 4085
rect 31450 4035 31500 4065
rect 31450 4015 31465 4035
rect 31485 4015 31500 4035
rect 31450 3985 31500 4015
rect 31450 3965 31465 3985
rect 31485 3965 31500 3985
rect 31450 3935 31500 3965
rect 31450 3915 31465 3935
rect 31485 3915 31500 3935
rect 31450 3885 31500 3915
rect 31450 3865 31465 3885
rect 31485 3865 31500 3885
rect 31450 3835 31500 3865
rect 31450 3815 31465 3835
rect 31485 3815 31500 3835
rect 31450 3785 31500 3815
rect 31450 3765 31465 3785
rect 31485 3765 31500 3785
rect 31450 3735 31500 3765
rect 31450 3715 31465 3735
rect 31485 3715 31500 3735
rect 31450 3700 31500 3715
rect 32050 4185 32100 4200
rect 32050 4165 32065 4185
rect 32085 4165 32100 4185
rect 32050 4135 32100 4165
rect 32050 4115 32065 4135
rect 32085 4115 32100 4135
rect 32050 4085 32100 4115
rect 32050 4065 32065 4085
rect 32085 4065 32100 4085
rect 32050 4035 32100 4065
rect 32050 4015 32065 4035
rect 32085 4015 32100 4035
rect 32050 3985 32100 4015
rect 32050 3965 32065 3985
rect 32085 3965 32100 3985
rect 32050 3935 32100 3965
rect 32050 3915 32065 3935
rect 32085 3915 32100 3935
rect 32050 3885 32100 3915
rect 32050 3865 32065 3885
rect 32085 3865 32100 3885
rect 32050 3835 32100 3865
rect 32050 3815 32065 3835
rect 32085 3815 32100 3835
rect 32050 3785 32100 3815
rect 32050 3765 32065 3785
rect 32085 3765 32100 3785
rect 32050 3735 32100 3765
rect 32050 3715 32065 3735
rect 32085 3715 32100 3735
rect 32050 3700 32100 3715
rect -600 3635 -350 3650
rect -600 3615 -585 3635
rect -565 3615 -535 3635
rect -515 3615 -485 3635
rect -465 3615 -435 3635
rect -415 3615 -385 3635
rect -365 3615 -350 3635
rect -600 3600 -350 3615
rect -300 3635 -50 3650
rect -300 3615 -285 3635
rect -265 3615 -235 3635
rect -215 3615 -185 3635
rect -165 3615 -135 3635
rect -115 3615 -85 3635
rect -65 3615 -50 3635
rect -300 3600 -50 3615
rect 0 3635 250 3650
rect 0 3615 15 3635
rect 35 3615 65 3635
rect 85 3615 115 3635
rect 135 3615 165 3635
rect 185 3615 215 3635
rect 235 3615 250 3635
rect 0 3600 250 3615
rect 300 3635 550 3650
rect 300 3615 315 3635
rect 335 3615 365 3635
rect 385 3615 415 3635
rect 435 3615 465 3635
rect 485 3615 515 3635
rect 535 3615 550 3635
rect 300 3600 550 3615
rect 600 3635 850 3650
rect 600 3615 615 3635
rect 635 3615 665 3635
rect 685 3615 715 3635
rect 735 3615 765 3635
rect 785 3615 815 3635
rect 835 3615 850 3635
rect 600 3600 850 3615
rect 900 3635 1150 3650
rect 900 3615 915 3635
rect 935 3615 965 3635
rect 985 3615 1015 3635
rect 1035 3615 1065 3635
rect 1085 3615 1115 3635
rect 1135 3615 1150 3635
rect 900 3600 1150 3615
rect 1200 3635 1450 3650
rect 1200 3615 1215 3635
rect 1235 3615 1265 3635
rect 1285 3615 1315 3635
rect 1335 3615 1365 3635
rect 1385 3615 1415 3635
rect 1435 3615 1450 3635
rect 1200 3600 1450 3615
rect 1500 3635 1750 3650
rect 1500 3615 1515 3635
rect 1535 3615 1565 3635
rect 1585 3615 1615 3635
rect 1635 3615 1665 3635
rect 1685 3615 1715 3635
rect 1735 3615 1750 3635
rect 1500 3600 1750 3615
rect 1800 3635 2050 3650
rect 1800 3615 1815 3635
rect 1835 3615 1865 3635
rect 1885 3615 1915 3635
rect 1935 3615 1965 3635
rect 1985 3615 2015 3635
rect 2035 3615 2050 3635
rect 1800 3600 2050 3615
rect 2100 3635 2350 3650
rect 2100 3615 2115 3635
rect 2135 3615 2165 3635
rect 2185 3615 2215 3635
rect 2235 3615 2265 3635
rect 2285 3615 2315 3635
rect 2335 3615 2350 3635
rect 2100 3600 2350 3615
rect 2400 3635 2650 3650
rect 2400 3615 2415 3635
rect 2435 3615 2465 3635
rect 2485 3615 2515 3635
rect 2535 3615 2565 3635
rect 2585 3615 2615 3635
rect 2635 3615 2650 3635
rect 2400 3600 2650 3615
rect 2700 3635 2950 3650
rect 2700 3615 2715 3635
rect 2735 3615 2765 3635
rect 2785 3615 2815 3635
rect 2835 3615 2865 3635
rect 2885 3615 2915 3635
rect 2935 3615 2950 3635
rect 2700 3600 2950 3615
rect 3000 3635 3250 3650
rect 3000 3615 3015 3635
rect 3035 3615 3065 3635
rect 3085 3615 3115 3635
rect 3135 3615 3165 3635
rect 3185 3615 3215 3635
rect 3235 3615 3250 3635
rect 3000 3600 3250 3615
rect 3300 3635 3550 3650
rect 3300 3615 3315 3635
rect 3335 3615 3365 3635
rect 3385 3615 3415 3635
rect 3435 3615 3465 3635
rect 3485 3615 3515 3635
rect 3535 3615 3550 3635
rect 3300 3600 3550 3615
rect 3600 3635 3850 3650
rect 3600 3615 3615 3635
rect 3635 3615 3665 3635
rect 3685 3615 3715 3635
rect 3735 3615 3765 3635
rect 3785 3615 3815 3635
rect 3835 3615 3850 3635
rect 3600 3600 3850 3615
rect 3900 3635 4150 3650
rect 3900 3615 3915 3635
rect 3935 3615 3965 3635
rect 3985 3615 4015 3635
rect 4035 3615 4065 3635
rect 4085 3615 4115 3635
rect 4135 3615 4150 3635
rect 3900 3600 4150 3615
rect 4200 3635 4450 3650
rect 4200 3615 4215 3635
rect 4235 3615 4265 3635
rect 4285 3615 4315 3635
rect 4335 3615 4365 3635
rect 4385 3615 4415 3635
rect 4435 3615 4450 3635
rect 4200 3600 4450 3615
rect 4500 3635 4750 3650
rect 4500 3615 4515 3635
rect 4535 3615 4565 3635
rect 4585 3615 4615 3635
rect 4635 3615 4665 3635
rect 4685 3615 4715 3635
rect 4735 3615 4750 3635
rect 4500 3600 4750 3615
rect 4800 3635 5050 3650
rect 4800 3615 4815 3635
rect 4835 3615 4865 3635
rect 4885 3615 4915 3635
rect 4935 3615 4965 3635
rect 4985 3615 5015 3635
rect 5035 3615 5050 3635
rect 4800 3600 5050 3615
rect 5100 3635 5350 3650
rect 5100 3615 5115 3635
rect 5135 3615 5165 3635
rect 5185 3615 5215 3635
rect 5235 3615 5265 3635
rect 5285 3615 5315 3635
rect 5335 3615 5350 3635
rect 5100 3600 5350 3615
rect 5400 3635 5650 3650
rect 5400 3615 5415 3635
rect 5435 3615 5465 3635
rect 5485 3615 5515 3635
rect 5535 3615 5565 3635
rect 5585 3615 5615 3635
rect 5635 3615 5650 3635
rect 5400 3600 5650 3615
rect 5700 3635 5950 3650
rect 5700 3615 5715 3635
rect 5735 3615 5765 3635
rect 5785 3615 5815 3635
rect 5835 3615 5865 3635
rect 5885 3615 5915 3635
rect 5935 3615 5950 3635
rect 5700 3600 5950 3615
rect 6000 3635 6250 3650
rect 6000 3615 6015 3635
rect 6035 3615 6065 3635
rect 6085 3615 6115 3635
rect 6135 3615 6165 3635
rect 6185 3615 6215 3635
rect 6235 3615 6250 3635
rect 6000 3600 6250 3615
rect 6300 3635 6550 3650
rect 6300 3615 6315 3635
rect 6335 3615 6365 3635
rect 6385 3615 6415 3635
rect 6435 3615 6465 3635
rect 6485 3615 6515 3635
rect 6535 3615 6550 3635
rect 6300 3600 6550 3615
rect 6600 3635 6850 3650
rect 6600 3615 6615 3635
rect 6635 3615 6665 3635
rect 6685 3615 6715 3635
rect 6735 3615 6765 3635
rect 6785 3615 6815 3635
rect 6835 3615 6850 3635
rect 6600 3600 6850 3615
rect 6900 3635 7150 3650
rect 6900 3615 6915 3635
rect 6935 3615 6965 3635
rect 6985 3615 7015 3635
rect 7035 3615 7065 3635
rect 7085 3615 7115 3635
rect 7135 3615 7150 3635
rect 6900 3600 7150 3615
rect 7200 3635 7450 3650
rect 7200 3615 7215 3635
rect 7235 3615 7265 3635
rect 7285 3615 7315 3635
rect 7335 3615 7365 3635
rect 7385 3615 7415 3635
rect 7435 3615 7450 3635
rect 7200 3600 7450 3615
rect 7500 3635 7750 3650
rect 7500 3615 7515 3635
rect 7535 3615 7565 3635
rect 7585 3615 7615 3635
rect 7635 3615 7665 3635
rect 7685 3615 7715 3635
rect 7735 3615 7750 3635
rect 7500 3600 7750 3615
rect 7800 3635 8050 3650
rect 7800 3615 7815 3635
rect 7835 3615 7865 3635
rect 7885 3615 7915 3635
rect 7935 3615 7965 3635
rect 7985 3615 8015 3635
rect 8035 3615 8050 3635
rect 7800 3600 8050 3615
rect 8100 3635 8350 3650
rect 8100 3615 8115 3635
rect 8135 3615 8165 3635
rect 8185 3615 8215 3635
rect 8235 3615 8265 3635
rect 8285 3615 8315 3635
rect 8335 3615 8350 3635
rect 8100 3600 8350 3615
rect 8400 3635 10750 3650
rect 8400 3615 8415 3635
rect 8435 3615 8465 3635
rect 8485 3615 8515 3635
rect 8535 3615 8565 3635
rect 8585 3615 8615 3635
rect 8635 3615 8715 3635
rect 8735 3615 8765 3635
rect 8785 3615 8815 3635
rect 8835 3615 8865 3635
rect 8885 3615 8915 3635
rect 8935 3615 9015 3635
rect 9035 3615 9065 3635
rect 9085 3615 9115 3635
rect 9135 3615 9165 3635
rect 9185 3615 9215 3635
rect 9235 3615 9315 3635
rect 9335 3615 9365 3635
rect 9385 3615 9415 3635
rect 9435 3615 9465 3635
rect 9485 3615 9515 3635
rect 9535 3615 9615 3635
rect 9635 3615 9665 3635
rect 9685 3615 9715 3635
rect 9735 3615 9765 3635
rect 9785 3615 9815 3635
rect 9835 3615 9915 3635
rect 9935 3615 9965 3635
rect 9985 3615 10015 3635
rect 10035 3615 10065 3635
rect 10085 3615 10115 3635
rect 10135 3615 10215 3635
rect 10235 3615 10265 3635
rect 10285 3615 10315 3635
rect 10335 3615 10365 3635
rect 10385 3615 10415 3635
rect 10435 3615 10515 3635
rect 10535 3615 10565 3635
rect 10585 3615 10615 3635
rect 10635 3615 10665 3635
rect 10685 3615 10715 3635
rect 10735 3615 10750 3635
rect 8400 3600 10750 3615
rect 10800 3635 11050 3650
rect 10800 3615 10815 3635
rect 10835 3615 10865 3635
rect 10885 3615 10915 3635
rect 10935 3615 10965 3635
rect 10985 3615 11015 3635
rect 11035 3615 11050 3635
rect 10800 3600 11050 3615
rect 11100 3635 11350 3650
rect 11100 3615 11115 3635
rect 11135 3615 11165 3635
rect 11185 3615 11215 3635
rect 11235 3615 11265 3635
rect 11285 3615 11315 3635
rect 11335 3615 11350 3635
rect 11100 3600 11350 3615
rect 11400 3635 11650 3650
rect 11400 3615 11415 3635
rect 11435 3615 11465 3635
rect 11485 3615 11515 3635
rect 11535 3615 11565 3635
rect 11585 3615 11615 3635
rect 11635 3615 11650 3635
rect 11400 3600 11650 3615
rect 11700 3635 11950 3650
rect 11700 3615 11715 3635
rect 11735 3615 11765 3635
rect 11785 3615 11815 3635
rect 11835 3615 11865 3635
rect 11885 3615 11915 3635
rect 11935 3615 11950 3635
rect 11700 3600 11950 3615
rect 12000 3635 12250 3650
rect 12000 3615 12015 3635
rect 12035 3615 12065 3635
rect 12085 3615 12115 3635
rect 12135 3615 12165 3635
rect 12185 3615 12215 3635
rect 12235 3615 12250 3635
rect 12000 3600 12250 3615
rect 12300 3635 12550 3650
rect 12300 3615 12315 3635
rect 12335 3615 12365 3635
rect 12385 3615 12415 3635
rect 12435 3615 12465 3635
rect 12485 3615 12515 3635
rect 12535 3615 12550 3635
rect 12300 3600 12550 3615
rect 12600 3635 12850 3650
rect 12600 3615 12615 3635
rect 12635 3615 12665 3635
rect 12685 3615 12715 3635
rect 12735 3615 12765 3635
rect 12785 3615 12815 3635
rect 12835 3615 12850 3635
rect 12600 3600 12850 3615
rect 12900 3635 13150 3650
rect 12900 3615 12915 3635
rect 12935 3615 12965 3635
rect 12985 3615 13015 3635
rect 13035 3615 13065 3635
rect 13085 3615 13115 3635
rect 13135 3615 13150 3635
rect 12900 3600 13150 3615
rect 13200 3635 13450 3650
rect 13200 3615 13215 3635
rect 13235 3615 13265 3635
rect 13285 3615 13315 3635
rect 13335 3615 13365 3635
rect 13385 3615 13415 3635
rect 13435 3615 13450 3635
rect 13200 3600 13450 3615
rect 13500 3635 13750 3650
rect 13500 3615 13515 3635
rect 13535 3615 13565 3635
rect 13585 3615 13615 3635
rect 13635 3615 13665 3635
rect 13685 3615 13715 3635
rect 13735 3615 13750 3635
rect 13500 3600 13750 3615
rect 13800 3635 14050 3650
rect 13800 3615 13815 3635
rect 13835 3615 13865 3635
rect 13885 3615 13915 3635
rect 13935 3615 13965 3635
rect 13985 3615 14015 3635
rect 14035 3615 14050 3635
rect 13800 3600 14050 3615
rect 14100 3635 14350 3650
rect 14100 3615 14115 3635
rect 14135 3615 14165 3635
rect 14185 3615 14215 3635
rect 14235 3615 14265 3635
rect 14285 3615 14315 3635
rect 14335 3615 14350 3635
rect 14100 3600 14350 3615
rect 14400 3635 14650 3650
rect 14400 3615 14415 3635
rect 14435 3615 14465 3635
rect 14485 3615 14515 3635
rect 14535 3615 14565 3635
rect 14585 3615 14615 3635
rect 14635 3615 14650 3635
rect 14400 3600 14650 3615
rect 14700 3635 14950 3650
rect 14700 3615 14715 3635
rect 14735 3615 14765 3635
rect 14785 3615 14815 3635
rect 14835 3615 14865 3635
rect 14885 3615 14915 3635
rect 14935 3615 14950 3635
rect 14700 3600 14950 3615
rect 15000 3635 15250 3650
rect 15000 3615 15015 3635
rect 15035 3615 15065 3635
rect 15085 3615 15115 3635
rect 15135 3615 15165 3635
rect 15185 3615 15215 3635
rect 15235 3615 15250 3635
rect 15000 3600 15250 3615
rect 15300 3635 15550 3650
rect 15300 3615 15315 3635
rect 15335 3615 15365 3635
rect 15385 3615 15415 3635
rect 15435 3615 15465 3635
rect 15485 3615 15515 3635
rect 15535 3615 15550 3635
rect 15300 3600 15550 3615
rect 15600 3635 15850 3650
rect 15600 3615 15615 3635
rect 15635 3615 15665 3635
rect 15685 3615 15715 3635
rect 15735 3615 15765 3635
rect 15785 3615 15815 3635
rect 15835 3615 15850 3635
rect 15600 3600 15850 3615
rect 15900 3635 16150 3650
rect 15900 3615 15915 3635
rect 15935 3615 15965 3635
rect 15985 3615 16015 3635
rect 16035 3615 16065 3635
rect 16085 3615 16115 3635
rect 16135 3615 16150 3635
rect 15900 3600 16150 3615
rect 16200 3635 16450 3650
rect 16200 3615 16215 3635
rect 16235 3615 16265 3635
rect 16285 3615 16315 3635
rect 16335 3615 16365 3635
rect 16385 3615 16415 3635
rect 16435 3615 16450 3635
rect 16200 3600 16450 3615
rect 16500 3635 16750 3650
rect 16500 3615 16515 3635
rect 16535 3615 16565 3635
rect 16585 3615 16615 3635
rect 16635 3615 16665 3635
rect 16685 3615 16715 3635
rect 16735 3615 16750 3635
rect 16500 3600 16750 3615
rect 16800 3635 17050 3650
rect 16800 3615 16815 3635
rect 16835 3615 16865 3635
rect 16885 3615 16915 3635
rect 16935 3615 16965 3635
rect 16985 3615 17015 3635
rect 17035 3615 17050 3635
rect 16800 3600 17050 3615
rect 17100 3635 17350 3650
rect 17100 3615 17115 3635
rect 17135 3615 17165 3635
rect 17185 3615 17215 3635
rect 17235 3615 17265 3635
rect 17285 3615 17315 3635
rect 17335 3615 17350 3635
rect 17100 3600 17350 3615
rect 17400 3635 17650 3650
rect 17400 3615 17415 3635
rect 17435 3615 17465 3635
rect 17485 3615 17515 3635
rect 17535 3615 17565 3635
rect 17585 3615 17615 3635
rect 17635 3615 17650 3635
rect 17400 3600 17650 3615
rect 17700 3635 17950 3650
rect 17700 3615 17715 3635
rect 17735 3615 17765 3635
rect 17785 3615 17815 3635
rect 17835 3615 17865 3635
rect 17885 3615 17915 3635
rect 17935 3615 17950 3635
rect 17700 3600 17950 3615
rect 18000 3635 18250 3650
rect 18000 3615 18015 3635
rect 18035 3615 18065 3635
rect 18085 3615 18115 3635
rect 18135 3615 18165 3635
rect 18185 3615 18215 3635
rect 18235 3615 18250 3635
rect 18000 3600 18250 3615
rect 18300 3635 18550 3650
rect 18300 3615 18315 3635
rect 18335 3615 18365 3635
rect 18385 3615 18415 3635
rect 18435 3615 18465 3635
rect 18485 3615 18515 3635
rect 18535 3615 18550 3635
rect 18300 3600 18550 3615
rect 18600 3635 18850 3650
rect 18600 3615 18615 3635
rect 18635 3615 18665 3635
rect 18685 3615 18715 3635
rect 18735 3615 18765 3635
rect 18785 3615 18815 3635
rect 18835 3615 18850 3635
rect 18600 3600 18850 3615
rect 18900 3635 19150 3650
rect 18900 3615 18915 3635
rect 18935 3615 18965 3635
rect 18985 3615 19015 3635
rect 19035 3615 19065 3635
rect 19085 3615 19115 3635
rect 19135 3615 19150 3635
rect 18900 3600 19150 3615
rect 19200 3635 19450 3650
rect 19200 3615 19215 3635
rect 19235 3615 19265 3635
rect 19285 3615 19315 3635
rect 19335 3615 19365 3635
rect 19385 3615 19415 3635
rect 19435 3615 19450 3635
rect 19200 3600 19450 3615
rect 19500 3635 19750 3650
rect 19500 3615 19515 3635
rect 19535 3615 19565 3635
rect 19585 3615 19615 3635
rect 19635 3615 19665 3635
rect 19685 3615 19715 3635
rect 19735 3615 19750 3635
rect 19500 3600 19750 3615
rect 19800 3635 20050 3650
rect 19800 3615 19815 3635
rect 19835 3615 19865 3635
rect 19885 3615 19915 3635
rect 19935 3615 19965 3635
rect 19985 3615 20015 3635
rect 20035 3615 20050 3635
rect 19800 3600 20050 3615
rect 20100 3635 20350 3650
rect 20100 3615 20115 3635
rect 20135 3615 20165 3635
rect 20185 3615 20215 3635
rect 20235 3615 20265 3635
rect 20285 3615 20315 3635
rect 20335 3615 20350 3635
rect 20100 3600 20350 3615
rect 20400 3635 20650 3650
rect 20400 3615 20415 3635
rect 20435 3615 20465 3635
rect 20485 3615 20515 3635
rect 20535 3615 20565 3635
rect 20585 3615 20615 3635
rect 20635 3615 20650 3635
rect 20400 3600 20650 3615
rect 20700 3635 20950 3650
rect 20700 3615 20715 3635
rect 20735 3615 20765 3635
rect 20785 3615 20815 3635
rect 20835 3615 20865 3635
rect 20885 3615 20915 3635
rect 20935 3615 20950 3635
rect 20700 3600 20950 3615
rect 21000 3635 21400 3650
rect 21000 3615 21015 3635
rect 21035 3615 21065 3635
rect 21085 3615 21115 3635
rect 21135 3615 21165 3635
rect 21185 3615 21215 3635
rect 21235 3615 21265 3635
rect 21285 3615 21315 3635
rect 21335 3615 21365 3635
rect 21385 3615 21400 3635
rect 21000 3600 21400 3615
rect 21450 3635 21850 3650
rect 21450 3615 21465 3635
rect 21485 3615 21515 3635
rect 21535 3615 21565 3635
rect 21585 3615 21615 3635
rect 21635 3615 21665 3635
rect 21685 3615 21715 3635
rect 21735 3615 21765 3635
rect 21785 3615 21815 3635
rect 21835 3615 21850 3635
rect 21450 3600 21850 3615
rect 21900 3635 22150 3650
rect 21900 3615 21915 3635
rect 21935 3615 21965 3635
rect 21985 3615 22015 3635
rect 22035 3615 22065 3635
rect 22085 3615 22115 3635
rect 22135 3615 22150 3635
rect 21900 3600 22150 3615
rect 22200 3635 22450 3650
rect 22200 3615 22215 3635
rect 22235 3615 22265 3635
rect 22285 3615 22315 3635
rect 22335 3615 22365 3635
rect 22385 3615 22415 3635
rect 22435 3615 22450 3635
rect 22200 3600 22450 3615
rect 22500 3635 22750 3650
rect 22500 3615 22515 3635
rect 22535 3615 22565 3635
rect 22585 3615 22615 3635
rect 22635 3615 22665 3635
rect 22685 3615 22715 3635
rect 22735 3615 22750 3635
rect 22500 3600 22750 3615
rect 22800 3635 23050 3650
rect 22800 3615 22815 3635
rect 22835 3615 22865 3635
rect 22885 3615 22915 3635
rect 22935 3615 22965 3635
rect 22985 3615 23015 3635
rect 23035 3615 23050 3635
rect 22800 3600 23050 3615
rect 23100 3635 23500 3650
rect 23100 3615 23115 3635
rect 23135 3615 23165 3635
rect 23185 3615 23215 3635
rect 23235 3615 23265 3635
rect 23285 3615 23315 3635
rect 23335 3615 23365 3635
rect 23385 3615 23415 3635
rect 23435 3615 23465 3635
rect 23485 3615 23500 3635
rect 23100 3600 23500 3615
rect 23550 3635 23950 3650
rect 23550 3615 23565 3635
rect 23585 3615 23615 3635
rect 23635 3615 23665 3635
rect 23685 3615 23715 3635
rect 23735 3615 23765 3635
rect 23785 3615 23815 3635
rect 23835 3615 23865 3635
rect 23885 3615 23915 3635
rect 23935 3615 23950 3635
rect 23550 3600 23950 3615
rect 24000 3635 24250 3650
rect 24000 3615 24015 3635
rect 24035 3615 24065 3635
rect 24085 3615 24115 3635
rect 24135 3615 24165 3635
rect 24185 3615 24215 3635
rect 24235 3615 24250 3635
rect 24000 3600 24250 3615
rect 24300 3635 24550 3650
rect 24300 3615 24315 3635
rect 24335 3615 24365 3635
rect 24385 3615 24415 3635
rect 24435 3615 24465 3635
rect 24485 3615 24515 3635
rect 24535 3615 24550 3635
rect 24300 3600 24550 3615
rect 24600 3635 24850 3650
rect 24600 3615 24615 3635
rect 24635 3615 24665 3635
rect 24685 3615 24715 3635
rect 24735 3615 24765 3635
rect 24785 3615 24815 3635
rect 24835 3615 24850 3635
rect 24600 3600 24850 3615
rect 24900 3635 25150 3650
rect 24900 3615 24915 3635
rect 24935 3615 24965 3635
rect 24985 3615 25015 3635
rect 25035 3615 25065 3635
rect 25085 3615 25115 3635
rect 25135 3615 25150 3635
rect 24900 3600 25150 3615
rect 25200 3635 25600 3650
rect 25200 3615 25215 3635
rect 25235 3615 25265 3635
rect 25285 3615 25315 3635
rect 25335 3615 25365 3635
rect 25385 3615 25415 3635
rect 25435 3615 25465 3635
rect 25485 3615 25515 3635
rect 25535 3615 25565 3635
rect 25585 3615 25600 3635
rect 25200 3600 25600 3615
rect 25650 3635 26050 3650
rect 25650 3615 25665 3635
rect 25685 3615 25715 3635
rect 25735 3615 25765 3635
rect 25785 3615 25815 3635
rect 25835 3615 25865 3635
rect 25885 3615 25915 3635
rect 25935 3615 25965 3635
rect 25985 3615 26015 3635
rect 26035 3615 26050 3635
rect 25650 3600 26050 3615
rect 26100 3635 26350 3650
rect 26100 3615 26115 3635
rect 26135 3615 26165 3635
rect 26185 3615 26215 3635
rect 26235 3615 26265 3635
rect 26285 3615 26315 3635
rect 26335 3615 26350 3635
rect 26100 3600 26350 3615
rect 26400 3635 26650 3650
rect 26400 3615 26415 3635
rect 26435 3615 26465 3635
rect 26485 3615 26515 3635
rect 26535 3615 26565 3635
rect 26585 3615 26615 3635
rect 26635 3615 26650 3635
rect 26400 3600 26650 3615
rect 26700 3635 26950 3650
rect 26700 3615 26715 3635
rect 26735 3615 26765 3635
rect 26785 3615 26815 3635
rect 26835 3615 26865 3635
rect 26885 3615 26915 3635
rect 26935 3615 26950 3635
rect 26700 3600 26950 3615
rect 27000 3635 27250 3650
rect 27000 3615 27015 3635
rect 27035 3615 27065 3635
rect 27085 3615 27115 3635
rect 27135 3615 27165 3635
rect 27185 3615 27215 3635
rect 27235 3615 27250 3635
rect 27000 3600 27250 3615
rect 27300 3635 27700 3650
rect 27300 3615 27315 3635
rect 27335 3615 27365 3635
rect 27385 3615 27415 3635
rect 27435 3615 27465 3635
rect 27485 3615 27515 3635
rect 27535 3615 27565 3635
rect 27585 3615 27615 3635
rect 27635 3615 27665 3635
rect 27685 3615 27700 3635
rect 27300 3600 27700 3615
rect 27750 3635 28150 3650
rect 27750 3615 27765 3635
rect 27785 3615 27815 3635
rect 27835 3615 27865 3635
rect 27885 3615 27915 3635
rect 27935 3615 27965 3635
rect 27985 3615 28015 3635
rect 28035 3615 28065 3635
rect 28085 3615 28115 3635
rect 28135 3615 28150 3635
rect 27750 3600 28150 3615
rect 28200 3635 28450 3650
rect 28200 3615 28215 3635
rect 28235 3615 28265 3635
rect 28285 3615 28315 3635
rect 28335 3615 28365 3635
rect 28385 3615 28415 3635
rect 28435 3615 28450 3635
rect 28200 3600 28450 3615
rect 28500 3635 28750 3650
rect 28500 3615 28515 3635
rect 28535 3615 28565 3635
rect 28585 3615 28615 3635
rect 28635 3615 28665 3635
rect 28685 3615 28715 3635
rect 28735 3615 28750 3635
rect 28500 3600 28750 3615
rect 28800 3635 29050 3650
rect 28800 3615 28815 3635
rect 28835 3615 28865 3635
rect 28885 3615 28915 3635
rect 28935 3615 28965 3635
rect 28985 3615 29015 3635
rect 29035 3615 29050 3635
rect 28800 3600 29050 3615
rect 29100 3635 29350 3650
rect 29100 3615 29115 3635
rect 29135 3615 29165 3635
rect 29185 3615 29215 3635
rect 29235 3615 29265 3635
rect 29285 3615 29315 3635
rect 29335 3615 29350 3635
rect 29100 3600 29350 3615
rect 29400 3635 29800 3650
rect 29400 3615 29415 3635
rect 29435 3615 29465 3635
rect 29485 3615 29515 3635
rect 29535 3615 29565 3635
rect 29585 3615 29615 3635
rect 29635 3615 29665 3635
rect 29685 3615 29715 3635
rect 29735 3615 29765 3635
rect 29785 3615 29800 3635
rect 29400 3600 29800 3615
rect 29850 3635 30100 3650
rect 29850 3615 29865 3635
rect 29885 3615 29915 3635
rect 29935 3615 29965 3635
rect 29985 3615 30015 3635
rect 30035 3615 30065 3635
rect 30085 3615 30100 3635
rect 29850 3600 30100 3615
rect 30150 3635 30400 3650
rect 30150 3615 30165 3635
rect 30185 3615 30215 3635
rect 30235 3615 30265 3635
rect 30285 3615 30315 3635
rect 30335 3615 30365 3635
rect 30385 3615 30400 3635
rect 30150 3600 30400 3615
rect 30450 3635 30700 3650
rect 30450 3615 30465 3635
rect 30485 3615 30515 3635
rect 30535 3615 30565 3635
rect 30585 3615 30615 3635
rect 30635 3615 30665 3635
rect 30685 3615 30700 3635
rect 30450 3600 30700 3615
rect 30750 3635 31000 3650
rect 30750 3615 30765 3635
rect 30785 3615 30815 3635
rect 30835 3615 30865 3635
rect 30885 3615 30915 3635
rect 30935 3615 30965 3635
rect 30985 3615 31000 3635
rect 30750 3600 31000 3615
rect 31050 3635 31450 3650
rect 31050 3615 31065 3635
rect 31085 3615 31115 3635
rect 31135 3615 31165 3635
rect 31185 3615 31215 3635
rect 31235 3615 31265 3635
rect 31285 3615 31315 3635
rect 31335 3615 31365 3635
rect 31385 3615 31415 3635
rect 31435 3615 31450 3635
rect 31050 3600 31450 3615
rect 31500 3635 31750 3650
rect 31500 3615 31515 3635
rect 31535 3615 31565 3635
rect 31585 3615 31615 3635
rect 31635 3615 31665 3635
rect 31685 3615 31715 3635
rect 31735 3615 31750 3635
rect 31500 3600 31750 3615
rect 31800 3635 32050 3650
rect 31800 3615 31815 3635
rect 31835 3615 31865 3635
rect 31885 3615 31915 3635
rect 31935 3615 31965 3635
rect 31985 3615 32015 3635
rect 32035 3615 32050 3635
rect 31800 3600 32050 3615
rect -650 3535 -600 3550
rect -650 3515 -635 3535
rect -615 3515 -600 3535
rect -650 3485 -600 3515
rect -650 3465 -635 3485
rect -615 3465 -600 3485
rect -650 3435 -600 3465
rect -650 3415 -635 3435
rect -615 3415 -600 3435
rect -650 3385 -600 3415
rect -650 3365 -635 3385
rect -615 3365 -600 3385
rect -650 3335 -600 3365
rect -650 3315 -635 3335
rect -615 3315 -600 3335
rect -650 3285 -600 3315
rect -650 3265 -635 3285
rect -615 3265 -600 3285
rect -650 3235 -600 3265
rect -650 3215 -635 3235
rect -615 3215 -600 3235
rect -650 3185 -600 3215
rect -650 3165 -635 3185
rect -615 3165 -600 3185
rect -650 3135 -600 3165
rect -650 3115 -635 3135
rect -615 3115 -600 3135
rect -650 3085 -600 3115
rect -650 3065 -635 3085
rect -615 3065 -600 3085
rect -650 3050 -600 3065
rect -500 3535 -450 3550
rect -500 3515 -485 3535
rect -465 3515 -450 3535
rect -500 3485 -450 3515
rect -500 3465 -485 3485
rect -465 3465 -450 3485
rect -500 3435 -450 3465
rect -500 3415 -485 3435
rect -465 3415 -450 3435
rect -500 3385 -450 3415
rect -500 3365 -485 3385
rect -465 3365 -450 3385
rect -500 3335 -450 3365
rect -500 3315 -485 3335
rect -465 3315 -450 3335
rect -500 3285 -450 3315
rect -500 3265 -485 3285
rect -465 3265 -450 3285
rect -500 3235 -450 3265
rect -500 3215 -485 3235
rect -465 3215 -450 3235
rect -500 3185 -450 3215
rect -500 3165 -485 3185
rect -465 3165 -450 3185
rect -500 3135 -450 3165
rect -500 3115 -485 3135
rect -465 3115 -450 3135
rect -500 3085 -450 3115
rect -500 3065 -485 3085
rect -465 3065 -450 3085
rect -500 3050 -450 3065
rect -350 3535 -300 3550
rect -350 3515 -335 3535
rect -315 3515 -300 3535
rect -350 3485 -300 3515
rect -350 3465 -335 3485
rect -315 3465 -300 3485
rect -350 3435 -300 3465
rect -350 3415 -335 3435
rect -315 3415 -300 3435
rect -350 3385 -300 3415
rect -350 3365 -335 3385
rect -315 3365 -300 3385
rect -350 3335 -300 3365
rect -350 3315 -335 3335
rect -315 3315 -300 3335
rect -350 3285 -300 3315
rect -350 3265 -335 3285
rect -315 3265 -300 3285
rect -350 3235 -300 3265
rect -350 3215 -335 3235
rect -315 3215 -300 3235
rect -350 3185 -300 3215
rect -350 3165 -335 3185
rect -315 3165 -300 3185
rect -350 3135 -300 3165
rect -350 3115 -335 3135
rect -315 3115 -300 3135
rect -350 3085 -300 3115
rect -350 3065 -335 3085
rect -315 3065 -300 3085
rect -350 3050 -300 3065
rect -200 3535 -150 3550
rect -200 3515 -185 3535
rect -165 3515 -150 3535
rect -200 3485 -150 3515
rect -200 3465 -185 3485
rect -165 3465 -150 3485
rect -200 3435 -150 3465
rect -200 3415 -185 3435
rect -165 3415 -150 3435
rect -200 3385 -150 3415
rect -200 3365 -185 3385
rect -165 3365 -150 3385
rect -200 3335 -150 3365
rect -200 3315 -185 3335
rect -165 3315 -150 3335
rect -200 3285 -150 3315
rect -200 3265 -185 3285
rect -165 3265 -150 3285
rect -200 3235 -150 3265
rect -200 3215 -185 3235
rect -165 3215 -150 3235
rect -200 3185 -150 3215
rect -200 3165 -185 3185
rect -165 3165 -150 3185
rect -200 3135 -150 3165
rect -200 3115 -185 3135
rect -165 3115 -150 3135
rect -200 3085 -150 3115
rect -200 3065 -185 3085
rect -165 3065 -150 3085
rect -200 3050 -150 3065
rect -50 3535 0 3550
rect -50 3515 -35 3535
rect -15 3515 0 3535
rect -50 3485 0 3515
rect -50 3465 -35 3485
rect -15 3465 0 3485
rect -50 3435 0 3465
rect -50 3415 -35 3435
rect -15 3415 0 3435
rect -50 3385 0 3415
rect -50 3365 -35 3385
rect -15 3365 0 3385
rect -50 3335 0 3365
rect -50 3315 -35 3335
rect -15 3315 0 3335
rect -50 3285 0 3315
rect -50 3265 -35 3285
rect -15 3265 0 3285
rect -50 3235 0 3265
rect -50 3215 -35 3235
rect -15 3215 0 3235
rect -50 3185 0 3215
rect -50 3165 -35 3185
rect -15 3165 0 3185
rect -50 3135 0 3165
rect -50 3115 -35 3135
rect -15 3115 0 3135
rect -50 3085 0 3115
rect -50 3065 -35 3085
rect -15 3065 0 3085
rect -50 3050 0 3065
rect 550 3535 600 3550
rect 550 3515 565 3535
rect 585 3515 600 3535
rect 550 3485 600 3515
rect 550 3465 565 3485
rect 585 3465 600 3485
rect 550 3435 600 3465
rect 550 3415 565 3435
rect 585 3415 600 3435
rect 550 3385 600 3415
rect 550 3365 565 3385
rect 585 3365 600 3385
rect 550 3335 600 3365
rect 550 3315 565 3335
rect 585 3315 600 3335
rect 550 3285 600 3315
rect 550 3265 565 3285
rect 585 3265 600 3285
rect 550 3235 600 3265
rect 550 3215 565 3235
rect 585 3215 600 3235
rect 550 3185 600 3215
rect 550 3165 565 3185
rect 585 3165 600 3185
rect 550 3135 600 3165
rect 550 3115 565 3135
rect 585 3115 600 3135
rect 550 3085 600 3115
rect 550 3065 565 3085
rect 585 3065 600 3085
rect 550 3050 600 3065
rect 700 3535 750 3550
rect 700 3515 715 3535
rect 735 3515 750 3535
rect 700 3485 750 3515
rect 700 3465 715 3485
rect 735 3465 750 3485
rect 700 3435 750 3465
rect 700 3415 715 3435
rect 735 3415 750 3435
rect 700 3385 750 3415
rect 700 3365 715 3385
rect 735 3365 750 3385
rect 700 3335 750 3365
rect 700 3315 715 3335
rect 735 3315 750 3335
rect 700 3285 750 3315
rect 700 3265 715 3285
rect 735 3265 750 3285
rect 700 3235 750 3265
rect 700 3215 715 3235
rect 735 3215 750 3235
rect 700 3185 750 3215
rect 700 3165 715 3185
rect 735 3165 750 3185
rect 700 3135 750 3165
rect 700 3115 715 3135
rect 735 3115 750 3135
rect 700 3085 750 3115
rect 700 3065 715 3085
rect 735 3065 750 3085
rect 700 3050 750 3065
rect 850 3535 900 3550
rect 850 3515 865 3535
rect 885 3515 900 3535
rect 850 3485 900 3515
rect 850 3465 865 3485
rect 885 3465 900 3485
rect 850 3435 900 3465
rect 850 3415 865 3435
rect 885 3415 900 3435
rect 850 3385 900 3415
rect 850 3365 865 3385
rect 885 3365 900 3385
rect 850 3335 900 3365
rect 850 3315 865 3335
rect 885 3315 900 3335
rect 850 3285 900 3315
rect 850 3265 865 3285
rect 885 3265 900 3285
rect 850 3235 900 3265
rect 850 3215 865 3235
rect 885 3215 900 3235
rect 850 3185 900 3215
rect 850 3165 865 3185
rect 885 3165 900 3185
rect 850 3135 900 3165
rect 850 3115 865 3135
rect 885 3115 900 3135
rect 850 3085 900 3115
rect 850 3065 865 3085
rect 885 3065 900 3085
rect 850 3050 900 3065
rect 1000 3535 1050 3550
rect 1000 3515 1015 3535
rect 1035 3515 1050 3535
rect 1000 3485 1050 3515
rect 1000 3465 1015 3485
rect 1035 3465 1050 3485
rect 1000 3435 1050 3465
rect 1000 3415 1015 3435
rect 1035 3415 1050 3435
rect 1000 3385 1050 3415
rect 1000 3365 1015 3385
rect 1035 3365 1050 3385
rect 1000 3335 1050 3365
rect 1000 3315 1015 3335
rect 1035 3315 1050 3335
rect 1000 3285 1050 3315
rect 1000 3265 1015 3285
rect 1035 3265 1050 3285
rect 1000 3235 1050 3265
rect 1000 3215 1015 3235
rect 1035 3215 1050 3235
rect 1000 3185 1050 3215
rect 1000 3165 1015 3185
rect 1035 3165 1050 3185
rect 1000 3135 1050 3165
rect 1000 3115 1015 3135
rect 1035 3115 1050 3135
rect 1000 3085 1050 3115
rect 1000 3065 1015 3085
rect 1035 3065 1050 3085
rect 1000 3050 1050 3065
rect 1150 3535 1200 3550
rect 1150 3515 1165 3535
rect 1185 3515 1200 3535
rect 1150 3485 1200 3515
rect 1150 3465 1165 3485
rect 1185 3465 1200 3485
rect 1150 3435 1200 3465
rect 1150 3415 1165 3435
rect 1185 3415 1200 3435
rect 1150 3385 1200 3415
rect 1150 3365 1165 3385
rect 1185 3365 1200 3385
rect 1150 3335 1200 3365
rect 1150 3315 1165 3335
rect 1185 3315 1200 3335
rect 1150 3285 1200 3315
rect 1150 3265 1165 3285
rect 1185 3265 1200 3285
rect 1150 3235 1200 3265
rect 1150 3215 1165 3235
rect 1185 3215 1200 3235
rect 1150 3185 1200 3215
rect 1150 3165 1165 3185
rect 1185 3165 1200 3185
rect 1150 3135 1200 3165
rect 1150 3115 1165 3135
rect 1185 3115 1200 3135
rect 1150 3085 1200 3115
rect 1150 3065 1165 3085
rect 1185 3065 1200 3085
rect 1150 3050 1200 3065
rect 1300 3535 1350 3550
rect 1300 3515 1315 3535
rect 1335 3515 1350 3535
rect 1300 3485 1350 3515
rect 1300 3465 1315 3485
rect 1335 3465 1350 3485
rect 1300 3435 1350 3465
rect 1300 3415 1315 3435
rect 1335 3415 1350 3435
rect 1300 3385 1350 3415
rect 1300 3365 1315 3385
rect 1335 3365 1350 3385
rect 1300 3335 1350 3365
rect 1300 3315 1315 3335
rect 1335 3315 1350 3335
rect 1300 3285 1350 3315
rect 1300 3265 1315 3285
rect 1335 3265 1350 3285
rect 1300 3235 1350 3265
rect 1300 3215 1315 3235
rect 1335 3215 1350 3235
rect 1300 3185 1350 3215
rect 1300 3165 1315 3185
rect 1335 3165 1350 3185
rect 1300 3135 1350 3165
rect 1300 3115 1315 3135
rect 1335 3115 1350 3135
rect 1300 3085 1350 3115
rect 1300 3065 1315 3085
rect 1335 3065 1350 3085
rect 1300 3050 1350 3065
rect 1450 3535 1500 3550
rect 1450 3515 1465 3535
rect 1485 3515 1500 3535
rect 1450 3485 1500 3515
rect 1450 3465 1465 3485
rect 1485 3465 1500 3485
rect 1450 3435 1500 3465
rect 1450 3415 1465 3435
rect 1485 3415 1500 3435
rect 1450 3385 1500 3415
rect 1450 3365 1465 3385
rect 1485 3365 1500 3385
rect 1450 3335 1500 3365
rect 1450 3315 1465 3335
rect 1485 3315 1500 3335
rect 1450 3285 1500 3315
rect 1450 3265 1465 3285
rect 1485 3265 1500 3285
rect 1450 3235 1500 3265
rect 1450 3215 1465 3235
rect 1485 3215 1500 3235
rect 1450 3185 1500 3215
rect 1450 3165 1465 3185
rect 1485 3165 1500 3185
rect 1450 3135 1500 3165
rect 1450 3115 1465 3135
rect 1485 3115 1500 3135
rect 1450 3085 1500 3115
rect 1450 3065 1465 3085
rect 1485 3065 1500 3085
rect 1450 3050 1500 3065
rect 1600 3535 1650 3550
rect 1600 3515 1615 3535
rect 1635 3515 1650 3535
rect 1600 3485 1650 3515
rect 1600 3465 1615 3485
rect 1635 3465 1650 3485
rect 1600 3435 1650 3465
rect 1600 3415 1615 3435
rect 1635 3415 1650 3435
rect 1600 3385 1650 3415
rect 1600 3365 1615 3385
rect 1635 3365 1650 3385
rect 1600 3335 1650 3365
rect 1600 3315 1615 3335
rect 1635 3315 1650 3335
rect 1600 3285 1650 3315
rect 1600 3265 1615 3285
rect 1635 3265 1650 3285
rect 1600 3235 1650 3265
rect 1600 3215 1615 3235
rect 1635 3215 1650 3235
rect 1600 3185 1650 3215
rect 1600 3165 1615 3185
rect 1635 3165 1650 3185
rect 1600 3135 1650 3165
rect 1600 3115 1615 3135
rect 1635 3115 1650 3135
rect 1600 3085 1650 3115
rect 1600 3065 1615 3085
rect 1635 3065 1650 3085
rect 1600 3050 1650 3065
rect 1750 3535 1800 3550
rect 1750 3515 1765 3535
rect 1785 3515 1800 3535
rect 1750 3485 1800 3515
rect 1750 3465 1765 3485
rect 1785 3465 1800 3485
rect 1750 3435 1800 3465
rect 1750 3415 1765 3435
rect 1785 3415 1800 3435
rect 1750 3385 1800 3415
rect 1750 3365 1765 3385
rect 1785 3365 1800 3385
rect 1750 3335 1800 3365
rect 1750 3315 1765 3335
rect 1785 3315 1800 3335
rect 1750 3285 1800 3315
rect 1750 3265 1765 3285
rect 1785 3265 1800 3285
rect 1750 3235 1800 3265
rect 1750 3215 1765 3235
rect 1785 3215 1800 3235
rect 1750 3185 1800 3215
rect 1750 3165 1765 3185
rect 1785 3165 1800 3185
rect 1750 3135 1800 3165
rect 1750 3115 1765 3135
rect 1785 3115 1800 3135
rect 1750 3085 1800 3115
rect 1750 3065 1765 3085
rect 1785 3065 1800 3085
rect 1750 3050 1800 3065
rect 1900 3535 1950 3550
rect 1900 3515 1915 3535
rect 1935 3515 1950 3535
rect 1900 3485 1950 3515
rect 1900 3465 1915 3485
rect 1935 3465 1950 3485
rect 1900 3435 1950 3465
rect 1900 3415 1915 3435
rect 1935 3415 1950 3435
rect 1900 3385 1950 3415
rect 1900 3365 1915 3385
rect 1935 3365 1950 3385
rect 1900 3335 1950 3365
rect 1900 3315 1915 3335
rect 1935 3315 1950 3335
rect 1900 3285 1950 3315
rect 1900 3265 1915 3285
rect 1935 3265 1950 3285
rect 1900 3235 1950 3265
rect 1900 3215 1915 3235
rect 1935 3215 1950 3235
rect 1900 3185 1950 3215
rect 1900 3165 1915 3185
rect 1935 3165 1950 3185
rect 1900 3135 1950 3165
rect 1900 3115 1915 3135
rect 1935 3115 1950 3135
rect 1900 3085 1950 3115
rect 1900 3065 1915 3085
rect 1935 3065 1950 3085
rect 1900 3050 1950 3065
rect 2050 3535 2100 3550
rect 2050 3515 2065 3535
rect 2085 3515 2100 3535
rect 2050 3485 2100 3515
rect 2050 3465 2065 3485
rect 2085 3465 2100 3485
rect 2050 3435 2100 3465
rect 2050 3415 2065 3435
rect 2085 3415 2100 3435
rect 2050 3385 2100 3415
rect 2050 3365 2065 3385
rect 2085 3365 2100 3385
rect 2050 3335 2100 3365
rect 2050 3315 2065 3335
rect 2085 3315 2100 3335
rect 2050 3285 2100 3315
rect 2050 3265 2065 3285
rect 2085 3265 2100 3285
rect 2050 3235 2100 3265
rect 2050 3215 2065 3235
rect 2085 3215 2100 3235
rect 2050 3185 2100 3215
rect 2050 3165 2065 3185
rect 2085 3165 2100 3185
rect 2050 3135 2100 3165
rect 2050 3115 2065 3135
rect 2085 3115 2100 3135
rect 2050 3085 2100 3115
rect 2050 3065 2065 3085
rect 2085 3065 2100 3085
rect 2050 3050 2100 3065
rect 2200 3535 2250 3550
rect 2200 3515 2215 3535
rect 2235 3515 2250 3535
rect 2200 3485 2250 3515
rect 2200 3465 2215 3485
rect 2235 3465 2250 3485
rect 2200 3435 2250 3465
rect 2200 3415 2215 3435
rect 2235 3415 2250 3435
rect 2200 3385 2250 3415
rect 2200 3365 2215 3385
rect 2235 3365 2250 3385
rect 2200 3335 2250 3365
rect 2200 3315 2215 3335
rect 2235 3315 2250 3335
rect 2200 3285 2250 3315
rect 2200 3265 2215 3285
rect 2235 3265 2250 3285
rect 2200 3235 2250 3265
rect 2200 3215 2215 3235
rect 2235 3215 2250 3235
rect 2200 3185 2250 3215
rect 2200 3165 2215 3185
rect 2235 3165 2250 3185
rect 2200 3135 2250 3165
rect 2200 3115 2215 3135
rect 2235 3115 2250 3135
rect 2200 3085 2250 3115
rect 2200 3065 2215 3085
rect 2235 3065 2250 3085
rect 2200 3050 2250 3065
rect 2350 3535 2400 3550
rect 2350 3515 2365 3535
rect 2385 3515 2400 3535
rect 2350 3485 2400 3515
rect 2350 3465 2365 3485
rect 2385 3465 2400 3485
rect 2350 3435 2400 3465
rect 2350 3415 2365 3435
rect 2385 3415 2400 3435
rect 2350 3385 2400 3415
rect 2350 3365 2365 3385
rect 2385 3365 2400 3385
rect 2350 3335 2400 3365
rect 2350 3315 2365 3335
rect 2385 3315 2400 3335
rect 2350 3285 2400 3315
rect 2350 3265 2365 3285
rect 2385 3265 2400 3285
rect 2350 3235 2400 3265
rect 2350 3215 2365 3235
rect 2385 3215 2400 3235
rect 2350 3185 2400 3215
rect 2350 3165 2365 3185
rect 2385 3165 2400 3185
rect 2350 3135 2400 3165
rect 2350 3115 2365 3135
rect 2385 3115 2400 3135
rect 2350 3085 2400 3115
rect 2350 3065 2365 3085
rect 2385 3065 2400 3085
rect 2350 3050 2400 3065
rect 2500 3535 2550 3550
rect 2500 3515 2515 3535
rect 2535 3515 2550 3535
rect 2500 3485 2550 3515
rect 2500 3465 2515 3485
rect 2535 3465 2550 3485
rect 2500 3435 2550 3465
rect 2500 3415 2515 3435
rect 2535 3415 2550 3435
rect 2500 3385 2550 3415
rect 2500 3365 2515 3385
rect 2535 3365 2550 3385
rect 2500 3335 2550 3365
rect 2500 3315 2515 3335
rect 2535 3315 2550 3335
rect 2500 3285 2550 3315
rect 2500 3265 2515 3285
rect 2535 3265 2550 3285
rect 2500 3235 2550 3265
rect 2500 3215 2515 3235
rect 2535 3215 2550 3235
rect 2500 3185 2550 3215
rect 2500 3165 2515 3185
rect 2535 3165 2550 3185
rect 2500 3135 2550 3165
rect 2500 3115 2515 3135
rect 2535 3115 2550 3135
rect 2500 3085 2550 3115
rect 2500 3065 2515 3085
rect 2535 3065 2550 3085
rect 2500 3050 2550 3065
rect 2650 3535 2700 3550
rect 2650 3515 2665 3535
rect 2685 3515 2700 3535
rect 2650 3485 2700 3515
rect 2650 3465 2665 3485
rect 2685 3465 2700 3485
rect 2650 3435 2700 3465
rect 2650 3415 2665 3435
rect 2685 3415 2700 3435
rect 2650 3385 2700 3415
rect 2650 3365 2665 3385
rect 2685 3365 2700 3385
rect 2650 3335 2700 3365
rect 2650 3315 2665 3335
rect 2685 3315 2700 3335
rect 2650 3285 2700 3315
rect 2650 3265 2665 3285
rect 2685 3265 2700 3285
rect 2650 3235 2700 3265
rect 2650 3215 2665 3235
rect 2685 3215 2700 3235
rect 2650 3185 2700 3215
rect 2650 3165 2665 3185
rect 2685 3165 2700 3185
rect 2650 3135 2700 3165
rect 2650 3115 2665 3135
rect 2685 3115 2700 3135
rect 2650 3085 2700 3115
rect 2650 3065 2665 3085
rect 2685 3065 2700 3085
rect 2650 3050 2700 3065
rect 2800 3535 2850 3550
rect 2800 3515 2815 3535
rect 2835 3515 2850 3535
rect 2800 3485 2850 3515
rect 2800 3465 2815 3485
rect 2835 3465 2850 3485
rect 2800 3435 2850 3465
rect 2800 3415 2815 3435
rect 2835 3415 2850 3435
rect 2800 3385 2850 3415
rect 2800 3365 2815 3385
rect 2835 3365 2850 3385
rect 2800 3335 2850 3365
rect 2800 3315 2815 3335
rect 2835 3315 2850 3335
rect 2800 3285 2850 3315
rect 2800 3265 2815 3285
rect 2835 3265 2850 3285
rect 2800 3235 2850 3265
rect 2800 3215 2815 3235
rect 2835 3215 2850 3235
rect 2800 3185 2850 3215
rect 2800 3165 2815 3185
rect 2835 3165 2850 3185
rect 2800 3135 2850 3165
rect 2800 3115 2815 3135
rect 2835 3115 2850 3135
rect 2800 3085 2850 3115
rect 2800 3065 2815 3085
rect 2835 3065 2850 3085
rect 2800 3050 2850 3065
rect 2950 3535 3000 3550
rect 2950 3515 2965 3535
rect 2985 3515 3000 3535
rect 2950 3485 3000 3515
rect 2950 3465 2965 3485
rect 2985 3465 3000 3485
rect 2950 3435 3000 3465
rect 2950 3415 2965 3435
rect 2985 3415 3000 3435
rect 2950 3385 3000 3415
rect 2950 3365 2965 3385
rect 2985 3365 3000 3385
rect 2950 3335 3000 3365
rect 2950 3315 2965 3335
rect 2985 3315 3000 3335
rect 2950 3285 3000 3315
rect 2950 3265 2965 3285
rect 2985 3265 3000 3285
rect 2950 3235 3000 3265
rect 2950 3215 2965 3235
rect 2985 3215 3000 3235
rect 2950 3185 3000 3215
rect 2950 3165 2965 3185
rect 2985 3165 3000 3185
rect 2950 3135 3000 3165
rect 2950 3115 2965 3135
rect 2985 3115 3000 3135
rect 2950 3085 3000 3115
rect 2950 3065 2965 3085
rect 2985 3065 3000 3085
rect 2950 3050 3000 3065
rect 3100 3535 3150 3550
rect 3100 3515 3115 3535
rect 3135 3515 3150 3535
rect 3100 3485 3150 3515
rect 3100 3465 3115 3485
rect 3135 3465 3150 3485
rect 3100 3435 3150 3465
rect 3100 3415 3115 3435
rect 3135 3415 3150 3435
rect 3100 3385 3150 3415
rect 3100 3365 3115 3385
rect 3135 3365 3150 3385
rect 3100 3335 3150 3365
rect 3100 3315 3115 3335
rect 3135 3315 3150 3335
rect 3100 3285 3150 3315
rect 3100 3265 3115 3285
rect 3135 3265 3150 3285
rect 3100 3235 3150 3265
rect 3100 3215 3115 3235
rect 3135 3215 3150 3235
rect 3100 3185 3150 3215
rect 3100 3165 3115 3185
rect 3135 3165 3150 3185
rect 3100 3135 3150 3165
rect 3100 3115 3115 3135
rect 3135 3115 3150 3135
rect 3100 3085 3150 3115
rect 3100 3065 3115 3085
rect 3135 3065 3150 3085
rect 3100 3050 3150 3065
rect 3250 3535 3300 3550
rect 3250 3515 3265 3535
rect 3285 3515 3300 3535
rect 3250 3485 3300 3515
rect 3250 3465 3265 3485
rect 3285 3465 3300 3485
rect 3250 3435 3300 3465
rect 3250 3415 3265 3435
rect 3285 3415 3300 3435
rect 3250 3385 3300 3415
rect 3250 3365 3265 3385
rect 3285 3365 3300 3385
rect 3250 3335 3300 3365
rect 3250 3315 3265 3335
rect 3285 3315 3300 3335
rect 3250 3285 3300 3315
rect 3250 3265 3265 3285
rect 3285 3265 3300 3285
rect 3250 3235 3300 3265
rect 3250 3215 3265 3235
rect 3285 3215 3300 3235
rect 3250 3185 3300 3215
rect 3250 3165 3265 3185
rect 3285 3165 3300 3185
rect 3250 3135 3300 3165
rect 3250 3115 3265 3135
rect 3285 3115 3300 3135
rect 3250 3085 3300 3115
rect 3250 3065 3265 3085
rect 3285 3065 3300 3085
rect 3250 3050 3300 3065
rect 3400 3535 3450 3550
rect 3400 3515 3415 3535
rect 3435 3515 3450 3535
rect 3400 3485 3450 3515
rect 3400 3465 3415 3485
rect 3435 3465 3450 3485
rect 3400 3435 3450 3465
rect 3400 3415 3415 3435
rect 3435 3415 3450 3435
rect 3400 3385 3450 3415
rect 3400 3365 3415 3385
rect 3435 3365 3450 3385
rect 3400 3335 3450 3365
rect 3400 3315 3415 3335
rect 3435 3315 3450 3335
rect 3400 3285 3450 3315
rect 3400 3265 3415 3285
rect 3435 3265 3450 3285
rect 3400 3235 3450 3265
rect 3400 3215 3415 3235
rect 3435 3215 3450 3235
rect 3400 3185 3450 3215
rect 3400 3165 3415 3185
rect 3435 3165 3450 3185
rect 3400 3135 3450 3165
rect 3400 3115 3415 3135
rect 3435 3115 3450 3135
rect 3400 3085 3450 3115
rect 3400 3065 3415 3085
rect 3435 3065 3450 3085
rect 3400 3050 3450 3065
rect 3550 3535 3600 3550
rect 3550 3515 3565 3535
rect 3585 3515 3600 3535
rect 3550 3485 3600 3515
rect 3550 3465 3565 3485
rect 3585 3465 3600 3485
rect 3550 3435 3600 3465
rect 3550 3415 3565 3435
rect 3585 3415 3600 3435
rect 3550 3385 3600 3415
rect 3550 3365 3565 3385
rect 3585 3365 3600 3385
rect 3550 3335 3600 3365
rect 3550 3315 3565 3335
rect 3585 3315 3600 3335
rect 3550 3285 3600 3315
rect 3550 3265 3565 3285
rect 3585 3265 3600 3285
rect 3550 3235 3600 3265
rect 3550 3215 3565 3235
rect 3585 3215 3600 3235
rect 3550 3185 3600 3215
rect 3550 3165 3565 3185
rect 3585 3165 3600 3185
rect 3550 3135 3600 3165
rect 3550 3115 3565 3135
rect 3585 3115 3600 3135
rect 3550 3085 3600 3115
rect 3550 3065 3565 3085
rect 3585 3065 3600 3085
rect 3550 3050 3600 3065
rect 4150 3535 4200 3550
rect 4150 3515 4165 3535
rect 4185 3515 4200 3535
rect 4150 3485 4200 3515
rect 4150 3465 4165 3485
rect 4185 3465 4200 3485
rect 4150 3435 4200 3465
rect 4150 3415 4165 3435
rect 4185 3415 4200 3435
rect 4150 3385 4200 3415
rect 4150 3365 4165 3385
rect 4185 3365 4200 3385
rect 4150 3335 4200 3365
rect 4150 3315 4165 3335
rect 4185 3315 4200 3335
rect 4150 3285 4200 3315
rect 4150 3265 4165 3285
rect 4185 3265 4200 3285
rect 4150 3235 4200 3265
rect 4150 3215 4165 3235
rect 4185 3215 4200 3235
rect 4150 3185 4200 3215
rect 4150 3165 4165 3185
rect 4185 3165 4200 3185
rect 4150 3135 4200 3165
rect 4150 3115 4165 3135
rect 4185 3115 4200 3135
rect 4150 3085 4200 3115
rect 4150 3065 4165 3085
rect 4185 3065 4200 3085
rect 4150 3050 4200 3065
rect 4750 3535 4800 3550
rect 4750 3515 4765 3535
rect 4785 3515 4800 3535
rect 4750 3485 4800 3515
rect 4750 3465 4765 3485
rect 4785 3465 4800 3485
rect 4750 3435 4800 3465
rect 4750 3415 4765 3435
rect 4785 3415 4800 3435
rect 4750 3385 4800 3415
rect 4750 3365 4765 3385
rect 4785 3365 4800 3385
rect 4750 3335 4800 3365
rect 4750 3315 4765 3335
rect 4785 3315 4800 3335
rect 4750 3285 4800 3315
rect 4750 3265 4765 3285
rect 4785 3265 4800 3285
rect 4750 3235 4800 3265
rect 4750 3215 4765 3235
rect 4785 3215 4800 3235
rect 4750 3185 4800 3215
rect 4750 3165 4765 3185
rect 4785 3165 4800 3185
rect 4750 3135 4800 3165
rect 4750 3115 4765 3135
rect 4785 3115 4800 3135
rect 4750 3085 4800 3115
rect 4750 3065 4765 3085
rect 4785 3065 4800 3085
rect 4750 3050 4800 3065
rect 4900 3535 4950 3550
rect 4900 3515 4915 3535
rect 4935 3515 4950 3535
rect 4900 3485 4950 3515
rect 4900 3465 4915 3485
rect 4935 3465 4950 3485
rect 4900 3435 4950 3465
rect 4900 3415 4915 3435
rect 4935 3415 4950 3435
rect 4900 3385 4950 3415
rect 4900 3365 4915 3385
rect 4935 3365 4950 3385
rect 4900 3335 4950 3365
rect 4900 3315 4915 3335
rect 4935 3315 4950 3335
rect 4900 3285 4950 3315
rect 4900 3265 4915 3285
rect 4935 3265 4950 3285
rect 4900 3235 4950 3265
rect 4900 3215 4915 3235
rect 4935 3215 4950 3235
rect 4900 3185 4950 3215
rect 4900 3165 4915 3185
rect 4935 3165 4950 3185
rect 4900 3135 4950 3165
rect 4900 3115 4915 3135
rect 4935 3115 4950 3135
rect 4900 3085 4950 3115
rect 4900 3065 4915 3085
rect 4935 3065 4950 3085
rect 4900 3050 4950 3065
rect 5050 3535 5100 3550
rect 5050 3515 5065 3535
rect 5085 3515 5100 3535
rect 5050 3485 5100 3515
rect 5050 3465 5065 3485
rect 5085 3465 5100 3485
rect 5050 3435 5100 3465
rect 5050 3415 5065 3435
rect 5085 3415 5100 3435
rect 5050 3385 5100 3415
rect 5050 3365 5065 3385
rect 5085 3365 5100 3385
rect 5050 3335 5100 3365
rect 5050 3315 5065 3335
rect 5085 3315 5100 3335
rect 5050 3285 5100 3315
rect 5050 3265 5065 3285
rect 5085 3265 5100 3285
rect 5050 3235 5100 3265
rect 5050 3215 5065 3235
rect 5085 3215 5100 3235
rect 5050 3185 5100 3215
rect 5050 3165 5065 3185
rect 5085 3165 5100 3185
rect 5050 3135 5100 3165
rect 5050 3115 5065 3135
rect 5085 3115 5100 3135
rect 5050 3085 5100 3115
rect 5050 3065 5065 3085
rect 5085 3065 5100 3085
rect 5050 3050 5100 3065
rect 5200 3535 5250 3550
rect 5200 3515 5215 3535
rect 5235 3515 5250 3535
rect 5200 3485 5250 3515
rect 5200 3465 5215 3485
rect 5235 3465 5250 3485
rect 5200 3435 5250 3465
rect 5200 3415 5215 3435
rect 5235 3415 5250 3435
rect 5200 3385 5250 3415
rect 5200 3365 5215 3385
rect 5235 3365 5250 3385
rect 5200 3335 5250 3365
rect 5200 3315 5215 3335
rect 5235 3315 5250 3335
rect 5200 3285 5250 3315
rect 5200 3265 5215 3285
rect 5235 3265 5250 3285
rect 5200 3235 5250 3265
rect 5200 3215 5215 3235
rect 5235 3215 5250 3235
rect 5200 3185 5250 3215
rect 5200 3165 5215 3185
rect 5235 3165 5250 3185
rect 5200 3135 5250 3165
rect 5200 3115 5215 3135
rect 5235 3115 5250 3135
rect 5200 3085 5250 3115
rect 5200 3065 5215 3085
rect 5235 3065 5250 3085
rect 5200 3050 5250 3065
rect 5350 3535 5400 3550
rect 5350 3515 5365 3535
rect 5385 3515 5400 3535
rect 5350 3485 5400 3515
rect 5350 3465 5365 3485
rect 5385 3465 5400 3485
rect 5350 3435 5400 3465
rect 5350 3415 5365 3435
rect 5385 3415 5400 3435
rect 5350 3385 5400 3415
rect 5350 3365 5365 3385
rect 5385 3365 5400 3385
rect 5350 3335 5400 3365
rect 5350 3315 5365 3335
rect 5385 3315 5400 3335
rect 5350 3285 5400 3315
rect 5350 3265 5365 3285
rect 5385 3265 5400 3285
rect 5350 3235 5400 3265
rect 5350 3215 5365 3235
rect 5385 3215 5400 3235
rect 5350 3185 5400 3215
rect 5350 3165 5365 3185
rect 5385 3165 5400 3185
rect 5350 3135 5400 3165
rect 5350 3115 5365 3135
rect 5385 3115 5400 3135
rect 5350 3085 5400 3115
rect 5350 3065 5365 3085
rect 5385 3065 5400 3085
rect 5350 3050 5400 3065
rect 5500 3535 5550 3550
rect 5500 3515 5515 3535
rect 5535 3515 5550 3535
rect 5500 3485 5550 3515
rect 5500 3465 5515 3485
rect 5535 3465 5550 3485
rect 5500 3435 5550 3465
rect 5500 3415 5515 3435
rect 5535 3415 5550 3435
rect 5500 3385 5550 3415
rect 5500 3365 5515 3385
rect 5535 3365 5550 3385
rect 5500 3335 5550 3365
rect 5500 3315 5515 3335
rect 5535 3315 5550 3335
rect 5500 3285 5550 3315
rect 5500 3265 5515 3285
rect 5535 3265 5550 3285
rect 5500 3235 5550 3265
rect 5500 3215 5515 3235
rect 5535 3215 5550 3235
rect 5500 3185 5550 3215
rect 5500 3165 5515 3185
rect 5535 3165 5550 3185
rect 5500 3135 5550 3165
rect 5500 3115 5515 3135
rect 5535 3115 5550 3135
rect 5500 3085 5550 3115
rect 5500 3065 5515 3085
rect 5535 3065 5550 3085
rect 5500 3050 5550 3065
rect 5650 3535 5700 3550
rect 5650 3515 5665 3535
rect 5685 3515 5700 3535
rect 5650 3485 5700 3515
rect 5650 3465 5665 3485
rect 5685 3465 5700 3485
rect 5650 3435 5700 3465
rect 5650 3415 5665 3435
rect 5685 3415 5700 3435
rect 5650 3385 5700 3415
rect 5650 3365 5665 3385
rect 5685 3365 5700 3385
rect 5650 3335 5700 3365
rect 5650 3315 5665 3335
rect 5685 3315 5700 3335
rect 5650 3285 5700 3315
rect 5650 3265 5665 3285
rect 5685 3265 5700 3285
rect 5650 3235 5700 3265
rect 5650 3215 5665 3235
rect 5685 3215 5700 3235
rect 5650 3185 5700 3215
rect 5650 3165 5665 3185
rect 5685 3165 5700 3185
rect 5650 3135 5700 3165
rect 5650 3115 5665 3135
rect 5685 3115 5700 3135
rect 5650 3085 5700 3115
rect 5650 3065 5665 3085
rect 5685 3065 5700 3085
rect 5650 3050 5700 3065
rect 5800 3535 5850 3550
rect 5800 3515 5815 3535
rect 5835 3515 5850 3535
rect 5800 3485 5850 3515
rect 5800 3465 5815 3485
rect 5835 3465 5850 3485
rect 5800 3435 5850 3465
rect 5800 3415 5815 3435
rect 5835 3415 5850 3435
rect 5800 3385 5850 3415
rect 5800 3365 5815 3385
rect 5835 3365 5850 3385
rect 5800 3335 5850 3365
rect 5800 3315 5815 3335
rect 5835 3315 5850 3335
rect 5800 3285 5850 3315
rect 5800 3265 5815 3285
rect 5835 3265 5850 3285
rect 5800 3235 5850 3265
rect 5800 3215 5815 3235
rect 5835 3215 5850 3235
rect 5800 3185 5850 3215
rect 5800 3165 5815 3185
rect 5835 3165 5850 3185
rect 5800 3135 5850 3165
rect 5800 3115 5815 3135
rect 5835 3115 5850 3135
rect 5800 3085 5850 3115
rect 5800 3065 5815 3085
rect 5835 3065 5850 3085
rect 5800 3050 5850 3065
rect 5950 3535 6000 3550
rect 5950 3515 5965 3535
rect 5985 3515 6000 3535
rect 5950 3485 6000 3515
rect 5950 3465 5965 3485
rect 5985 3465 6000 3485
rect 5950 3435 6000 3465
rect 5950 3415 5965 3435
rect 5985 3415 6000 3435
rect 5950 3385 6000 3415
rect 5950 3365 5965 3385
rect 5985 3365 6000 3385
rect 5950 3335 6000 3365
rect 5950 3315 5965 3335
rect 5985 3315 6000 3335
rect 5950 3285 6000 3315
rect 5950 3265 5965 3285
rect 5985 3265 6000 3285
rect 5950 3235 6000 3265
rect 5950 3215 5965 3235
rect 5985 3215 6000 3235
rect 5950 3185 6000 3215
rect 5950 3165 5965 3185
rect 5985 3165 6000 3185
rect 5950 3135 6000 3165
rect 5950 3115 5965 3135
rect 5985 3115 6000 3135
rect 5950 3085 6000 3115
rect 5950 3065 5965 3085
rect 5985 3065 6000 3085
rect 5950 3050 6000 3065
rect 6100 3535 6150 3550
rect 6100 3515 6115 3535
rect 6135 3515 6150 3535
rect 6100 3485 6150 3515
rect 6100 3465 6115 3485
rect 6135 3465 6150 3485
rect 6100 3435 6150 3465
rect 6100 3415 6115 3435
rect 6135 3415 6150 3435
rect 6100 3385 6150 3415
rect 6100 3365 6115 3385
rect 6135 3365 6150 3385
rect 6100 3335 6150 3365
rect 6100 3315 6115 3335
rect 6135 3315 6150 3335
rect 6100 3285 6150 3315
rect 6100 3265 6115 3285
rect 6135 3265 6150 3285
rect 6100 3235 6150 3265
rect 6100 3215 6115 3235
rect 6135 3215 6150 3235
rect 6100 3185 6150 3215
rect 6100 3165 6115 3185
rect 6135 3165 6150 3185
rect 6100 3135 6150 3165
rect 6100 3115 6115 3135
rect 6135 3115 6150 3135
rect 6100 3085 6150 3115
rect 6100 3065 6115 3085
rect 6135 3065 6150 3085
rect 6100 3050 6150 3065
rect 6250 3535 6300 3550
rect 6250 3515 6265 3535
rect 6285 3515 6300 3535
rect 6250 3485 6300 3515
rect 6250 3465 6265 3485
rect 6285 3465 6300 3485
rect 6250 3435 6300 3465
rect 6250 3415 6265 3435
rect 6285 3415 6300 3435
rect 6250 3385 6300 3415
rect 6250 3365 6265 3385
rect 6285 3365 6300 3385
rect 6250 3335 6300 3365
rect 6250 3315 6265 3335
rect 6285 3315 6300 3335
rect 6250 3285 6300 3315
rect 6250 3265 6265 3285
rect 6285 3265 6300 3285
rect 6250 3235 6300 3265
rect 6250 3215 6265 3235
rect 6285 3215 6300 3235
rect 6250 3185 6300 3215
rect 6250 3165 6265 3185
rect 6285 3165 6300 3185
rect 6250 3135 6300 3165
rect 6250 3115 6265 3135
rect 6285 3115 6300 3135
rect 6250 3085 6300 3115
rect 6250 3065 6265 3085
rect 6285 3065 6300 3085
rect 6250 3050 6300 3065
rect 6400 3535 6450 3550
rect 6400 3515 6415 3535
rect 6435 3515 6450 3535
rect 6400 3485 6450 3515
rect 6400 3465 6415 3485
rect 6435 3465 6450 3485
rect 6400 3435 6450 3465
rect 6400 3415 6415 3435
rect 6435 3415 6450 3435
rect 6400 3385 6450 3415
rect 6400 3365 6415 3385
rect 6435 3365 6450 3385
rect 6400 3335 6450 3365
rect 6400 3315 6415 3335
rect 6435 3315 6450 3335
rect 6400 3285 6450 3315
rect 6400 3265 6415 3285
rect 6435 3265 6450 3285
rect 6400 3235 6450 3265
rect 6400 3215 6415 3235
rect 6435 3215 6450 3235
rect 6400 3185 6450 3215
rect 6400 3165 6415 3185
rect 6435 3165 6450 3185
rect 6400 3135 6450 3165
rect 6400 3115 6415 3135
rect 6435 3115 6450 3135
rect 6400 3085 6450 3115
rect 6400 3065 6415 3085
rect 6435 3065 6450 3085
rect 6400 3050 6450 3065
rect 6550 3535 6600 3550
rect 6550 3515 6565 3535
rect 6585 3515 6600 3535
rect 6550 3485 6600 3515
rect 6550 3465 6565 3485
rect 6585 3465 6600 3485
rect 6550 3435 6600 3465
rect 6550 3415 6565 3435
rect 6585 3415 6600 3435
rect 6550 3385 6600 3415
rect 6550 3365 6565 3385
rect 6585 3365 6600 3385
rect 6550 3335 6600 3365
rect 6550 3315 6565 3335
rect 6585 3315 6600 3335
rect 6550 3285 6600 3315
rect 6550 3265 6565 3285
rect 6585 3265 6600 3285
rect 6550 3235 6600 3265
rect 6550 3215 6565 3235
rect 6585 3215 6600 3235
rect 6550 3185 6600 3215
rect 6550 3165 6565 3185
rect 6585 3165 6600 3185
rect 6550 3135 6600 3165
rect 6550 3115 6565 3135
rect 6585 3115 6600 3135
rect 6550 3085 6600 3115
rect 6550 3065 6565 3085
rect 6585 3065 6600 3085
rect 6550 3050 6600 3065
rect 6700 3535 6750 3550
rect 6700 3515 6715 3535
rect 6735 3515 6750 3535
rect 6700 3485 6750 3515
rect 6700 3465 6715 3485
rect 6735 3465 6750 3485
rect 6700 3435 6750 3465
rect 6700 3415 6715 3435
rect 6735 3415 6750 3435
rect 6700 3385 6750 3415
rect 6700 3365 6715 3385
rect 6735 3365 6750 3385
rect 6700 3335 6750 3365
rect 6700 3315 6715 3335
rect 6735 3315 6750 3335
rect 6700 3285 6750 3315
rect 6700 3265 6715 3285
rect 6735 3265 6750 3285
rect 6700 3235 6750 3265
rect 6700 3215 6715 3235
rect 6735 3215 6750 3235
rect 6700 3185 6750 3215
rect 6700 3165 6715 3185
rect 6735 3165 6750 3185
rect 6700 3135 6750 3165
rect 6700 3115 6715 3135
rect 6735 3115 6750 3135
rect 6700 3085 6750 3115
rect 6700 3065 6715 3085
rect 6735 3065 6750 3085
rect 6700 3050 6750 3065
rect 6850 3535 6900 3550
rect 6850 3515 6865 3535
rect 6885 3515 6900 3535
rect 6850 3485 6900 3515
rect 6850 3465 6865 3485
rect 6885 3465 6900 3485
rect 6850 3435 6900 3465
rect 6850 3415 6865 3435
rect 6885 3415 6900 3435
rect 6850 3385 6900 3415
rect 6850 3365 6865 3385
rect 6885 3365 6900 3385
rect 6850 3335 6900 3365
rect 6850 3315 6865 3335
rect 6885 3315 6900 3335
rect 6850 3285 6900 3315
rect 6850 3265 6865 3285
rect 6885 3265 6900 3285
rect 6850 3235 6900 3265
rect 6850 3215 6865 3235
rect 6885 3215 6900 3235
rect 6850 3185 6900 3215
rect 6850 3165 6865 3185
rect 6885 3165 6900 3185
rect 6850 3135 6900 3165
rect 6850 3115 6865 3135
rect 6885 3115 6900 3135
rect 6850 3085 6900 3115
rect 6850 3065 6865 3085
rect 6885 3065 6900 3085
rect 6850 3050 6900 3065
rect 7000 3535 7050 3550
rect 7000 3515 7015 3535
rect 7035 3515 7050 3535
rect 7000 3485 7050 3515
rect 7000 3465 7015 3485
rect 7035 3465 7050 3485
rect 7000 3435 7050 3465
rect 7000 3415 7015 3435
rect 7035 3415 7050 3435
rect 7000 3385 7050 3415
rect 7000 3365 7015 3385
rect 7035 3365 7050 3385
rect 7000 3335 7050 3365
rect 7000 3315 7015 3335
rect 7035 3315 7050 3335
rect 7000 3285 7050 3315
rect 7000 3265 7015 3285
rect 7035 3265 7050 3285
rect 7000 3235 7050 3265
rect 7000 3215 7015 3235
rect 7035 3215 7050 3235
rect 7000 3185 7050 3215
rect 7000 3165 7015 3185
rect 7035 3165 7050 3185
rect 7000 3135 7050 3165
rect 7000 3115 7015 3135
rect 7035 3115 7050 3135
rect 7000 3085 7050 3115
rect 7000 3065 7015 3085
rect 7035 3065 7050 3085
rect 7000 3050 7050 3065
rect 7150 3535 7200 3550
rect 7150 3515 7165 3535
rect 7185 3515 7200 3535
rect 7150 3485 7200 3515
rect 7150 3465 7165 3485
rect 7185 3465 7200 3485
rect 7150 3435 7200 3465
rect 7150 3415 7165 3435
rect 7185 3415 7200 3435
rect 7150 3385 7200 3415
rect 7150 3365 7165 3385
rect 7185 3365 7200 3385
rect 7150 3335 7200 3365
rect 7150 3315 7165 3335
rect 7185 3315 7200 3335
rect 7150 3285 7200 3315
rect 7150 3265 7165 3285
rect 7185 3265 7200 3285
rect 7150 3235 7200 3265
rect 7150 3215 7165 3235
rect 7185 3215 7200 3235
rect 7150 3185 7200 3215
rect 7150 3165 7165 3185
rect 7185 3165 7200 3185
rect 7150 3135 7200 3165
rect 7150 3115 7165 3135
rect 7185 3115 7200 3135
rect 7150 3085 7200 3115
rect 7150 3065 7165 3085
rect 7185 3065 7200 3085
rect 7150 3050 7200 3065
rect 7300 3535 7350 3550
rect 7300 3515 7315 3535
rect 7335 3515 7350 3535
rect 7300 3485 7350 3515
rect 7300 3465 7315 3485
rect 7335 3465 7350 3485
rect 7300 3435 7350 3465
rect 7300 3415 7315 3435
rect 7335 3415 7350 3435
rect 7300 3385 7350 3415
rect 7300 3365 7315 3385
rect 7335 3365 7350 3385
rect 7300 3335 7350 3365
rect 7300 3315 7315 3335
rect 7335 3315 7350 3335
rect 7300 3285 7350 3315
rect 7300 3265 7315 3285
rect 7335 3265 7350 3285
rect 7300 3235 7350 3265
rect 7300 3215 7315 3235
rect 7335 3215 7350 3235
rect 7300 3185 7350 3215
rect 7300 3165 7315 3185
rect 7335 3165 7350 3185
rect 7300 3135 7350 3165
rect 7300 3115 7315 3135
rect 7335 3115 7350 3135
rect 7300 3085 7350 3115
rect 7300 3065 7315 3085
rect 7335 3065 7350 3085
rect 7300 3050 7350 3065
rect 7450 3535 7500 3550
rect 7450 3515 7465 3535
rect 7485 3515 7500 3535
rect 7450 3485 7500 3515
rect 7450 3465 7465 3485
rect 7485 3465 7500 3485
rect 7450 3435 7500 3465
rect 7450 3415 7465 3435
rect 7485 3415 7500 3435
rect 7450 3385 7500 3415
rect 7450 3365 7465 3385
rect 7485 3365 7500 3385
rect 7450 3335 7500 3365
rect 7450 3315 7465 3335
rect 7485 3315 7500 3335
rect 7450 3285 7500 3315
rect 7450 3265 7465 3285
rect 7485 3265 7500 3285
rect 7450 3235 7500 3265
rect 7450 3215 7465 3235
rect 7485 3215 7500 3235
rect 7450 3185 7500 3215
rect 7450 3165 7465 3185
rect 7485 3165 7500 3185
rect 7450 3135 7500 3165
rect 7450 3115 7465 3135
rect 7485 3115 7500 3135
rect 7450 3085 7500 3115
rect 7450 3065 7465 3085
rect 7485 3065 7500 3085
rect 7450 3050 7500 3065
rect 7600 3535 7650 3550
rect 7600 3515 7615 3535
rect 7635 3515 7650 3535
rect 7600 3485 7650 3515
rect 7600 3465 7615 3485
rect 7635 3465 7650 3485
rect 7600 3435 7650 3465
rect 7600 3415 7615 3435
rect 7635 3415 7650 3435
rect 7600 3385 7650 3415
rect 7600 3365 7615 3385
rect 7635 3365 7650 3385
rect 7600 3335 7650 3365
rect 7600 3315 7615 3335
rect 7635 3315 7650 3335
rect 7600 3285 7650 3315
rect 7600 3265 7615 3285
rect 7635 3265 7650 3285
rect 7600 3235 7650 3265
rect 7600 3215 7615 3235
rect 7635 3215 7650 3235
rect 7600 3185 7650 3215
rect 7600 3165 7615 3185
rect 7635 3165 7650 3185
rect 7600 3135 7650 3165
rect 7600 3115 7615 3135
rect 7635 3115 7650 3135
rect 7600 3085 7650 3115
rect 7600 3065 7615 3085
rect 7635 3065 7650 3085
rect 7600 3050 7650 3065
rect 7750 3535 7800 3550
rect 7750 3515 7765 3535
rect 7785 3515 7800 3535
rect 7750 3485 7800 3515
rect 7750 3465 7765 3485
rect 7785 3465 7800 3485
rect 7750 3435 7800 3465
rect 7750 3415 7765 3435
rect 7785 3415 7800 3435
rect 7750 3385 7800 3415
rect 7750 3365 7765 3385
rect 7785 3365 7800 3385
rect 7750 3335 7800 3365
rect 7750 3315 7765 3335
rect 7785 3315 7800 3335
rect 7750 3285 7800 3315
rect 7750 3265 7765 3285
rect 7785 3265 7800 3285
rect 7750 3235 7800 3265
rect 7750 3215 7765 3235
rect 7785 3215 7800 3235
rect 7750 3185 7800 3215
rect 7750 3165 7765 3185
rect 7785 3165 7800 3185
rect 7750 3135 7800 3165
rect 7750 3115 7765 3135
rect 7785 3115 7800 3135
rect 7750 3085 7800 3115
rect 7750 3065 7765 3085
rect 7785 3065 7800 3085
rect 7750 3050 7800 3065
rect 8350 3535 8400 3550
rect 8350 3515 8365 3535
rect 8385 3515 8400 3535
rect 8350 3485 8400 3515
rect 8350 3465 8365 3485
rect 8385 3465 8400 3485
rect 8350 3435 8400 3465
rect 8350 3415 8365 3435
rect 8385 3415 8400 3435
rect 8350 3385 8400 3415
rect 8350 3365 8365 3385
rect 8385 3365 8400 3385
rect 8350 3335 8400 3365
rect 8350 3315 8365 3335
rect 8385 3315 8400 3335
rect 8350 3285 8400 3315
rect 8350 3265 8365 3285
rect 8385 3265 8400 3285
rect 8350 3235 8400 3265
rect 8350 3215 8365 3235
rect 8385 3215 8400 3235
rect 8350 3185 8400 3215
rect 8350 3165 8365 3185
rect 8385 3165 8400 3185
rect 8350 3135 8400 3165
rect 8350 3115 8365 3135
rect 8385 3115 8400 3135
rect 8350 3085 8400 3115
rect 8350 3065 8365 3085
rect 8385 3065 8400 3085
rect 8350 3050 8400 3065
rect 8500 3535 8550 3600
rect 8500 3515 8515 3535
rect 8535 3515 8550 3535
rect 8500 3485 8550 3515
rect 8500 3465 8515 3485
rect 8535 3465 8550 3485
rect 8500 3435 8550 3465
rect 8500 3415 8515 3435
rect 8535 3415 8550 3435
rect 8500 3385 8550 3415
rect 8500 3365 8515 3385
rect 8535 3365 8550 3385
rect 8500 3335 8550 3365
rect 8500 3315 8515 3335
rect 8535 3315 8550 3335
rect 8500 3285 8550 3315
rect 8500 3265 8515 3285
rect 8535 3265 8550 3285
rect 8500 3235 8550 3265
rect 8500 3215 8515 3235
rect 8535 3215 8550 3235
rect 8500 3185 8550 3215
rect 8500 3165 8515 3185
rect 8535 3165 8550 3185
rect 8500 3135 8550 3165
rect 8500 3115 8515 3135
rect 8535 3115 8550 3135
rect 8500 3085 8550 3115
rect 8500 3065 8515 3085
rect 8535 3065 8550 3085
rect 8500 3050 8550 3065
rect 8650 3535 8700 3550
rect 8650 3515 8665 3535
rect 8685 3515 8700 3535
rect 8650 3485 8700 3515
rect 8650 3465 8665 3485
rect 8685 3465 8700 3485
rect 8650 3435 8700 3465
rect 8650 3415 8665 3435
rect 8685 3415 8700 3435
rect 8650 3385 8700 3415
rect 8650 3365 8665 3385
rect 8685 3365 8700 3385
rect 8650 3335 8700 3365
rect 8650 3315 8665 3335
rect 8685 3315 8700 3335
rect 8650 3285 8700 3315
rect 8650 3265 8665 3285
rect 8685 3265 8700 3285
rect 8650 3235 8700 3265
rect 8650 3215 8665 3235
rect 8685 3215 8700 3235
rect 8650 3185 8700 3215
rect 8650 3165 8665 3185
rect 8685 3165 8700 3185
rect 8650 3135 8700 3165
rect 8650 3115 8665 3135
rect 8685 3115 8700 3135
rect 8650 3085 8700 3115
rect 8650 3065 8665 3085
rect 8685 3065 8700 3085
rect 8650 3050 8700 3065
rect 8800 3535 8850 3600
rect 8800 3515 8815 3535
rect 8835 3515 8850 3535
rect 8800 3485 8850 3515
rect 8800 3465 8815 3485
rect 8835 3465 8850 3485
rect 8800 3435 8850 3465
rect 8800 3415 8815 3435
rect 8835 3415 8850 3435
rect 8800 3385 8850 3415
rect 8800 3365 8815 3385
rect 8835 3365 8850 3385
rect 8800 3335 8850 3365
rect 8800 3315 8815 3335
rect 8835 3315 8850 3335
rect 8800 3285 8850 3315
rect 8800 3265 8815 3285
rect 8835 3265 8850 3285
rect 8800 3235 8850 3265
rect 8800 3215 8815 3235
rect 8835 3215 8850 3235
rect 8800 3185 8850 3215
rect 8800 3165 8815 3185
rect 8835 3165 8850 3185
rect 8800 3135 8850 3165
rect 8800 3115 8815 3135
rect 8835 3115 8850 3135
rect 8800 3085 8850 3115
rect 8800 3065 8815 3085
rect 8835 3065 8850 3085
rect 8800 3050 8850 3065
rect 8950 3535 9000 3550
rect 8950 3515 8965 3535
rect 8985 3515 9000 3535
rect 8950 3485 9000 3515
rect 8950 3465 8965 3485
rect 8985 3465 9000 3485
rect 8950 3435 9000 3465
rect 8950 3415 8965 3435
rect 8985 3415 9000 3435
rect 8950 3385 9000 3415
rect 8950 3365 8965 3385
rect 8985 3365 9000 3385
rect 8950 3335 9000 3365
rect 8950 3315 8965 3335
rect 8985 3315 9000 3335
rect 8950 3285 9000 3315
rect 8950 3265 8965 3285
rect 8985 3265 9000 3285
rect 8950 3235 9000 3265
rect 8950 3215 8965 3235
rect 8985 3215 9000 3235
rect 8950 3185 9000 3215
rect 8950 3165 8965 3185
rect 8985 3165 9000 3185
rect 8950 3135 9000 3165
rect 8950 3115 8965 3135
rect 8985 3115 9000 3135
rect 8950 3085 9000 3115
rect 8950 3065 8965 3085
rect 8985 3065 9000 3085
rect 8950 3050 9000 3065
rect 9100 3535 9150 3600
rect 9100 3515 9115 3535
rect 9135 3515 9150 3535
rect 9100 3485 9150 3515
rect 9100 3465 9115 3485
rect 9135 3465 9150 3485
rect 9100 3435 9150 3465
rect 9100 3415 9115 3435
rect 9135 3415 9150 3435
rect 9100 3385 9150 3415
rect 9100 3365 9115 3385
rect 9135 3365 9150 3385
rect 9100 3335 9150 3365
rect 9100 3315 9115 3335
rect 9135 3315 9150 3335
rect 9100 3285 9150 3315
rect 9100 3265 9115 3285
rect 9135 3265 9150 3285
rect 9100 3235 9150 3265
rect 9100 3215 9115 3235
rect 9135 3215 9150 3235
rect 9100 3185 9150 3215
rect 9100 3165 9115 3185
rect 9135 3165 9150 3185
rect 9100 3135 9150 3165
rect 9100 3115 9115 3135
rect 9135 3115 9150 3135
rect 9100 3085 9150 3115
rect 9100 3065 9115 3085
rect 9135 3065 9150 3085
rect 9100 3050 9150 3065
rect 9250 3535 9300 3550
rect 9250 3515 9265 3535
rect 9285 3515 9300 3535
rect 9250 3485 9300 3515
rect 9250 3465 9265 3485
rect 9285 3465 9300 3485
rect 9250 3435 9300 3465
rect 9250 3415 9265 3435
rect 9285 3415 9300 3435
rect 9250 3385 9300 3415
rect 9250 3365 9265 3385
rect 9285 3365 9300 3385
rect 9250 3335 9300 3365
rect 9250 3315 9265 3335
rect 9285 3315 9300 3335
rect 9250 3285 9300 3315
rect 9250 3265 9265 3285
rect 9285 3265 9300 3285
rect 9250 3235 9300 3265
rect 9250 3215 9265 3235
rect 9285 3215 9300 3235
rect 9250 3185 9300 3215
rect 9250 3165 9265 3185
rect 9285 3165 9300 3185
rect 9250 3135 9300 3165
rect 9250 3115 9265 3135
rect 9285 3115 9300 3135
rect 9250 3085 9300 3115
rect 9250 3065 9265 3085
rect 9285 3065 9300 3085
rect 9250 3050 9300 3065
rect 9400 3535 9450 3600
rect 9400 3515 9415 3535
rect 9435 3515 9450 3535
rect 9400 3485 9450 3515
rect 9400 3465 9415 3485
rect 9435 3465 9450 3485
rect 9400 3435 9450 3465
rect 9400 3415 9415 3435
rect 9435 3415 9450 3435
rect 9400 3385 9450 3415
rect 9400 3365 9415 3385
rect 9435 3365 9450 3385
rect 9400 3335 9450 3365
rect 9400 3315 9415 3335
rect 9435 3315 9450 3335
rect 9400 3285 9450 3315
rect 9400 3265 9415 3285
rect 9435 3265 9450 3285
rect 9400 3235 9450 3265
rect 9400 3215 9415 3235
rect 9435 3215 9450 3235
rect 9400 3185 9450 3215
rect 9400 3165 9415 3185
rect 9435 3165 9450 3185
rect 9400 3135 9450 3165
rect 9400 3115 9415 3135
rect 9435 3115 9450 3135
rect 9400 3085 9450 3115
rect 9400 3065 9415 3085
rect 9435 3065 9450 3085
rect 9400 3050 9450 3065
rect 9550 3535 9600 3550
rect 9550 3515 9565 3535
rect 9585 3515 9600 3535
rect 9550 3485 9600 3515
rect 9550 3465 9565 3485
rect 9585 3465 9600 3485
rect 9550 3435 9600 3465
rect 9550 3415 9565 3435
rect 9585 3415 9600 3435
rect 9550 3385 9600 3415
rect 9550 3365 9565 3385
rect 9585 3365 9600 3385
rect 9550 3335 9600 3365
rect 9550 3315 9565 3335
rect 9585 3315 9600 3335
rect 9550 3285 9600 3315
rect 9550 3265 9565 3285
rect 9585 3265 9600 3285
rect 9550 3235 9600 3265
rect 9550 3215 9565 3235
rect 9585 3215 9600 3235
rect 9550 3185 9600 3215
rect 9550 3165 9565 3185
rect 9585 3165 9600 3185
rect 9550 3135 9600 3165
rect 9550 3115 9565 3135
rect 9585 3115 9600 3135
rect 9550 3085 9600 3115
rect 9550 3065 9565 3085
rect 9585 3065 9600 3085
rect 9550 3050 9600 3065
rect 9700 3535 9750 3600
rect 9700 3515 9715 3535
rect 9735 3515 9750 3535
rect 9700 3485 9750 3515
rect 9700 3465 9715 3485
rect 9735 3465 9750 3485
rect 9700 3435 9750 3465
rect 9700 3415 9715 3435
rect 9735 3415 9750 3435
rect 9700 3385 9750 3415
rect 9700 3365 9715 3385
rect 9735 3365 9750 3385
rect 9700 3335 9750 3365
rect 9700 3315 9715 3335
rect 9735 3315 9750 3335
rect 9700 3285 9750 3315
rect 9700 3265 9715 3285
rect 9735 3265 9750 3285
rect 9700 3235 9750 3265
rect 9700 3215 9715 3235
rect 9735 3215 9750 3235
rect 9700 3185 9750 3215
rect 9700 3165 9715 3185
rect 9735 3165 9750 3185
rect 9700 3135 9750 3165
rect 9700 3115 9715 3135
rect 9735 3115 9750 3135
rect 9700 3085 9750 3115
rect 9700 3065 9715 3085
rect 9735 3065 9750 3085
rect 9700 3050 9750 3065
rect 9850 3535 9900 3550
rect 9850 3515 9865 3535
rect 9885 3515 9900 3535
rect 9850 3485 9900 3515
rect 9850 3465 9865 3485
rect 9885 3465 9900 3485
rect 9850 3435 9900 3465
rect 9850 3415 9865 3435
rect 9885 3415 9900 3435
rect 9850 3385 9900 3415
rect 9850 3365 9865 3385
rect 9885 3365 9900 3385
rect 9850 3335 9900 3365
rect 9850 3315 9865 3335
rect 9885 3315 9900 3335
rect 9850 3285 9900 3315
rect 9850 3265 9865 3285
rect 9885 3265 9900 3285
rect 9850 3235 9900 3265
rect 9850 3215 9865 3235
rect 9885 3215 9900 3235
rect 9850 3185 9900 3215
rect 9850 3165 9865 3185
rect 9885 3165 9900 3185
rect 9850 3135 9900 3165
rect 9850 3115 9865 3135
rect 9885 3115 9900 3135
rect 9850 3085 9900 3115
rect 9850 3065 9865 3085
rect 9885 3065 9900 3085
rect 9850 3050 9900 3065
rect 10000 3535 10050 3600
rect 10000 3515 10015 3535
rect 10035 3515 10050 3535
rect 10000 3485 10050 3515
rect 10000 3465 10015 3485
rect 10035 3465 10050 3485
rect 10000 3435 10050 3465
rect 10000 3415 10015 3435
rect 10035 3415 10050 3435
rect 10000 3385 10050 3415
rect 10000 3365 10015 3385
rect 10035 3365 10050 3385
rect 10000 3335 10050 3365
rect 10000 3315 10015 3335
rect 10035 3315 10050 3335
rect 10000 3285 10050 3315
rect 10000 3265 10015 3285
rect 10035 3265 10050 3285
rect 10000 3235 10050 3265
rect 10000 3215 10015 3235
rect 10035 3215 10050 3235
rect 10000 3185 10050 3215
rect 10000 3165 10015 3185
rect 10035 3165 10050 3185
rect 10000 3135 10050 3165
rect 10000 3115 10015 3135
rect 10035 3115 10050 3135
rect 10000 3085 10050 3115
rect 10000 3065 10015 3085
rect 10035 3065 10050 3085
rect 10000 3050 10050 3065
rect 10150 3535 10200 3550
rect 10150 3515 10165 3535
rect 10185 3515 10200 3535
rect 10150 3485 10200 3515
rect 10150 3465 10165 3485
rect 10185 3465 10200 3485
rect 10150 3435 10200 3465
rect 10150 3415 10165 3435
rect 10185 3415 10200 3435
rect 10150 3385 10200 3415
rect 10150 3365 10165 3385
rect 10185 3365 10200 3385
rect 10150 3335 10200 3365
rect 10150 3315 10165 3335
rect 10185 3315 10200 3335
rect 10150 3285 10200 3315
rect 10150 3265 10165 3285
rect 10185 3265 10200 3285
rect 10150 3235 10200 3265
rect 10150 3215 10165 3235
rect 10185 3215 10200 3235
rect 10150 3185 10200 3215
rect 10150 3165 10165 3185
rect 10185 3165 10200 3185
rect 10150 3135 10200 3165
rect 10150 3115 10165 3135
rect 10185 3115 10200 3135
rect 10150 3085 10200 3115
rect 10150 3065 10165 3085
rect 10185 3065 10200 3085
rect 10150 3050 10200 3065
rect 10300 3535 10350 3600
rect 10300 3515 10315 3535
rect 10335 3515 10350 3535
rect 10300 3485 10350 3515
rect 10300 3465 10315 3485
rect 10335 3465 10350 3485
rect 10300 3435 10350 3465
rect 10300 3415 10315 3435
rect 10335 3415 10350 3435
rect 10300 3385 10350 3415
rect 10300 3365 10315 3385
rect 10335 3365 10350 3385
rect 10300 3335 10350 3365
rect 10300 3315 10315 3335
rect 10335 3315 10350 3335
rect 10300 3285 10350 3315
rect 10300 3265 10315 3285
rect 10335 3265 10350 3285
rect 10300 3235 10350 3265
rect 10300 3215 10315 3235
rect 10335 3215 10350 3235
rect 10300 3185 10350 3215
rect 10300 3165 10315 3185
rect 10335 3165 10350 3185
rect 10300 3135 10350 3165
rect 10300 3115 10315 3135
rect 10335 3115 10350 3135
rect 10300 3085 10350 3115
rect 10300 3065 10315 3085
rect 10335 3065 10350 3085
rect 10300 3050 10350 3065
rect 10450 3535 10500 3550
rect 10450 3515 10465 3535
rect 10485 3515 10500 3535
rect 10450 3485 10500 3515
rect 10450 3465 10465 3485
rect 10485 3465 10500 3485
rect 10450 3435 10500 3465
rect 10450 3415 10465 3435
rect 10485 3415 10500 3435
rect 10450 3385 10500 3415
rect 10450 3365 10465 3385
rect 10485 3365 10500 3385
rect 10450 3335 10500 3365
rect 10450 3315 10465 3335
rect 10485 3315 10500 3335
rect 10450 3285 10500 3315
rect 10450 3265 10465 3285
rect 10485 3265 10500 3285
rect 10450 3235 10500 3265
rect 10450 3215 10465 3235
rect 10485 3215 10500 3235
rect 10450 3185 10500 3215
rect 10450 3165 10465 3185
rect 10485 3165 10500 3185
rect 10450 3135 10500 3165
rect 10450 3115 10465 3135
rect 10485 3115 10500 3135
rect 10450 3085 10500 3115
rect 10450 3065 10465 3085
rect 10485 3065 10500 3085
rect 10450 3050 10500 3065
rect 10600 3535 10650 3600
rect 10600 3515 10615 3535
rect 10635 3515 10650 3535
rect 10600 3485 10650 3515
rect 10600 3465 10615 3485
rect 10635 3465 10650 3485
rect 10600 3435 10650 3465
rect 10600 3415 10615 3435
rect 10635 3415 10650 3435
rect 10600 3385 10650 3415
rect 10600 3365 10615 3385
rect 10635 3365 10650 3385
rect 10600 3335 10650 3365
rect 10600 3315 10615 3335
rect 10635 3315 10650 3335
rect 10600 3285 10650 3315
rect 10600 3265 10615 3285
rect 10635 3265 10650 3285
rect 10600 3235 10650 3265
rect 10600 3215 10615 3235
rect 10635 3215 10650 3235
rect 10600 3185 10650 3215
rect 10600 3165 10615 3185
rect 10635 3165 10650 3185
rect 10600 3135 10650 3165
rect 10600 3115 10615 3135
rect 10635 3115 10650 3135
rect 10600 3085 10650 3115
rect 10600 3065 10615 3085
rect 10635 3065 10650 3085
rect 10600 3050 10650 3065
rect 10750 3535 10800 3550
rect 10750 3515 10765 3535
rect 10785 3515 10800 3535
rect 10750 3485 10800 3515
rect 10750 3465 10765 3485
rect 10785 3465 10800 3485
rect 10750 3435 10800 3465
rect 10750 3415 10765 3435
rect 10785 3415 10800 3435
rect 10750 3385 10800 3415
rect 10750 3365 10765 3385
rect 10785 3365 10800 3385
rect 10750 3335 10800 3365
rect 10750 3315 10765 3335
rect 10785 3315 10800 3335
rect 10750 3285 10800 3315
rect 10750 3265 10765 3285
rect 10785 3265 10800 3285
rect 10750 3235 10800 3265
rect 10750 3215 10765 3235
rect 10785 3215 10800 3235
rect 10750 3185 10800 3215
rect 10750 3165 10765 3185
rect 10785 3165 10800 3185
rect 10750 3135 10800 3165
rect 10750 3115 10765 3135
rect 10785 3115 10800 3135
rect 10750 3085 10800 3115
rect 10750 3065 10765 3085
rect 10785 3065 10800 3085
rect 10750 3050 10800 3065
rect 11350 3535 11400 3550
rect 11350 3515 11365 3535
rect 11385 3515 11400 3535
rect 11350 3485 11400 3515
rect 11350 3465 11365 3485
rect 11385 3465 11400 3485
rect 11350 3435 11400 3465
rect 11350 3415 11365 3435
rect 11385 3415 11400 3435
rect 11350 3385 11400 3415
rect 11350 3365 11365 3385
rect 11385 3365 11400 3385
rect 11350 3335 11400 3365
rect 11350 3315 11365 3335
rect 11385 3315 11400 3335
rect 11350 3285 11400 3315
rect 11350 3265 11365 3285
rect 11385 3265 11400 3285
rect 11350 3235 11400 3265
rect 11350 3215 11365 3235
rect 11385 3215 11400 3235
rect 11350 3185 11400 3215
rect 11350 3165 11365 3185
rect 11385 3165 11400 3185
rect 11350 3135 11400 3165
rect 11350 3115 11365 3135
rect 11385 3115 11400 3135
rect 11350 3085 11400 3115
rect 11350 3065 11365 3085
rect 11385 3065 11400 3085
rect 11350 3050 11400 3065
rect 11950 3535 12000 3550
rect 11950 3515 11965 3535
rect 11985 3515 12000 3535
rect 11950 3485 12000 3515
rect 11950 3465 11965 3485
rect 11985 3465 12000 3485
rect 11950 3435 12000 3465
rect 11950 3415 11965 3435
rect 11985 3415 12000 3435
rect 11950 3385 12000 3415
rect 11950 3365 11965 3385
rect 11985 3365 12000 3385
rect 11950 3335 12000 3365
rect 11950 3315 11965 3335
rect 11985 3315 12000 3335
rect 11950 3285 12000 3315
rect 11950 3265 11965 3285
rect 11985 3265 12000 3285
rect 11950 3235 12000 3265
rect 11950 3215 11965 3235
rect 11985 3215 12000 3235
rect 11950 3185 12000 3215
rect 11950 3165 11965 3185
rect 11985 3165 12000 3185
rect 11950 3135 12000 3165
rect 11950 3115 11965 3135
rect 11985 3115 12000 3135
rect 11950 3085 12000 3115
rect 11950 3065 11965 3085
rect 11985 3065 12000 3085
rect 11950 3050 12000 3065
rect 12550 3535 12600 3550
rect 12550 3515 12565 3535
rect 12585 3515 12600 3535
rect 12550 3485 12600 3515
rect 12550 3465 12565 3485
rect 12585 3465 12600 3485
rect 12550 3435 12600 3465
rect 12550 3415 12565 3435
rect 12585 3415 12600 3435
rect 12550 3385 12600 3415
rect 12550 3365 12565 3385
rect 12585 3365 12600 3385
rect 12550 3335 12600 3365
rect 12550 3315 12565 3335
rect 12585 3315 12600 3335
rect 12550 3285 12600 3315
rect 12550 3265 12565 3285
rect 12585 3265 12600 3285
rect 12550 3235 12600 3265
rect 12550 3215 12565 3235
rect 12585 3215 12600 3235
rect 12550 3185 12600 3215
rect 12550 3165 12565 3185
rect 12585 3165 12600 3185
rect 12550 3135 12600 3165
rect 12550 3115 12565 3135
rect 12585 3115 12600 3135
rect 12550 3085 12600 3115
rect 12550 3065 12565 3085
rect 12585 3065 12600 3085
rect 12550 3050 12600 3065
rect 13150 3535 13200 3550
rect 13150 3515 13165 3535
rect 13185 3515 13200 3535
rect 13150 3485 13200 3515
rect 13150 3465 13165 3485
rect 13185 3465 13200 3485
rect 13150 3435 13200 3465
rect 13150 3415 13165 3435
rect 13185 3415 13200 3435
rect 13150 3385 13200 3415
rect 13150 3365 13165 3385
rect 13185 3365 13200 3385
rect 13150 3335 13200 3365
rect 13150 3315 13165 3335
rect 13185 3315 13200 3335
rect 13150 3285 13200 3315
rect 13150 3265 13165 3285
rect 13185 3265 13200 3285
rect 13150 3235 13200 3265
rect 13150 3215 13165 3235
rect 13185 3215 13200 3235
rect 13150 3185 13200 3215
rect 13150 3165 13165 3185
rect 13185 3165 13200 3185
rect 13150 3135 13200 3165
rect 13150 3115 13165 3135
rect 13185 3115 13200 3135
rect 13150 3085 13200 3115
rect 13150 3065 13165 3085
rect 13185 3065 13200 3085
rect 13150 3050 13200 3065
rect 13750 3535 13800 3550
rect 13750 3515 13765 3535
rect 13785 3515 13800 3535
rect 13750 3485 13800 3515
rect 13750 3465 13765 3485
rect 13785 3465 13800 3485
rect 13750 3435 13800 3465
rect 13750 3415 13765 3435
rect 13785 3415 13800 3435
rect 13750 3385 13800 3415
rect 13750 3365 13765 3385
rect 13785 3365 13800 3385
rect 13750 3335 13800 3365
rect 13750 3315 13765 3335
rect 13785 3315 13800 3335
rect 13750 3285 13800 3315
rect 13750 3265 13765 3285
rect 13785 3265 13800 3285
rect 13750 3235 13800 3265
rect 13750 3215 13765 3235
rect 13785 3215 13800 3235
rect 13750 3185 13800 3215
rect 13750 3165 13765 3185
rect 13785 3165 13800 3185
rect 13750 3135 13800 3165
rect 13750 3115 13765 3135
rect 13785 3115 13800 3135
rect 13750 3085 13800 3115
rect 13750 3065 13765 3085
rect 13785 3065 13800 3085
rect 13750 3050 13800 3065
rect 14350 3535 14400 3550
rect 14350 3515 14365 3535
rect 14385 3515 14400 3535
rect 14350 3485 14400 3515
rect 14350 3465 14365 3485
rect 14385 3465 14400 3485
rect 14350 3435 14400 3465
rect 14350 3415 14365 3435
rect 14385 3415 14400 3435
rect 14350 3385 14400 3415
rect 14350 3365 14365 3385
rect 14385 3365 14400 3385
rect 14350 3335 14400 3365
rect 14350 3315 14365 3335
rect 14385 3315 14400 3335
rect 14350 3285 14400 3315
rect 14350 3265 14365 3285
rect 14385 3265 14400 3285
rect 14350 3235 14400 3265
rect 14350 3215 14365 3235
rect 14385 3215 14400 3235
rect 14350 3185 14400 3215
rect 14350 3165 14365 3185
rect 14385 3165 14400 3185
rect 14350 3135 14400 3165
rect 14350 3115 14365 3135
rect 14385 3115 14400 3135
rect 14350 3085 14400 3115
rect 14350 3065 14365 3085
rect 14385 3065 14400 3085
rect 14350 3050 14400 3065
rect 14950 3535 15000 3550
rect 14950 3515 14965 3535
rect 14985 3515 15000 3535
rect 14950 3485 15000 3515
rect 14950 3465 14965 3485
rect 14985 3465 15000 3485
rect 14950 3435 15000 3465
rect 14950 3415 14965 3435
rect 14985 3415 15000 3435
rect 14950 3385 15000 3415
rect 14950 3365 14965 3385
rect 14985 3365 15000 3385
rect 14950 3335 15000 3365
rect 14950 3315 14965 3335
rect 14985 3315 15000 3335
rect 14950 3285 15000 3315
rect 14950 3265 14965 3285
rect 14985 3265 15000 3285
rect 14950 3235 15000 3265
rect 14950 3215 14965 3235
rect 14985 3215 15000 3235
rect 14950 3185 15000 3215
rect 14950 3165 14965 3185
rect 14985 3165 15000 3185
rect 14950 3135 15000 3165
rect 14950 3115 14965 3135
rect 14985 3115 15000 3135
rect 14950 3085 15000 3115
rect 14950 3065 14965 3085
rect 14985 3065 15000 3085
rect 14950 3050 15000 3065
rect 15550 3535 15600 3550
rect 15550 3515 15565 3535
rect 15585 3515 15600 3535
rect 15550 3485 15600 3515
rect 15550 3465 15565 3485
rect 15585 3465 15600 3485
rect 15550 3435 15600 3465
rect 15550 3415 15565 3435
rect 15585 3415 15600 3435
rect 15550 3385 15600 3415
rect 15550 3365 15565 3385
rect 15585 3365 15600 3385
rect 15550 3335 15600 3365
rect 15550 3315 15565 3335
rect 15585 3315 15600 3335
rect 15550 3285 15600 3315
rect 15550 3265 15565 3285
rect 15585 3265 15600 3285
rect 15550 3235 15600 3265
rect 15550 3215 15565 3235
rect 15585 3215 15600 3235
rect 15550 3185 15600 3215
rect 15550 3165 15565 3185
rect 15585 3165 15600 3185
rect 15550 3135 15600 3165
rect 15550 3115 15565 3135
rect 15585 3115 15600 3135
rect 15550 3085 15600 3115
rect 15550 3065 15565 3085
rect 15585 3065 15600 3085
rect 15550 3050 15600 3065
rect 16150 3535 16200 3550
rect 16150 3515 16165 3535
rect 16185 3515 16200 3535
rect 16150 3485 16200 3515
rect 16150 3465 16165 3485
rect 16185 3465 16200 3485
rect 16150 3435 16200 3465
rect 16150 3415 16165 3435
rect 16185 3415 16200 3435
rect 16150 3385 16200 3415
rect 16150 3365 16165 3385
rect 16185 3365 16200 3385
rect 16150 3335 16200 3365
rect 16150 3315 16165 3335
rect 16185 3315 16200 3335
rect 16150 3285 16200 3315
rect 16150 3265 16165 3285
rect 16185 3265 16200 3285
rect 16150 3235 16200 3265
rect 16150 3215 16165 3235
rect 16185 3215 16200 3235
rect 16150 3185 16200 3215
rect 16150 3165 16165 3185
rect 16185 3165 16200 3185
rect 16150 3135 16200 3165
rect 16150 3115 16165 3135
rect 16185 3115 16200 3135
rect 16150 3085 16200 3115
rect 16150 3065 16165 3085
rect 16185 3065 16200 3085
rect 16150 3050 16200 3065
rect 16300 3535 16350 3550
rect 16300 3515 16315 3535
rect 16335 3515 16350 3535
rect 16300 3485 16350 3515
rect 16300 3465 16315 3485
rect 16335 3465 16350 3485
rect 16300 3435 16350 3465
rect 16300 3415 16315 3435
rect 16335 3415 16350 3435
rect 16300 3385 16350 3415
rect 16300 3365 16315 3385
rect 16335 3365 16350 3385
rect 16300 3335 16350 3365
rect 16300 3315 16315 3335
rect 16335 3315 16350 3335
rect 16300 3285 16350 3315
rect 16300 3265 16315 3285
rect 16335 3265 16350 3285
rect 16300 3235 16350 3265
rect 16300 3215 16315 3235
rect 16335 3215 16350 3235
rect 16300 3185 16350 3215
rect 16300 3165 16315 3185
rect 16335 3165 16350 3185
rect 16300 3135 16350 3165
rect 16300 3115 16315 3135
rect 16335 3115 16350 3135
rect 16300 3085 16350 3115
rect 16300 3065 16315 3085
rect 16335 3065 16350 3085
rect 16300 3050 16350 3065
rect 16450 3535 16500 3550
rect 16450 3515 16465 3535
rect 16485 3515 16500 3535
rect 16450 3485 16500 3515
rect 16450 3465 16465 3485
rect 16485 3465 16500 3485
rect 16450 3435 16500 3465
rect 16450 3415 16465 3435
rect 16485 3415 16500 3435
rect 16450 3385 16500 3415
rect 16450 3365 16465 3385
rect 16485 3365 16500 3385
rect 16450 3335 16500 3365
rect 16450 3315 16465 3335
rect 16485 3315 16500 3335
rect 16450 3285 16500 3315
rect 16450 3265 16465 3285
rect 16485 3265 16500 3285
rect 16450 3235 16500 3265
rect 16450 3215 16465 3235
rect 16485 3215 16500 3235
rect 16450 3185 16500 3215
rect 16450 3165 16465 3185
rect 16485 3165 16500 3185
rect 16450 3135 16500 3165
rect 16450 3115 16465 3135
rect 16485 3115 16500 3135
rect 16450 3085 16500 3115
rect 16450 3065 16465 3085
rect 16485 3065 16500 3085
rect 16450 3050 16500 3065
rect 16600 3535 16650 3550
rect 16600 3515 16615 3535
rect 16635 3515 16650 3535
rect 16600 3485 16650 3515
rect 16600 3465 16615 3485
rect 16635 3465 16650 3485
rect 16600 3435 16650 3465
rect 16600 3415 16615 3435
rect 16635 3415 16650 3435
rect 16600 3385 16650 3415
rect 16600 3365 16615 3385
rect 16635 3365 16650 3385
rect 16600 3335 16650 3365
rect 16600 3315 16615 3335
rect 16635 3315 16650 3335
rect 16600 3285 16650 3315
rect 16600 3265 16615 3285
rect 16635 3265 16650 3285
rect 16600 3235 16650 3265
rect 16600 3215 16615 3235
rect 16635 3215 16650 3235
rect 16600 3185 16650 3215
rect 16600 3165 16615 3185
rect 16635 3165 16650 3185
rect 16600 3135 16650 3165
rect 16600 3115 16615 3135
rect 16635 3115 16650 3135
rect 16600 3085 16650 3115
rect 16600 3065 16615 3085
rect 16635 3065 16650 3085
rect 16600 3050 16650 3065
rect 16750 3535 16800 3550
rect 16750 3515 16765 3535
rect 16785 3515 16800 3535
rect 16750 3485 16800 3515
rect 16750 3465 16765 3485
rect 16785 3465 16800 3485
rect 16750 3435 16800 3465
rect 16750 3415 16765 3435
rect 16785 3415 16800 3435
rect 16750 3385 16800 3415
rect 16750 3365 16765 3385
rect 16785 3365 16800 3385
rect 16750 3335 16800 3365
rect 16750 3315 16765 3335
rect 16785 3315 16800 3335
rect 16750 3285 16800 3315
rect 16750 3265 16765 3285
rect 16785 3265 16800 3285
rect 16750 3235 16800 3265
rect 16750 3215 16765 3235
rect 16785 3215 16800 3235
rect 16750 3185 16800 3215
rect 16750 3165 16765 3185
rect 16785 3165 16800 3185
rect 16750 3135 16800 3165
rect 16750 3115 16765 3135
rect 16785 3115 16800 3135
rect 16750 3085 16800 3115
rect 16750 3065 16765 3085
rect 16785 3065 16800 3085
rect 16750 3050 16800 3065
rect 16900 3535 16950 3550
rect 16900 3515 16915 3535
rect 16935 3515 16950 3535
rect 16900 3485 16950 3515
rect 16900 3465 16915 3485
rect 16935 3465 16950 3485
rect 16900 3435 16950 3465
rect 16900 3415 16915 3435
rect 16935 3415 16950 3435
rect 16900 3385 16950 3415
rect 16900 3365 16915 3385
rect 16935 3365 16950 3385
rect 16900 3335 16950 3365
rect 16900 3315 16915 3335
rect 16935 3315 16950 3335
rect 16900 3285 16950 3315
rect 16900 3265 16915 3285
rect 16935 3265 16950 3285
rect 16900 3235 16950 3265
rect 16900 3215 16915 3235
rect 16935 3215 16950 3235
rect 16900 3185 16950 3215
rect 16900 3165 16915 3185
rect 16935 3165 16950 3185
rect 16900 3135 16950 3165
rect 16900 3115 16915 3135
rect 16935 3115 16950 3135
rect 16900 3085 16950 3115
rect 16900 3065 16915 3085
rect 16935 3065 16950 3085
rect 16900 3050 16950 3065
rect 17050 3535 17100 3550
rect 17050 3515 17065 3535
rect 17085 3515 17100 3535
rect 17050 3485 17100 3515
rect 17050 3465 17065 3485
rect 17085 3465 17100 3485
rect 17050 3435 17100 3465
rect 17050 3415 17065 3435
rect 17085 3415 17100 3435
rect 17050 3385 17100 3415
rect 17050 3365 17065 3385
rect 17085 3365 17100 3385
rect 17050 3335 17100 3365
rect 17050 3315 17065 3335
rect 17085 3315 17100 3335
rect 17050 3285 17100 3315
rect 17050 3265 17065 3285
rect 17085 3265 17100 3285
rect 17050 3235 17100 3265
rect 17050 3215 17065 3235
rect 17085 3215 17100 3235
rect 17050 3185 17100 3215
rect 17050 3165 17065 3185
rect 17085 3165 17100 3185
rect 17050 3135 17100 3165
rect 17050 3115 17065 3135
rect 17085 3115 17100 3135
rect 17050 3085 17100 3115
rect 17050 3065 17065 3085
rect 17085 3065 17100 3085
rect 17050 3050 17100 3065
rect 17200 3535 17250 3550
rect 17200 3515 17215 3535
rect 17235 3515 17250 3535
rect 17200 3485 17250 3515
rect 17200 3465 17215 3485
rect 17235 3465 17250 3485
rect 17200 3435 17250 3465
rect 17200 3415 17215 3435
rect 17235 3415 17250 3435
rect 17200 3385 17250 3415
rect 17200 3365 17215 3385
rect 17235 3365 17250 3385
rect 17200 3335 17250 3365
rect 17200 3315 17215 3335
rect 17235 3315 17250 3335
rect 17200 3285 17250 3315
rect 17200 3265 17215 3285
rect 17235 3265 17250 3285
rect 17200 3235 17250 3265
rect 17200 3215 17215 3235
rect 17235 3215 17250 3235
rect 17200 3185 17250 3215
rect 17200 3165 17215 3185
rect 17235 3165 17250 3185
rect 17200 3135 17250 3165
rect 17200 3115 17215 3135
rect 17235 3115 17250 3135
rect 17200 3085 17250 3115
rect 17200 3065 17215 3085
rect 17235 3065 17250 3085
rect 17200 3050 17250 3065
rect 17350 3535 17400 3550
rect 17350 3515 17365 3535
rect 17385 3515 17400 3535
rect 17350 3485 17400 3515
rect 17350 3465 17365 3485
rect 17385 3465 17400 3485
rect 17350 3435 17400 3465
rect 17350 3415 17365 3435
rect 17385 3415 17400 3435
rect 17350 3385 17400 3415
rect 17350 3365 17365 3385
rect 17385 3365 17400 3385
rect 17350 3335 17400 3365
rect 17350 3315 17365 3335
rect 17385 3315 17400 3335
rect 17350 3285 17400 3315
rect 17350 3265 17365 3285
rect 17385 3265 17400 3285
rect 17350 3235 17400 3265
rect 17350 3215 17365 3235
rect 17385 3215 17400 3235
rect 17350 3185 17400 3215
rect 17350 3165 17365 3185
rect 17385 3165 17400 3185
rect 17350 3135 17400 3165
rect 17350 3115 17365 3135
rect 17385 3115 17400 3135
rect 17350 3085 17400 3115
rect 17350 3065 17365 3085
rect 17385 3065 17400 3085
rect 17350 3050 17400 3065
rect 17950 3535 18000 3550
rect 17950 3515 17965 3535
rect 17985 3515 18000 3535
rect 17950 3485 18000 3515
rect 17950 3465 17965 3485
rect 17985 3465 18000 3485
rect 17950 3435 18000 3465
rect 17950 3415 17965 3435
rect 17985 3415 18000 3435
rect 17950 3385 18000 3415
rect 17950 3365 17965 3385
rect 17985 3365 18000 3385
rect 17950 3335 18000 3365
rect 17950 3315 17965 3335
rect 17985 3315 18000 3335
rect 17950 3285 18000 3315
rect 17950 3265 17965 3285
rect 17985 3265 18000 3285
rect 17950 3235 18000 3265
rect 17950 3215 17965 3235
rect 17985 3215 18000 3235
rect 17950 3185 18000 3215
rect 17950 3165 17965 3185
rect 17985 3165 18000 3185
rect 17950 3135 18000 3165
rect 17950 3115 17965 3135
rect 17985 3115 18000 3135
rect 17950 3085 18000 3115
rect 17950 3065 17965 3085
rect 17985 3065 18000 3085
rect 17950 3050 18000 3065
rect 18550 3535 18600 3550
rect 18550 3515 18565 3535
rect 18585 3515 18600 3535
rect 18550 3485 18600 3515
rect 18550 3465 18565 3485
rect 18585 3465 18600 3485
rect 18550 3435 18600 3465
rect 18550 3415 18565 3435
rect 18585 3415 18600 3435
rect 18550 3385 18600 3415
rect 18550 3365 18565 3385
rect 18585 3365 18600 3385
rect 18550 3335 18600 3365
rect 18550 3315 18565 3335
rect 18585 3315 18600 3335
rect 18550 3285 18600 3315
rect 18550 3265 18565 3285
rect 18585 3265 18600 3285
rect 18550 3235 18600 3265
rect 18550 3215 18565 3235
rect 18585 3215 18600 3235
rect 18550 3185 18600 3215
rect 18550 3165 18565 3185
rect 18585 3165 18600 3185
rect 18550 3135 18600 3165
rect 18550 3115 18565 3135
rect 18585 3115 18600 3135
rect 18550 3085 18600 3115
rect 18550 3065 18565 3085
rect 18585 3065 18600 3085
rect 18550 3050 18600 3065
rect 18700 3535 18750 3550
rect 18700 3515 18715 3535
rect 18735 3515 18750 3535
rect 18700 3485 18750 3515
rect 18700 3465 18715 3485
rect 18735 3465 18750 3485
rect 18700 3435 18750 3465
rect 18700 3415 18715 3435
rect 18735 3415 18750 3435
rect 18700 3385 18750 3415
rect 18700 3365 18715 3385
rect 18735 3365 18750 3385
rect 18700 3335 18750 3365
rect 18700 3315 18715 3335
rect 18735 3315 18750 3335
rect 18700 3285 18750 3315
rect 18700 3265 18715 3285
rect 18735 3265 18750 3285
rect 18700 3235 18750 3265
rect 18700 3215 18715 3235
rect 18735 3215 18750 3235
rect 18700 3185 18750 3215
rect 18700 3165 18715 3185
rect 18735 3165 18750 3185
rect 18700 3135 18750 3165
rect 18700 3115 18715 3135
rect 18735 3115 18750 3135
rect 18700 3085 18750 3115
rect 18700 3065 18715 3085
rect 18735 3065 18750 3085
rect 18700 3050 18750 3065
rect 18850 3535 18900 3550
rect 18850 3515 18865 3535
rect 18885 3515 18900 3535
rect 18850 3485 18900 3515
rect 18850 3465 18865 3485
rect 18885 3465 18900 3485
rect 18850 3435 18900 3465
rect 18850 3415 18865 3435
rect 18885 3415 18900 3435
rect 18850 3385 18900 3415
rect 18850 3365 18865 3385
rect 18885 3365 18900 3385
rect 18850 3335 18900 3365
rect 18850 3315 18865 3335
rect 18885 3315 18900 3335
rect 18850 3285 18900 3315
rect 18850 3265 18865 3285
rect 18885 3265 18900 3285
rect 18850 3235 18900 3265
rect 18850 3215 18865 3235
rect 18885 3215 18900 3235
rect 18850 3185 18900 3215
rect 18850 3165 18865 3185
rect 18885 3165 18900 3185
rect 18850 3135 18900 3165
rect 18850 3115 18865 3135
rect 18885 3115 18900 3135
rect 18850 3085 18900 3115
rect 18850 3065 18865 3085
rect 18885 3065 18900 3085
rect 18850 3050 18900 3065
rect 19000 3535 19050 3550
rect 19000 3515 19015 3535
rect 19035 3515 19050 3535
rect 19000 3485 19050 3515
rect 19000 3465 19015 3485
rect 19035 3465 19050 3485
rect 19000 3435 19050 3465
rect 19000 3415 19015 3435
rect 19035 3415 19050 3435
rect 19000 3385 19050 3415
rect 19000 3365 19015 3385
rect 19035 3365 19050 3385
rect 19000 3335 19050 3365
rect 19000 3315 19015 3335
rect 19035 3315 19050 3335
rect 19000 3285 19050 3315
rect 19000 3265 19015 3285
rect 19035 3265 19050 3285
rect 19000 3235 19050 3265
rect 19000 3215 19015 3235
rect 19035 3215 19050 3235
rect 19000 3185 19050 3215
rect 19000 3165 19015 3185
rect 19035 3165 19050 3185
rect 19000 3135 19050 3165
rect 19000 3115 19015 3135
rect 19035 3115 19050 3135
rect 19000 3085 19050 3115
rect 19000 3065 19015 3085
rect 19035 3065 19050 3085
rect 19000 3050 19050 3065
rect 19150 3535 19200 3550
rect 19150 3515 19165 3535
rect 19185 3515 19200 3535
rect 19150 3485 19200 3515
rect 19150 3465 19165 3485
rect 19185 3465 19200 3485
rect 19150 3435 19200 3465
rect 19150 3415 19165 3435
rect 19185 3415 19200 3435
rect 19150 3385 19200 3415
rect 19150 3365 19165 3385
rect 19185 3365 19200 3385
rect 19150 3335 19200 3365
rect 19150 3315 19165 3335
rect 19185 3315 19200 3335
rect 19150 3285 19200 3315
rect 19150 3265 19165 3285
rect 19185 3265 19200 3285
rect 19150 3235 19200 3265
rect 19150 3215 19165 3235
rect 19185 3215 19200 3235
rect 19150 3185 19200 3215
rect 19150 3165 19165 3185
rect 19185 3165 19200 3185
rect 19150 3135 19200 3165
rect 19150 3115 19165 3135
rect 19185 3115 19200 3135
rect 19150 3085 19200 3115
rect 19150 3065 19165 3085
rect 19185 3065 19200 3085
rect 19150 3050 19200 3065
rect 19300 3535 19350 3550
rect 19300 3515 19315 3535
rect 19335 3515 19350 3535
rect 19300 3485 19350 3515
rect 19300 3465 19315 3485
rect 19335 3465 19350 3485
rect 19300 3435 19350 3465
rect 19300 3415 19315 3435
rect 19335 3415 19350 3435
rect 19300 3385 19350 3415
rect 19300 3365 19315 3385
rect 19335 3365 19350 3385
rect 19300 3335 19350 3365
rect 19300 3315 19315 3335
rect 19335 3315 19350 3335
rect 19300 3285 19350 3315
rect 19300 3265 19315 3285
rect 19335 3265 19350 3285
rect 19300 3235 19350 3265
rect 19300 3215 19315 3235
rect 19335 3215 19350 3235
rect 19300 3185 19350 3215
rect 19300 3165 19315 3185
rect 19335 3165 19350 3185
rect 19300 3135 19350 3165
rect 19300 3115 19315 3135
rect 19335 3115 19350 3135
rect 19300 3085 19350 3115
rect 19300 3065 19315 3085
rect 19335 3065 19350 3085
rect 19300 3050 19350 3065
rect 19450 3535 19500 3550
rect 19450 3515 19465 3535
rect 19485 3515 19500 3535
rect 19450 3485 19500 3515
rect 19450 3465 19465 3485
rect 19485 3465 19500 3485
rect 19450 3435 19500 3465
rect 19450 3415 19465 3435
rect 19485 3415 19500 3435
rect 19450 3385 19500 3415
rect 19450 3365 19465 3385
rect 19485 3365 19500 3385
rect 19450 3335 19500 3365
rect 19450 3315 19465 3335
rect 19485 3315 19500 3335
rect 19450 3285 19500 3315
rect 19450 3265 19465 3285
rect 19485 3265 19500 3285
rect 19450 3235 19500 3265
rect 19450 3215 19465 3235
rect 19485 3215 19500 3235
rect 19450 3185 19500 3215
rect 19450 3165 19465 3185
rect 19485 3165 19500 3185
rect 19450 3135 19500 3165
rect 19450 3115 19465 3135
rect 19485 3115 19500 3135
rect 19450 3085 19500 3115
rect 19450 3065 19465 3085
rect 19485 3065 19500 3085
rect 19450 3050 19500 3065
rect 19600 3535 19650 3550
rect 19600 3515 19615 3535
rect 19635 3515 19650 3535
rect 19600 3485 19650 3515
rect 19600 3465 19615 3485
rect 19635 3465 19650 3485
rect 19600 3435 19650 3465
rect 19600 3415 19615 3435
rect 19635 3415 19650 3435
rect 19600 3385 19650 3415
rect 19600 3365 19615 3385
rect 19635 3365 19650 3385
rect 19600 3335 19650 3365
rect 19600 3315 19615 3335
rect 19635 3315 19650 3335
rect 19600 3285 19650 3315
rect 19600 3265 19615 3285
rect 19635 3265 19650 3285
rect 19600 3235 19650 3265
rect 19600 3215 19615 3235
rect 19635 3215 19650 3235
rect 19600 3185 19650 3215
rect 19600 3165 19615 3185
rect 19635 3165 19650 3185
rect 19600 3135 19650 3165
rect 19600 3115 19615 3135
rect 19635 3115 19650 3135
rect 19600 3085 19650 3115
rect 19600 3065 19615 3085
rect 19635 3065 19650 3085
rect 19600 3050 19650 3065
rect 19750 3535 19800 3550
rect 19750 3515 19765 3535
rect 19785 3515 19800 3535
rect 19750 3485 19800 3515
rect 19750 3465 19765 3485
rect 19785 3465 19800 3485
rect 19750 3435 19800 3465
rect 19750 3415 19765 3435
rect 19785 3415 19800 3435
rect 19750 3385 19800 3415
rect 19750 3365 19765 3385
rect 19785 3365 19800 3385
rect 19750 3335 19800 3365
rect 19750 3315 19765 3335
rect 19785 3315 19800 3335
rect 19750 3285 19800 3315
rect 19750 3265 19765 3285
rect 19785 3265 19800 3285
rect 19750 3235 19800 3265
rect 19750 3215 19765 3235
rect 19785 3215 19800 3235
rect 19750 3185 19800 3215
rect 19750 3165 19765 3185
rect 19785 3165 19800 3185
rect 19750 3135 19800 3165
rect 19750 3115 19765 3135
rect 19785 3115 19800 3135
rect 19750 3085 19800 3115
rect 19750 3065 19765 3085
rect 19785 3065 19800 3085
rect 19750 3050 19800 3065
rect 20350 3535 20400 3550
rect 20350 3515 20365 3535
rect 20385 3515 20400 3535
rect 20350 3485 20400 3515
rect 20350 3465 20365 3485
rect 20385 3465 20400 3485
rect 20350 3435 20400 3465
rect 20350 3415 20365 3435
rect 20385 3415 20400 3435
rect 20350 3385 20400 3415
rect 20350 3365 20365 3385
rect 20385 3365 20400 3385
rect 20350 3335 20400 3365
rect 20350 3315 20365 3335
rect 20385 3315 20400 3335
rect 20350 3285 20400 3315
rect 20350 3265 20365 3285
rect 20385 3265 20400 3285
rect 20350 3235 20400 3265
rect 20350 3215 20365 3235
rect 20385 3215 20400 3235
rect 20350 3185 20400 3215
rect 20350 3165 20365 3185
rect 20385 3165 20400 3185
rect 20350 3135 20400 3165
rect 20350 3115 20365 3135
rect 20385 3115 20400 3135
rect 20350 3085 20400 3115
rect 20350 3065 20365 3085
rect 20385 3065 20400 3085
rect 20350 3050 20400 3065
rect 20950 3535 21000 3550
rect 20950 3515 20965 3535
rect 20985 3515 21000 3535
rect 20950 3485 21000 3515
rect 20950 3465 20965 3485
rect 20985 3465 21000 3485
rect 20950 3435 21000 3465
rect 20950 3415 20965 3435
rect 20985 3415 21000 3435
rect 20950 3385 21000 3415
rect 20950 3365 20965 3385
rect 20985 3365 21000 3385
rect 20950 3335 21000 3365
rect 20950 3315 20965 3335
rect 20985 3315 21000 3335
rect 20950 3285 21000 3315
rect 20950 3265 20965 3285
rect 20985 3265 21000 3285
rect 20950 3235 21000 3265
rect 20950 3215 20965 3235
rect 20985 3215 21000 3235
rect 20950 3185 21000 3215
rect 20950 3165 20965 3185
rect 20985 3165 21000 3185
rect 20950 3135 21000 3165
rect 20950 3115 20965 3135
rect 20985 3115 21000 3135
rect 20950 3085 21000 3115
rect 20950 3065 20965 3085
rect 20985 3065 21000 3085
rect 20950 3050 21000 3065
rect 21400 3535 21450 3550
rect 21400 3515 21415 3535
rect 21435 3515 21450 3535
rect 21400 3485 21450 3515
rect 21400 3465 21415 3485
rect 21435 3465 21450 3485
rect 21400 3435 21450 3465
rect 21400 3415 21415 3435
rect 21435 3415 21450 3435
rect 21400 3385 21450 3415
rect 21400 3365 21415 3385
rect 21435 3365 21450 3385
rect 21400 3335 21450 3365
rect 21400 3315 21415 3335
rect 21435 3315 21450 3335
rect 21400 3285 21450 3315
rect 21400 3265 21415 3285
rect 21435 3265 21450 3285
rect 21400 3235 21450 3265
rect 21400 3215 21415 3235
rect 21435 3215 21450 3235
rect 21400 3185 21450 3215
rect 21400 3165 21415 3185
rect 21435 3165 21450 3185
rect 21400 3135 21450 3165
rect 21400 3115 21415 3135
rect 21435 3115 21450 3135
rect 21400 3085 21450 3115
rect 21400 3065 21415 3085
rect 21435 3065 21450 3085
rect 21400 3050 21450 3065
rect 21850 3535 21900 3550
rect 21850 3515 21865 3535
rect 21885 3515 21900 3535
rect 21850 3485 21900 3515
rect 21850 3465 21865 3485
rect 21885 3465 21900 3485
rect 21850 3435 21900 3465
rect 21850 3415 21865 3435
rect 21885 3415 21900 3435
rect 21850 3385 21900 3415
rect 21850 3365 21865 3385
rect 21885 3365 21900 3385
rect 21850 3335 21900 3365
rect 21850 3315 21865 3335
rect 21885 3315 21900 3335
rect 21850 3285 21900 3315
rect 21850 3265 21865 3285
rect 21885 3265 21900 3285
rect 21850 3235 21900 3265
rect 21850 3215 21865 3235
rect 21885 3215 21900 3235
rect 21850 3185 21900 3215
rect 21850 3165 21865 3185
rect 21885 3165 21900 3185
rect 21850 3135 21900 3165
rect 21850 3115 21865 3135
rect 21885 3115 21900 3135
rect 21850 3085 21900 3115
rect 21850 3065 21865 3085
rect 21885 3065 21900 3085
rect 21850 3050 21900 3065
rect 22450 3535 22500 3550
rect 22450 3515 22465 3535
rect 22485 3515 22500 3535
rect 22450 3485 22500 3515
rect 22450 3465 22465 3485
rect 22485 3465 22500 3485
rect 22450 3435 22500 3465
rect 22450 3415 22465 3435
rect 22485 3415 22500 3435
rect 22450 3385 22500 3415
rect 22450 3365 22465 3385
rect 22485 3365 22500 3385
rect 22450 3335 22500 3365
rect 22450 3315 22465 3335
rect 22485 3315 22500 3335
rect 22450 3285 22500 3315
rect 22450 3265 22465 3285
rect 22485 3265 22500 3285
rect 22450 3235 22500 3265
rect 22450 3215 22465 3235
rect 22485 3215 22500 3235
rect 22450 3185 22500 3215
rect 22450 3165 22465 3185
rect 22485 3165 22500 3185
rect 22450 3135 22500 3165
rect 22450 3115 22465 3135
rect 22485 3115 22500 3135
rect 22450 3085 22500 3115
rect 22450 3065 22465 3085
rect 22485 3065 22500 3085
rect 22450 3050 22500 3065
rect 23050 3535 23100 3550
rect 23050 3515 23065 3535
rect 23085 3515 23100 3535
rect 23050 3485 23100 3515
rect 23050 3465 23065 3485
rect 23085 3465 23100 3485
rect 23050 3435 23100 3465
rect 23050 3415 23065 3435
rect 23085 3415 23100 3435
rect 23050 3385 23100 3415
rect 23050 3365 23065 3385
rect 23085 3365 23100 3385
rect 23050 3335 23100 3365
rect 23050 3315 23065 3335
rect 23085 3315 23100 3335
rect 23050 3285 23100 3315
rect 23050 3265 23065 3285
rect 23085 3265 23100 3285
rect 23050 3235 23100 3265
rect 23050 3215 23065 3235
rect 23085 3215 23100 3235
rect 23050 3185 23100 3215
rect 23050 3165 23065 3185
rect 23085 3165 23100 3185
rect 23050 3135 23100 3165
rect 23050 3115 23065 3135
rect 23085 3115 23100 3135
rect 23050 3085 23100 3115
rect 23050 3065 23065 3085
rect 23085 3065 23100 3085
rect 23050 3050 23100 3065
rect 23500 3535 23550 3550
rect 23500 3515 23515 3535
rect 23535 3515 23550 3535
rect 23500 3485 23550 3515
rect 23500 3465 23515 3485
rect 23535 3465 23550 3485
rect 23500 3435 23550 3465
rect 23500 3415 23515 3435
rect 23535 3415 23550 3435
rect 23500 3385 23550 3415
rect 23500 3365 23515 3385
rect 23535 3365 23550 3385
rect 23500 3335 23550 3365
rect 23500 3315 23515 3335
rect 23535 3315 23550 3335
rect 23500 3285 23550 3315
rect 23500 3265 23515 3285
rect 23535 3265 23550 3285
rect 23500 3235 23550 3265
rect 23500 3215 23515 3235
rect 23535 3215 23550 3235
rect 23500 3185 23550 3215
rect 23500 3165 23515 3185
rect 23535 3165 23550 3185
rect 23500 3135 23550 3165
rect 23500 3115 23515 3135
rect 23535 3115 23550 3135
rect 23500 3085 23550 3115
rect 23500 3065 23515 3085
rect 23535 3065 23550 3085
rect 23500 3050 23550 3065
rect 23950 3535 24000 3550
rect 23950 3515 23965 3535
rect 23985 3515 24000 3535
rect 23950 3485 24000 3515
rect 23950 3465 23965 3485
rect 23985 3465 24000 3485
rect 23950 3435 24000 3465
rect 23950 3415 23965 3435
rect 23985 3415 24000 3435
rect 23950 3385 24000 3415
rect 23950 3365 23965 3385
rect 23985 3365 24000 3385
rect 23950 3335 24000 3365
rect 23950 3315 23965 3335
rect 23985 3315 24000 3335
rect 23950 3285 24000 3315
rect 23950 3265 23965 3285
rect 23985 3265 24000 3285
rect 23950 3235 24000 3265
rect 23950 3215 23965 3235
rect 23985 3215 24000 3235
rect 23950 3185 24000 3215
rect 23950 3165 23965 3185
rect 23985 3165 24000 3185
rect 23950 3135 24000 3165
rect 23950 3115 23965 3135
rect 23985 3115 24000 3135
rect 23950 3085 24000 3115
rect 23950 3065 23965 3085
rect 23985 3065 24000 3085
rect 23950 3050 24000 3065
rect 24550 3535 24600 3550
rect 24550 3515 24565 3535
rect 24585 3515 24600 3535
rect 24550 3485 24600 3515
rect 24550 3465 24565 3485
rect 24585 3465 24600 3485
rect 24550 3435 24600 3465
rect 24550 3415 24565 3435
rect 24585 3415 24600 3435
rect 24550 3385 24600 3415
rect 24550 3365 24565 3385
rect 24585 3365 24600 3385
rect 24550 3335 24600 3365
rect 24550 3315 24565 3335
rect 24585 3315 24600 3335
rect 24550 3285 24600 3315
rect 24550 3265 24565 3285
rect 24585 3265 24600 3285
rect 24550 3235 24600 3265
rect 24550 3215 24565 3235
rect 24585 3215 24600 3235
rect 24550 3185 24600 3215
rect 24550 3165 24565 3185
rect 24585 3165 24600 3185
rect 24550 3135 24600 3165
rect 24550 3115 24565 3135
rect 24585 3115 24600 3135
rect 24550 3085 24600 3115
rect 24550 3065 24565 3085
rect 24585 3065 24600 3085
rect 24550 3050 24600 3065
rect 25150 3535 25200 3550
rect 25150 3515 25165 3535
rect 25185 3515 25200 3535
rect 25150 3485 25200 3515
rect 25150 3465 25165 3485
rect 25185 3465 25200 3485
rect 25150 3435 25200 3465
rect 25150 3415 25165 3435
rect 25185 3415 25200 3435
rect 25150 3385 25200 3415
rect 25150 3365 25165 3385
rect 25185 3365 25200 3385
rect 25150 3335 25200 3365
rect 25150 3315 25165 3335
rect 25185 3315 25200 3335
rect 25150 3285 25200 3315
rect 25150 3265 25165 3285
rect 25185 3265 25200 3285
rect 25150 3235 25200 3265
rect 25150 3215 25165 3235
rect 25185 3215 25200 3235
rect 25150 3185 25200 3215
rect 25150 3165 25165 3185
rect 25185 3165 25200 3185
rect 25150 3135 25200 3165
rect 25150 3115 25165 3135
rect 25185 3115 25200 3135
rect 25150 3085 25200 3115
rect 25150 3065 25165 3085
rect 25185 3065 25200 3085
rect 25150 3050 25200 3065
rect 25600 3535 25650 3550
rect 25600 3515 25615 3535
rect 25635 3515 25650 3535
rect 25600 3485 25650 3515
rect 25600 3465 25615 3485
rect 25635 3465 25650 3485
rect 25600 3435 25650 3465
rect 25600 3415 25615 3435
rect 25635 3415 25650 3435
rect 25600 3385 25650 3415
rect 25600 3365 25615 3385
rect 25635 3365 25650 3385
rect 25600 3335 25650 3365
rect 25600 3315 25615 3335
rect 25635 3315 25650 3335
rect 25600 3285 25650 3315
rect 25600 3265 25615 3285
rect 25635 3265 25650 3285
rect 25600 3235 25650 3265
rect 25600 3215 25615 3235
rect 25635 3215 25650 3235
rect 25600 3185 25650 3215
rect 25600 3165 25615 3185
rect 25635 3165 25650 3185
rect 25600 3135 25650 3165
rect 25600 3115 25615 3135
rect 25635 3115 25650 3135
rect 25600 3085 25650 3115
rect 25600 3065 25615 3085
rect 25635 3065 25650 3085
rect 25600 3050 25650 3065
rect 26050 3535 26100 3550
rect 26050 3515 26065 3535
rect 26085 3515 26100 3535
rect 26050 3485 26100 3515
rect 26050 3465 26065 3485
rect 26085 3465 26100 3485
rect 26050 3435 26100 3465
rect 26050 3415 26065 3435
rect 26085 3415 26100 3435
rect 26050 3385 26100 3415
rect 26050 3365 26065 3385
rect 26085 3365 26100 3385
rect 26050 3335 26100 3365
rect 26050 3315 26065 3335
rect 26085 3315 26100 3335
rect 26050 3285 26100 3315
rect 26050 3265 26065 3285
rect 26085 3265 26100 3285
rect 26050 3235 26100 3265
rect 26050 3215 26065 3235
rect 26085 3215 26100 3235
rect 26050 3185 26100 3215
rect 26050 3165 26065 3185
rect 26085 3165 26100 3185
rect 26050 3135 26100 3165
rect 26050 3115 26065 3135
rect 26085 3115 26100 3135
rect 26050 3085 26100 3115
rect 26050 3065 26065 3085
rect 26085 3065 26100 3085
rect 26050 3050 26100 3065
rect 26650 3535 26700 3550
rect 26650 3515 26665 3535
rect 26685 3515 26700 3535
rect 26650 3485 26700 3515
rect 26650 3465 26665 3485
rect 26685 3465 26700 3485
rect 26650 3435 26700 3465
rect 26650 3415 26665 3435
rect 26685 3415 26700 3435
rect 26650 3385 26700 3415
rect 26650 3365 26665 3385
rect 26685 3365 26700 3385
rect 26650 3335 26700 3365
rect 26650 3315 26665 3335
rect 26685 3315 26700 3335
rect 26650 3285 26700 3315
rect 26650 3265 26665 3285
rect 26685 3265 26700 3285
rect 26650 3235 26700 3265
rect 26650 3215 26665 3235
rect 26685 3215 26700 3235
rect 26650 3185 26700 3215
rect 26650 3165 26665 3185
rect 26685 3165 26700 3185
rect 26650 3135 26700 3165
rect 26650 3115 26665 3135
rect 26685 3115 26700 3135
rect 26650 3085 26700 3115
rect 26650 3065 26665 3085
rect 26685 3065 26700 3085
rect 26650 3050 26700 3065
rect 27250 3535 27300 3550
rect 27250 3515 27265 3535
rect 27285 3515 27300 3535
rect 27250 3485 27300 3515
rect 27250 3465 27265 3485
rect 27285 3465 27300 3485
rect 27250 3435 27300 3465
rect 27250 3415 27265 3435
rect 27285 3415 27300 3435
rect 27250 3385 27300 3415
rect 27250 3365 27265 3385
rect 27285 3365 27300 3385
rect 27250 3335 27300 3365
rect 27250 3315 27265 3335
rect 27285 3315 27300 3335
rect 27250 3285 27300 3315
rect 27250 3265 27265 3285
rect 27285 3265 27300 3285
rect 27250 3235 27300 3265
rect 27250 3215 27265 3235
rect 27285 3215 27300 3235
rect 27250 3185 27300 3215
rect 27250 3165 27265 3185
rect 27285 3165 27300 3185
rect 27250 3135 27300 3165
rect 27250 3115 27265 3135
rect 27285 3115 27300 3135
rect 27250 3085 27300 3115
rect 27250 3065 27265 3085
rect 27285 3065 27300 3085
rect 27250 3050 27300 3065
rect 27700 3535 27750 3550
rect 27700 3515 27715 3535
rect 27735 3515 27750 3535
rect 27700 3485 27750 3515
rect 27700 3465 27715 3485
rect 27735 3465 27750 3485
rect 27700 3435 27750 3465
rect 27700 3415 27715 3435
rect 27735 3415 27750 3435
rect 27700 3385 27750 3415
rect 27700 3365 27715 3385
rect 27735 3365 27750 3385
rect 27700 3335 27750 3365
rect 27700 3315 27715 3335
rect 27735 3315 27750 3335
rect 27700 3285 27750 3315
rect 27700 3265 27715 3285
rect 27735 3265 27750 3285
rect 27700 3235 27750 3265
rect 27700 3215 27715 3235
rect 27735 3215 27750 3235
rect 27700 3185 27750 3215
rect 27700 3165 27715 3185
rect 27735 3165 27750 3185
rect 27700 3135 27750 3165
rect 27700 3115 27715 3135
rect 27735 3115 27750 3135
rect 27700 3085 27750 3115
rect 27700 3065 27715 3085
rect 27735 3065 27750 3085
rect 27700 3050 27750 3065
rect 28150 3535 28200 3550
rect 28150 3515 28165 3535
rect 28185 3515 28200 3535
rect 28150 3485 28200 3515
rect 28150 3465 28165 3485
rect 28185 3465 28200 3485
rect 28150 3435 28200 3465
rect 28150 3415 28165 3435
rect 28185 3415 28200 3435
rect 28150 3385 28200 3415
rect 28150 3365 28165 3385
rect 28185 3365 28200 3385
rect 28150 3335 28200 3365
rect 28150 3315 28165 3335
rect 28185 3315 28200 3335
rect 28150 3285 28200 3315
rect 28150 3265 28165 3285
rect 28185 3265 28200 3285
rect 28150 3235 28200 3265
rect 28150 3215 28165 3235
rect 28185 3215 28200 3235
rect 28150 3185 28200 3215
rect 28150 3165 28165 3185
rect 28185 3165 28200 3185
rect 28150 3135 28200 3165
rect 28150 3115 28165 3135
rect 28185 3115 28200 3135
rect 28150 3085 28200 3115
rect 28150 3065 28165 3085
rect 28185 3065 28200 3085
rect 28150 3050 28200 3065
rect 28750 3535 28800 3550
rect 28750 3515 28765 3535
rect 28785 3515 28800 3535
rect 28750 3485 28800 3515
rect 28750 3465 28765 3485
rect 28785 3465 28800 3485
rect 28750 3435 28800 3465
rect 28750 3415 28765 3435
rect 28785 3415 28800 3435
rect 28750 3385 28800 3415
rect 28750 3365 28765 3385
rect 28785 3365 28800 3385
rect 28750 3335 28800 3365
rect 28750 3315 28765 3335
rect 28785 3315 28800 3335
rect 28750 3285 28800 3315
rect 28750 3265 28765 3285
rect 28785 3265 28800 3285
rect 28750 3235 28800 3265
rect 28750 3215 28765 3235
rect 28785 3215 28800 3235
rect 28750 3185 28800 3215
rect 28750 3165 28765 3185
rect 28785 3165 28800 3185
rect 28750 3135 28800 3165
rect 28750 3115 28765 3135
rect 28785 3115 28800 3135
rect 28750 3085 28800 3115
rect 28750 3065 28765 3085
rect 28785 3065 28800 3085
rect 28750 3050 28800 3065
rect 29350 3535 29400 3550
rect 29350 3515 29365 3535
rect 29385 3515 29400 3535
rect 29350 3485 29400 3515
rect 29350 3465 29365 3485
rect 29385 3465 29400 3485
rect 29350 3435 29400 3465
rect 29350 3415 29365 3435
rect 29385 3415 29400 3435
rect 29350 3385 29400 3415
rect 29350 3365 29365 3385
rect 29385 3365 29400 3385
rect 29350 3335 29400 3365
rect 29350 3315 29365 3335
rect 29385 3315 29400 3335
rect 29350 3285 29400 3315
rect 29350 3265 29365 3285
rect 29385 3265 29400 3285
rect 29350 3235 29400 3265
rect 29350 3215 29365 3235
rect 29385 3215 29400 3235
rect 29350 3185 29400 3215
rect 29350 3165 29365 3185
rect 29385 3165 29400 3185
rect 29350 3135 29400 3165
rect 29350 3115 29365 3135
rect 29385 3115 29400 3135
rect 29350 3085 29400 3115
rect 29350 3065 29365 3085
rect 29385 3065 29400 3085
rect 29350 3050 29400 3065
rect 29500 3535 29550 3550
rect 29500 3515 29515 3535
rect 29535 3515 29550 3535
rect 29500 3485 29550 3515
rect 29500 3465 29515 3485
rect 29535 3465 29550 3485
rect 29500 3435 29550 3465
rect 29500 3415 29515 3435
rect 29535 3415 29550 3435
rect 29500 3385 29550 3415
rect 29500 3365 29515 3385
rect 29535 3365 29550 3385
rect 29500 3335 29550 3365
rect 29500 3315 29515 3335
rect 29535 3315 29550 3335
rect 29500 3285 29550 3315
rect 29500 3265 29515 3285
rect 29535 3265 29550 3285
rect 29500 3235 29550 3265
rect 29500 3215 29515 3235
rect 29535 3215 29550 3235
rect 29500 3185 29550 3215
rect 29500 3165 29515 3185
rect 29535 3165 29550 3185
rect 29500 3135 29550 3165
rect 29500 3115 29515 3135
rect 29535 3115 29550 3135
rect 29500 3085 29550 3115
rect 29500 3065 29515 3085
rect 29535 3065 29550 3085
rect 29500 3050 29550 3065
rect 29650 3535 29700 3550
rect 29650 3515 29665 3535
rect 29685 3515 29700 3535
rect 29650 3485 29700 3515
rect 29650 3465 29665 3485
rect 29685 3465 29700 3485
rect 29650 3435 29700 3465
rect 29650 3415 29665 3435
rect 29685 3415 29700 3435
rect 29650 3385 29700 3415
rect 29650 3365 29665 3385
rect 29685 3365 29700 3385
rect 29650 3335 29700 3365
rect 29650 3315 29665 3335
rect 29685 3315 29700 3335
rect 29650 3285 29700 3315
rect 29650 3265 29665 3285
rect 29685 3265 29700 3285
rect 29650 3235 29700 3265
rect 29650 3215 29665 3235
rect 29685 3215 29700 3235
rect 29650 3185 29700 3215
rect 29650 3165 29665 3185
rect 29685 3165 29700 3185
rect 29650 3135 29700 3165
rect 29650 3115 29665 3135
rect 29685 3115 29700 3135
rect 29650 3085 29700 3115
rect 29650 3065 29665 3085
rect 29685 3065 29700 3085
rect 29650 3050 29700 3065
rect 29800 3535 29850 3550
rect 29800 3515 29815 3535
rect 29835 3515 29850 3535
rect 29800 3485 29850 3515
rect 29800 3465 29815 3485
rect 29835 3465 29850 3485
rect 29800 3435 29850 3465
rect 29800 3415 29815 3435
rect 29835 3415 29850 3435
rect 29800 3385 29850 3415
rect 29800 3365 29815 3385
rect 29835 3365 29850 3385
rect 29800 3335 29850 3365
rect 29800 3315 29815 3335
rect 29835 3315 29850 3335
rect 29800 3285 29850 3315
rect 29800 3265 29815 3285
rect 29835 3265 29850 3285
rect 29800 3235 29850 3265
rect 29800 3215 29815 3235
rect 29835 3215 29850 3235
rect 29800 3185 29850 3215
rect 29800 3165 29815 3185
rect 29835 3165 29850 3185
rect 29800 3135 29850 3165
rect 29800 3115 29815 3135
rect 29835 3115 29850 3135
rect 29800 3085 29850 3115
rect 29800 3065 29815 3085
rect 29835 3065 29850 3085
rect 29800 3050 29850 3065
rect 29950 3535 30000 3550
rect 29950 3515 29965 3535
rect 29985 3515 30000 3535
rect 29950 3485 30000 3515
rect 29950 3465 29965 3485
rect 29985 3465 30000 3485
rect 29950 3435 30000 3465
rect 29950 3415 29965 3435
rect 29985 3415 30000 3435
rect 29950 3385 30000 3415
rect 29950 3365 29965 3385
rect 29985 3365 30000 3385
rect 29950 3335 30000 3365
rect 29950 3315 29965 3335
rect 29985 3315 30000 3335
rect 29950 3285 30000 3315
rect 29950 3265 29965 3285
rect 29985 3265 30000 3285
rect 29950 3235 30000 3265
rect 29950 3215 29965 3235
rect 29985 3215 30000 3235
rect 29950 3185 30000 3215
rect 29950 3165 29965 3185
rect 29985 3165 30000 3185
rect 29950 3135 30000 3165
rect 29950 3115 29965 3135
rect 29985 3115 30000 3135
rect 29950 3085 30000 3115
rect 29950 3065 29965 3085
rect 29985 3065 30000 3085
rect 29950 3050 30000 3065
rect 30100 3535 30150 3550
rect 30100 3515 30115 3535
rect 30135 3515 30150 3535
rect 30100 3485 30150 3515
rect 30100 3465 30115 3485
rect 30135 3465 30150 3485
rect 30100 3435 30150 3465
rect 30100 3415 30115 3435
rect 30135 3415 30150 3435
rect 30100 3385 30150 3415
rect 30100 3365 30115 3385
rect 30135 3365 30150 3385
rect 30100 3335 30150 3365
rect 30100 3315 30115 3335
rect 30135 3315 30150 3335
rect 30100 3285 30150 3315
rect 30100 3265 30115 3285
rect 30135 3265 30150 3285
rect 30100 3235 30150 3265
rect 30100 3215 30115 3235
rect 30135 3215 30150 3235
rect 30100 3185 30150 3215
rect 30100 3165 30115 3185
rect 30135 3165 30150 3185
rect 30100 3135 30150 3165
rect 30100 3115 30115 3135
rect 30135 3115 30150 3135
rect 30100 3085 30150 3115
rect 30100 3065 30115 3085
rect 30135 3065 30150 3085
rect 30100 3050 30150 3065
rect 30250 3535 30300 3550
rect 30250 3515 30265 3535
rect 30285 3515 30300 3535
rect 30250 3485 30300 3515
rect 30250 3465 30265 3485
rect 30285 3465 30300 3485
rect 30250 3435 30300 3465
rect 30250 3415 30265 3435
rect 30285 3415 30300 3435
rect 30250 3385 30300 3415
rect 30250 3365 30265 3385
rect 30285 3365 30300 3385
rect 30250 3335 30300 3365
rect 30250 3315 30265 3335
rect 30285 3315 30300 3335
rect 30250 3285 30300 3315
rect 30250 3265 30265 3285
rect 30285 3265 30300 3285
rect 30250 3235 30300 3265
rect 30250 3215 30265 3235
rect 30285 3215 30300 3235
rect 30250 3185 30300 3215
rect 30250 3165 30265 3185
rect 30285 3165 30300 3185
rect 30250 3135 30300 3165
rect 30250 3115 30265 3135
rect 30285 3115 30300 3135
rect 30250 3085 30300 3115
rect 30250 3065 30265 3085
rect 30285 3065 30300 3085
rect 30250 3050 30300 3065
rect 30400 3535 30450 3550
rect 30400 3515 30415 3535
rect 30435 3515 30450 3535
rect 30400 3485 30450 3515
rect 30400 3465 30415 3485
rect 30435 3465 30450 3485
rect 30400 3435 30450 3465
rect 30400 3415 30415 3435
rect 30435 3415 30450 3435
rect 30400 3385 30450 3415
rect 30400 3365 30415 3385
rect 30435 3365 30450 3385
rect 30400 3335 30450 3365
rect 30400 3315 30415 3335
rect 30435 3315 30450 3335
rect 30400 3285 30450 3315
rect 30400 3265 30415 3285
rect 30435 3265 30450 3285
rect 30400 3235 30450 3265
rect 30400 3215 30415 3235
rect 30435 3215 30450 3235
rect 30400 3185 30450 3215
rect 30400 3165 30415 3185
rect 30435 3165 30450 3185
rect 30400 3135 30450 3165
rect 30400 3115 30415 3135
rect 30435 3115 30450 3135
rect 30400 3085 30450 3115
rect 30400 3065 30415 3085
rect 30435 3065 30450 3085
rect 30400 3050 30450 3065
rect 30550 3535 30600 3550
rect 30550 3515 30565 3535
rect 30585 3515 30600 3535
rect 30550 3485 30600 3515
rect 30550 3465 30565 3485
rect 30585 3465 30600 3485
rect 30550 3435 30600 3465
rect 30550 3415 30565 3435
rect 30585 3415 30600 3435
rect 30550 3385 30600 3415
rect 30550 3365 30565 3385
rect 30585 3365 30600 3385
rect 30550 3335 30600 3365
rect 30550 3315 30565 3335
rect 30585 3315 30600 3335
rect 30550 3285 30600 3315
rect 30550 3265 30565 3285
rect 30585 3265 30600 3285
rect 30550 3235 30600 3265
rect 30550 3215 30565 3235
rect 30585 3215 30600 3235
rect 30550 3185 30600 3215
rect 30550 3165 30565 3185
rect 30585 3165 30600 3185
rect 30550 3135 30600 3165
rect 30550 3115 30565 3135
rect 30585 3115 30600 3135
rect 30550 3085 30600 3115
rect 30550 3065 30565 3085
rect 30585 3065 30600 3085
rect 30550 3050 30600 3065
rect 30700 3535 30750 3550
rect 30700 3515 30715 3535
rect 30735 3515 30750 3535
rect 30700 3485 30750 3515
rect 30700 3465 30715 3485
rect 30735 3465 30750 3485
rect 30700 3435 30750 3465
rect 30700 3415 30715 3435
rect 30735 3415 30750 3435
rect 30700 3385 30750 3415
rect 30700 3365 30715 3385
rect 30735 3365 30750 3385
rect 30700 3335 30750 3365
rect 30700 3315 30715 3335
rect 30735 3315 30750 3335
rect 30700 3285 30750 3315
rect 30700 3265 30715 3285
rect 30735 3265 30750 3285
rect 30700 3235 30750 3265
rect 30700 3215 30715 3235
rect 30735 3215 30750 3235
rect 30700 3185 30750 3215
rect 30700 3165 30715 3185
rect 30735 3165 30750 3185
rect 30700 3135 30750 3165
rect 30700 3115 30715 3135
rect 30735 3115 30750 3135
rect 30700 3085 30750 3115
rect 30700 3065 30715 3085
rect 30735 3065 30750 3085
rect 30700 3050 30750 3065
rect 30850 3535 30900 3550
rect 30850 3515 30865 3535
rect 30885 3515 30900 3535
rect 30850 3485 30900 3515
rect 30850 3465 30865 3485
rect 30885 3465 30900 3485
rect 30850 3435 30900 3465
rect 30850 3415 30865 3435
rect 30885 3415 30900 3435
rect 30850 3385 30900 3415
rect 30850 3365 30865 3385
rect 30885 3365 30900 3385
rect 30850 3335 30900 3365
rect 30850 3315 30865 3335
rect 30885 3315 30900 3335
rect 30850 3285 30900 3315
rect 30850 3265 30865 3285
rect 30885 3265 30900 3285
rect 30850 3235 30900 3265
rect 30850 3215 30865 3235
rect 30885 3215 30900 3235
rect 30850 3185 30900 3215
rect 30850 3165 30865 3185
rect 30885 3165 30900 3185
rect 30850 3135 30900 3165
rect 30850 3115 30865 3135
rect 30885 3115 30900 3135
rect 30850 3085 30900 3115
rect 30850 3065 30865 3085
rect 30885 3065 30900 3085
rect 30850 3050 30900 3065
rect 31000 3535 31050 3550
rect 31000 3515 31015 3535
rect 31035 3515 31050 3535
rect 31000 3485 31050 3515
rect 31000 3465 31015 3485
rect 31035 3465 31050 3485
rect 31000 3435 31050 3465
rect 31000 3415 31015 3435
rect 31035 3415 31050 3435
rect 31000 3385 31050 3415
rect 31000 3365 31015 3385
rect 31035 3365 31050 3385
rect 31000 3335 31050 3365
rect 31000 3315 31015 3335
rect 31035 3315 31050 3335
rect 31000 3285 31050 3315
rect 31000 3265 31015 3285
rect 31035 3265 31050 3285
rect 31000 3235 31050 3265
rect 31000 3215 31015 3235
rect 31035 3215 31050 3235
rect 31000 3185 31050 3215
rect 31000 3165 31015 3185
rect 31035 3165 31050 3185
rect 31000 3135 31050 3165
rect 31000 3115 31015 3135
rect 31035 3115 31050 3135
rect 31000 3085 31050 3115
rect 31000 3065 31015 3085
rect 31035 3065 31050 3085
rect 31000 3050 31050 3065
rect 31150 3535 31200 3550
rect 31150 3515 31165 3535
rect 31185 3515 31200 3535
rect 31150 3485 31200 3515
rect 31150 3465 31165 3485
rect 31185 3465 31200 3485
rect 31150 3435 31200 3465
rect 31150 3415 31165 3435
rect 31185 3415 31200 3435
rect 31150 3385 31200 3415
rect 31150 3365 31165 3385
rect 31185 3365 31200 3385
rect 31150 3335 31200 3365
rect 31150 3315 31165 3335
rect 31185 3315 31200 3335
rect 31150 3285 31200 3315
rect 31150 3265 31165 3285
rect 31185 3265 31200 3285
rect 31150 3235 31200 3265
rect 31150 3215 31165 3235
rect 31185 3215 31200 3235
rect 31150 3185 31200 3215
rect 31150 3165 31165 3185
rect 31185 3165 31200 3185
rect 31150 3135 31200 3165
rect 31150 3115 31165 3135
rect 31185 3115 31200 3135
rect 31150 3085 31200 3115
rect 31150 3065 31165 3085
rect 31185 3065 31200 3085
rect 31150 3050 31200 3065
rect 31300 3535 31350 3550
rect 31300 3515 31315 3535
rect 31335 3515 31350 3535
rect 31300 3485 31350 3515
rect 31300 3465 31315 3485
rect 31335 3465 31350 3485
rect 31300 3435 31350 3465
rect 31300 3415 31315 3435
rect 31335 3415 31350 3435
rect 31300 3385 31350 3415
rect 31300 3365 31315 3385
rect 31335 3365 31350 3385
rect 31300 3335 31350 3365
rect 31300 3315 31315 3335
rect 31335 3315 31350 3335
rect 31300 3285 31350 3315
rect 31300 3265 31315 3285
rect 31335 3265 31350 3285
rect 31300 3235 31350 3265
rect 31300 3215 31315 3235
rect 31335 3215 31350 3235
rect 31300 3185 31350 3215
rect 31300 3165 31315 3185
rect 31335 3165 31350 3185
rect 31300 3135 31350 3165
rect 31300 3115 31315 3135
rect 31335 3115 31350 3135
rect 31300 3085 31350 3115
rect 31300 3065 31315 3085
rect 31335 3065 31350 3085
rect 31300 3050 31350 3065
rect 31450 3535 31500 3550
rect 31450 3515 31465 3535
rect 31485 3515 31500 3535
rect 31450 3485 31500 3515
rect 31450 3465 31465 3485
rect 31485 3465 31500 3485
rect 31450 3435 31500 3465
rect 31450 3415 31465 3435
rect 31485 3415 31500 3435
rect 31450 3385 31500 3415
rect 31450 3365 31465 3385
rect 31485 3365 31500 3385
rect 31450 3335 31500 3365
rect 31450 3315 31465 3335
rect 31485 3315 31500 3335
rect 31450 3285 31500 3315
rect 31450 3265 31465 3285
rect 31485 3265 31500 3285
rect 31450 3235 31500 3265
rect 31450 3215 31465 3235
rect 31485 3215 31500 3235
rect 31450 3185 31500 3215
rect 31450 3165 31465 3185
rect 31485 3165 31500 3185
rect 31450 3135 31500 3165
rect 31450 3115 31465 3135
rect 31485 3115 31500 3135
rect 31450 3085 31500 3115
rect 31450 3065 31465 3085
rect 31485 3065 31500 3085
rect 31450 3050 31500 3065
rect 32050 3535 32100 3550
rect 32050 3515 32065 3535
rect 32085 3515 32100 3535
rect 32050 3485 32100 3515
rect 32050 3465 32065 3485
rect 32085 3465 32100 3485
rect 32050 3435 32100 3465
rect 32050 3415 32065 3435
rect 32085 3415 32100 3435
rect 32050 3385 32100 3415
rect 32050 3365 32065 3385
rect 32085 3365 32100 3385
rect 32050 3335 32100 3365
rect 32050 3315 32065 3335
rect 32085 3315 32100 3335
rect 32050 3285 32100 3315
rect 32050 3265 32065 3285
rect 32085 3265 32100 3285
rect 32050 3235 32100 3265
rect 32050 3215 32065 3235
rect 32085 3215 32100 3235
rect 32050 3185 32100 3215
rect 32050 3165 32065 3185
rect 32085 3165 32100 3185
rect 32050 3135 32100 3165
rect 32050 3115 32065 3135
rect 32085 3115 32100 3135
rect 32050 3085 32100 3115
rect 32050 3065 32065 3085
rect 32085 3065 32100 3085
rect 32050 3050 32100 3065
rect -650 2985 32100 3000
rect -650 2965 -635 2985
rect -615 2965 -585 2985
rect -565 2965 -535 2985
rect -515 2965 -485 2985
rect -465 2965 -435 2985
rect -415 2965 -385 2985
rect -365 2965 -335 2985
rect -315 2965 -285 2985
rect -265 2965 -235 2985
rect -215 2965 -185 2985
rect -165 2965 -135 2985
rect -115 2965 -85 2985
rect -65 2965 -35 2985
rect -15 2965 15 2985
rect 35 2965 65 2985
rect 85 2965 115 2985
rect 135 2965 165 2985
rect 185 2965 215 2985
rect 235 2965 265 2985
rect 285 2965 315 2985
rect 335 2965 365 2985
rect 385 2965 415 2985
rect 435 2965 465 2985
rect 485 2965 515 2985
rect 535 2965 565 2985
rect 585 2965 615 2985
rect 635 2965 665 2985
rect 685 2965 715 2985
rect 735 2965 765 2985
rect 785 2965 815 2985
rect 835 2965 865 2985
rect 885 2965 915 2985
rect 935 2965 965 2985
rect 985 2965 1015 2985
rect 1035 2965 1065 2985
rect 1085 2965 1115 2985
rect 1135 2965 1165 2985
rect 1185 2965 1215 2985
rect 1235 2965 1265 2985
rect 1285 2965 1315 2985
rect 1335 2965 1365 2985
rect 1385 2965 1415 2985
rect 1435 2965 1465 2985
rect 1485 2965 1515 2985
rect 1535 2965 1565 2985
rect 1585 2965 1615 2985
rect 1635 2965 1665 2985
rect 1685 2965 1715 2985
rect 1735 2965 1765 2985
rect 1785 2965 1815 2985
rect 1835 2965 1865 2985
rect 1885 2965 1915 2985
rect 1935 2965 1965 2985
rect 1985 2965 2015 2985
rect 2035 2965 2065 2985
rect 2085 2965 2115 2985
rect 2135 2965 2165 2985
rect 2185 2965 2215 2985
rect 2235 2965 2265 2985
rect 2285 2965 2315 2985
rect 2335 2965 2365 2985
rect 2385 2965 2415 2985
rect 2435 2965 2465 2985
rect 2485 2965 2515 2985
rect 2535 2965 2565 2985
rect 2585 2965 2615 2985
rect 2635 2965 2665 2985
rect 2685 2965 2715 2985
rect 2735 2965 2765 2985
rect 2785 2965 2815 2985
rect 2835 2965 2865 2985
rect 2885 2965 2915 2985
rect 2935 2965 2965 2985
rect 2985 2965 3015 2985
rect 3035 2965 3065 2985
rect 3085 2965 3115 2985
rect 3135 2965 3165 2985
rect 3185 2965 3215 2985
rect 3235 2965 3265 2985
rect 3285 2965 3315 2985
rect 3335 2965 3365 2985
rect 3385 2965 3415 2985
rect 3435 2965 3465 2985
rect 3485 2965 3515 2985
rect 3535 2965 3565 2985
rect 3585 2965 3615 2985
rect 3635 2965 3665 2985
rect 3685 2965 3715 2985
rect 3735 2965 3765 2985
rect 3785 2965 3815 2985
rect 3835 2965 3865 2985
rect 3885 2965 3915 2985
rect 3935 2965 3965 2985
rect 3985 2965 4015 2985
rect 4035 2965 4065 2985
rect 4085 2965 4115 2985
rect 4135 2965 4165 2985
rect 4185 2965 4215 2985
rect 4235 2965 4265 2985
rect 4285 2965 4315 2985
rect 4335 2965 4365 2985
rect 4385 2965 4415 2985
rect 4435 2965 4465 2985
rect 4485 2965 4515 2985
rect 4535 2965 4565 2985
rect 4585 2965 4615 2985
rect 4635 2965 4665 2985
rect 4685 2965 4715 2985
rect 4735 2965 4765 2985
rect 4785 2965 4815 2985
rect 4835 2965 4865 2985
rect 4885 2965 4915 2985
rect 4935 2965 4965 2985
rect 4985 2965 5015 2985
rect 5035 2965 5065 2985
rect 5085 2965 5115 2985
rect 5135 2965 5165 2985
rect 5185 2965 5215 2985
rect 5235 2965 5265 2985
rect 5285 2965 5315 2985
rect 5335 2965 5365 2985
rect 5385 2965 5415 2985
rect 5435 2965 5465 2985
rect 5485 2965 5515 2985
rect 5535 2965 5565 2985
rect 5585 2965 5615 2985
rect 5635 2965 5665 2985
rect 5685 2965 5715 2985
rect 5735 2965 5765 2985
rect 5785 2965 5815 2985
rect 5835 2965 5865 2985
rect 5885 2965 5915 2985
rect 5935 2965 5965 2985
rect 5985 2965 6015 2985
rect 6035 2965 6065 2985
rect 6085 2965 6115 2985
rect 6135 2965 6165 2985
rect 6185 2965 6215 2985
rect 6235 2965 6265 2985
rect 6285 2965 6315 2985
rect 6335 2965 6365 2985
rect 6385 2965 6415 2985
rect 6435 2965 6465 2985
rect 6485 2965 6515 2985
rect 6535 2965 6565 2985
rect 6585 2965 6615 2985
rect 6635 2965 6665 2985
rect 6685 2965 6715 2985
rect 6735 2965 6765 2985
rect 6785 2965 6815 2985
rect 6835 2965 6865 2985
rect 6885 2965 6915 2985
rect 6935 2965 6965 2985
rect 6985 2965 7015 2985
rect 7035 2965 7065 2985
rect 7085 2965 7115 2985
rect 7135 2965 7165 2985
rect 7185 2965 7215 2985
rect 7235 2965 7265 2985
rect 7285 2965 7315 2985
rect 7335 2965 7365 2985
rect 7385 2965 7415 2985
rect 7435 2965 7465 2985
rect 7485 2965 7515 2985
rect 7535 2965 7565 2985
rect 7585 2965 7615 2985
rect 7635 2965 7665 2985
rect 7685 2965 7715 2985
rect 7735 2965 7765 2985
rect 7785 2965 7815 2985
rect 7835 2965 7865 2985
rect 7885 2965 7915 2985
rect 7935 2965 7965 2985
rect 7985 2965 8015 2985
rect 8035 2965 8065 2985
rect 8085 2965 8115 2985
rect 8135 2965 8165 2985
rect 8185 2965 8215 2985
rect 8235 2965 8265 2985
rect 8285 2965 8315 2985
rect 8335 2965 8365 2985
rect 8385 2965 8415 2985
rect 8435 2965 8465 2985
rect 8485 2965 8515 2985
rect 8535 2965 8565 2985
rect 8585 2965 8615 2985
rect 8635 2965 8665 2985
rect 8685 2965 8715 2985
rect 8735 2965 8765 2985
rect 8785 2965 8815 2985
rect 8835 2965 8865 2985
rect 8885 2965 8915 2985
rect 8935 2965 8965 2985
rect 8985 2965 9015 2985
rect 9035 2965 9065 2985
rect 9085 2965 9115 2985
rect 9135 2965 9165 2985
rect 9185 2965 9215 2985
rect 9235 2965 9265 2985
rect 9285 2965 9315 2985
rect 9335 2965 9365 2985
rect 9385 2965 9415 2985
rect 9435 2965 9465 2985
rect 9485 2965 9515 2985
rect 9535 2965 9565 2985
rect 9585 2965 9615 2985
rect 9635 2965 9665 2985
rect 9685 2965 9715 2985
rect 9735 2965 9765 2985
rect 9785 2965 9815 2985
rect 9835 2965 9865 2985
rect 9885 2965 9915 2985
rect 9935 2965 9965 2985
rect 9985 2965 10015 2985
rect 10035 2965 10065 2985
rect 10085 2965 10115 2985
rect 10135 2965 10165 2985
rect 10185 2965 10215 2985
rect 10235 2965 10265 2985
rect 10285 2965 10315 2985
rect 10335 2965 10365 2985
rect 10385 2965 10415 2985
rect 10435 2965 10465 2985
rect 10485 2965 10515 2985
rect 10535 2965 10565 2985
rect 10585 2965 10615 2985
rect 10635 2965 10665 2985
rect 10685 2965 10715 2985
rect 10735 2965 10765 2985
rect 10785 2965 10815 2985
rect 10835 2965 10865 2985
rect 10885 2965 10915 2985
rect 10935 2965 10965 2985
rect 10985 2965 11015 2985
rect 11035 2965 11065 2985
rect 11085 2965 11115 2985
rect 11135 2965 11165 2985
rect 11185 2965 11215 2985
rect 11235 2965 11265 2985
rect 11285 2965 11315 2985
rect 11335 2965 11365 2985
rect 11385 2965 11415 2985
rect 11435 2965 11465 2985
rect 11485 2965 11515 2985
rect 11535 2965 11565 2985
rect 11585 2965 11615 2985
rect 11635 2965 11665 2985
rect 11685 2965 11715 2985
rect 11735 2965 11765 2985
rect 11785 2965 11815 2985
rect 11835 2965 11865 2985
rect 11885 2965 11915 2985
rect 11935 2965 11965 2985
rect 11985 2965 12015 2985
rect 12035 2965 12065 2985
rect 12085 2965 12115 2985
rect 12135 2965 12165 2985
rect 12185 2965 12215 2985
rect 12235 2965 12265 2985
rect 12285 2965 12315 2985
rect 12335 2965 12365 2985
rect 12385 2965 12415 2985
rect 12435 2965 12465 2985
rect 12485 2965 12515 2985
rect 12535 2965 12565 2985
rect 12585 2965 12615 2985
rect 12635 2965 12665 2985
rect 12685 2965 12715 2985
rect 12735 2965 12765 2985
rect 12785 2965 12815 2985
rect 12835 2965 12865 2985
rect 12885 2965 12915 2985
rect 12935 2965 12965 2985
rect 12985 2965 13015 2985
rect 13035 2965 13065 2985
rect 13085 2965 13115 2985
rect 13135 2965 13165 2985
rect 13185 2965 13215 2985
rect 13235 2965 13265 2985
rect 13285 2965 13315 2985
rect 13335 2965 13365 2985
rect 13385 2965 13415 2985
rect 13435 2965 13465 2985
rect 13485 2965 13515 2985
rect 13535 2965 13565 2985
rect 13585 2965 13615 2985
rect 13635 2965 13665 2985
rect 13685 2965 13715 2985
rect 13735 2965 13765 2985
rect 13785 2965 13815 2985
rect 13835 2965 13865 2985
rect 13885 2965 13915 2985
rect 13935 2965 13965 2985
rect 13985 2965 14015 2985
rect 14035 2965 14065 2985
rect 14085 2965 14115 2985
rect 14135 2965 14165 2985
rect 14185 2965 14215 2985
rect 14235 2965 14265 2985
rect 14285 2965 14315 2985
rect 14335 2965 14365 2985
rect 14385 2965 14415 2985
rect 14435 2965 14465 2985
rect 14485 2965 14515 2985
rect 14535 2965 14565 2985
rect 14585 2965 14615 2985
rect 14635 2965 14665 2985
rect 14685 2965 14715 2985
rect 14735 2965 14765 2985
rect 14785 2965 14815 2985
rect 14835 2965 14865 2985
rect 14885 2965 14915 2985
rect 14935 2965 14965 2985
rect 14985 2965 15015 2985
rect 15035 2965 15065 2985
rect 15085 2965 15115 2985
rect 15135 2965 15165 2985
rect 15185 2965 15215 2985
rect 15235 2965 15265 2985
rect 15285 2965 15315 2985
rect 15335 2965 15365 2985
rect 15385 2965 15415 2985
rect 15435 2965 15465 2985
rect 15485 2965 15515 2985
rect 15535 2965 15565 2985
rect 15585 2965 15615 2985
rect 15635 2965 15665 2985
rect 15685 2965 15715 2985
rect 15735 2965 15765 2985
rect 15785 2965 15815 2985
rect 15835 2965 15865 2985
rect 15885 2965 15915 2985
rect 15935 2965 15965 2985
rect 15985 2965 16015 2985
rect 16035 2965 16065 2985
rect 16085 2965 16115 2985
rect 16135 2965 16165 2985
rect 16185 2965 16215 2985
rect 16235 2965 16265 2985
rect 16285 2965 16315 2985
rect 16335 2965 16365 2985
rect 16385 2965 16415 2985
rect 16435 2965 16465 2985
rect 16485 2965 16515 2985
rect 16535 2965 16565 2985
rect 16585 2965 16615 2985
rect 16635 2965 16665 2985
rect 16685 2965 16715 2985
rect 16735 2965 16765 2985
rect 16785 2965 16815 2985
rect 16835 2965 16865 2985
rect 16885 2965 16915 2985
rect 16935 2965 16965 2985
rect 16985 2965 17015 2985
rect 17035 2965 17065 2985
rect 17085 2965 17115 2985
rect 17135 2965 17165 2985
rect 17185 2965 17215 2985
rect 17235 2965 17265 2985
rect 17285 2965 17315 2985
rect 17335 2965 17365 2985
rect 17385 2965 17415 2985
rect 17435 2965 17465 2985
rect 17485 2965 17515 2985
rect 17535 2965 17565 2985
rect 17585 2965 17615 2985
rect 17635 2965 17665 2985
rect 17685 2965 17715 2985
rect 17735 2965 17765 2985
rect 17785 2965 17815 2985
rect 17835 2965 17865 2985
rect 17885 2965 17915 2985
rect 17935 2965 17965 2985
rect 17985 2965 18015 2985
rect 18035 2965 18065 2985
rect 18085 2965 18115 2985
rect 18135 2965 18165 2985
rect 18185 2965 18215 2985
rect 18235 2965 18265 2985
rect 18285 2965 18315 2985
rect 18335 2965 18365 2985
rect 18385 2965 18415 2985
rect 18435 2965 18465 2985
rect 18485 2965 18515 2985
rect 18535 2965 18565 2985
rect 18585 2965 18615 2985
rect 18635 2965 18665 2985
rect 18685 2965 18715 2985
rect 18735 2965 18765 2985
rect 18785 2965 18815 2985
rect 18835 2965 18865 2985
rect 18885 2965 18915 2985
rect 18935 2965 18965 2985
rect 18985 2965 19015 2985
rect 19035 2965 19065 2985
rect 19085 2965 19115 2985
rect 19135 2965 19165 2985
rect 19185 2965 19215 2985
rect 19235 2965 19265 2985
rect 19285 2965 19315 2985
rect 19335 2965 19365 2985
rect 19385 2965 19415 2985
rect 19435 2965 19465 2985
rect 19485 2965 19515 2985
rect 19535 2965 19565 2985
rect 19585 2965 19615 2985
rect 19635 2965 19665 2985
rect 19685 2965 19715 2985
rect 19735 2965 19765 2985
rect 19785 2965 19815 2985
rect 19835 2965 19865 2985
rect 19885 2965 19915 2985
rect 19935 2965 19965 2985
rect 19985 2965 20015 2985
rect 20035 2965 20065 2985
rect 20085 2965 20115 2985
rect 20135 2965 20165 2985
rect 20185 2965 20215 2985
rect 20235 2965 20265 2985
rect 20285 2965 20315 2985
rect 20335 2965 20365 2985
rect 20385 2965 20415 2985
rect 20435 2965 20465 2985
rect 20485 2965 20515 2985
rect 20535 2965 20565 2985
rect 20585 2965 20615 2985
rect 20635 2965 20665 2985
rect 20685 2965 20715 2985
rect 20735 2965 20765 2985
rect 20785 2965 20815 2985
rect 20835 2965 20865 2985
rect 20885 2965 20915 2985
rect 20935 2965 20965 2985
rect 20985 2965 21015 2985
rect 21035 2965 21065 2985
rect 21085 2965 21115 2985
rect 21135 2965 21165 2985
rect 21185 2965 21215 2985
rect 21235 2965 21265 2985
rect 21285 2965 21315 2985
rect 21335 2965 21365 2985
rect 21385 2965 21415 2985
rect 21435 2965 21465 2985
rect 21485 2965 21515 2985
rect 21535 2965 21565 2985
rect 21585 2965 21615 2985
rect 21635 2965 21665 2985
rect 21685 2965 21715 2985
rect 21735 2965 21765 2985
rect 21785 2965 21815 2985
rect 21835 2965 21865 2985
rect 21885 2965 21915 2985
rect 21935 2965 21965 2985
rect 21985 2965 22015 2985
rect 22035 2965 22065 2985
rect 22085 2965 22115 2985
rect 22135 2965 22165 2985
rect 22185 2965 22215 2985
rect 22235 2965 22265 2985
rect 22285 2965 22315 2985
rect 22335 2965 22365 2985
rect 22385 2965 22415 2985
rect 22435 2965 22465 2985
rect 22485 2965 22515 2985
rect 22535 2965 22565 2985
rect 22585 2965 22615 2985
rect 22635 2965 22665 2985
rect 22685 2965 22715 2985
rect 22735 2965 22765 2985
rect 22785 2965 22815 2985
rect 22835 2965 22865 2985
rect 22885 2965 22915 2985
rect 22935 2965 22965 2985
rect 22985 2965 23015 2985
rect 23035 2965 23065 2985
rect 23085 2965 23115 2985
rect 23135 2965 23165 2985
rect 23185 2965 23215 2985
rect 23235 2965 23265 2985
rect 23285 2965 23315 2985
rect 23335 2965 23365 2985
rect 23385 2965 23415 2985
rect 23435 2965 23465 2985
rect 23485 2965 23515 2985
rect 23535 2965 23565 2985
rect 23585 2965 23615 2985
rect 23635 2965 23665 2985
rect 23685 2965 23715 2985
rect 23735 2965 23765 2985
rect 23785 2965 23815 2985
rect 23835 2965 23865 2985
rect 23885 2965 23915 2985
rect 23935 2965 23965 2985
rect 23985 2965 24015 2985
rect 24035 2965 24065 2985
rect 24085 2965 24115 2985
rect 24135 2965 24165 2985
rect 24185 2965 24215 2985
rect 24235 2965 24265 2985
rect 24285 2965 24315 2985
rect 24335 2965 24365 2985
rect 24385 2965 24415 2985
rect 24435 2965 24465 2985
rect 24485 2965 24515 2985
rect 24535 2965 24565 2985
rect 24585 2965 24615 2985
rect 24635 2965 24665 2985
rect 24685 2965 24715 2985
rect 24735 2965 24765 2985
rect 24785 2965 24815 2985
rect 24835 2965 24865 2985
rect 24885 2965 24915 2985
rect 24935 2965 24965 2985
rect 24985 2965 25015 2985
rect 25035 2965 25065 2985
rect 25085 2965 25115 2985
rect 25135 2965 25165 2985
rect 25185 2965 25215 2985
rect 25235 2965 25265 2985
rect 25285 2965 25315 2985
rect 25335 2965 25365 2985
rect 25385 2965 25415 2985
rect 25435 2965 25465 2985
rect 25485 2965 25515 2985
rect 25535 2965 25565 2985
rect 25585 2965 25615 2985
rect 25635 2965 25665 2985
rect 25685 2965 25715 2985
rect 25735 2965 25765 2985
rect 25785 2965 25815 2985
rect 25835 2965 25865 2985
rect 25885 2965 25915 2985
rect 25935 2965 25965 2985
rect 25985 2965 26015 2985
rect 26035 2965 26065 2985
rect 26085 2965 26115 2985
rect 26135 2965 26165 2985
rect 26185 2965 26215 2985
rect 26235 2965 26265 2985
rect 26285 2965 26315 2985
rect 26335 2965 26365 2985
rect 26385 2965 26415 2985
rect 26435 2965 26465 2985
rect 26485 2965 26515 2985
rect 26535 2965 26565 2985
rect 26585 2965 26615 2985
rect 26635 2965 26665 2985
rect 26685 2965 26715 2985
rect 26735 2965 26765 2985
rect 26785 2965 26815 2985
rect 26835 2965 26865 2985
rect 26885 2965 26915 2985
rect 26935 2965 26965 2985
rect 26985 2965 27015 2985
rect 27035 2965 27065 2985
rect 27085 2965 27115 2985
rect 27135 2965 27165 2985
rect 27185 2965 27215 2985
rect 27235 2965 27265 2985
rect 27285 2965 27315 2985
rect 27335 2965 27365 2985
rect 27385 2965 27415 2985
rect 27435 2965 27465 2985
rect 27485 2965 27515 2985
rect 27535 2965 27565 2985
rect 27585 2965 27615 2985
rect 27635 2965 27665 2985
rect 27685 2965 27715 2985
rect 27735 2965 27765 2985
rect 27785 2965 27815 2985
rect 27835 2965 27865 2985
rect 27885 2965 27915 2985
rect 27935 2965 27965 2985
rect 27985 2965 28015 2985
rect 28035 2965 28065 2985
rect 28085 2965 28115 2985
rect 28135 2965 28165 2985
rect 28185 2965 28215 2985
rect 28235 2965 28265 2985
rect 28285 2965 28315 2985
rect 28335 2965 28365 2985
rect 28385 2965 28415 2985
rect 28435 2965 28465 2985
rect 28485 2965 28515 2985
rect 28535 2965 28565 2985
rect 28585 2965 28615 2985
rect 28635 2965 28665 2985
rect 28685 2965 28715 2985
rect 28735 2965 28765 2985
rect 28785 2965 28815 2985
rect 28835 2965 28865 2985
rect 28885 2965 28915 2985
rect 28935 2965 28965 2985
rect 28985 2965 29015 2985
rect 29035 2965 29065 2985
rect 29085 2965 29115 2985
rect 29135 2965 29165 2985
rect 29185 2965 29215 2985
rect 29235 2965 29265 2985
rect 29285 2965 29315 2985
rect 29335 2965 29365 2985
rect 29385 2965 29415 2985
rect 29435 2965 29465 2985
rect 29485 2965 29515 2985
rect 29535 2965 29565 2985
rect 29585 2965 29615 2985
rect 29635 2965 29665 2985
rect 29685 2965 29715 2985
rect 29735 2965 29765 2985
rect 29785 2965 29815 2985
rect 29835 2965 29865 2985
rect 29885 2965 29915 2985
rect 29935 2965 29965 2985
rect 29985 2965 30015 2985
rect 30035 2965 30065 2985
rect 30085 2965 30115 2985
rect 30135 2965 30165 2985
rect 30185 2965 30215 2985
rect 30235 2965 30265 2985
rect 30285 2965 30315 2985
rect 30335 2965 30365 2985
rect 30385 2965 30415 2985
rect 30435 2965 30465 2985
rect 30485 2965 30515 2985
rect 30535 2965 30565 2985
rect 30585 2965 30615 2985
rect 30635 2965 30665 2985
rect 30685 2965 30715 2985
rect 30735 2965 30765 2985
rect 30785 2965 30815 2985
rect 30835 2965 30865 2985
rect 30885 2965 30915 2985
rect 30935 2965 30965 2985
rect 30985 2965 31015 2985
rect 31035 2965 31065 2985
rect 31085 2965 31115 2985
rect 31135 2965 31165 2985
rect 31185 2965 31215 2985
rect 31235 2965 31265 2985
rect 31285 2965 31315 2985
rect 31335 2965 31365 2985
rect 31385 2965 31415 2985
rect 31435 2965 31465 2985
rect 31485 2965 31515 2985
rect 31535 2965 31565 2985
rect 31585 2965 31615 2985
rect 31635 2965 31665 2985
rect 31685 2965 31715 2985
rect 31735 2965 31765 2985
rect 31785 2965 31815 2985
rect 31835 2965 31865 2985
rect 31885 2965 31915 2985
rect 31935 2965 31965 2985
rect 31985 2965 32015 2985
rect 32035 2965 32065 2985
rect 32085 2965 32100 2985
rect -650 2950 32100 2965
rect -900 2835 32100 2850
rect -900 2815 -885 2835
rect -865 2815 -835 2835
rect -815 2815 -785 2835
rect -765 2815 -735 2835
rect -715 2815 -685 2835
rect -665 2815 -635 2835
rect -615 2815 -585 2835
rect -565 2815 -535 2835
rect -515 2815 -485 2835
rect -465 2815 -435 2835
rect -415 2815 -385 2835
rect -365 2815 -335 2835
rect -315 2815 -285 2835
rect -265 2815 -235 2835
rect -215 2815 -185 2835
rect -165 2815 -135 2835
rect -115 2815 -85 2835
rect -65 2815 -35 2835
rect -15 2815 15 2835
rect 35 2815 65 2835
rect 85 2815 115 2835
rect 135 2815 165 2835
rect 185 2815 215 2835
rect 235 2815 265 2835
rect 285 2815 315 2835
rect 335 2815 365 2835
rect 385 2815 415 2835
rect 435 2815 465 2835
rect 485 2815 515 2835
rect 535 2815 565 2835
rect 585 2815 615 2835
rect 635 2815 665 2835
rect 685 2815 715 2835
rect 735 2815 765 2835
rect 785 2815 815 2835
rect 835 2815 865 2835
rect 885 2815 915 2835
rect 935 2815 965 2835
rect 985 2815 1015 2835
rect 1035 2815 1065 2835
rect 1085 2815 1115 2835
rect 1135 2815 1165 2835
rect 1185 2815 1215 2835
rect 1235 2815 1265 2835
rect 1285 2815 1315 2835
rect 1335 2815 1365 2835
rect 1385 2815 1415 2835
rect 1435 2815 1465 2835
rect 1485 2815 1515 2835
rect 1535 2815 1565 2835
rect 1585 2815 1615 2835
rect 1635 2815 1665 2835
rect 1685 2815 1715 2835
rect 1735 2815 1765 2835
rect 1785 2815 1815 2835
rect 1835 2815 1865 2835
rect 1885 2815 1915 2835
rect 1935 2815 1965 2835
rect 1985 2815 2015 2835
rect 2035 2815 2065 2835
rect 2085 2815 2115 2835
rect 2135 2815 2165 2835
rect 2185 2815 2215 2835
rect 2235 2815 2265 2835
rect 2285 2815 2315 2835
rect 2335 2815 2365 2835
rect 2385 2815 2415 2835
rect 2435 2815 2465 2835
rect 2485 2815 2515 2835
rect 2535 2815 2565 2835
rect 2585 2815 2615 2835
rect 2635 2815 2665 2835
rect 2685 2815 2715 2835
rect 2735 2815 2765 2835
rect 2785 2815 2815 2835
rect 2835 2815 2865 2835
rect 2885 2815 2915 2835
rect 2935 2815 2965 2835
rect 2985 2815 3015 2835
rect 3035 2815 3065 2835
rect 3085 2815 3115 2835
rect 3135 2815 3165 2835
rect 3185 2815 3215 2835
rect 3235 2815 3265 2835
rect 3285 2815 3315 2835
rect 3335 2815 3365 2835
rect 3385 2815 3415 2835
rect 3435 2815 3465 2835
rect 3485 2815 3515 2835
rect 3535 2815 3565 2835
rect 3585 2815 3615 2835
rect 3635 2815 3665 2835
rect 3685 2815 3715 2835
rect 3735 2815 3765 2835
rect 3785 2815 3815 2835
rect 3835 2815 3865 2835
rect 3885 2815 3915 2835
rect 3935 2815 3965 2835
rect 3985 2815 4015 2835
rect 4035 2815 4065 2835
rect 4085 2815 4115 2835
rect 4135 2815 4165 2835
rect 4185 2815 4215 2835
rect 4235 2815 4265 2835
rect 4285 2815 4315 2835
rect 4335 2815 4365 2835
rect 4385 2815 4415 2835
rect 4435 2815 4465 2835
rect 4485 2815 4515 2835
rect 4535 2815 4565 2835
rect 4585 2815 4615 2835
rect 4635 2815 4665 2835
rect 4685 2815 4715 2835
rect 4735 2815 4765 2835
rect 4785 2815 4815 2835
rect 4835 2815 4865 2835
rect 4885 2815 4915 2835
rect 4935 2815 4965 2835
rect 4985 2815 5015 2835
rect 5035 2815 5065 2835
rect 5085 2815 5115 2835
rect 5135 2815 5165 2835
rect 5185 2815 5215 2835
rect 5235 2815 5265 2835
rect 5285 2815 5315 2835
rect 5335 2815 5365 2835
rect 5385 2815 5415 2835
rect 5435 2815 5465 2835
rect 5485 2815 5515 2835
rect 5535 2815 5565 2835
rect 5585 2815 5615 2835
rect 5635 2815 5665 2835
rect 5685 2815 5715 2835
rect 5735 2815 5765 2835
rect 5785 2815 5815 2835
rect 5835 2815 5865 2835
rect 5885 2815 5915 2835
rect 5935 2815 5965 2835
rect 5985 2815 6015 2835
rect 6035 2815 6065 2835
rect 6085 2815 6115 2835
rect 6135 2815 6165 2835
rect 6185 2815 6215 2835
rect 6235 2815 6265 2835
rect 6285 2815 6315 2835
rect 6335 2815 6365 2835
rect 6385 2815 6415 2835
rect 6435 2815 6465 2835
rect 6485 2815 6515 2835
rect 6535 2815 6565 2835
rect 6585 2815 6615 2835
rect 6635 2815 6665 2835
rect 6685 2815 6715 2835
rect 6735 2815 6765 2835
rect 6785 2815 6815 2835
rect 6835 2815 6865 2835
rect 6885 2815 6915 2835
rect 6935 2815 6965 2835
rect 6985 2815 7015 2835
rect 7035 2815 7065 2835
rect 7085 2815 7115 2835
rect 7135 2815 7165 2835
rect 7185 2815 7215 2835
rect 7235 2815 7265 2835
rect 7285 2815 7315 2835
rect 7335 2815 7365 2835
rect 7385 2815 7415 2835
rect 7435 2815 7465 2835
rect 7485 2815 7515 2835
rect 7535 2815 7565 2835
rect 7585 2815 7615 2835
rect 7635 2815 7665 2835
rect 7685 2815 7715 2835
rect 7735 2815 7765 2835
rect 7785 2815 7815 2835
rect 7835 2815 7865 2835
rect 7885 2815 7915 2835
rect 7935 2815 7965 2835
rect 7985 2815 8015 2835
rect 8035 2815 8065 2835
rect 8085 2815 8115 2835
rect 8135 2815 8165 2835
rect 8185 2815 8215 2835
rect 8235 2815 8265 2835
rect 8285 2815 8315 2835
rect 8335 2815 8365 2835
rect 8385 2815 8415 2835
rect 8435 2815 8465 2835
rect 8485 2815 8515 2835
rect 8535 2815 8565 2835
rect 8585 2815 8615 2835
rect 8635 2815 8665 2835
rect 8685 2815 8715 2835
rect 8735 2815 8765 2835
rect 8785 2815 8815 2835
rect 8835 2815 8865 2835
rect 8885 2815 8915 2835
rect 8935 2815 8965 2835
rect 8985 2815 9015 2835
rect 9035 2815 9065 2835
rect 9085 2815 9115 2835
rect 9135 2815 9165 2835
rect 9185 2815 9215 2835
rect 9235 2815 9265 2835
rect 9285 2815 9315 2835
rect 9335 2815 9365 2835
rect 9385 2815 9415 2835
rect 9435 2815 9465 2835
rect 9485 2815 9515 2835
rect 9535 2815 9565 2835
rect 9585 2815 9615 2835
rect 9635 2815 9665 2835
rect 9685 2815 9715 2835
rect 9735 2815 9765 2835
rect 9785 2815 9815 2835
rect 9835 2815 9865 2835
rect 9885 2815 9915 2835
rect 9935 2815 9965 2835
rect 9985 2815 10015 2835
rect 10035 2815 10065 2835
rect 10085 2815 10115 2835
rect 10135 2815 10165 2835
rect 10185 2815 10215 2835
rect 10235 2815 10265 2835
rect 10285 2815 10315 2835
rect 10335 2815 10365 2835
rect 10385 2815 10415 2835
rect 10435 2815 10465 2835
rect 10485 2815 10515 2835
rect 10535 2815 10565 2835
rect 10585 2815 10615 2835
rect 10635 2815 10665 2835
rect 10685 2815 10715 2835
rect 10735 2815 10765 2835
rect 10785 2815 10815 2835
rect 10835 2815 10865 2835
rect 10885 2815 10915 2835
rect 10935 2815 10965 2835
rect 10985 2815 11015 2835
rect 11035 2815 11065 2835
rect 11085 2815 11115 2835
rect 11135 2815 11165 2835
rect 11185 2815 11215 2835
rect 11235 2815 11265 2835
rect 11285 2815 11315 2835
rect 11335 2815 11365 2835
rect 11385 2815 11415 2835
rect 11435 2815 11465 2835
rect 11485 2815 11515 2835
rect 11535 2815 11565 2835
rect 11585 2815 11615 2835
rect 11635 2815 11665 2835
rect 11685 2815 11715 2835
rect 11735 2815 11765 2835
rect 11785 2815 11815 2835
rect 11835 2815 11865 2835
rect 11885 2815 11915 2835
rect 11935 2815 11965 2835
rect 11985 2815 12015 2835
rect 12035 2815 12065 2835
rect 12085 2815 12115 2835
rect 12135 2815 12165 2835
rect 12185 2815 12215 2835
rect 12235 2815 12265 2835
rect 12285 2815 12315 2835
rect 12335 2815 12365 2835
rect 12385 2815 12415 2835
rect 12435 2815 12465 2835
rect 12485 2815 12515 2835
rect 12535 2815 12565 2835
rect 12585 2815 12615 2835
rect 12635 2815 12665 2835
rect 12685 2815 12715 2835
rect 12735 2815 12765 2835
rect 12785 2815 12815 2835
rect 12835 2815 12865 2835
rect 12885 2815 12915 2835
rect 12935 2815 12965 2835
rect 12985 2815 13015 2835
rect 13035 2815 13065 2835
rect 13085 2815 13115 2835
rect 13135 2815 13165 2835
rect 13185 2815 13215 2835
rect 13235 2815 13265 2835
rect 13285 2815 13315 2835
rect 13335 2815 13365 2835
rect 13385 2815 13415 2835
rect 13435 2815 13465 2835
rect 13485 2815 13515 2835
rect 13535 2815 13565 2835
rect 13585 2815 13615 2835
rect 13635 2815 13665 2835
rect 13685 2815 13715 2835
rect 13735 2815 13765 2835
rect 13785 2815 13815 2835
rect 13835 2815 13865 2835
rect 13885 2815 13915 2835
rect 13935 2815 13965 2835
rect 13985 2815 14015 2835
rect 14035 2815 14065 2835
rect 14085 2815 14115 2835
rect 14135 2815 14165 2835
rect 14185 2815 14215 2835
rect 14235 2815 14265 2835
rect 14285 2815 14315 2835
rect 14335 2815 14365 2835
rect 14385 2815 14415 2835
rect 14435 2815 14465 2835
rect 14485 2815 14515 2835
rect 14535 2815 14565 2835
rect 14585 2815 14615 2835
rect 14635 2815 14665 2835
rect 14685 2815 14715 2835
rect 14735 2815 14765 2835
rect 14785 2815 14815 2835
rect 14835 2815 14865 2835
rect 14885 2815 14915 2835
rect 14935 2815 14965 2835
rect 14985 2815 15015 2835
rect 15035 2815 15065 2835
rect 15085 2815 15115 2835
rect 15135 2815 15165 2835
rect 15185 2815 15215 2835
rect 15235 2815 15265 2835
rect 15285 2815 15315 2835
rect 15335 2815 15365 2835
rect 15385 2815 15415 2835
rect 15435 2815 15465 2835
rect 15485 2815 15515 2835
rect 15535 2815 15565 2835
rect 15585 2815 15615 2835
rect 15635 2815 15665 2835
rect 15685 2815 15715 2835
rect 15735 2815 15765 2835
rect 15785 2815 15815 2835
rect 15835 2815 15865 2835
rect 15885 2815 15915 2835
rect 15935 2815 15965 2835
rect 15985 2815 16015 2835
rect 16035 2815 16065 2835
rect 16085 2815 16115 2835
rect 16135 2815 16165 2835
rect 16185 2815 16215 2835
rect 16235 2815 16265 2835
rect 16285 2815 16315 2835
rect 16335 2815 16365 2835
rect 16385 2815 16415 2835
rect 16435 2815 16465 2835
rect 16485 2815 16515 2835
rect 16535 2815 16565 2835
rect 16585 2815 16615 2835
rect 16635 2815 16665 2835
rect 16685 2815 16715 2835
rect 16735 2815 16765 2835
rect 16785 2815 16815 2835
rect 16835 2815 16865 2835
rect 16885 2815 16915 2835
rect 16935 2815 16965 2835
rect 16985 2815 17015 2835
rect 17035 2815 17065 2835
rect 17085 2815 17115 2835
rect 17135 2815 17165 2835
rect 17185 2815 17215 2835
rect 17235 2815 17265 2835
rect 17285 2815 17315 2835
rect 17335 2815 17365 2835
rect 17385 2815 17415 2835
rect 17435 2815 17465 2835
rect 17485 2815 17515 2835
rect 17535 2815 17565 2835
rect 17585 2815 17615 2835
rect 17635 2815 17665 2835
rect 17685 2815 17715 2835
rect 17735 2815 17765 2835
rect 17785 2815 17815 2835
rect 17835 2815 17865 2835
rect 17885 2815 17915 2835
rect 17935 2815 17965 2835
rect 17985 2815 18015 2835
rect 18035 2815 18065 2835
rect 18085 2815 18115 2835
rect 18135 2815 18165 2835
rect 18185 2815 18215 2835
rect 18235 2815 18265 2835
rect 18285 2815 18315 2835
rect 18335 2815 18365 2835
rect 18385 2815 18415 2835
rect 18435 2815 18465 2835
rect 18485 2815 18515 2835
rect 18535 2815 18565 2835
rect 18585 2815 18615 2835
rect 18635 2815 18665 2835
rect 18685 2815 18715 2835
rect 18735 2815 18765 2835
rect 18785 2815 18815 2835
rect 18835 2815 18865 2835
rect 18885 2815 18915 2835
rect 18935 2815 18965 2835
rect 18985 2815 19015 2835
rect 19035 2815 19065 2835
rect 19085 2815 19115 2835
rect 19135 2815 19165 2835
rect 19185 2815 19215 2835
rect 19235 2815 19265 2835
rect 19285 2815 19315 2835
rect 19335 2815 19365 2835
rect 19385 2815 19415 2835
rect 19435 2815 19465 2835
rect 19485 2815 19515 2835
rect 19535 2815 19565 2835
rect 19585 2815 19615 2835
rect 19635 2815 19665 2835
rect 19685 2815 19715 2835
rect 19735 2815 19765 2835
rect 19785 2815 19815 2835
rect 19835 2815 19865 2835
rect 19885 2815 19915 2835
rect 19935 2815 19965 2835
rect 19985 2815 20015 2835
rect 20035 2815 20065 2835
rect 20085 2815 20115 2835
rect 20135 2815 20165 2835
rect 20185 2815 20215 2835
rect 20235 2815 20265 2835
rect 20285 2815 20315 2835
rect 20335 2815 20365 2835
rect 20385 2815 20415 2835
rect 20435 2815 20465 2835
rect 20485 2815 20515 2835
rect 20535 2815 20565 2835
rect 20585 2815 20615 2835
rect 20635 2815 20665 2835
rect 20685 2815 20715 2835
rect 20735 2815 20765 2835
rect 20785 2815 20815 2835
rect 20835 2815 20865 2835
rect 20885 2815 20915 2835
rect 20935 2815 20965 2835
rect 20985 2815 21015 2835
rect 21035 2815 21065 2835
rect 21085 2815 21115 2835
rect 21135 2815 21165 2835
rect 21185 2815 21215 2835
rect 21235 2815 21265 2835
rect 21285 2815 21315 2835
rect 21335 2815 21365 2835
rect 21385 2815 21415 2835
rect 21435 2815 21465 2835
rect 21485 2815 21515 2835
rect 21535 2815 21565 2835
rect 21585 2815 21615 2835
rect 21635 2815 21665 2835
rect 21685 2815 21715 2835
rect 21735 2815 21765 2835
rect 21785 2815 21815 2835
rect 21835 2815 21865 2835
rect 21885 2815 21915 2835
rect 21935 2815 21965 2835
rect 21985 2815 22015 2835
rect 22035 2815 22065 2835
rect 22085 2815 22115 2835
rect 22135 2815 22165 2835
rect 22185 2815 22215 2835
rect 22235 2815 22265 2835
rect 22285 2815 22315 2835
rect 22335 2815 22365 2835
rect 22385 2815 22415 2835
rect 22435 2815 22465 2835
rect 22485 2815 22515 2835
rect 22535 2815 22565 2835
rect 22585 2815 22615 2835
rect 22635 2815 22665 2835
rect 22685 2815 22715 2835
rect 22735 2815 22765 2835
rect 22785 2815 22815 2835
rect 22835 2815 22865 2835
rect 22885 2815 22915 2835
rect 22935 2815 22965 2835
rect 22985 2815 23015 2835
rect 23035 2815 23065 2835
rect 23085 2815 23115 2835
rect 23135 2815 23165 2835
rect 23185 2815 23215 2835
rect 23235 2815 23265 2835
rect 23285 2815 23315 2835
rect 23335 2815 23365 2835
rect 23385 2815 23415 2835
rect 23435 2815 23465 2835
rect 23485 2815 23515 2835
rect 23535 2815 23565 2835
rect 23585 2815 23615 2835
rect 23635 2815 23665 2835
rect 23685 2815 23715 2835
rect 23735 2815 23765 2835
rect 23785 2815 23815 2835
rect 23835 2815 23865 2835
rect 23885 2815 23915 2835
rect 23935 2815 23965 2835
rect 23985 2815 24015 2835
rect 24035 2815 24065 2835
rect 24085 2815 24115 2835
rect 24135 2815 24165 2835
rect 24185 2815 24215 2835
rect 24235 2815 24265 2835
rect 24285 2815 24315 2835
rect 24335 2815 24365 2835
rect 24385 2815 24415 2835
rect 24435 2815 24465 2835
rect 24485 2815 24515 2835
rect 24535 2815 24565 2835
rect 24585 2815 24615 2835
rect 24635 2815 24665 2835
rect 24685 2815 24715 2835
rect 24735 2815 24765 2835
rect 24785 2815 24815 2835
rect 24835 2815 24865 2835
rect 24885 2815 24915 2835
rect 24935 2815 24965 2835
rect 24985 2815 25015 2835
rect 25035 2815 25065 2835
rect 25085 2815 25115 2835
rect 25135 2815 25165 2835
rect 25185 2815 25215 2835
rect 25235 2815 25265 2835
rect 25285 2815 25315 2835
rect 25335 2815 25365 2835
rect 25385 2815 25415 2835
rect 25435 2815 25465 2835
rect 25485 2815 25515 2835
rect 25535 2815 25565 2835
rect 25585 2815 25615 2835
rect 25635 2815 25665 2835
rect 25685 2815 25715 2835
rect 25735 2815 25765 2835
rect 25785 2815 25815 2835
rect 25835 2815 25865 2835
rect 25885 2815 25915 2835
rect 25935 2815 25965 2835
rect 25985 2815 26015 2835
rect 26035 2815 26065 2835
rect 26085 2815 26115 2835
rect 26135 2815 26165 2835
rect 26185 2815 26215 2835
rect 26235 2815 26265 2835
rect 26285 2815 26315 2835
rect 26335 2815 26365 2835
rect 26385 2815 26415 2835
rect 26435 2815 26465 2835
rect 26485 2815 26515 2835
rect 26535 2815 26565 2835
rect 26585 2815 26615 2835
rect 26635 2815 26665 2835
rect 26685 2815 26715 2835
rect 26735 2815 26765 2835
rect 26785 2815 26815 2835
rect 26835 2815 26865 2835
rect 26885 2815 26915 2835
rect 26935 2815 26965 2835
rect 26985 2815 27015 2835
rect 27035 2815 27065 2835
rect 27085 2815 27115 2835
rect 27135 2815 27165 2835
rect 27185 2815 27215 2835
rect 27235 2815 27265 2835
rect 27285 2815 27315 2835
rect 27335 2815 27365 2835
rect 27385 2815 27415 2835
rect 27435 2815 27465 2835
rect 27485 2815 27515 2835
rect 27535 2815 27565 2835
rect 27585 2815 27615 2835
rect 27635 2815 27665 2835
rect 27685 2815 27715 2835
rect 27735 2815 27765 2835
rect 27785 2815 27815 2835
rect 27835 2815 27865 2835
rect 27885 2815 27915 2835
rect 27935 2815 27965 2835
rect 27985 2815 28015 2835
rect 28035 2815 28065 2835
rect 28085 2815 28115 2835
rect 28135 2815 28165 2835
rect 28185 2815 28215 2835
rect 28235 2815 28265 2835
rect 28285 2815 28315 2835
rect 28335 2815 28365 2835
rect 28385 2815 28415 2835
rect 28435 2815 28465 2835
rect 28485 2815 28515 2835
rect 28535 2815 28565 2835
rect 28585 2815 28615 2835
rect 28635 2815 28665 2835
rect 28685 2815 28715 2835
rect 28735 2815 28765 2835
rect 28785 2815 28815 2835
rect 28835 2815 28865 2835
rect 28885 2815 28915 2835
rect 28935 2815 28965 2835
rect 28985 2815 29015 2835
rect 29035 2815 29065 2835
rect 29085 2815 29115 2835
rect 29135 2815 29165 2835
rect 29185 2815 29215 2835
rect 29235 2815 29265 2835
rect 29285 2815 29315 2835
rect 29335 2815 29365 2835
rect 29385 2815 29415 2835
rect 29435 2815 29465 2835
rect 29485 2815 29515 2835
rect 29535 2815 29565 2835
rect 29585 2815 29615 2835
rect 29635 2815 29665 2835
rect 29685 2815 29715 2835
rect 29735 2815 29765 2835
rect 29785 2815 29815 2835
rect 29835 2815 29865 2835
rect 29885 2815 29915 2835
rect 29935 2815 29965 2835
rect 29985 2815 30015 2835
rect 30035 2815 30065 2835
rect 30085 2815 30115 2835
rect 30135 2815 30165 2835
rect 30185 2815 30215 2835
rect 30235 2815 30265 2835
rect 30285 2815 30315 2835
rect 30335 2815 30365 2835
rect 30385 2815 30415 2835
rect 30435 2815 30465 2835
rect 30485 2815 30515 2835
rect 30535 2815 30565 2835
rect 30585 2815 30615 2835
rect 30635 2815 30665 2835
rect 30685 2815 30715 2835
rect 30735 2815 30765 2835
rect 30785 2815 30815 2835
rect 30835 2815 30865 2835
rect 30885 2815 30915 2835
rect 30935 2815 30965 2835
rect 30985 2815 31015 2835
rect 31035 2815 31065 2835
rect 31085 2815 31115 2835
rect 31135 2815 31165 2835
rect 31185 2815 31215 2835
rect 31235 2815 31265 2835
rect 31285 2815 31315 2835
rect 31335 2815 31365 2835
rect 31385 2815 31415 2835
rect 31435 2815 31465 2835
rect 31485 2815 31515 2835
rect 31535 2815 31565 2835
rect 31585 2815 31615 2835
rect 31635 2815 31665 2835
rect 31685 2815 31715 2835
rect 31735 2815 31765 2835
rect 31785 2815 31815 2835
rect 31835 2815 31865 2835
rect 31885 2815 31915 2835
rect 31935 2815 31965 2835
rect 31985 2815 32015 2835
rect 32035 2815 32065 2835
rect 32085 2815 32100 2835
rect -900 2800 32100 2815
rect -900 2035 28800 2050
rect -900 2015 -885 2035
rect -865 2015 -835 2035
rect -815 2015 -785 2035
rect -765 2015 -735 2035
rect -715 2015 -685 2035
rect -665 2015 -635 2035
rect -615 2015 -585 2035
rect -565 2015 -535 2035
rect -515 2015 -485 2035
rect -465 2015 -435 2035
rect -415 2015 -385 2035
rect -365 2015 -335 2035
rect -315 2015 -285 2035
rect -265 2015 -235 2035
rect -215 2015 -185 2035
rect -165 2015 -135 2035
rect -115 2015 -85 2035
rect -65 2015 -35 2035
rect -15 2015 15 2035
rect 35 2015 65 2035
rect 85 2015 115 2035
rect 135 2015 165 2035
rect 185 2015 215 2035
rect 235 2015 265 2035
rect 285 2015 315 2035
rect 335 2015 365 2035
rect 385 2015 415 2035
rect 435 2015 465 2035
rect 485 2015 515 2035
rect 535 2015 565 2035
rect 585 2015 615 2035
rect 635 2015 665 2035
rect 685 2015 715 2035
rect 735 2015 765 2035
rect 785 2015 815 2035
rect 835 2015 865 2035
rect 885 2015 915 2035
rect 935 2015 965 2035
rect 985 2015 1015 2035
rect 1035 2015 1065 2035
rect 1085 2015 1115 2035
rect 1135 2015 1165 2035
rect 1185 2015 1215 2035
rect 1235 2015 1265 2035
rect 1285 2015 1315 2035
rect 1335 2015 1365 2035
rect 1385 2015 1415 2035
rect 1435 2015 1465 2035
rect 1485 2015 1515 2035
rect 1535 2015 1565 2035
rect 1585 2015 1615 2035
rect 1635 2015 1665 2035
rect 1685 2015 1715 2035
rect 1735 2015 1765 2035
rect 1785 2015 1815 2035
rect 1835 2015 1865 2035
rect 1885 2015 1915 2035
rect 1935 2015 1965 2035
rect 1985 2015 2015 2035
rect 2035 2015 2065 2035
rect 2085 2015 2115 2035
rect 2135 2015 2165 2035
rect 2185 2015 2215 2035
rect 2235 2015 2265 2035
rect 2285 2015 2315 2035
rect 2335 2015 2365 2035
rect 2385 2015 2415 2035
rect 2435 2015 2465 2035
rect 2485 2015 2515 2035
rect 2535 2015 2565 2035
rect 2585 2015 2615 2035
rect 2635 2015 2665 2035
rect 2685 2015 2715 2035
rect 2735 2015 2765 2035
rect 2785 2015 2815 2035
rect 2835 2015 2865 2035
rect 2885 2015 2915 2035
rect 2935 2015 2965 2035
rect 2985 2015 3015 2035
rect 3035 2015 3065 2035
rect 3085 2015 3115 2035
rect 3135 2015 3165 2035
rect 3185 2015 3215 2035
rect 3235 2015 3265 2035
rect 3285 2015 3315 2035
rect 3335 2015 3365 2035
rect 3385 2015 3415 2035
rect 3435 2015 3465 2035
rect 3485 2015 3515 2035
rect 3535 2015 3565 2035
rect 3585 2015 3615 2035
rect 3635 2015 3665 2035
rect 3685 2015 3715 2035
rect 3735 2015 3765 2035
rect 3785 2015 3815 2035
rect 3835 2015 3865 2035
rect 3885 2015 3915 2035
rect 3935 2015 3965 2035
rect 3985 2015 4015 2035
rect 4035 2015 4065 2035
rect 4085 2015 4115 2035
rect 4135 2015 4165 2035
rect 4185 2015 4215 2035
rect 4235 2015 4265 2035
rect 4285 2015 4315 2035
rect 4335 2015 4365 2035
rect 4385 2015 4415 2035
rect 4435 2015 4465 2035
rect 4485 2015 4515 2035
rect 4535 2015 4565 2035
rect 4585 2015 4615 2035
rect 4635 2015 4665 2035
rect 4685 2015 4715 2035
rect 4735 2015 4765 2035
rect 4785 2015 4815 2035
rect 4835 2015 4865 2035
rect 4885 2015 4915 2035
rect 4935 2015 4965 2035
rect 4985 2015 5015 2035
rect 5035 2015 5065 2035
rect 5085 2015 5115 2035
rect 5135 2015 5165 2035
rect 5185 2015 5215 2035
rect 5235 2015 5265 2035
rect 5285 2015 5315 2035
rect 5335 2015 5365 2035
rect 5385 2015 5415 2035
rect 5435 2015 5465 2035
rect 5485 2015 5515 2035
rect 5535 2015 5565 2035
rect 5585 2015 5615 2035
rect 5635 2015 5665 2035
rect 5685 2015 5715 2035
rect 5735 2015 5765 2035
rect 5785 2015 5815 2035
rect 5835 2015 5865 2035
rect 5885 2015 5915 2035
rect 5935 2015 5965 2035
rect 5985 2015 6015 2035
rect 6035 2015 6065 2035
rect 6085 2015 6115 2035
rect 6135 2015 6165 2035
rect 6185 2015 6215 2035
rect 6235 2015 6265 2035
rect 6285 2015 6315 2035
rect 6335 2015 6365 2035
rect 6385 2015 6415 2035
rect 6435 2015 6465 2035
rect 6485 2015 6515 2035
rect 6535 2015 6565 2035
rect 6585 2015 6615 2035
rect 6635 2015 6665 2035
rect 6685 2015 6715 2035
rect 6735 2015 6765 2035
rect 6785 2015 6815 2035
rect 6835 2015 6865 2035
rect 6885 2015 6915 2035
rect 6935 2015 6965 2035
rect 6985 2015 7015 2035
rect 7035 2015 7065 2035
rect 7085 2015 7115 2035
rect 7135 2015 7165 2035
rect 7185 2015 7215 2035
rect 7235 2015 7265 2035
rect 7285 2015 7315 2035
rect 7335 2015 7365 2035
rect 7385 2015 7415 2035
rect 7435 2015 7465 2035
rect 7485 2015 7515 2035
rect 7535 2015 7565 2035
rect 7585 2015 7615 2035
rect 7635 2015 7665 2035
rect 7685 2015 7715 2035
rect 7735 2015 7765 2035
rect 7785 2015 7815 2035
rect 7835 2015 7865 2035
rect 7885 2015 7915 2035
rect 7935 2015 7965 2035
rect 7985 2015 8015 2035
rect 8035 2015 8065 2035
rect 8085 2015 8115 2035
rect 8135 2015 8165 2035
rect 8185 2015 8215 2035
rect 8235 2015 8265 2035
rect 8285 2015 8315 2035
rect 8335 2015 8365 2035
rect 8385 2015 8415 2035
rect 8435 2015 8465 2035
rect 8485 2015 8515 2035
rect 8535 2015 8565 2035
rect 8585 2015 8615 2035
rect 8635 2015 8665 2035
rect 8685 2015 8715 2035
rect 8735 2015 8765 2035
rect 8785 2015 8815 2035
rect 8835 2015 8865 2035
rect 8885 2015 8915 2035
rect 8935 2015 8965 2035
rect 8985 2015 9015 2035
rect 9035 2015 9065 2035
rect 9085 2015 9115 2035
rect 9135 2015 9165 2035
rect 9185 2015 9215 2035
rect 9235 2015 9265 2035
rect 9285 2015 9315 2035
rect 9335 2015 9365 2035
rect 9385 2015 9415 2035
rect 9435 2015 9465 2035
rect 9485 2015 9515 2035
rect 9535 2015 9565 2035
rect 9585 2015 9615 2035
rect 9635 2015 9665 2035
rect 9685 2015 9715 2035
rect 9735 2015 9765 2035
rect 9785 2015 9815 2035
rect 9835 2015 9865 2035
rect 9885 2015 9915 2035
rect 9935 2015 9965 2035
rect 9985 2015 10015 2035
rect 10035 2015 10065 2035
rect 10085 2015 10115 2035
rect 10135 2015 10165 2035
rect 10185 2015 10215 2035
rect 10235 2015 10265 2035
rect 10285 2015 10315 2035
rect 10335 2015 10365 2035
rect 10385 2015 10415 2035
rect 10435 2015 10465 2035
rect 10485 2015 10515 2035
rect 10535 2015 10565 2035
rect 10585 2015 10615 2035
rect 10635 2015 10665 2035
rect 10685 2015 10715 2035
rect 10735 2015 10765 2035
rect 10785 2015 10815 2035
rect 10835 2015 10865 2035
rect 10885 2015 10915 2035
rect 10935 2015 10965 2035
rect 10985 2015 11015 2035
rect 11035 2015 11065 2035
rect 11085 2015 11115 2035
rect 11135 2015 11165 2035
rect 11185 2015 11215 2035
rect 11235 2015 11265 2035
rect 11285 2015 11315 2035
rect 11335 2015 11365 2035
rect 11385 2015 11415 2035
rect 11435 2015 11465 2035
rect 11485 2015 11515 2035
rect 11535 2015 11565 2035
rect 11585 2015 11615 2035
rect 11635 2015 11665 2035
rect 11685 2015 11715 2035
rect 11735 2015 11765 2035
rect 11785 2015 11815 2035
rect 11835 2015 11865 2035
rect 11885 2015 11915 2035
rect 11935 2015 11965 2035
rect 11985 2015 12015 2035
rect 12035 2015 12065 2035
rect 12085 2015 12115 2035
rect 12135 2015 12165 2035
rect 12185 2015 12215 2035
rect 12235 2015 12265 2035
rect 12285 2015 12315 2035
rect 12335 2015 12365 2035
rect 12385 2015 12415 2035
rect 12435 2015 12465 2035
rect 12485 2015 12515 2035
rect 12535 2015 12565 2035
rect 12585 2015 12615 2035
rect 12635 2015 12665 2035
rect 12685 2015 12715 2035
rect 12735 2015 12765 2035
rect 12785 2015 12815 2035
rect 12835 2015 12865 2035
rect 12885 2015 12915 2035
rect 12935 2015 12965 2035
rect 12985 2015 13015 2035
rect 13035 2015 13065 2035
rect 13085 2015 13115 2035
rect 13135 2015 13165 2035
rect 13185 2015 13215 2035
rect 13235 2015 13265 2035
rect 13285 2015 13315 2035
rect 13335 2015 13365 2035
rect 13385 2015 13415 2035
rect 13435 2015 13465 2035
rect 13485 2015 13515 2035
rect 13535 2015 13565 2035
rect 13585 2015 13615 2035
rect 13635 2015 13665 2035
rect 13685 2015 13715 2035
rect 13735 2015 13765 2035
rect 13785 2015 13815 2035
rect 13835 2015 13865 2035
rect 13885 2015 13915 2035
rect 13935 2015 13965 2035
rect 13985 2015 14015 2035
rect 14035 2015 14065 2035
rect 14085 2015 14115 2035
rect 14135 2015 14165 2035
rect 14185 2015 14215 2035
rect 14235 2015 14265 2035
rect 14285 2015 14315 2035
rect 14335 2015 14365 2035
rect 14385 2015 14415 2035
rect 14435 2015 14465 2035
rect 14485 2015 14515 2035
rect 14535 2015 14565 2035
rect 14585 2015 14615 2035
rect 14635 2015 14665 2035
rect 14685 2015 14715 2035
rect 14735 2015 14765 2035
rect 14785 2015 14815 2035
rect 14835 2015 14865 2035
rect 14885 2015 14915 2035
rect 14935 2015 14965 2035
rect 14985 2015 15015 2035
rect 15035 2015 15065 2035
rect 15085 2015 15115 2035
rect 15135 2015 15165 2035
rect 15185 2015 15215 2035
rect 15235 2015 15265 2035
rect 15285 2015 15315 2035
rect 15335 2015 15365 2035
rect 15385 2015 15415 2035
rect 15435 2015 15465 2035
rect 15485 2015 15515 2035
rect 15535 2015 15565 2035
rect 15585 2015 15615 2035
rect 15635 2015 15665 2035
rect 15685 2015 15715 2035
rect 15735 2015 15765 2035
rect 15785 2015 15815 2035
rect 15835 2015 15865 2035
rect 15885 2015 15915 2035
rect 15935 2015 15965 2035
rect 15985 2015 16015 2035
rect 16035 2015 16065 2035
rect 16085 2015 16115 2035
rect 16135 2015 16165 2035
rect 16185 2015 16215 2035
rect 16235 2015 16265 2035
rect 16285 2015 16315 2035
rect 16335 2015 16365 2035
rect 16385 2015 16415 2035
rect 16435 2015 16465 2035
rect 16485 2015 16515 2035
rect 16535 2015 16565 2035
rect 16585 2015 16615 2035
rect 16635 2015 16665 2035
rect 16685 2015 16715 2035
rect 16735 2015 16765 2035
rect 16785 2015 16815 2035
rect 16835 2015 16865 2035
rect 16885 2015 16915 2035
rect 16935 2015 16965 2035
rect 16985 2015 17015 2035
rect 17035 2015 17065 2035
rect 17085 2015 17115 2035
rect 17135 2015 17165 2035
rect 17185 2015 17215 2035
rect 17235 2015 17265 2035
rect 17285 2015 17315 2035
rect 17335 2015 17365 2035
rect 17385 2015 17415 2035
rect 17435 2015 17465 2035
rect 17485 2015 17515 2035
rect 17535 2015 17565 2035
rect 17585 2015 17615 2035
rect 17635 2015 17665 2035
rect 17685 2015 17715 2035
rect 17735 2015 17765 2035
rect 17785 2015 17815 2035
rect 17835 2015 17865 2035
rect 17885 2015 17915 2035
rect 17935 2015 17965 2035
rect 17985 2015 18015 2035
rect 18035 2015 18065 2035
rect 18085 2015 18115 2035
rect 18135 2015 18165 2035
rect 18185 2015 18215 2035
rect 18235 2015 18265 2035
rect 18285 2015 18315 2035
rect 18335 2015 18365 2035
rect 18385 2015 18415 2035
rect 18435 2015 18465 2035
rect 18485 2015 18515 2035
rect 18535 2015 18565 2035
rect 18585 2015 18615 2035
rect 18635 2015 18665 2035
rect 18685 2015 18715 2035
rect 18735 2015 18765 2035
rect 18785 2015 18815 2035
rect 18835 2015 18865 2035
rect 18885 2015 18915 2035
rect 18935 2015 18965 2035
rect 18985 2015 19015 2035
rect 19035 2015 19065 2035
rect 19085 2015 19115 2035
rect 19135 2015 19165 2035
rect 19185 2015 19215 2035
rect 19235 2015 19265 2035
rect 19285 2015 19315 2035
rect 19335 2015 19365 2035
rect 19385 2015 19415 2035
rect 19435 2015 19465 2035
rect 19485 2015 19515 2035
rect 19535 2015 19565 2035
rect 19585 2015 19615 2035
rect 19635 2015 19665 2035
rect 19685 2015 19715 2035
rect 19735 2015 19765 2035
rect 19785 2015 19815 2035
rect 19835 2015 19865 2035
rect 19885 2015 19915 2035
rect 19935 2015 19965 2035
rect 19985 2015 20015 2035
rect 20035 2015 20065 2035
rect 20085 2015 20115 2035
rect 20135 2015 20165 2035
rect 20185 2015 20215 2035
rect 20235 2015 20265 2035
rect 20285 2015 20315 2035
rect 20335 2015 20365 2035
rect 20385 2015 20415 2035
rect 20435 2015 20465 2035
rect 20485 2015 20515 2035
rect 20535 2015 20565 2035
rect 20585 2015 20615 2035
rect 20635 2015 20665 2035
rect 20685 2015 20715 2035
rect 20735 2015 20765 2035
rect 20785 2015 20815 2035
rect 20835 2015 20865 2035
rect 20885 2015 20915 2035
rect 20935 2015 20965 2035
rect 20985 2015 21015 2035
rect 21035 2015 21065 2035
rect 21085 2015 21115 2035
rect 21135 2015 21165 2035
rect 21185 2015 21215 2035
rect 21235 2015 21265 2035
rect 21285 2015 21315 2035
rect 21335 2015 21365 2035
rect 21385 2015 21415 2035
rect 21435 2015 21465 2035
rect 21485 2015 21515 2035
rect 21535 2015 21565 2035
rect 21585 2015 21615 2035
rect 21635 2015 21665 2035
rect 21685 2015 21715 2035
rect 21735 2015 21765 2035
rect 21785 2015 21815 2035
rect 21835 2015 21865 2035
rect 21885 2015 21915 2035
rect 21935 2015 21965 2035
rect 21985 2015 22015 2035
rect 22035 2015 22065 2035
rect 22085 2015 22115 2035
rect 22135 2015 22165 2035
rect 22185 2015 22215 2035
rect 22235 2015 22265 2035
rect 22285 2015 22315 2035
rect 22335 2015 22365 2035
rect 22385 2015 22415 2035
rect 22435 2015 22465 2035
rect 22485 2015 22515 2035
rect 22535 2015 22565 2035
rect 22585 2015 22615 2035
rect 22635 2015 22665 2035
rect 22685 2015 22715 2035
rect 22735 2015 22765 2035
rect 22785 2015 22815 2035
rect 22835 2015 22865 2035
rect 22885 2015 22915 2035
rect 22935 2015 22965 2035
rect 22985 2015 23015 2035
rect 23035 2015 23065 2035
rect 23085 2015 23115 2035
rect 23135 2015 23165 2035
rect 23185 2015 23215 2035
rect 23235 2015 23265 2035
rect 23285 2015 23315 2035
rect 23335 2015 23365 2035
rect 23385 2015 23415 2035
rect 23435 2015 23465 2035
rect 23485 2015 23515 2035
rect 23535 2015 23565 2035
rect 23585 2015 23615 2035
rect 23635 2015 23665 2035
rect 23685 2015 23715 2035
rect 23735 2015 23765 2035
rect 23785 2015 23815 2035
rect 23835 2015 23865 2035
rect 23885 2015 23915 2035
rect 23935 2015 23965 2035
rect 23985 2015 24015 2035
rect 24035 2015 24065 2035
rect 24085 2015 24115 2035
rect 24135 2015 24165 2035
rect 24185 2015 24215 2035
rect 24235 2015 24265 2035
rect 24285 2015 24315 2035
rect 24335 2015 24365 2035
rect 24385 2015 24415 2035
rect 24435 2015 24465 2035
rect 24485 2015 24515 2035
rect 24535 2015 24565 2035
rect 24585 2015 24615 2035
rect 24635 2015 24665 2035
rect 24685 2015 24715 2035
rect 24735 2015 24765 2035
rect 24785 2015 24815 2035
rect 24835 2015 24865 2035
rect 24885 2015 24915 2035
rect 24935 2015 24965 2035
rect 24985 2015 25015 2035
rect 25035 2015 25065 2035
rect 25085 2015 25115 2035
rect 25135 2015 25165 2035
rect 25185 2015 25215 2035
rect 25235 2015 25265 2035
rect 25285 2015 25315 2035
rect 25335 2015 25365 2035
rect 25385 2015 25415 2035
rect 25435 2015 25465 2035
rect 25485 2015 25515 2035
rect 25535 2015 25565 2035
rect 25585 2015 25615 2035
rect 25635 2015 25665 2035
rect 25685 2015 25715 2035
rect 25735 2015 25765 2035
rect 25785 2015 25815 2035
rect 25835 2015 25865 2035
rect 25885 2015 25915 2035
rect 25935 2015 25965 2035
rect 25985 2015 26015 2035
rect 26035 2015 26065 2035
rect 26085 2015 26115 2035
rect 26135 2015 26165 2035
rect 26185 2015 26215 2035
rect 26235 2015 26265 2035
rect 26285 2015 26315 2035
rect 26335 2015 26365 2035
rect 26385 2015 26415 2035
rect 26435 2015 26465 2035
rect 26485 2015 26515 2035
rect 26535 2015 26565 2035
rect 26585 2015 26615 2035
rect 26635 2015 26665 2035
rect 26685 2015 26715 2035
rect 26735 2015 26765 2035
rect 26785 2015 26815 2035
rect 26835 2015 26865 2035
rect 26885 2015 26915 2035
rect 26935 2015 26965 2035
rect 26985 2015 27015 2035
rect 27035 2015 27065 2035
rect 27085 2015 27115 2035
rect 27135 2015 27165 2035
rect 27185 2015 27215 2035
rect 27235 2015 27265 2035
rect 27285 2015 27315 2035
rect 27335 2015 27365 2035
rect 27385 2015 27415 2035
rect 27435 2015 27465 2035
rect 27485 2015 27515 2035
rect 27535 2015 27565 2035
rect 27585 2015 27615 2035
rect 27635 2015 27665 2035
rect 27685 2015 27715 2035
rect 27735 2015 27765 2035
rect 27785 2015 27815 2035
rect 27835 2015 27865 2035
rect 27885 2015 27915 2035
rect 27935 2015 27965 2035
rect 27985 2015 28015 2035
rect 28035 2015 28065 2035
rect 28085 2015 28115 2035
rect 28135 2015 28165 2035
rect 28185 2015 28215 2035
rect 28235 2015 28265 2035
rect 28285 2015 28315 2035
rect 28335 2015 28365 2035
rect 28385 2015 28415 2035
rect 28435 2015 28465 2035
rect 28485 2015 28515 2035
rect 28535 2015 28565 2035
rect 28585 2015 28615 2035
rect 28635 2015 28665 2035
rect 28685 2015 28715 2035
rect 28735 2015 28765 2035
rect 28785 2015 28800 2035
rect -900 2000 28800 2015
rect -650 1835 28800 1850
rect -650 1815 -635 1835
rect -615 1815 -585 1835
rect -565 1815 -535 1835
rect -515 1815 -485 1835
rect -465 1815 -435 1835
rect -415 1815 -385 1835
rect -365 1815 -335 1835
rect -315 1815 -285 1835
rect -265 1815 -235 1835
rect -215 1815 -185 1835
rect -165 1815 -135 1835
rect -115 1815 -85 1835
rect -65 1815 -35 1835
rect -15 1815 15 1835
rect 35 1815 65 1835
rect 85 1815 115 1835
rect 135 1815 165 1835
rect 185 1815 215 1835
rect 235 1815 265 1835
rect 285 1815 315 1835
rect 335 1815 365 1835
rect 385 1815 415 1835
rect 435 1815 465 1835
rect 485 1815 515 1835
rect 535 1815 565 1835
rect 585 1815 615 1835
rect 635 1815 665 1835
rect 685 1815 715 1835
rect 735 1815 765 1835
rect 785 1815 815 1835
rect 835 1815 865 1835
rect 885 1815 915 1835
rect 935 1815 965 1835
rect 985 1815 1015 1835
rect 1035 1815 1065 1835
rect 1085 1815 1115 1835
rect 1135 1815 1165 1835
rect 1185 1815 1215 1835
rect 1235 1815 1265 1835
rect 1285 1815 1315 1835
rect 1335 1815 1365 1835
rect 1385 1815 1415 1835
rect 1435 1815 1465 1835
rect 1485 1815 1515 1835
rect 1535 1815 1565 1835
rect 1585 1815 1615 1835
rect 1635 1815 1665 1835
rect 1685 1815 1715 1835
rect 1735 1815 1765 1835
rect 1785 1815 1815 1835
rect 1835 1815 1865 1835
rect 1885 1815 1915 1835
rect 1935 1815 1965 1835
rect 1985 1815 2015 1835
rect 2035 1815 2065 1835
rect 2085 1815 2115 1835
rect 2135 1815 2165 1835
rect 2185 1815 2215 1835
rect 2235 1815 2265 1835
rect 2285 1815 2315 1835
rect 2335 1815 2365 1835
rect 2385 1815 2415 1835
rect 2435 1815 2465 1835
rect 2485 1815 2515 1835
rect 2535 1815 2565 1835
rect 2585 1815 2615 1835
rect 2635 1815 2665 1835
rect 2685 1815 2715 1835
rect 2735 1815 2765 1835
rect 2785 1815 2815 1835
rect 2835 1815 2865 1835
rect 2885 1815 2915 1835
rect 2935 1815 2965 1835
rect 2985 1815 3015 1835
rect 3035 1815 3065 1835
rect 3085 1815 3115 1835
rect 3135 1815 3165 1835
rect 3185 1815 3215 1835
rect 3235 1815 3265 1835
rect 3285 1815 3315 1835
rect 3335 1815 3365 1835
rect 3385 1815 3415 1835
rect 3435 1815 3465 1835
rect 3485 1815 3515 1835
rect 3535 1815 3565 1835
rect 3585 1815 3615 1835
rect 3635 1815 3665 1835
rect 3685 1815 3715 1835
rect 3735 1815 3765 1835
rect 3785 1815 3815 1835
rect 3835 1815 3865 1835
rect 3885 1815 3915 1835
rect 3935 1815 3965 1835
rect 3985 1815 4015 1835
rect 4035 1815 4065 1835
rect 4085 1815 4115 1835
rect 4135 1815 4165 1835
rect 4185 1815 4215 1835
rect 4235 1815 4265 1835
rect 4285 1815 4315 1835
rect 4335 1815 4365 1835
rect 4385 1815 4415 1835
rect 4435 1815 4465 1835
rect 4485 1815 4515 1835
rect 4535 1815 4565 1835
rect 4585 1815 4615 1835
rect 4635 1815 4665 1835
rect 4685 1815 4715 1835
rect 4735 1815 4765 1835
rect 4785 1815 4815 1835
rect 4835 1815 4865 1835
rect 4885 1815 4915 1835
rect 4935 1815 4965 1835
rect 4985 1815 5015 1835
rect 5035 1815 5065 1835
rect 5085 1815 5115 1835
rect 5135 1815 5165 1835
rect 5185 1815 5215 1835
rect 5235 1815 5265 1835
rect 5285 1815 5315 1835
rect 5335 1815 5365 1835
rect 5385 1815 5415 1835
rect 5435 1815 5465 1835
rect 5485 1815 5515 1835
rect 5535 1815 5565 1835
rect 5585 1815 5615 1835
rect 5635 1815 5665 1835
rect 5685 1815 5715 1835
rect 5735 1815 5765 1835
rect 5785 1815 5815 1835
rect 5835 1815 5865 1835
rect 5885 1815 5915 1835
rect 5935 1815 5965 1835
rect 5985 1815 6015 1835
rect 6035 1815 6065 1835
rect 6085 1815 6115 1835
rect 6135 1815 6165 1835
rect 6185 1815 6215 1835
rect 6235 1815 6265 1835
rect 6285 1815 6315 1835
rect 6335 1815 6365 1835
rect 6385 1815 6415 1835
rect 6435 1815 6465 1835
rect 6485 1815 6515 1835
rect 6535 1815 6565 1835
rect 6585 1815 6615 1835
rect 6635 1815 6665 1835
rect 6685 1815 6715 1835
rect 6735 1815 6765 1835
rect 6785 1815 6815 1835
rect 6835 1815 6865 1835
rect 6885 1815 6915 1835
rect 6935 1815 6965 1835
rect 6985 1815 7015 1835
rect 7035 1815 7065 1835
rect 7085 1815 7115 1835
rect 7135 1815 7165 1835
rect 7185 1815 7215 1835
rect 7235 1815 7265 1835
rect 7285 1815 7315 1835
rect 7335 1815 7365 1835
rect 7385 1815 7415 1835
rect 7435 1815 7465 1835
rect 7485 1815 7515 1835
rect 7535 1815 7565 1835
rect 7585 1815 7615 1835
rect 7635 1815 7665 1835
rect 7685 1815 7715 1835
rect 7735 1815 7765 1835
rect 7785 1815 7815 1835
rect 7835 1815 7865 1835
rect 7885 1815 7915 1835
rect 7935 1815 7965 1835
rect 7985 1815 8015 1835
rect 8035 1815 8065 1835
rect 8085 1815 8115 1835
rect 8135 1815 8165 1835
rect 8185 1815 8215 1835
rect 8235 1815 8265 1835
rect 8285 1815 8315 1835
rect 8335 1815 8365 1835
rect 8385 1815 8415 1835
rect 8435 1815 8465 1835
rect 8485 1815 8515 1835
rect 8535 1815 8565 1835
rect 8585 1815 8615 1835
rect 8635 1815 8665 1835
rect 8685 1815 8715 1835
rect 8735 1815 8765 1835
rect 8785 1815 8815 1835
rect 8835 1815 8865 1835
rect 8885 1815 8915 1835
rect 8935 1815 8965 1835
rect 8985 1815 9015 1835
rect 9035 1815 9065 1835
rect 9085 1815 9115 1835
rect 9135 1815 9165 1835
rect 9185 1815 9215 1835
rect 9235 1815 9265 1835
rect 9285 1815 9315 1835
rect 9335 1815 9365 1835
rect 9385 1815 9415 1835
rect 9435 1815 9465 1835
rect 9485 1815 9515 1835
rect 9535 1815 9565 1835
rect 9585 1815 9615 1835
rect 9635 1815 9665 1835
rect 9685 1815 9715 1835
rect 9735 1815 9765 1835
rect 9785 1815 9815 1835
rect 9835 1815 9865 1835
rect 9885 1815 9915 1835
rect 9935 1815 9965 1835
rect 9985 1815 10015 1835
rect 10035 1815 10065 1835
rect 10085 1815 10115 1835
rect 10135 1815 10165 1835
rect 10185 1815 10215 1835
rect 10235 1815 10265 1835
rect 10285 1815 10315 1835
rect 10335 1815 10365 1835
rect 10385 1815 10415 1835
rect 10435 1815 10465 1835
rect 10485 1815 10515 1835
rect 10535 1815 10565 1835
rect 10585 1815 10615 1835
rect 10635 1815 10665 1835
rect 10685 1815 10715 1835
rect 10735 1815 10765 1835
rect 10785 1815 10815 1835
rect 10835 1815 10865 1835
rect 10885 1815 10915 1835
rect 10935 1815 10965 1835
rect 10985 1815 11015 1835
rect 11035 1815 11065 1835
rect 11085 1815 11115 1835
rect 11135 1815 11165 1835
rect 11185 1815 11215 1835
rect 11235 1815 11265 1835
rect 11285 1815 11315 1835
rect 11335 1815 11365 1835
rect 11385 1815 11415 1835
rect 11435 1815 11465 1835
rect 11485 1815 11515 1835
rect 11535 1815 11565 1835
rect 11585 1815 11615 1835
rect 11635 1815 11665 1835
rect 11685 1815 11715 1835
rect 11735 1815 11765 1835
rect 11785 1815 11815 1835
rect 11835 1815 11865 1835
rect 11885 1815 11915 1835
rect 11935 1815 11965 1835
rect 11985 1815 12015 1835
rect 12035 1815 12065 1835
rect 12085 1815 12115 1835
rect 12135 1815 12165 1835
rect 12185 1815 12215 1835
rect 12235 1815 12265 1835
rect 12285 1815 12315 1835
rect 12335 1815 12365 1835
rect 12385 1815 12415 1835
rect 12435 1815 12465 1835
rect 12485 1815 12515 1835
rect 12535 1815 12565 1835
rect 12585 1815 12615 1835
rect 12635 1815 12665 1835
rect 12685 1815 12715 1835
rect 12735 1815 12765 1835
rect 12785 1815 12815 1835
rect 12835 1815 12865 1835
rect 12885 1815 12915 1835
rect 12935 1815 12965 1835
rect 12985 1815 13015 1835
rect 13035 1815 13065 1835
rect 13085 1815 13115 1835
rect 13135 1815 13165 1835
rect 13185 1815 13215 1835
rect 13235 1815 13265 1835
rect 13285 1815 13315 1835
rect 13335 1815 13365 1835
rect 13385 1815 13415 1835
rect 13435 1815 13465 1835
rect 13485 1815 13515 1835
rect 13535 1815 13565 1835
rect 13585 1815 13615 1835
rect 13635 1815 13665 1835
rect 13685 1815 13715 1835
rect 13735 1815 13765 1835
rect 13785 1815 13815 1835
rect 13835 1815 13865 1835
rect 13885 1815 13915 1835
rect 13935 1815 13965 1835
rect 13985 1815 14015 1835
rect 14035 1815 14065 1835
rect 14085 1815 14115 1835
rect 14135 1815 14165 1835
rect 14185 1815 14215 1835
rect 14235 1815 14265 1835
rect 14285 1815 14315 1835
rect 14335 1815 14365 1835
rect 14385 1815 14415 1835
rect 14435 1815 14465 1835
rect 14485 1815 14515 1835
rect 14535 1815 14565 1835
rect 14585 1815 14615 1835
rect 14635 1815 14665 1835
rect 14685 1815 14715 1835
rect 14735 1815 14765 1835
rect 14785 1815 14815 1835
rect 14835 1815 14865 1835
rect 14885 1815 14915 1835
rect 14935 1815 14965 1835
rect 14985 1815 15015 1835
rect 15035 1815 15065 1835
rect 15085 1815 15115 1835
rect 15135 1815 15165 1835
rect 15185 1815 15215 1835
rect 15235 1815 15265 1835
rect 15285 1815 15315 1835
rect 15335 1815 15365 1835
rect 15385 1815 15415 1835
rect 15435 1815 15465 1835
rect 15485 1815 15515 1835
rect 15535 1815 15565 1835
rect 15585 1815 15615 1835
rect 15635 1815 15665 1835
rect 15685 1815 15715 1835
rect 15735 1815 15765 1835
rect 15785 1815 15815 1835
rect 15835 1815 15865 1835
rect 15885 1815 15915 1835
rect 15935 1815 15965 1835
rect 15985 1815 16015 1835
rect 16035 1815 16065 1835
rect 16085 1815 16115 1835
rect 16135 1815 16165 1835
rect 16185 1815 16215 1835
rect 16235 1815 16265 1835
rect 16285 1815 16315 1835
rect 16335 1815 16365 1835
rect 16385 1815 16415 1835
rect 16435 1815 16465 1835
rect 16485 1815 16515 1835
rect 16535 1815 16565 1835
rect 16585 1815 16615 1835
rect 16635 1815 16665 1835
rect 16685 1815 16715 1835
rect 16735 1815 16765 1835
rect 16785 1815 16815 1835
rect 16835 1815 16865 1835
rect 16885 1815 16915 1835
rect 16935 1815 16965 1835
rect 16985 1815 17015 1835
rect 17035 1815 17065 1835
rect 17085 1815 17115 1835
rect 17135 1815 17165 1835
rect 17185 1815 17215 1835
rect 17235 1815 17265 1835
rect 17285 1815 17315 1835
rect 17335 1815 17365 1835
rect 17385 1815 17415 1835
rect 17435 1815 17465 1835
rect 17485 1815 17515 1835
rect 17535 1815 17565 1835
rect 17585 1815 17615 1835
rect 17635 1815 17665 1835
rect 17685 1815 17715 1835
rect 17735 1815 17765 1835
rect 17785 1815 17815 1835
rect 17835 1815 17865 1835
rect 17885 1815 17915 1835
rect 17935 1815 17965 1835
rect 17985 1815 18015 1835
rect 18035 1815 18065 1835
rect 18085 1815 18115 1835
rect 18135 1815 18165 1835
rect 18185 1815 18215 1835
rect 18235 1815 18265 1835
rect 18285 1815 18315 1835
rect 18335 1815 18365 1835
rect 18385 1815 18415 1835
rect 18435 1815 18465 1835
rect 18485 1815 18515 1835
rect 18535 1815 18565 1835
rect 18585 1815 18615 1835
rect 18635 1815 18665 1835
rect 18685 1815 18715 1835
rect 18735 1815 18765 1835
rect 18785 1815 18815 1835
rect 18835 1815 18865 1835
rect 18885 1815 18915 1835
rect 18935 1815 18965 1835
rect 18985 1815 19015 1835
rect 19035 1815 19065 1835
rect 19085 1815 19115 1835
rect 19135 1815 19165 1835
rect 19185 1815 19215 1835
rect 19235 1815 19265 1835
rect 19285 1815 19315 1835
rect 19335 1815 19365 1835
rect 19385 1815 19415 1835
rect 19435 1815 19465 1835
rect 19485 1815 19515 1835
rect 19535 1815 19565 1835
rect 19585 1815 19615 1835
rect 19635 1815 19665 1835
rect 19685 1815 19715 1835
rect 19735 1815 19765 1835
rect 19785 1815 19815 1835
rect 19835 1815 19865 1835
rect 19885 1815 19915 1835
rect 19935 1815 19965 1835
rect 19985 1815 20015 1835
rect 20035 1815 20065 1835
rect 20085 1815 20115 1835
rect 20135 1815 20165 1835
rect 20185 1815 20215 1835
rect 20235 1815 20265 1835
rect 20285 1815 20315 1835
rect 20335 1815 20365 1835
rect 20385 1815 20415 1835
rect 20435 1815 20465 1835
rect 20485 1815 20515 1835
rect 20535 1815 20565 1835
rect 20585 1815 20615 1835
rect 20635 1815 20665 1835
rect 20685 1815 20715 1835
rect 20735 1815 20765 1835
rect 20785 1815 20815 1835
rect 20835 1815 20865 1835
rect 20885 1815 20915 1835
rect 20935 1815 20965 1835
rect 20985 1815 21015 1835
rect 21035 1815 21065 1835
rect 21085 1815 21115 1835
rect 21135 1815 21165 1835
rect 21185 1815 21215 1835
rect 21235 1815 21265 1835
rect 21285 1815 21315 1835
rect 21335 1815 21365 1835
rect 21385 1815 21415 1835
rect 21435 1815 21465 1835
rect 21485 1815 21515 1835
rect 21535 1815 21565 1835
rect 21585 1815 21615 1835
rect 21635 1815 21665 1835
rect 21685 1815 21715 1835
rect 21735 1815 21765 1835
rect 21785 1815 21815 1835
rect 21835 1815 21865 1835
rect 21885 1815 21915 1835
rect 21935 1815 21965 1835
rect 21985 1815 22015 1835
rect 22035 1815 22065 1835
rect 22085 1815 22115 1835
rect 22135 1815 22165 1835
rect 22185 1815 22215 1835
rect 22235 1815 22265 1835
rect 22285 1815 22315 1835
rect 22335 1815 22365 1835
rect 22385 1815 22415 1835
rect 22435 1815 22465 1835
rect 22485 1815 22515 1835
rect 22535 1815 22565 1835
rect 22585 1815 22615 1835
rect 22635 1815 22665 1835
rect 22685 1815 22715 1835
rect 22735 1815 22765 1835
rect 22785 1815 22815 1835
rect 22835 1815 22865 1835
rect 22885 1815 22915 1835
rect 22935 1815 22965 1835
rect 22985 1815 23015 1835
rect 23035 1815 23065 1835
rect 23085 1815 23115 1835
rect 23135 1815 23165 1835
rect 23185 1815 23215 1835
rect 23235 1815 23265 1835
rect 23285 1815 23315 1835
rect 23335 1815 23365 1835
rect 23385 1815 23415 1835
rect 23435 1815 23465 1835
rect 23485 1815 23515 1835
rect 23535 1815 23565 1835
rect 23585 1815 23615 1835
rect 23635 1815 23665 1835
rect 23685 1815 23715 1835
rect 23735 1815 23765 1835
rect 23785 1815 23815 1835
rect 23835 1815 23865 1835
rect 23885 1815 23915 1835
rect 23935 1815 23965 1835
rect 23985 1815 24015 1835
rect 24035 1815 24065 1835
rect 24085 1815 24115 1835
rect 24135 1815 24165 1835
rect 24185 1815 24215 1835
rect 24235 1815 24265 1835
rect 24285 1815 24315 1835
rect 24335 1815 24365 1835
rect 24385 1815 24415 1835
rect 24435 1815 24465 1835
rect 24485 1815 24515 1835
rect 24535 1815 24565 1835
rect 24585 1815 24615 1835
rect 24635 1815 24665 1835
rect 24685 1815 24715 1835
rect 24735 1815 24765 1835
rect 24785 1815 24815 1835
rect 24835 1815 24865 1835
rect 24885 1815 24915 1835
rect 24935 1815 24965 1835
rect 24985 1815 25015 1835
rect 25035 1815 25065 1835
rect 25085 1815 25115 1835
rect 25135 1815 25165 1835
rect 25185 1815 25215 1835
rect 25235 1815 25265 1835
rect 25285 1815 25315 1835
rect 25335 1815 25365 1835
rect 25385 1815 25415 1835
rect 25435 1815 25465 1835
rect 25485 1815 25515 1835
rect 25535 1815 25565 1835
rect 25585 1815 25615 1835
rect 25635 1815 25665 1835
rect 25685 1815 25715 1835
rect 25735 1815 25765 1835
rect 25785 1815 25815 1835
rect 25835 1815 25865 1835
rect 25885 1815 25915 1835
rect 25935 1815 25965 1835
rect 25985 1815 26015 1835
rect 26035 1815 26065 1835
rect 26085 1815 26115 1835
rect 26135 1815 26165 1835
rect 26185 1815 26215 1835
rect 26235 1815 26265 1835
rect 26285 1815 26315 1835
rect 26335 1815 26365 1835
rect 26385 1815 26415 1835
rect 26435 1815 26465 1835
rect 26485 1815 26515 1835
rect 26535 1815 26565 1835
rect 26585 1815 26615 1835
rect 26635 1815 26665 1835
rect 26685 1815 26715 1835
rect 26735 1815 26765 1835
rect 26785 1815 26815 1835
rect 26835 1815 26865 1835
rect 26885 1815 26915 1835
rect 26935 1815 26965 1835
rect 26985 1815 27015 1835
rect 27035 1815 27065 1835
rect 27085 1815 27115 1835
rect 27135 1815 27165 1835
rect 27185 1815 27215 1835
rect 27235 1815 27265 1835
rect 27285 1815 27315 1835
rect 27335 1815 27365 1835
rect 27385 1815 27415 1835
rect 27435 1815 27465 1835
rect 27485 1815 27515 1835
rect 27535 1815 27565 1835
rect 27585 1815 27615 1835
rect 27635 1815 27665 1835
rect 27685 1815 27715 1835
rect 27735 1815 27765 1835
rect 27785 1815 27815 1835
rect 27835 1815 27865 1835
rect 27885 1815 27915 1835
rect 27935 1815 27965 1835
rect 27985 1815 28015 1835
rect 28035 1815 28065 1835
rect 28085 1815 28115 1835
rect 28135 1815 28165 1835
rect 28185 1815 28215 1835
rect 28235 1815 28265 1835
rect 28285 1815 28315 1835
rect 28335 1815 28365 1835
rect 28385 1815 28415 1835
rect 28435 1815 28465 1835
rect 28485 1815 28515 1835
rect 28535 1815 28565 1835
rect 28585 1815 28615 1835
rect 28635 1815 28665 1835
rect 28685 1815 28715 1835
rect 28735 1815 28765 1835
rect 28785 1815 28800 1835
rect -650 1800 28800 1815
rect -650 1685 28800 1700
rect -650 1665 -635 1685
rect -615 1665 -585 1685
rect -565 1665 -535 1685
rect -515 1665 -485 1685
rect -465 1665 -435 1685
rect -415 1665 -385 1685
rect -365 1665 -335 1685
rect -315 1665 -285 1685
rect -265 1665 -235 1685
rect -215 1665 -185 1685
rect -165 1665 -135 1685
rect -115 1665 -85 1685
rect -65 1665 -35 1685
rect -15 1665 15 1685
rect 35 1665 65 1685
rect 85 1665 115 1685
rect 135 1665 165 1685
rect 185 1665 215 1685
rect 235 1665 265 1685
rect 285 1665 315 1685
rect 335 1665 365 1685
rect 385 1665 415 1685
rect 435 1665 465 1685
rect 485 1665 515 1685
rect 535 1665 565 1685
rect 585 1665 615 1685
rect 635 1665 665 1685
rect 685 1665 715 1685
rect 735 1665 765 1685
rect 785 1665 815 1685
rect 835 1665 865 1685
rect 885 1665 915 1685
rect 935 1665 965 1685
rect 985 1665 1015 1685
rect 1035 1665 1065 1685
rect 1085 1665 1115 1685
rect 1135 1665 1165 1685
rect 1185 1665 1215 1685
rect 1235 1665 1265 1685
rect 1285 1665 1315 1685
rect 1335 1665 1365 1685
rect 1385 1665 1415 1685
rect 1435 1665 1465 1685
rect 1485 1665 1515 1685
rect 1535 1665 1565 1685
rect 1585 1665 1615 1685
rect 1635 1665 1665 1685
rect 1685 1665 1715 1685
rect 1735 1665 1765 1685
rect 1785 1665 1815 1685
rect 1835 1665 1865 1685
rect 1885 1665 1915 1685
rect 1935 1665 1965 1685
rect 1985 1665 2015 1685
rect 2035 1665 2065 1685
rect 2085 1665 2115 1685
rect 2135 1665 2165 1685
rect 2185 1665 2215 1685
rect 2235 1665 2265 1685
rect 2285 1665 2315 1685
rect 2335 1665 2365 1685
rect 2385 1665 2415 1685
rect 2435 1665 2465 1685
rect 2485 1665 2515 1685
rect 2535 1665 2565 1685
rect 2585 1665 2615 1685
rect 2635 1665 2665 1685
rect 2685 1665 2715 1685
rect 2735 1665 2765 1685
rect 2785 1665 2815 1685
rect 2835 1665 2865 1685
rect 2885 1665 2915 1685
rect 2935 1665 2965 1685
rect 2985 1665 3015 1685
rect 3035 1665 3065 1685
rect 3085 1665 3115 1685
rect 3135 1665 3165 1685
rect 3185 1665 3215 1685
rect 3235 1665 3265 1685
rect 3285 1665 3315 1685
rect 3335 1665 3365 1685
rect 3385 1665 3415 1685
rect 3435 1665 3465 1685
rect 3485 1665 3515 1685
rect 3535 1665 3565 1685
rect 3585 1665 3615 1685
rect 3635 1665 3665 1685
rect 3685 1665 3715 1685
rect 3735 1665 3765 1685
rect 3785 1665 3815 1685
rect 3835 1665 3865 1685
rect 3885 1665 3915 1685
rect 3935 1665 3965 1685
rect 3985 1665 4015 1685
rect 4035 1665 4065 1685
rect 4085 1665 4115 1685
rect 4135 1665 4165 1685
rect 4185 1665 4215 1685
rect 4235 1665 4265 1685
rect 4285 1665 4315 1685
rect 4335 1665 4365 1685
rect 4385 1665 4415 1685
rect 4435 1665 4465 1685
rect 4485 1665 4515 1685
rect 4535 1665 4565 1685
rect 4585 1665 4615 1685
rect 4635 1665 4665 1685
rect 4685 1665 4715 1685
rect 4735 1665 4765 1685
rect 4785 1665 4815 1685
rect 4835 1665 4865 1685
rect 4885 1665 4915 1685
rect 4935 1665 4965 1685
rect 4985 1665 5015 1685
rect 5035 1665 5065 1685
rect 5085 1665 5115 1685
rect 5135 1665 5165 1685
rect 5185 1665 5215 1685
rect 5235 1665 5265 1685
rect 5285 1665 5315 1685
rect 5335 1665 5365 1685
rect 5385 1665 5415 1685
rect 5435 1665 5465 1685
rect 5485 1665 5515 1685
rect 5535 1665 5565 1685
rect 5585 1665 5615 1685
rect 5635 1665 5665 1685
rect 5685 1665 5715 1685
rect 5735 1665 5765 1685
rect 5785 1665 5815 1685
rect 5835 1665 5865 1685
rect 5885 1665 5915 1685
rect 5935 1665 5965 1685
rect 5985 1665 6015 1685
rect 6035 1665 6065 1685
rect 6085 1665 6115 1685
rect 6135 1665 6165 1685
rect 6185 1665 6215 1685
rect 6235 1665 6265 1685
rect 6285 1665 6315 1685
rect 6335 1665 6365 1685
rect 6385 1665 6415 1685
rect 6435 1665 6465 1685
rect 6485 1665 6515 1685
rect 6535 1665 6565 1685
rect 6585 1665 6615 1685
rect 6635 1665 6665 1685
rect 6685 1665 6715 1685
rect 6735 1665 6765 1685
rect 6785 1665 6815 1685
rect 6835 1665 6865 1685
rect 6885 1665 6915 1685
rect 6935 1665 6965 1685
rect 6985 1665 7015 1685
rect 7035 1665 7065 1685
rect 7085 1665 7115 1685
rect 7135 1665 7165 1685
rect 7185 1665 7215 1685
rect 7235 1665 7265 1685
rect 7285 1665 7315 1685
rect 7335 1665 7365 1685
rect 7385 1665 7415 1685
rect 7435 1665 7465 1685
rect 7485 1665 7515 1685
rect 7535 1665 7565 1685
rect 7585 1665 7615 1685
rect 7635 1665 7665 1685
rect 7685 1665 7715 1685
rect 7735 1665 7765 1685
rect 7785 1665 7815 1685
rect 7835 1665 7865 1685
rect 7885 1665 7915 1685
rect 7935 1665 7965 1685
rect 7985 1665 8015 1685
rect 8035 1665 8065 1685
rect 8085 1665 8115 1685
rect 8135 1665 8165 1685
rect 8185 1665 8215 1685
rect 8235 1665 8265 1685
rect 8285 1665 8315 1685
rect 8335 1665 8365 1685
rect 8385 1665 8415 1685
rect 8435 1665 8465 1685
rect 8485 1665 8515 1685
rect 8535 1665 8565 1685
rect 8585 1665 8615 1685
rect 8635 1665 8665 1685
rect 8685 1665 8715 1685
rect 8735 1665 8765 1685
rect 8785 1665 8815 1685
rect 8835 1665 8865 1685
rect 8885 1665 8915 1685
rect 8935 1665 8965 1685
rect 8985 1665 9015 1685
rect 9035 1665 9065 1685
rect 9085 1665 9115 1685
rect 9135 1665 9165 1685
rect 9185 1665 9215 1685
rect 9235 1665 9265 1685
rect 9285 1665 9315 1685
rect 9335 1665 9365 1685
rect 9385 1665 9415 1685
rect 9435 1665 9465 1685
rect 9485 1665 9515 1685
rect 9535 1665 9565 1685
rect 9585 1665 9615 1685
rect 9635 1665 9665 1685
rect 9685 1665 9715 1685
rect 9735 1665 9765 1685
rect 9785 1665 9815 1685
rect 9835 1665 9865 1685
rect 9885 1665 9915 1685
rect 9935 1665 9965 1685
rect 9985 1665 10015 1685
rect 10035 1665 10065 1685
rect 10085 1665 10115 1685
rect 10135 1665 10165 1685
rect 10185 1665 10215 1685
rect 10235 1665 10265 1685
rect 10285 1665 10315 1685
rect 10335 1665 10365 1685
rect 10385 1665 10415 1685
rect 10435 1665 10465 1685
rect 10485 1665 10515 1685
rect 10535 1665 10565 1685
rect 10585 1665 10615 1685
rect 10635 1665 10665 1685
rect 10685 1665 10715 1685
rect 10735 1665 10765 1685
rect 10785 1665 10815 1685
rect 10835 1665 10865 1685
rect 10885 1665 10915 1685
rect 10935 1665 10965 1685
rect 10985 1665 11015 1685
rect 11035 1665 11065 1685
rect 11085 1665 11115 1685
rect 11135 1665 11165 1685
rect 11185 1665 11215 1685
rect 11235 1665 11265 1685
rect 11285 1665 11315 1685
rect 11335 1665 11365 1685
rect 11385 1665 11415 1685
rect 11435 1665 11465 1685
rect 11485 1665 11515 1685
rect 11535 1665 11565 1685
rect 11585 1665 11615 1685
rect 11635 1665 11665 1685
rect 11685 1665 11715 1685
rect 11735 1665 11765 1685
rect 11785 1665 11815 1685
rect 11835 1665 11865 1685
rect 11885 1665 11915 1685
rect 11935 1665 11965 1685
rect 11985 1665 12015 1685
rect 12035 1665 12065 1685
rect 12085 1665 12115 1685
rect 12135 1665 12165 1685
rect 12185 1665 12215 1685
rect 12235 1665 12265 1685
rect 12285 1665 12315 1685
rect 12335 1665 12365 1685
rect 12385 1665 12415 1685
rect 12435 1665 12465 1685
rect 12485 1665 12515 1685
rect 12535 1665 12565 1685
rect 12585 1665 12615 1685
rect 12635 1665 12665 1685
rect 12685 1665 12715 1685
rect 12735 1665 12765 1685
rect 12785 1665 12815 1685
rect 12835 1665 12865 1685
rect 12885 1665 12915 1685
rect 12935 1665 12965 1685
rect 12985 1665 13015 1685
rect 13035 1665 13065 1685
rect 13085 1665 13115 1685
rect 13135 1665 13165 1685
rect 13185 1665 13215 1685
rect 13235 1665 13265 1685
rect 13285 1665 13315 1685
rect 13335 1665 13365 1685
rect 13385 1665 13415 1685
rect 13435 1665 13465 1685
rect 13485 1665 13515 1685
rect 13535 1665 13565 1685
rect 13585 1665 13615 1685
rect 13635 1665 13665 1685
rect 13685 1665 13715 1685
rect 13735 1665 13765 1685
rect 13785 1665 13815 1685
rect 13835 1665 13865 1685
rect 13885 1665 13915 1685
rect 13935 1665 13965 1685
rect 13985 1665 14015 1685
rect 14035 1665 14065 1685
rect 14085 1665 14115 1685
rect 14135 1665 14165 1685
rect 14185 1665 14215 1685
rect 14235 1665 14265 1685
rect 14285 1665 14315 1685
rect 14335 1665 14365 1685
rect 14385 1665 14415 1685
rect 14435 1665 14465 1685
rect 14485 1665 14515 1685
rect 14535 1665 14565 1685
rect 14585 1665 14615 1685
rect 14635 1665 14665 1685
rect 14685 1665 14715 1685
rect 14735 1665 14765 1685
rect 14785 1665 14815 1685
rect 14835 1665 14865 1685
rect 14885 1665 14915 1685
rect 14935 1665 14965 1685
rect 14985 1665 15015 1685
rect 15035 1665 15065 1685
rect 15085 1665 15115 1685
rect 15135 1665 15165 1685
rect 15185 1665 15215 1685
rect 15235 1665 15265 1685
rect 15285 1665 15315 1685
rect 15335 1665 15365 1685
rect 15385 1665 15415 1685
rect 15435 1665 15465 1685
rect 15485 1665 15515 1685
rect 15535 1665 15565 1685
rect 15585 1665 15615 1685
rect 15635 1665 15665 1685
rect 15685 1665 15715 1685
rect 15735 1665 15765 1685
rect 15785 1665 15815 1685
rect 15835 1665 15865 1685
rect 15885 1665 15915 1685
rect 15935 1665 15965 1685
rect 15985 1665 16015 1685
rect 16035 1665 16065 1685
rect 16085 1665 16115 1685
rect 16135 1665 16165 1685
rect 16185 1665 16215 1685
rect 16235 1665 16265 1685
rect 16285 1665 16315 1685
rect 16335 1665 16365 1685
rect 16385 1665 16415 1685
rect 16435 1665 16465 1685
rect 16485 1665 16515 1685
rect 16535 1665 16565 1685
rect 16585 1665 16615 1685
rect 16635 1665 16665 1685
rect 16685 1665 16715 1685
rect 16735 1665 16765 1685
rect 16785 1665 16815 1685
rect 16835 1665 16865 1685
rect 16885 1665 16915 1685
rect 16935 1665 16965 1685
rect 16985 1665 17015 1685
rect 17035 1665 17065 1685
rect 17085 1665 17115 1685
rect 17135 1665 17165 1685
rect 17185 1665 17215 1685
rect 17235 1665 17265 1685
rect 17285 1665 17315 1685
rect 17335 1665 17365 1685
rect 17385 1665 17415 1685
rect 17435 1665 17465 1685
rect 17485 1665 17515 1685
rect 17535 1665 17565 1685
rect 17585 1665 17615 1685
rect 17635 1665 17665 1685
rect 17685 1665 17715 1685
rect 17735 1665 17765 1685
rect 17785 1665 17815 1685
rect 17835 1665 17865 1685
rect 17885 1665 17915 1685
rect 17935 1665 17965 1685
rect 17985 1665 18015 1685
rect 18035 1665 18065 1685
rect 18085 1665 18115 1685
rect 18135 1665 18165 1685
rect 18185 1665 18215 1685
rect 18235 1665 18265 1685
rect 18285 1665 18315 1685
rect 18335 1665 18365 1685
rect 18385 1665 18415 1685
rect 18435 1665 18465 1685
rect 18485 1665 18515 1685
rect 18535 1665 18565 1685
rect 18585 1665 18615 1685
rect 18635 1665 18665 1685
rect 18685 1665 18715 1685
rect 18735 1665 18765 1685
rect 18785 1665 18815 1685
rect 18835 1665 18865 1685
rect 18885 1665 18915 1685
rect 18935 1665 18965 1685
rect 18985 1665 19015 1685
rect 19035 1665 19065 1685
rect 19085 1665 19115 1685
rect 19135 1665 19165 1685
rect 19185 1665 19215 1685
rect 19235 1665 19265 1685
rect 19285 1665 19315 1685
rect 19335 1665 19365 1685
rect 19385 1665 19415 1685
rect 19435 1665 19465 1685
rect 19485 1665 19515 1685
rect 19535 1665 19565 1685
rect 19585 1665 19615 1685
rect 19635 1665 19665 1685
rect 19685 1665 19715 1685
rect 19735 1665 19765 1685
rect 19785 1665 19815 1685
rect 19835 1665 19865 1685
rect 19885 1665 19915 1685
rect 19935 1665 19965 1685
rect 19985 1665 20015 1685
rect 20035 1665 20065 1685
rect 20085 1665 20115 1685
rect 20135 1665 20165 1685
rect 20185 1665 20215 1685
rect 20235 1665 20265 1685
rect 20285 1665 20315 1685
rect 20335 1665 20365 1685
rect 20385 1665 20415 1685
rect 20435 1665 20465 1685
rect 20485 1665 20515 1685
rect 20535 1665 20565 1685
rect 20585 1665 20615 1685
rect 20635 1665 20665 1685
rect 20685 1665 20715 1685
rect 20735 1665 20765 1685
rect 20785 1665 20815 1685
rect 20835 1665 20865 1685
rect 20885 1665 20915 1685
rect 20935 1665 20965 1685
rect 20985 1665 21015 1685
rect 21035 1665 21065 1685
rect 21085 1665 21115 1685
rect 21135 1665 21165 1685
rect 21185 1665 21215 1685
rect 21235 1665 21265 1685
rect 21285 1665 21315 1685
rect 21335 1665 21365 1685
rect 21385 1665 21415 1685
rect 21435 1665 21465 1685
rect 21485 1665 21515 1685
rect 21535 1665 21565 1685
rect 21585 1665 21615 1685
rect 21635 1665 21665 1685
rect 21685 1665 21715 1685
rect 21735 1665 21765 1685
rect 21785 1665 21815 1685
rect 21835 1665 21865 1685
rect 21885 1665 21915 1685
rect 21935 1665 21965 1685
rect 21985 1665 22015 1685
rect 22035 1665 22065 1685
rect 22085 1665 22115 1685
rect 22135 1665 22165 1685
rect 22185 1665 22215 1685
rect 22235 1665 22265 1685
rect 22285 1665 22315 1685
rect 22335 1665 22365 1685
rect 22385 1665 22415 1685
rect 22435 1665 22465 1685
rect 22485 1665 22515 1685
rect 22535 1665 22565 1685
rect 22585 1665 22615 1685
rect 22635 1665 22665 1685
rect 22685 1665 22715 1685
rect 22735 1665 22765 1685
rect 22785 1665 22815 1685
rect 22835 1665 22865 1685
rect 22885 1665 22915 1685
rect 22935 1665 22965 1685
rect 22985 1665 23015 1685
rect 23035 1665 23065 1685
rect 23085 1665 23115 1685
rect 23135 1665 23165 1685
rect 23185 1665 23215 1685
rect 23235 1665 23265 1685
rect 23285 1665 23315 1685
rect 23335 1665 23365 1685
rect 23385 1665 23415 1685
rect 23435 1665 23465 1685
rect 23485 1665 23515 1685
rect 23535 1665 23565 1685
rect 23585 1665 23615 1685
rect 23635 1665 23665 1685
rect 23685 1665 23715 1685
rect 23735 1665 23765 1685
rect 23785 1665 23815 1685
rect 23835 1665 23865 1685
rect 23885 1665 23915 1685
rect 23935 1665 23965 1685
rect 23985 1665 24015 1685
rect 24035 1665 24065 1685
rect 24085 1665 24115 1685
rect 24135 1665 24165 1685
rect 24185 1665 24215 1685
rect 24235 1665 24265 1685
rect 24285 1665 24315 1685
rect 24335 1665 24365 1685
rect 24385 1665 24415 1685
rect 24435 1665 24465 1685
rect 24485 1665 24515 1685
rect 24535 1665 24565 1685
rect 24585 1665 24615 1685
rect 24635 1665 24665 1685
rect 24685 1665 24715 1685
rect 24735 1665 24765 1685
rect 24785 1665 24815 1685
rect 24835 1665 24865 1685
rect 24885 1665 24915 1685
rect 24935 1665 24965 1685
rect 24985 1665 25015 1685
rect 25035 1665 25065 1685
rect 25085 1665 25115 1685
rect 25135 1665 25165 1685
rect 25185 1665 25215 1685
rect 25235 1665 25265 1685
rect 25285 1665 25315 1685
rect 25335 1665 25365 1685
rect 25385 1665 25415 1685
rect 25435 1665 25465 1685
rect 25485 1665 25515 1685
rect 25535 1665 25565 1685
rect 25585 1665 25615 1685
rect 25635 1665 25665 1685
rect 25685 1665 25715 1685
rect 25735 1665 25765 1685
rect 25785 1665 25815 1685
rect 25835 1665 25865 1685
rect 25885 1665 25915 1685
rect 25935 1665 25965 1685
rect 25985 1665 26015 1685
rect 26035 1665 26065 1685
rect 26085 1665 26115 1685
rect 26135 1665 26165 1685
rect 26185 1665 26215 1685
rect 26235 1665 26265 1685
rect 26285 1665 26315 1685
rect 26335 1665 26365 1685
rect 26385 1665 26415 1685
rect 26435 1665 26465 1685
rect 26485 1665 26515 1685
rect 26535 1665 26565 1685
rect 26585 1665 26615 1685
rect 26635 1665 26665 1685
rect 26685 1665 26715 1685
rect 26735 1665 26765 1685
rect 26785 1665 26815 1685
rect 26835 1665 26865 1685
rect 26885 1665 26915 1685
rect 26935 1665 26965 1685
rect 26985 1665 27015 1685
rect 27035 1665 27065 1685
rect 27085 1665 27115 1685
rect 27135 1665 27165 1685
rect 27185 1665 27215 1685
rect 27235 1665 27265 1685
rect 27285 1665 27315 1685
rect 27335 1665 27365 1685
rect 27385 1665 27415 1685
rect 27435 1665 27465 1685
rect 27485 1665 27515 1685
rect 27535 1665 27565 1685
rect 27585 1665 27615 1685
rect 27635 1665 27665 1685
rect 27685 1665 27715 1685
rect 27735 1665 27765 1685
rect 27785 1665 27815 1685
rect 27835 1665 27865 1685
rect 27885 1665 27915 1685
rect 27935 1665 27965 1685
rect 27985 1665 28015 1685
rect 28035 1665 28065 1685
rect 28085 1665 28115 1685
rect 28135 1665 28165 1685
rect 28185 1665 28215 1685
rect 28235 1665 28265 1685
rect 28285 1665 28315 1685
rect 28335 1665 28365 1685
rect 28385 1665 28415 1685
rect 28435 1665 28465 1685
rect 28485 1665 28515 1685
rect 28535 1665 28565 1685
rect 28585 1665 28615 1685
rect 28635 1665 28665 1685
rect 28685 1665 28715 1685
rect 28735 1665 28765 1685
rect 28785 1665 28800 1685
rect -650 1650 28800 1665
rect -650 1585 -600 1600
rect -650 1565 -635 1585
rect -615 1565 -600 1585
rect -650 1535 -600 1565
rect -650 1515 -635 1535
rect -615 1515 -600 1535
rect -650 1485 -600 1515
rect -650 1465 -635 1485
rect -615 1465 -600 1485
rect -650 1435 -600 1465
rect -650 1415 -635 1435
rect -615 1415 -600 1435
rect -650 1385 -600 1415
rect -650 1365 -635 1385
rect -615 1365 -600 1385
rect -650 1335 -600 1365
rect -650 1315 -635 1335
rect -615 1315 -600 1335
rect -650 1285 -600 1315
rect -650 1265 -635 1285
rect -615 1265 -600 1285
rect -650 1235 -600 1265
rect -650 1215 -635 1235
rect -615 1215 -600 1235
rect -650 1185 -600 1215
rect -650 1165 -635 1185
rect -615 1165 -600 1185
rect -650 1135 -600 1165
rect -650 1115 -635 1135
rect -615 1115 -600 1135
rect -650 1085 -600 1115
rect -650 1065 -635 1085
rect -615 1065 -600 1085
rect -650 1035 -600 1065
rect -650 1015 -635 1035
rect -615 1015 -600 1035
rect -650 985 -600 1015
rect -650 965 -635 985
rect -615 965 -600 985
rect -650 935 -600 965
rect -650 915 -635 935
rect -615 915 -600 935
rect -650 900 -600 915
rect -500 1585 -450 1600
rect -500 1565 -485 1585
rect -465 1565 -450 1585
rect -500 1535 -450 1565
rect -500 1515 -485 1535
rect -465 1515 -450 1535
rect -500 1485 -450 1515
rect -500 1465 -485 1485
rect -465 1465 -450 1485
rect -500 1435 -450 1465
rect -500 1415 -485 1435
rect -465 1415 -450 1435
rect -500 1385 -450 1415
rect -500 1365 -485 1385
rect -465 1365 -450 1385
rect -500 1335 -450 1365
rect -500 1315 -485 1335
rect -465 1315 -450 1335
rect -500 1285 -450 1315
rect -500 1265 -485 1285
rect -465 1265 -450 1285
rect -500 1235 -450 1265
rect -500 1215 -485 1235
rect -465 1215 -450 1235
rect -500 1185 -450 1215
rect -500 1165 -485 1185
rect -465 1165 -450 1185
rect -500 1135 -450 1165
rect -500 1115 -485 1135
rect -465 1115 -450 1135
rect -500 1085 -450 1115
rect -500 1065 -485 1085
rect -465 1065 -450 1085
rect -500 1035 -450 1065
rect -500 1015 -485 1035
rect -465 1015 -450 1035
rect -500 985 -450 1015
rect -500 965 -485 985
rect -465 965 -450 985
rect -500 935 -450 965
rect -500 915 -485 935
rect -465 915 -450 935
rect -500 900 -450 915
rect -350 1585 -300 1600
rect -350 1565 -335 1585
rect -315 1565 -300 1585
rect -350 1535 -300 1565
rect -350 1515 -335 1535
rect -315 1515 -300 1535
rect -350 1485 -300 1515
rect -350 1465 -335 1485
rect -315 1465 -300 1485
rect -350 1435 -300 1465
rect -350 1415 -335 1435
rect -315 1415 -300 1435
rect -350 1385 -300 1415
rect -350 1365 -335 1385
rect -315 1365 -300 1385
rect -350 1335 -300 1365
rect -350 1315 -335 1335
rect -315 1315 -300 1335
rect -350 1285 -300 1315
rect -350 1265 -335 1285
rect -315 1265 -300 1285
rect -350 1235 -300 1265
rect -350 1215 -335 1235
rect -315 1215 -300 1235
rect -350 1185 -300 1215
rect -350 1165 -335 1185
rect -315 1165 -300 1185
rect -350 1135 -300 1165
rect -350 1115 -335 1135
rect -315 1115 -300 1135
rect -350 1085 -300 1115
rect -350 1065 -335 1085
rect -315 1065 -300 1085
rect -350 1035 -300 1065
rect -350 1015 -335 1035
rect -315 1015 -300 1035
rect -350 985 -300 1015
rect -350 965 -335 985
rect -315 965 -300 985
rect -350 935 -300 965
rect -350 915 -335 935
rect -315 915 -300 935
rect -350 900 -300 915
rect -200 1585 -150 1600
rect -200 1565 -185 1585
rect -165 1565 -150 1585
rect -200 1535 -150 1565
rect -200 1515 -185 1535
rect -165 1515 -150 1535
rect -200 1485 -150 1515
rect -200 1465 -185 1485
rect -165 1465 -150 1485
rect -200 1435 -150 1465
rect -200 1415 -185 1435
rect -165 1415 -150 1435
rect -200 1385 -150 1415
rect -200 1365 -185 1385
rect -165 1365 -150 1385
rect -200 1335 -150 1365
rect -200 1315 -185 1335
rect -165 1315 -150 1335
rect -200 1285 -150 1315
rect -200 1265 -185 1285
rect -165 1265 -150 1285
rect -200 1235 -150 1265
rect -200 1215 -185 1235
rect -165 1215 -150 1235
rect -200 1185 -150 1215
rect -200 1165 -185 1185
rect -165 1165 -150 1185
rect -200 1135 -150 1165
rect -200 1115 -185 1135
rect -165 1115 -150 1135
rect -200 1085 -150 1115
rect -200 1065 -185 1085
rect -165 1065 -150 1085
rect -200 1035 -150 1065
rect -200 1015 -185 1035
rect -165 1015 -150 1035
rect -200 985 -150 1015
rect -200 965 -185 985
rect -165 965 -150 985
rect -200 935 -150 965
rect -200 915 -185 935
rect -165 915 -150 935
rect -200 900 -150 915
rect -50 1585 0 1600
rect -50 1565 -35 1585
rect -15 1565 0 1585
rect -50 1535 0 1565
rect -50 1515 -35 1535
rect -15 1515 0 1535
rect -50 1485 0 1515
rect -50 1465 -35 1485
rect -15 1465 0 1485
rect -50 1435 0 1465
rect -50 1415 -35 1435
rect -15 1415 0 1435
rect -50 1385 0 1415
rect -50 1365 -35 1385
rect -15 1365 0 1385
rect -50 1335 0 1365
rect -50 1315 -35 1335
rect -15 1315 0 1335
rect -50 1285 0 1315
rect -50 1265 -35 1285
rect -15 1265 0 1285
rect -50 1235 0 1265
rect -50 1215 -35 1235
rect -15 1215 0 1235
rect -50 1185 0 1215
rect -50 1165 -35 1185
rect -15 1165 0 1185
rect -50 1135 0 1165
rect -50 1115 -35 1135
rect -15 1115 0 1135
rect -50 1085 0 1115
rect -50 1065 -35 1085
rect -15 1065 0 1085
rect -50 1035 0 1065
rect -50 1015 -35 1035
rect -15 1015 0 1035
rect -50 985 0 1015
rect -50 965 -35 985
rect -15 965 0 985
rect -50 935 0 965
rect -50 915 -35 935
rect -15 915 0 935
rect -50 900 0 915
rect 1150 1585 1200 1600
rect 1150 1565 1165 1585
rect 1185 1565 1200 1585
rect 1150 1535 1200 1565
rect 1150 1515 1165 1535
rect 1185 1515 1200 1535
rect 1150 1485 1200 1515
rect 1150 1465 1165 1485
rect 1185 1465 1200 1485
rect 1150 1435 1200 1465
rect 1150 1415 1165 1435
rect 1185 1415 1200 1435
rect 1150 1385 1200 1415
rect 1150 1365 1165 1385
rect 1185 1365 1200 1385
rect 1150 1335 1200 1365
rect 1150 1315 1165 1335
rect 1185 1315 1200 1335
rect 1150 1285 1200 1315
rect 1150 1265 1165 1285
rect 1185 1265 1200 1285
rect 1150 1235 1200 1265
rect 1150 1215 1165 1235
rect 1185 1215 1200 1235
rect 1150 1185 1200 1215
rect 1150 1165 1165 1185
rect 1185 1165 1200 1185
rect 1150 1135 1200 1165
rect 1150 1115 1165 1135
rect 1185 1115 1200 1135
rect 1150 1085 1200 1115
rect 1150 1065 1165 1085
rect 1185 1065 1200 1085
rect 1150 1035 1200 1065
rect 1150 1015 1165 1035
rect 1185 1015 1200 1035
rect 1150 985 1200 1015
rect 1150 965 1165 985
rect 1185 965 1200 985
rect 1150 935 1200 965
rect 1150 915 1165 935
rect 1185 915 1200 935
rect 1150 900 1200 915
rect 1450 1585 1500 1600
rect 1450 1565 1465 1585
rect 1485 1565 1500 1585
rect 1450 1535 1500 1565
rect 1450 1515 1465 1535
rect 1485 1515 1500 1535
rect 1450 1485 1500 1515
rect 1450 1465 1465 1485
rect 1485 1465 1500 1485
rect 1450 1435 1500 1465
rect 1450 1415 1465 1435
rect 1485 1415 1500 1435
rect 1450 1385 1500 1415
rect 1450 1365 1465 1385
rect 1485 1365 1500 1385
rect 1450 1335 1500 1365
rect 1450 1315 1465 1335
rect 1485 1315 1500 1335
rect 1450 1285 1500 1315
rect 1450 1265 1465 1285
rect 1485 1265 1500 1285
rect 1450 1235 1500 1265
rect 1450 1215 1465 1235
rect 1485 1215 1500 1235
rect 1450 1185 1500 1215
rect 1450 1165 1465 1185
rect 1485 1165 1500 1185
rect 1450 1135 1500 1165
rect 1450 1115 1465 1135
rect 1485 1115 1500 1135
rect 1450 1085 1500 1115
rect 1450 1065 1465 1085
rect 1485 1065 1500 1085
rect 1450 1035 1500 1065
rect 1450 1015 1465 1035
rect 1485 1015 1500 1035
rect 1450 985 1500 1015
rect 1450 965 1465 985
rect 1485 965 1500 985
rect 1450 935 1500 965
rect 1450 915 1465 935
rect 1485 915 1500 935
rect 1450 900 1500 915
rect 1750 1585 1800 1600
rect 1750 1565 1765 1585
rect 1785 1565 1800 1585
rect 1750 1535 1800 1565
rect 1750 1515 1765 1535
rect 1785 1515 1800 1535
rect 1750 1485 1800 1515
rect 1750 1465 1765 1485
rect 1785 1465 1800 1485
rect 1750 1435 1800 1465
rect 1750 1415 1765 1435
rect 1785 1415 1800 1435
rect 1750 1385 1800 1415
rect 1750 1365 1765 1385
rect 1785 1365 1800 1385
rect 1750 1335 1800 1365
rect 1750 1315 1765 1335
rect 1785 1315 1800 1335
rect 1750 1285 1800 1315
rect 1750 1265 1765 1285
rect 1785 1265 1800 1285
rect 1750 1235 1800 1265
rect 1750 1215 1765 1235
rect 1785 1215 1800 1235
rect 1750 1185 1800 1215
rect 1750 1165 1765 1185
rect 1785 1165 1800 1185
rect 1750 1135 1800 1165
rect 1750 1115 1765 1135
rect 1785 1115 1800 1135
rect 1750 1085 1800 1115
rect 1750 1065 1765 1085
rect 1785 1065 1800 1085
rect 1750 1035 1800 1065
rect 1750 1015 1765 1035
rect 1785 1015 1800 1035
rect 1750 985 1800 1015
rect 1750 965 1765 985
rect 1785 965 1800 985
rect 1750 935 1800 965
rect 1750 915 1765 935
rect 1785 915 1800 935
rect 1750 900 1800 915
rect 2050 1585 2100 1600
rect 2050 1565 2065 1585
rect 2085 1565 2100 1585
rect 2050 1535 2100 1565
rect 2050 1515 2065 1535
rect 2085 1515 2100 1535
rect 2050 1485 2100 1515
rect 2050 1465 2065 1485
rect 2085 1465 2100 1485
rect 2050 1435 2100 1465
rect 2050 1415 2065 1435
rect 2085 1415 2100 1435
rect 2050 1385 2100 1415
rect 2050 1365 2065 1385
rect 2085 1365 2100 1385
rect 2050 1335 2100 1365
rect 2050 1315 2065 1335
rect 2085 1315 2100 1335
rect 2050 1285 2100 1315
rect 2050 1265 2065 1285
rect 2085 1265 2100 1285
rect 2050 1235 2100 1265
rect 2050 1215 2065 1235
rect 2085 1215 2100 1235
rect 2050 1185 2100 1215
rect 2050 1165 2065 1185
rect 2085 1165 2100 1185
rect 2050 1135 2100 1165
rect 2050 1115 2065 1135
rect 2085 1115 2100 1135
rect 2050 1085 2100 1115
rect 2050 1065 2065 1085
rect 2085 1065 2100 1085
rect 2050 1035 2100 1065
rect 2050 1015 2065 1035
rect 2085 1015 2100 1035
rect 2050 985 2100 1015
rect 2050 965 2065 985
rect 2085 965 2100 985
rect 2050 935 2100 965
rect 2050 915 2065 935
rect 2085 915 2100 935
rect 2050 900 2100 915
rect 2350 1585 2400 1600
rect 2350 1565 2365 1585
rect 2385 1565 2400 1585
rect 2350 1535 2400 1565
rect 2350 1515 2365 1535
rect 2385 1515 2400 1535
rect 2350 1485 2400 1515
rect 2350 1465 2365 1485
rect 2385 1465 2400 1485
rect 2350 1435 2400 1465
rect 2350 1415 2365 1435
rect 2385 1415 2400 1435
rect 2350 1385 2400 1415
rect 2350 1365 2365 1385
rect 2385 1365 2400 1385
rect 2350 1335 2400 1365
rect 2350 1315 2365 1335
rect 2385 1315 2400 1335
rect 2350 1285 2400 1315
rect 2350 1265 2365 1285
rect 2385 1265 2400 1285
rect 2350 1235 2400 1265
rect 2350 1215 2365 1235
rect 2385 1215 2400 1235
rect 2350 1185 2400 1215
rect 2350 1165 2365 1185
rect 2385 1165 2400 1185
rect 2350 1135 2400 1165
rect 2350 1115 2365 1135
rect 2385 1115 2400 1135
rect 2350 1085 2400 1115
rect 2350 1065 2365 1085
rect 2385 1065 2400 1085
rect 2350 1035 2400 1065
rect 2350 1015 2365 1035
rect 2385 1015 2400 1035
rect 2350 985 2400 1015
rect 2350 965 2365 985
rect 2385 965 2400 985
rect 2350 935 2400 965
rect 2350 915 2365 935
rect 2385 915 2400 935
rect 2350 900 2400 915
rect 2650 1585 2700 1600
rect 2650 1565 2665 1585
rect 2685 1565 2700 1585
rect 2650 1535 2700 1565
rect 2650 1515 2665 1535
rect 2685 1515 2700 1535
rect 2650 1485 2700 1515
rect 2650 1465 2665 1485
rect 2685 1465 2700 1485
rect 2650 1435 2700 1465
rect 2650 1415 2665 1435
rect 2685 1415 2700 1435
rect 2650 1385 2700 1415
rect 2650 1365 2665 1385
rect 2685 1365 2700 1385
rect 2650 1335 2700 1365
rect 2650 1315 2665 1335
rect 2685 1315 2700 1335
rect 2650 1285 2700 1315
rect 2650 1265 2665 1285
rect 2685 1265 2700 1285
rect 2650 1235 2700 1265
rect 2650 1215 2665 1235
rect 2685 1215 2700 1235
rect 2650 1185 2700 1215
rect 2650 1165 2665 1185
rect 2685 1165 2700 1185
rect 2650 1135 2700 1165
rect 2650 1115 2665 1135
rect 2685 1115 2700 1135
rect 2650 1085 2700 1115
rect 2650 1065 2665 1085
rect 2685 1065 2700 1085
rect 2650 1035 2700 1065
rect 2650 1015 2665 1035
rect 2685 1015 2700 1035
rect 2650 985 2700 1015
rect 2650 965 2665 985
rect 2685 965 2700 985
rect 2650 935 2700 965
rect 2650 915 2665 935
rect 2685 915 2700 935
rect 2650 900 2700 915
rect 2950 1585 3000 1600
rect 2950 1565 2965 1585
rect 2985 1565 3000 1585
rect 2950 1535 3000 1565
rect 2950 1515 2965 1535
rect 2985 1515 3000 1535
rect 2950 1485 3000 1515
rect 2950 1465 2965 1485
rect 2985 1465 3000 1485
rect 2950 1435 3000 1465
rect 2950 1415 2965 1435
rect 2985 1415 3000 1435
rect 2950 1385 3000 1415
rect 2950 1365 2965 1385
rect 2985 1365 3000 1385
rect 2950 1335 3000 1365
rect 2950 1315 2965 1335
rect 2985 1315 3000 1335
rect 2950 1285 3000 1315
rect 2950 1265 2965 1285
rect 2985 1265 3000 1285
rect 2950 1235 3000 1265
rect 2950 1215 2965 1235
rect 2985 1215 3000 1235
rect 2950 1185 3000 1215
rect 2950 1165 2965 1185
rect 2985 1165 3000 1185
rect 2950 1135 3000 1165
rect 2950 1115 2965 1135
rect 2985 1115 3000 1135
rect 2950 1085 3000 1115
rect 2950 1065 2965 1085
rect 2985 1065 3000 1085
rect 2950 1035 3000 1065
rect 2950 1015 2965 1035
rect 2985 1015 3000 1035
rect 2950 985 3000 1015
rect 2950 965 2965 985
rect 2985 965 3000 985
rect 2950 935 3000 965
rect 2950 915 2965 935
rect 2985 915 3000 935
rect 2950 900 3000 915
rect 3250 1585 3300 1600
rect 3250 1565 3265 1585
rect 3285 1565 3300 1585
rect 3250 1535 3300 1565
rect 3250 1515 3265 1535
rect 3285 1515 3300 1535
rect 3250 1485 3300 1515
rect 3250 1465 3265 1485
rect 3285 1465 3300 1485
rect 3250 1435 3300 1465
rect 3250 1415 3265 1435
rect 3285 1415 3300 1435
rect 3250 1385 3300 1415
rect 3250 1365 3265 1385
rect 3285 1365 3300 1385
rect 3250 1335 3300 1365
rect 3250 1315 3265 1335
rect 3285 1315 3300 1335
rect 3250 1285 3300 1315
rect 3250 1265 3265 1285
rect 3285 1265 3300 1285
rect 3250 1235 3300 1265
rect 3250 1215 3265 1235
rect 3285 1215 3300 1235
rect 3250 1185 3300 1215
rect 3250 1165 3265 1185
rect 3285 1165 3300 1185
rect 3250 1135 3300 1165
rect 3250 1115 3265 1135
rect 3285 1115 3300 1135
rect 3250 1085 3300 1115
rect 3250 1065 3265 1085
rect 3285 1065 3300 1085
rect 3250 1035 3300 1065
rect 3250 1015 3265 1035
rect 3285 1015 3300 1035
rect 3250 985 3300 1015
rect 3250 965 3265 985
rect 3285 965 3300 985
rect 3250 935 3300 965
rect 3250 915 3265 935
rect 3285 915 3300 935
rect 3250 900 3300 915
rect 3550 1585 3600 1600
rect 3550 1565 3565 1585
rect 3585 1565 3600 1585
rect 3550 1535 3600 1565
rect 3550 1515 3565 1535
rect 3585 1515 3600 1535
rect 3550 1485 3600 1515
rect 3550 1465 3565 1485
rect 3585 1465 3600 1485
rect 3550 1435 3600 1465
rect 3550 1415 3565 1435
rect 3585 1415 3600 1435
rect 3550 1385 3600 1415
rect 3550 1365 3565 1385
rect 3585 1365 3600 1385
rect 3550 1335 3600 1365
rect 3550 1315 3565 1335
rect 3585 1315 3600 1335
rect 3550 1285 3600 1315
rect 3550 1265 3565 1285
rect 3585 1265 3600 1285
rect 3550 1235 3600 1265
rect 3550 1215 3565 1235
rect 3585 1215 3600 1235
rect 3550 1185 3600 1215
rect 3550 1165 3565 1185
rect 3585 1165 3600 1185
rect 3550 1135 3600 1165
rect 3550 1115 3565 1135
rect 3585 1115 3600 1135
rect 3550 1085 3600 1115
rect 3550 1065 3565 1085
rect 3585 1065 3600 1085
rect 3550 1035 3600 1065
rect 3550 1015 3565 1035
rect 3585 1015 3600 1035
rect 3550 985 3600 1015
rect 3550 965 3565 985
rect 3585 965 3600 985
rect 3550 935 3600 965
rect 3550 915 3565 935
rect 3585 915 3600 935
rect 3550 900 3600 915
rect 3700 1585 3750 1600
rect 3700 1565 3715 1585
rect 3735 1565 3750 1585
rect 3700 1535 3750 1565
rect 3700 1515 3715 1535
rect 3735 1515 3750 1535
rect 3700 1485 3750 1515
rect 3700 1465 3715 1485
rect 3735 1465 3750 1485
rect 3700 1435 3750 1465
rect 3700 1415 3715 1435
rect 3735 1415 3750 1435
rect 3700 1385 3750 1415
rect 3700 1365 3715 1385
rect 3735 1365 3750 1385
rect 3700 1335 3750 1365
rect 3700 1315 3715 1335
rect 3735 1315 3750 1335
rect 3700 1285 3750 1315
rect 3700 1265 3715 1285
rect 3735 1265 3750 1285
rect 3700 1235 3750 1265
rect 3700 1215 3715 1235
rect 3735 1215 3750 1235
rect 3700 1185 3750 1215
rect 3700 1165 3715 1185
rect 3735 1165 3750 1185
rect 3700 1135 3750 1165
rect 3700 1115 3715 1135
rect 3735 1115 3750 1135
rect 3700 1085 3750 1115
rect 3700 1065 3715 1085
rect 3735 1065 3750 1085
rect 3700 1035 3750 1065
rect 3700 1015 3715 1035
rect 3735 1015 3750 1035
rect 3700 985 3750 1015
rect 3700 965 3715 985
rect 3735 965 3750 985
rect 3700 935 3750 965
rect 3700 915 3715 935
rect 3735 915 3750 935
rect 3700 900 3750 915
rect 3850 1585 3900 1600
rect 3850 1565 3865 1585
rect 3885 1565 3900 1585
rect 3850 1535 3900 1565
rect 3850 1515 3865 1535
rect 3885 1515 3900 1535
rect 3850 1485 3900 1515
rect 3850 1465 3865 1485
rect 3885 1465 3900 1485
rect 3850 1435 3900 1465
rect 3850 1415 3865 1435
rect 3885 1415 3900 1435
rect 3850 1385 3900 1415
rect 3850 1365 3865 1385
rect 3885 1365 3900 1385
rect 3850 1335 3900 1365
rect 3850 1315 3865 1335
rect 3885 1315 3900 1335
rect 3850 1285 3900 1315
rect 3850 1265 3865 1285
rect 3885 1265 3900 1285
rect 3850 1235 3900 1265
rect 3850 1215 3865 1235
rect 3885 1215 3900 1235
rect 3850 1185 3900 1215
rect 3850 1165 3865 1185
rect 3885 1165 3900 1185
rect 3850 1135 3900 1165
rect 3850 1115 3865 1135
rect 3885 1115 3900 1135
rect 3850 1085 3900 1115
rect 3850 1065 3865 1085
rect 3885 1065 3900 1085
rect 3850 1035 3900 1065
rect 3850 1015 3865 1035
rect 3885 1015 3900 1035
rect 3850 985 3900 1015
rect 3850 965 3865 985
rect 3885 965 3900 985
rect 3850 935 3900 965
rect 3850 915 3865 935
rect 3885 915 3900 935
rect 3850 900 3900 915
rect 4000 1585 4050 1600
rect 4000 1565 4015 1585
rect 4035 1565 4050 1585
rect 4000 1535 4050 1565
rect 4000 1515 4015 1535
rect 4035 1515 4050 1535
rect 4000 1485 4050 1515
rect 4000 1465 4015 1485
rect 4035 1465 4050 1485
rect 4000 1435 4050 1465
rect 4000 1415 4015 1435
rect 4035 1415 4050 1435
rect 4000 1385 4050 1415
rect 4000 1365 4015 1385
rect 4035 1365 4050 1385
rect 4000 1335 4050 1365
rect 4000 1315 4015 1335
rect 4035 1315 4050 1335
rect 4000 1285 4050 1315
rect 4000 1265 4015 1285
rect 4035 1265 4050 1285
rect 4000 1235 4050 1265
rect 4000 1215 4015 1235
rect 4035 1215 4050 1235
rect 4000 1185 4050 1215
rect 4000 1165 4015 1185
rect 4035 1165 4050 1185
rect 4000 1135 4050 1165
rect 4000 1115 4015 1135
rect 4035 1115 4050 1135
rect 4000 1085 4050 1115
rect 4000 1065 4015 1085
rect 4035 1065 4050 1085
rect 4000 1035 4050 1065
rect 4000 1015 4015 1035
rect 4035 1015 4050 1035
rect 4000 985 4050 1015
rect 4000 965 4015 985
rect 4035 965 4050 985
rect 4000 935 4050 965
rect 4000 915 4015 935
rect 4035 915 4050 935
rect 4000 900 4050 915
rect 4150 1585 4200 1600
rect 4150 1565 4165 1585
rect 4185 1565 4200 1585
rect 4150 1535 4200 1565
rect 4150 1515 4165 1535
rect 4185 1515 4200 1535
rect 4150 1485 4200 1515
rect 4150 1465 4165 1485
rect 4185 1465 4200 1485
rect 4150 1435 4200 1465
rect 4150 1415 4165 1435
rect 4185 1415 4200 1435
rect 4150 1385 4200 1415
rect 4150 1365 4165 1385
rect 4185 1365 4200 1385
rect 4150 1335 4200 1365
rect 4150 1315 4165 1335
rect 4185 1315 4200 1335
rect 4150 1285 4200 1315
rect 4150 1265 4165 1285
rect 4185 1265 4200 1285
rect 4150 1235 4200 1265
rect 4150 1215 4165 1235
rect 4185 1215 4200 1235
rect 4150 1185 4200 1215
rect 4150 1165 4165 1185
rect 4185 1165 4200 1185
rect 4150 1135 4200 1165
rect 4150 1115 4165 1135
rect 4185 1115 4200 1135
rect 4150 1085 4200 1115
rect 4150 1065 4165 1085
rect 4185 1065 4200 1085
rect 4150 1035 4200 1065
rect 4150 1015 4165 1035
rect 4185 1015 4200 1035
rect 4150 985 4200 1015
rect 4150 965 4165 985
rect 4185 965 4200 985
rect 4150 935 4200 965
rect 4150 915 4165 935
rect 4185 915 4200 935
rect 4150 900 4200 915
rect 4300 1585 4350 1600
rect 4300 1565 4315 1585
rect 4335 1565 4350 1585
rect 4300 1535 4350 1565
rect 4300 1515 4315 1535
rect 4335 1515 4350 1535
rect 4300 1485 4350 1515
rect 4300 1465 4315 1485
rect 4335 1465 4350 1485
rect 4300 1435 4350 1465
rect 4300 1415 4315 1435
rect 4335 1415 4350 1435
rect 4300 1385 4350 1415
rect 4300 1365 4315 1385
rect 4335 1365 4350 1385
rect 4300 1335 4350 1365
rect 4300 1315 4315 1335
rect 4335 1315 4350 1335
rect 4300 1285 4350 1315
rect 4300 1265 4315 1285
rect 4335 1265 4350 1285
rect 4300 1235 4350 1265
rect 4300 1215 4315 1235
rect 4335 1215 4350 1235
rect 4300 1185 4350 1215
rect 4300 1165 4315 1185
rect 4335 1165 4350 1185
rect 4300 1135 4350 1165
rect 4300 1115 4315 1135
rect 4335 1115 4350 1135
rect 4300 1085 4350 1115
rect 4300 1065 4315 1085
rect 4335 1065 4350 1085
rect 4300 1035 4350 1065
rect 4300 1015 4315 1035
rect 4335 1015 4350 1035
rect 4300 985 4350 1015
rect 4300 965 4315 985
rect 4335 965 4350 985
rect 4300 935 4350 965
rect 4300 915 4315 935
rect 4335 915 4350 935
rect 4300 900 4350 915
rect 4450 1585 4500 1600
rect 4450 1565 4465 1585
rect 4485 1565 4500 1585
rect 4450 1535 4500 1565
rect 4450 1515 4465 1535
rect 4485 1515 4500 1535
rect 4450 1485 4500 1515
rect 4450 1465 4465 1485
rect 4485 1465 4500 1485
rect 4450 1435 4500 1465
rect 4450 1415 4465 1435
rect 4485 1415 4500 1435
rect 4450 1385 4500 1415
rect 4450 1365 4465 1385
rect 4485 1365 4500 1385
rect 4450 1335 4500 1365
rect 4450 1315 4465 1335
rect 4485 1315 4500 1335
rect 4450 1285 4500 1315
rect 4450 1265 4465 1285
rect 4485 1265 4500 1285
rect 4450 1235 4500 1265
rect 4450 1215 4465 1235
rect 4485 1215 4500 1235
rect 4450 1185 4500 1215
rect 4450 1165 4465 1185
rect 4485 1165 4500 1185
rect 4450 1135 4500 1165
rect 4450 1115 4465 1135
rect 4485 1115 4500 1135
rect 4450 1085 4500 1115
rect 4450 1065 4465 1085
rect 4485 1065 4500 1085
rect 4450 1035 4500 1065
rect 4450 1015 4465 1035
rect 4485 1015 4500 1035
rect 4450 985 4500 1015
rect 4450 965 4465 985
rect 4485 965 4500 985
rect 4450 935 4500 965
rect 4450 915 4465 935
rect 4485 915 4500 935
rect 4450 900 4500 915
rect 4600 1585 4650 1600
rect 4600 1565 4615 1585
rect 4635 1565 4650 1585
rect 4600 1535 4650 1565
rect 4600 1515 4615 1535
rect 4635 1515 4650 1535
rect 4600 1485 4650 1515
rect 4600 1465 4615 1485
rect 4635 1465 4650 1485
rect 4600 1435 4650 1465
rect 4600 1415 4615 1435
rect 4635 1415 4650 1435
rect 4600 1385 4650 1415
rect 4600 1365 4615 1385
rect 4635 1365 4650 1385
rect 4600 1335 4650 1365
rect 4600 1315 4615 1335
rect 4635 1315 4650 1335
rect 4600 1285 4650 1315
rect 4600 1265 4615 1285
rect 4635 1265 4650 1285
rect 4600 1235 4650 1265
rect 4600 1215 4615 1235
rect 4635 1215 4650 1235
rect 4600 1185 4650 1215
rect 4600 1165 4615 1185
rect 4635 1165 4650 1185
rect 4600 1135 4650 1165
rect 4600 1115 4615 1135
rect 4635 1115 4650 1135
rect 4600 1085 4650 1115
rect 4600 1065 4615 1085
rect 4635 1065 4650 1085
rect 4600 1035 4650 1065
rect 4600 1015 4615 1035
rect 4635 1015 4650 1035
rect 4600 985 4650 1015
rect 4600 965 4615 985
rect 4635 965 4650 985
rect 4600 935 4650 965
rect 4600 915 4615 935
rect 4635 915 4650 935
rect 4600 900 4650 915
rect 4750 1585 4800 1600
rect 4750 1565 4765 1585
rect 4785 1565 4800 1585
rect 4750 1535 4800 1565
rect 4750 1515 4765 1535
rect 4785 1515 4800 1535
rect 4750 1485 4800 1515
rect 4750 1465 4765 1485
rect 4785 1465 4800 1485
rect 4750 1435 4800 1465
rect 4750 1415 4765 1435
rect 4785 1415 4800 1435
rect 4750 1385 4800 1415
rect 4750 1365 4765 1385
rect 4785 1365 4800 1385
rect 4750 1335 4800 1365
rect 4750 1315 4765 1335
rect 4785 1315 4800 1335
rect 4750 1285 4800 1315
rect 4750 1265 4765 1285
rect 4785 1265 4800 1285
rect 4750 1235 4800 1265
rect 4750 1215 4765 1235
rect 4785 1215 4800 1235
rect 4750 1185 4800 1215
rect 4750 1165 4765 1185
rect 4785 1165 4800 1185
rect 4750 1135 4800 1165
rect 4750 1115 4765 1135
rect 4785 1115 4800 1135
rect 4750 1085 4800 1115
rect 4750 1065 4765 1085
rect 4785 1065 4800 1085
rect 4750 1035 4800 1065
rect 4750 1015 4765 1035
rect 4785 1015 4800 1035
rect 4750 985 4800 1015
rect 4750 965 4765 985
rect 4785 965 4800 985
rect 4750 935 4800 965
rect 4750 915 4765 935
rect 4785 915 4800 935
rect 4750 900 4800 915
rect 5050 1585 5100 1600
rect 5050 1565 5065 1585
rect 5085 1565 5100 1585
rect 5050 1535 5100 1565
rect 5050 1515 5065 1535
rect 5085 1515 5100 1535
rect 5050 1485 5100 1515
rect 5050 1465 5065 1485
rect 5085 1465 5100 1485
rect 5050 1435 5100 1465
rect 5050 1415 5065 1435
rect 5085 1415 5100 1435
rect 5050 1385 5100 1415
rect 5050 1365 5065 1385
rect 5085 1365 5100 1385
rect 5050 1335 5100 1365
rect 5050 1315 5065 1335
rect 5085 1315 5100 1335
rect 5050 1285 5100 1315
rect 5050 1265 5065 1285
rect 5085 1265 5100 1285
rect 5050 1235 5100 1265
rect 5050 1215 5065 1235
rect 5085 1215 5100 1235
rect 5050 1185 5100 1215
rect 5050 1165 5065 1185
rect 5085 1165 5100 1185
rect 5050 1135 5100 1165
rect 5050 1115 5065 1135
rect 5085 1115 5100 1135
rect 5050 1085 5100 1115
rect 5050 1065 5065 1085
rect 5085 1065 5100 1085
rect 5050 1035 5100 1065
rect 5050 1015 5065 1035
rect 5085 1015 5100 1035
rect 5050 985 5100 1015
rect 5050 965 5065 985
rect 5085 965 5100 985
rect 5050 935 5100 965
rect 5050 915 5065 935
rect 5085 915 5100 935
rect 5050 900 5100 915
rect 5350 1585 5400 1600
rect 5350 1565 5365 1585
rect 5385 1565 5400 1585
rect 5350 1535 5400 1565
rect 5350 1515 5365 1535
rect 5385 1515 5400 1535
rect 5350 1485 5400 1515
rect 5350 1465 5365 1485
rect 5385 1465 5400 1485
rect 5350 1435 5400 1465
rect 5350 1415 5365 1435
rect 5385 1415 5400 1435
rect 5350 1385 5400 1415
rect 5350 1365 5365 1385
rect 5385 1365 5400 1385
rect 5350 1335 5400 1365
rect 5350 1315 5365 1335
rect 5385 1315 5400 1335
rect 5350 1285 5400 1315
rect 5350 1265 5365 1285
rect 5385 1265 5400 1285
rect 5350 1235 5400 1265
rect 5350 1215 5365 1235
rect 5385 1215 5400 1235
rect 5350 1185 5400 1215
rect 5350 1165 5365 1185
rect 5385 1165 5400 1185
rect 5350 1135 5400 1165
rect 5350 1115 5365 1135
rect 5385 1115 5400 1135
rect 5350 1085 5400 1115
rect 5350 1065 5365 1085
rect 5385 1065 5400 1085
rect 5350 1035 5400 1065
rect 5350 1015 5365 1035
rect 5385 1015 5400 1035
rect 5350 985 5400 1015
rect 5350 965 5365 985
rect 5385 965 5400 985
rect 5350 935 5400 965
rect 5350 915 5365 935
rect 5385 915 5400 935
rect 5350 900 5400 915
rect 5650 1585 5700 1600
rect 5650 1565 5665 1585
rect 5685 1565 5700 1585
rect 5650 1535 5700 1565
rect 5650 1515 5665 1535
rect 5685 1515 5700 1535
rect 5650 1485 5700 1515
rect 5650 1465 5665 1485
rect 5685 1465 5700 1485
rect 5650 1435 5700 1465
rect 5650 1415 5665 1435
rect 5685 1415 5700 1435
rect 5650 1385 5700 1415
rect 5650 1365 5665 1385
rect 5685 1365 5700 1385
rect 5650 1335 5700 1365
rect 5650 1315 5665 1335
rect 5685 1315 5700 1335
rect 5650 1285 5700 1315
rect 5650 1265 5665 1285
rect 5685 1265 5700 1285
rect 5650 1235 5700 1265
rect 5650 1215 5665 1235
rect 5685 1215 5700 1235
rect 5650 1185 5700 1215
rect 5650 1165 5665 1185
rect 5685 1165 5700 1185
rect 5650 1135 5700 1165
rect 5650 1115 5665 1135
rect 5685 1115 5700 1135
rect 5650 1085 5700 1115
rect 5650 1065 5665 1085
rect 5685 1065 5700 1085
rect 5650 1035 5700 1065
rect 5650 1015 5665 1035
rect 5685 1015 5700 1035
rect 5650 985 5700 1015
rect 5650 965 5665 985
rect 5685 965 5700 985
rect 5650 935 5700 965
rect 5650 915 5665 935
rect 5685 915 5700 935
rect 5650 900 5700 915
rect 5950 1585 6000 1600
rect 5950 1565 5965 1585
rect 5985 1565 6000 1585
rect 5950 1535 6000 1565
rect 5950 1515 5965 1535
rect 5985 1515 6000 1535
rect 5950 1485 6000 1515
rect 5950 1465 5965 1485
rect 5985 1465 6000 1485
rect 5950 1435 6000 1465
rect 5950 1415 5965 1435
rect 5985 1415 6000 1435
rect 5950 1385 6000 1415
rect 5950 1365 5965 1385
rect 5985 1365 6000 1385
rect 5950 1335 6000 1365
rect 5950 1315 5965 1335
rect 5985 1315 6000 1335
rect 5950 1285 6000 1315
rect 5950 1265 5965 1285
rect 5985 1265 6000 1285
rect 5950 1235 6000 1265
rect 5950 1215 5965 1235
rect 5985 1215 6000 1235
rect 5950 1185 6000 1215
rect 5950 1165 5965 1185
rect 5985 1165 6000 1185
rect 5950 1135 6000 1165
rect 5950 1115 5965 1135
rect 5985 1115 6000 1135
rect 5950 1085 6000 1115
rect 5950 1065 5965 1085
rect 5985 1065 6000 1085
rect 5950 1035 6000 1065
rect 5950 1015 5965 1035
rect 5985 1015 6000 1035
rect 5950 985 6000 1015
rect 5950 965 5965 985
rect 5985 965 6000 985
rect 5950 935 6000 965
rect 5950 915 5965 935
rect 5985 915 6000 935
rect 5950 900 6000 915
rect 6250 1585 6300 1600
rect 6250 1565 6265 1585
rect 6285 1565 6300 1585
rect 6250 1535 6300 1565
rect 6250 1515 6265 1535
rect 6285 1515 6300 1535
rect 6250 1485 6300 1515
rect 6250 1465 6265 1485
rect 6285 1465 6300 1485
rect 6250 1435 6300 1465
rect 6250 1415 6265 1435
rect 6285 1415 6300 1435
rect 6250 1385 6300 1415
rect 6250 1365 6265 1385
rect 6285 1365 6300 1385
rect 6250 1335 6300 1365
rect 6250 1315 6265 1335
rect 6285 1315 6300 1335
rect 6250 1285 6300 1315
rect 6250 1265 6265 1285
rect 6285 1265 6300 1285
rect 6250 1235 6300 1265
rect 6250 1215 6265 1235
rect 6285 1215 6300 1235
rect 6250 1185 6300 1215
rect 6250 1165 6265 1185
rect 6285 1165 6300 1185
rect 6250 1135 6300 1165
rect 6250 1115 6265 1135
rect 6285 1115 6300 1135
rect 6250 1085 6300 1115
rect 6250 1065 6265 1085
rect 6285 1065 6300 1085
rect 6250 1035 6300 1065
rect 6250 1015 6265 1035
rect 6285 1015 6300 1035
rect 6250 985 6300 1015
rect 6250 965 6265 985
rect 6285 965 6300 985
rect 6250 935 6300 965
rect 6250 915 6265 935
rect 6285 915 6300 935
rect 6250 900 6300 915
rect 6550 1585 6600 1600
rect 6550 1565 6565 1585
rect 6585 1565 6600 1585
rect 6550 1535 6600 1565
rect 6550 1515 6565 1535
rect 6585 1515 6600 1535
rect 6550 1485 6600 1515
rect 6550 1465 6565 1485
rect 6585 1465 6600 1485
rect 6550 1435 6600 1465
rect 6550 1415 6565 1435
rect 6585 1415 6600 1435
rect 6550 1385 6600 1415
rect 6550 1365 6565 1385
rect 6585 1365 6600 1385
rect 6550 1335 6600 1365
rect 6550 1315 6565 1335
rect 6585 1315 6600 1335
rect 6550 1285 6600 1315
rect 6550 1265 6565 1285
rect 6585 1265 6600 1285
rect 6550 1235 6600 1265
rect 6550 1215 6565 1235
rect 6585 1215 6600 1235
rect 6550 1185 6600 1215
rect 6550 1165 6565 1185
rect 6585 1165 6600 1185
rect 6550 1135 6600 1165
rect 6550 1115 6565 1135
rect 6585 1115 6600 1135
rect 6550 1085 6600 1115
rect 6550 1065 6565 1085
rect 6585 1065 6600 1085
rect 6550 1035 6600 1065
rect 6550 1015 6565 1035
rect 6585 1015 6600 1035
rect 6550 985 6600 1015
rect 6550 965 6565 985
rect 6585 965 6600 985
rect 6550 935 6600 965
rect 6550 915 6565 935
rect 6585 915 6600 935
rect 6550 900 6600 915
rect 6850 1585 6900 1600
rect 6850 1565 6865 1585
rect 6885 1565 6900 1585
rect 6850 1535 6900 1565
rect 6850 1515 6865 1535
rect 6885 1515 6900 1535
rect 6850 1485 6900 1515
rect 6850 1465 6865 1485
rect 6885 1465 6900 1485
rect 6850 1435 6900 1465
rect 6850 1415 6865 1435
rect 6885 1415 6900 1435
rect 6850 1385 6900 1415
rect 6850 1365 6865 1385
rect 6885 1365 6900 1385
rect 6850 1335 6900 1365
rect 6850 1315 6865 1335
rect 6885 1315 6900 1335
rect 6850 1285 6900 1315
rect 6850 1265 6865 1285
rect 6885 1265 6900 1285
rect 6850 1235 6900 1265
rect 6850 1215 6865 1235
rect 6885 1215 6900 1235
rect 6850 1185 6900 1215
rect 6850 1165 6865 1185
rect 6885 1165 6900 1185
rect 6850 1135 6900 1165
rect 6850 1115 6865 1135
rect 6885 1115 6900 1135
rect 6850 1085 6900 1115
rect 6850 1065 6865 1085
rect 6885 1065 6900 1085
rect 6850 1035 6900 1065
rect 6850 1015 6865 1035
rect 6885 1015 6900 1035
rect 6850 985 6900 1015
rect 6850 965 6865 985
rect 6885 965 6900 985
rect 6850 935 6900 965
rect 6850 915 6865 935
rect 6885 915 6900 935
rect 6850 900 6900 915
rect 7150 1585 7200 1600
rect 7150 1565 7165 1585
rect 7185 1565 7200 1585
rect 7150 1535 7200 1565
rect 7150 1515 7165 1535
rect 7185 1515 7200 1535
rect 7150 1485 7200 1515
rect 7150 1465 7165 1485
rect 7185 1465 7200 1485
rect 7150 1435 7200 1465
rect 7150 1415 7165 1435
rect 7185 1415 7200 1435
rect 7150 1385 7200 1415
rect 7150 1365 7165 1385
rect 7185 1365 7200 1385
rect 7150 1335 7200 1365
rect 7150 1315 7165 1335
rect 7185 1315 7200 1335
rect 7150 1285 7200 1315
rect 7150 1265 7165 1285
rect 7185 1265 7200 1285
rect 7150 1235 7200 1265
rect 7150 1215 7165 1235
rect 7185 1215 7200 1235
rect 7150 1185 7200 1215
rect 7150 1165 7165 1185
rect 7185 1165 7200 1185
rect 7150 1135 7200 1165
rect 7150 1115 7165 1135
rect 7185 1115 7200 1135
rect 7150 1085 7200 1115
rect 7150 1065 7165 1085
rect 7185 1065 7200 1085
rect 7150 1035 7200 1065
rect 7150 1015 7165 1035
rect 7185 1015 7200 1035
rect 7150 985 7200 1015
rect 7150 965 7165 985
rect 7185 965 7200 985
rect 7150 935 7200 965
rect 7150 915 7165 935
rect 7185 915 7200 935
rect 7150 900 7200 915
rect 8350 1585 8400 1600
rect 8350 1565 8365 1585
rect 8385 1565 8400 1585
rect 8350 1535 8400 1565
rect 8350 1515 8365 1535
rect 8385 1515 8400 1535
rect 8350 1485 8400 1515
rect 8350 1465 8365 1485
rect 8385 1465 8400 1485
rect 8350 1435 8400 1465
rect 8350 1415 8365 1435
rect 8385 1415 8400 1435
rect 8350 1385 8400 1415
rect 8350 1365 8365 1385
rect 8385 1365 8400 1385
rect 8350 1335 8400 1365
rect 8350 1315 8365 1335
rect 8385 1315 8400 1335
rect 8350 1285 8400 1315
rect 8350 1265 8365 1285
rect 8385 1265 8400 1285
rect 8350 1235 8400 1265
rect 8350 1215 8365 1235
rect 8385 1215 8400 1235
rect 8350 1185 8400 1215
rect 8350 1165 8365 1185
rect 8385 1165 8400 1185
rect 8350 1135 8400 1165
rect 8350 1115 8365 1135
rect 8385 1115 8400 1135
rect 8350 1085 8400 1115
rect 8350 1065 8365 1085
rect 8385 1065 8400 1085
rect 8350 1035 8400 1065
rect 8350 1015 8365 1035
rect 8385 1015 8400 1035
rect 8350 985 8400 1015
rect 8350 965 8365 985
rect 8385 965 8400 985
rect 8350 935 8400 965
rect 8350 915 8365 935
rect 8385 915 8400 935
rect 8350 900 8400 915
rect 9550 1585 9600 1600
rect 9550 1565 9565 1585
rect 9585 1565 9600 1585
rect 9550 1535 9600 1565
rect 9550 1515 9565 1535
rect 9585 1515 9600 1535
rect 9550 1485 9600 1515
rect 9550 1465 9565 1485
rect 9585 1465 9600 1485
rect 9550 1435 9600 1465
rect 9550 1415 9565 1435
rect 9585 1415 9600 1435
rect 9550 1385 9600 1415
rect 9550 1365 9565 1385
rect 9585 1365 9600 1385
rect 9550 1335 9600 1365
rect 9550 1315 9565 1335
rect 9585 1315 9600 1335
rect 9550 1285 9600 1315
rect 9550 1265 9565 1285
rect 9585 1265 9600 1285
rect 9550 1235 9600 1265
rect 9550 1215 9565 1235
rect 9585 1215 9600 1235
rect 9550 1185 9600 1215
rect 9550 1165 9565 1185
rect 9585 1165 9600 1185
rect 9550 1135 9600 1165
rect 9550 1115 9565 1135
rect 9585 1115 9600 1135
rect 9550 1085 9600 1115
rect 9550 1065 9565 1085
rect 9585 1065 9600 1085
rect 9550 1035 9600 1065
rect 9550 1015 9565 1035
rect 9585 1015 9600 1035
rect 9550 985 9600 1015
rect 9550 965 9565 985
rect 9585 965 9600 985
rect 9550 935 9600 965
rect 9550 915 9565 935
rect 9585 915 9600 935
rect 9550 900 9600 915
rect 10750 1585 10800 1600
rect 10750 1565 10765 1585
rect 10785 1565 10800 1585
rect 10750 1535 10800 1565
rect 10750 1515 10765 1535
rect 10785 1515 10800 1535
rect 10750 1485 10800 1515
rect 10750 1465 10765 1485
rect 10785 1465 10800 1485
rect 10750 1435 10800 1465
rect 10750 1415 10765 1435
rect 10785 1415 10800 1435
rect 10750 1385 10800 1415
rect 10750 1365 10765 1385
rect 10785 1365 10800 1385
rect 10750 1335 10800 1365
rect 10750 1315 10765 1335
rect 10785 1315 10800 1335
rect 10750 1285 10800 1315
rect 10750 1265 10765 1285
rect 10785 1265 10800 1285
rect 10750 1235 10800 1265
rect 10750 1215 10765 1235
rect 10785 1215 10800 1235
rect 10750 1185 10800 1215
rect 10750 1165 10765 1185
rect 10785 1165 10800 1185
rect 10750 1135 10800 1165
rect 10750 1115 10765 1135
rect 10785 1115 10800 1135
rect 10750 1085 10800 1115
rect 10750 1065 10765 1085
rect 10785 1065 10800 1085
rect 10750 1035 10800 1065
rect 10750 1015 10765 1035
rect 10785 1015 10800 1035
rect 10750 985 10800 1015
rect 10750 965 10765 985
rect 10785 965 10800 985
rect 10750 935 10800 965
rect 10750 915 10765 935
rect 10785 915 10800 935
rect 10750 900 10800 915
rect 11950 1585 12000 1600
rect 11950 1565 11965 1585
rect 11985 1565 12000 1585
rect 11950 1535 12000 1565
rect 11950 1515 11965 1535
rect 11985 1515 12000 1535
rect 11950 1485 12000 1515
rect 11950 1465 11965 1485
rect 11985 1465 12000 1485
rect 11950 1435 12000 1465
rect 11950 1415 11965 1435
rect 11985 1415 12000 1435
rect 11950 1385 12000 1415
rect 11950 1365 11965 1385
rect 11985 1365 12000 1385
rect 11950 1335 12000 1365
rect 11950 1315 11965 1335
rect 11985 1315 12000 1335
rect 11950 1285 12000 1315
rect 11950 1265 11965 1285
rect 11985 1265 12000 1285
rect 11950 1235 12000 1265
rect 11950 1215 11965 1235
rect 11985 1215 12000 1235
rect 11950 1185 12000 1215
rect 11950 1165 11965 1185
rect 11985 1165 12000 1185
rect 11950 1135 12000 1165
rect 11950 1115 11965 1135
rect 11985 1115 12000 1135
rect 11950 1085 12000 1115
rect 11950 1065 11965 1085
rect 11985 1065 12000 1085
rect 11950 1035 12000 1065
rect 11950 1015 11965 1035
rect 11985 1015 12000 1035
rect 11950 985 12000 1015
rect 11950 965 11965 985
rect 11985 965 12000 985
rect 11950 935 12000 965
rect 11950 915 11965 935
rect 11985 915 12000 935
rect 11950 900 12000 915
rect 12250 1585 12300 1600
rect 12250 1565 12265 1585
rect 12285 1565 12300 1585
rect 12250 1535 12300 1565
rect 12250 1515 12265 1535
rect 12285 1515 12300 1535
rect 12250 1485 12300 1515
rect 12250 1465 12265 1485
rect 12285 1465 12300 1485
rect 12250 1435 12300 1465
rect 12250 1415 12265 1435
rect 12285 1415 12300 1435
rect 12250 1385 12300 1415
rect 12250 1365 12265 1385
rect 12285 1365 12300 1385
rect 12250 1335 12300 1365
rect 12250 1315 12265 1335
rect 12285 1315 12300 1335
rect 12250 1285 12300 1315
rect 12250 1265 12265 1285
rect 12285 1265 12300 1285
rect 12250 1235 12300 1265
rect 12250 1215 12265 1235
rect 12285 1215 12300 1235
rect 12250 1185 12300 1215
rect 12250 1165 12265 1185
rect 12285 1165 12300 1185
rect 12250 1135 12300 1165
rect 12250 1115 12265 1135
rect 12285 1115 12300 1135
rect 12250 1085 12300 1115
rect 12250 1065 12265 1085
rect 12285 1065 12300 1085
rect 12250 1035 12300 1065
rect 12250 1015 12265 1035
rect 12285 1015 12300 1035
rect 12250 985 12300 1015
rect 12250 965 12265 985
rect 12285 965 12300 985
rect 12250 935 12300 965
rect 12250 915 12265 935
rect 12285 915 12300 935
rect 12250 900 12300 915
rect 12550 1585 12600 1600
rect 12550 1565 12565 1585
rect 12585 1565 12600 1585
rect 12550 1535 12600 1565
rect 12550 1515 12565 1535
rect 12585 1515 12600 1535
rect 12550 1485 12600 1515
rect 12550 1465 12565 1485
rect 12585 1465 12600 1485
rect 12550 1435 12600 1465
rect 12550 1415 12565 1435
rect 12585 1415 12600 1435
rect 12550 1385 12600 1415
rect 12550 1365 12565 1385
rect 12585 1365 12600 1385
rect 12550 1335 12600 1365
rect 12550 1315 12565 1335
rect 12585 1315 12600 1335
rect 12550 1285 12600 1315
rect 12550 1265 12565 1285
rect 12585 1265 12600 1285
rect 12550 1235 12600 1265
rect 12550 1215 12565 1235
rect 12585 1215 12600 1235
rect 12550 1185 12600 1215
rect 12550 1165 12565 1185
rect 12585 1165 12600 1185
rect 12550 1135 12600 1165
rect 12550 1115 12565 1135
rect 12585 1115 12600 1135
rect 12550 1085 12600 1115
rect 12550 1065 12565 1085
rect 12585 1065 12600 1085
rect 12550 1035 12600 1065
rect 12550 1015 12565 1035
rect 12585 1015 12600 1035
rect 12550 985 12600 1015
rect 12550 965 12565 985
rect 12585 965 12600 985
rect 12550 935 12600 965
rect 12550 915 12565 935
rect 12585 915 12600 935
rect 12550 900 12600 915
rect 12850 1585 12900 1600
rect 12850 1565 12865 1585
rect 12885 1565 12900 1585
rect 12850 1535 12900 1565
rect 12850 1515 12865 1535
rect 12885 1515 12900 1535
rect 12850 1485 12900 1515
rect 12850 1465 12865 1485
rect 12885 1465 12900 1485
rect 12850 1435 12900 1465
rect 12850 1415 12865 1435
rect 12885 1415 12900 1435
rect 12850 1385 12900 1415
rect 12850 1365 12865 1385
rect 12885 1365 12900 1385
rect 12850 1335 12900 1365
rect 12850 1315 12865 1335
rect 12885 1315 12900 1335
rect 12850 1285 12900 1315
rect 12850 1265 12865 1285
rect 12885 1265 12900 1285
rect 12850 1235 12900 1265
rect 12850 1215 12865 1235
rect 12885 1215 12900 1235
rect 12850 1185 12900 1215
rect 12850 1165 12865 1185
rect 12885 1165 12900 1185
rect 12850 1135 12900 1165
rect 12850 1115 12865 1135
rect 12885 1115 12900 1135
rect 12850 1085 12900 1115
rect 12850 1065 12865 1085
rect 12885 1065 12900 1085
rect 12850 1035 12900 1065
rect 12850 1015 12865 1035
rect 12885 1015 12900 1035
rect 12850 985 12900 1015
rect 12850 965 12865 985
rect 12885 965 12900 985
rect 12850 935 12900 965
rect 12850 915 12865 935
rect 12885 915 12900 935
rect 12850 900 12900 915
rect 13150 1585 13200 1600
rect 13150 1565 13165 1585
rect 13185 1565 13200 1585
rect 13150 1535 13200 1565
rect 13150 1515 13165 1535
rect 13185 1515 13200 1535
rect 13150 1485 13200 1515
rect 13150 1465 13165 1485
rect 13185 1465 13200 1485
rect 13150 1435 13200 1465
rect 13150 1415 13165 1435
rect 13185 1415 13200 1435
rect 13150 1385 13200 1415
rect 13150 1365 13165 1385
rect 13185 1365 13200 1385
rect 13150 1335 13200 1365
rect 13150 1315 13165 1335
rect 13185 1315 13200 1335
rect 13150 1285 13200 1315
rect 13150 1265 13165 1285
rect 13185 1265 13200 1285
rect 13150 1235 13200 1265
rect 13150 1215 13165 1235
rect 13185 1215 13200 1235
rect 13150 1185 13200 1215
rect 13150 1165 13165 1185
rect 13185 1165 13200 1185
rect 13150 1135 13200 1165
rect 13150 1115 13165 1135
rect 13185 1115 13200 1135
rect 13150 1085 13200 1115
rect 13150 1065 13165 1085
rect 13185 1065 13200 1085
rect 13150 1035 13200 1065
rect 13150 1015 13165 1035
rect 13185 1015 13200 1035
rect 13150 985 13200 1015
rect 13150 965 13165 985
rect 13185 965 13200 985
rect 13150 935 13200 965
rect 13150 915 13165 935
rect 13185 915 13200 935
rect 13150 900 13200 915
rect 13450 1585 13500 1600
rect 13450 1565 13465 1585
rect 13485 1565 13500 1585
rect 13450 1535 13500 1565
rect 13450 1515 13465 1535
rect 13485 1515 13500 1535
rect 13450 1485 13500 1515
rect 13450 1465 13465 1485
rect 13485 1465 13500 1485
rect 13450 1435 13500 1465
rect 13450 1415 13465 1435
rect 13485 1415 13500 1435
rect 13450 1385 13500 1415
rect 13450 1365 13465 1385
rect 13485 1365 13500 1385
rect 13450 1335 13500 1365
rect 13450 1315 13465 1335
rect 13485 1315 13500 1335
rect 13450 1285 13500 1315
rect 13450 1265 13465 1285
rect 13485 1265 13500 1285
rect 13450 1235 13500 1265
rect 13450 1215 13465 1235
rect 13485 1215 13500 1235
rect 13450 1185 13500 1215
rect 13450 1165 13465 1185
rect 13485 1165 13500 1185
rect 13450 1135 13500 1165
rect 13450 1115 13465 1135
rect 13485 1115 13500 1135
rect 13450 1085 13500 1115
rect 13450 1065 13465 1085
rect 13485 1065 13500 1085
rect 13450 1035 13500 1065
rect 13450 1015 13465 1035
rect 13485 1015 13500 1035
rect 13450 985 13500 1015
rect 13450 965 13465 985
rect 13485 965 13500 985
rect 13450 935 13500 965
rect 13450 915 13465 935
rect 13485 915 13500 935
rect 13450 900 13500 915
rect 13750 1585 13800 1600
rect 13750 1565 13765 1585
rect 13785 1565 13800 1585
rect 13750 1535 13800 1565
rect 13750 1515 13765 1535
rect 13785 1515 13800 1535
rect 13750 1485 13800 1515
rect 13750 1465 13765 1485
rect 13785 1465 13800 1485
rect 13750 1435 13800 1465
rect 13750 1415 13765 1435
rect 13785 1415 13800 1435
rect 13750 1385 13800 1415
rect 13750 1365 13765 1385
rect 13785 1365 13800 1385
rect 13750 1335 13800 1365
rect 13750 1315 13765 1335
rect 13785 1315 13800 1335
rect 13750 1285 13800 1315
rect 13750 1265 13765 1285
rect 13785 1265 13800 1285
rect 13750 1235 13800 1265
rect 13750 1215 13765 1235
rect 13785 1215 13800 1235
rect 13750 1185 13800 1215
rect 13750 1165 13765 1185
rect 13785 1165 13800 1185
rect 13750 1135 13800 1165
rect 13750 1115 13765 1135
rect 13785 1115 13800 1135
rect 13750 1085 13800 1115
rect 13750 1065 13765 1085
rect 13785 1065 13800 1085
rect 13750 1035 13800 1065
rect 13750 1015 13765 1035
rect 13785 1015 13800 1035
rect 13750 985 13800 1015
rect 13750 965 13765 985
rect 13785 965 13800 985
rect 13750 935 13800 965
rect 13750 915 13765 935
rect 13785 915 13800 935
rect 13750 900 13800 915
rect 14050 1585 14100 1600
rect 14050 1565 14065 1585
rect 14085 1565 14100 1585
rect 14050 1535 14100 1565
rect 14050 1515 14065 1535
rect 14085 1515 14100 1535
rect 14050 1485 14100 1515
rect 14050 1465 14065 1485
rect 14085 1465 14100 1485
rect 14050 1435 14100 1465
rect 14050 1415 14065 1435
rect 14085 1415 14100 1435
rect 14050 1385 14100 1415
rect 14050 1365 14065 1385
rect 14085 1365 14100 1385
rect 14050 1335 14100 1365
rect 14050 1315 14065 1335
rect 14085 1315 14100 1335
rect 14050 1285 14100 1315
rect 14050 1265 14065 1285
rect 14085 1265 14100 1285
rect 14050 1235 14100 1265
rect 14050 1215 14065 1235
rect 14085 1215 14100 1235
rect 14050 1185 14100 1215
rect 14050 1165 14065 1185
rect 14085 1165 14100 1185
rect 14050 1135 14100 1165
rect 14050 1115 14065 1135
rect 14085 1115 14100 1135
rect 14050 1085 14100 1115
rect 14050 1065 14065 1085
rect 14085 1065 14100 1085
rect 14050 1035 14100 1065
rect 14050 1015 14065 1035
rect 14085 1015 14100 1035
rect 14050 985 14100 1015
rect 14050 965 14065 985
rect 14085 965 14100 985
rect 14050 935 14100 965
rect 14050 915 14065 935
rect 14085 915 14100 935
rect 14050 900 14100 915
rect 14350 1585 14400 1600
rect 14350 1565 14365 1585
rect 14385 1565 14400 1585
rect 14350 1535 14400 1565
rect 14350 1515 14365 1535
rect 14385 1515 14400 1535
rect 14350 1485 14400 1515
rect 14350 1465 14365 1485
rect 14385 1465 14400 1485
rect 14350 1435 14400 1465
rect 14350 1415 14365 1435
rect 14385 1415 14400 1435
rect 14350 1385 14400 1415
rect 14350 1365 14365 1385
rect 14385 1365 14400 1385
rect 14350 1335 14400 1365
rect 14350 1315 14365 1335
rect 14385 1315 14400 1335
rect 14350 1285 14400 1315
rect 14350 1265 14365 1285
rect 14385 1265 14400 1285
rect 14350 1235 14400 1265
rect 14350 1215 14365 1235
rect 14385 1215 14400 1235
rect 14350 1185 14400 1215
rect 14350 1165 14365 1185
rect 14385 1165 14400 1185
rect 14350 1135 14400 1165
rect 14350 1115 14365 1135
rect 14385 1115 14400 1135
rect 14350 1085 14400 1115
rect 14350 1065 14365 1085
rect 14385 1065 14400 1085
rect 14350 1035 14400 1065
rect 14350 1015 14365 1035
rect 14385 1015 14400 1035
rect 14350 985 14400 1015
rect 14350 965 14365 985
rect 14385 965 14400 985
rect 14350 935 14400 965
rect 14350 915 14365 935
rect 14385 915 14400 935
rect 14350 900 14400 915
rect 15550 1585 15600 1600
rect 15550 1565 15565 1585
rect 15585 1565 15600 1585
rect 15550 1535 15600 1565
rect 15550 1515 15565 1535
rect 15585 1515 15600 1535
rect 15550 1485 15600 1515
rect 15550 1465 15565 1485
rect 15585 1465 15600 1485
rect 15550 1435 15600 1465
rect 15550 1415 15565 1435
rect 15585 1415 15600 1435
rect 15550 1385 15600 1415
rect 15550 1365 15565 1385
rect 15585 1365 15600 1385
rect 15550 1335 15600 1365
rect 15550 1315 15565 1335
rect 15585 1315 15600 1335
rect 15550 1285 15600 1315
rect 15550 1265 15565 1285
rect 15585 1265 15600 1285
rect 15550 1235 15600 1265
rect 15550 1215 15565 1235
rect 15585 1215 15600 1235
rect 15550 1185 15600 1215
rect 15550 1165 15565 1185
rect 15585 1165 15600 1185
rect 15550 1135 15600 1165
rect 15550 1115 15565 1135
rect 15585 1115 15600 1135
rect 15550 1085 15600 1115
rect 15550 1065 15565 1085
rect 15585 1065 15600 1085
rect 15550 1035 15600 1065
rect 15550 1015 15565 1035
rect 15585 1015 15600 1035
rect 15550 985 15600 1015
rect 15550 965 15565 985
rect 15585 965 15600 985
rect 15550 935 15600 965
rect 15550 915 15565 935
rect 15585 915 15600 935
rect 15550 900 15600 915
rect 16750 1585 16800 1600
rect 16750 1565 16765 1585
rect 16785 1565 16800 1585
rect 16750 1535 16800 1565
rect 16750 1515 16765 1535
rect 16785 1515 16800 1535
rect 16750 1485 16800 1515
rect 16750 1465 16765 1485
rect 16785 1465 16800 1485
rect 16750 1435 16800 1465
rect 16750 1415 16765 1435
rect 16785 1415 16800 1435
rect 16750 1385 16800 1415
rect 16750 1365 16765 1385
rect 16785 1365 16800 1385
rect 16750 1335 16800 1365
rect 16750 1315 16765 1335
rect 16785 1315 16800 1335
rect 16750 1285 16800 1315
rect 16750 1265 16765 1285
rect 16785 1265 16800 1285
rect 16750 1235 16800 1265
rect 16750 1215 16765 1235
rect 16785 1215 16800 1235
rect 16750 1185 16800 1215
rect 16750 1165 16765 1185
rect 16785 1165 16800 1185
rect 16750 1135 16800 1165
rect 16750 1115 16765 1135
rect 16785 1115 16800 1135
rect 16750 1085 16800 1115
rect 16750 1065 16765 1085
rect 16785 1065 16800 1085
rect 16750 1035 16800 1065
rect 16750 1015 16765 1035
rect 16785 1015 16800 1035
rect 16750 985 16800 1015
rect 16750 965 16765 985
rect 16785 965 16800 985
rect 16750 935 16800 965
rect 16750 915 16765 935
rect 16785 915 16800 935
rect 16750 900 16800 915
rect 17950 1585 18000 1600
rect 17950 1565 17965 1585
rect 17985 1565 18000 1585
rect 17950 1535 18000 1565
rect 17950 1515 17965 1535
rect 17985 1515 18000 1535
rect 17950 1485 18000 1515
rect 17950 1465 17965 1485
rect 17985 1465 18000 1485
rect 17950 1435 18000 1465
rect 17950 1415 17965 1435
rect 17985 1415 18000 1435
rect 17950 1385 18000 1415
rect 17950 1365 17965 1385
rect 17985 1365 18000 1385
rect 17950 1335 18000 1365
rect 17950 1315 17965 1335
rect 17985 1315 18000 1335
rect 17950 1285 18000 1315
rect 17950 1265 17965 1285
rect 17985 1265 18000 1285
rect 17950 1235 18000 1265
rect 17950 1215 17965 1235
rect 17985 1215 18000 1235
rect 17950 1185 18000 1215
rect 17950 1165 17965 1185
rect 17985 1165 18000 1185
rect 17950 1135 18000 1165
rect 17950 1115 17965 1135
rect 17985 1115 18000 1135
rect 17950 1085 18000 1115
rect 17950 1065 17965 1085
rect 17985 1065 18000 1085
rect 17950 1035 18000 1065
rect 17950 1015 17965 1035
rect 17985 1015 18000 1035
rect 17950 985 18000 1015
rect 17950 965 17965 985
rect 17985 965 18000 985
rect 17950 935 18000 965
rect 17950 915 17965 935
rect 17985 915 18000 935
rect 17950 900 18000 915
rect 19150 1585 19200 1600
rect 19150 1565 19165 1585
rect 19185 1565 19200 1585
rect 19150 1535 19200 1565
rect 19150 1515 19165 1535
rect 19185 1515 19200 1535
rect 19150 1485 19200 1515
rect 19150 1465 19165 1485
rect 19185 1465 19200 1485
rect 19150 1435 19200 1465
rect 19150 1415 19165 1435
rect 19185 1415 19200 1435
rect 19150 1385 19200 1415
rect 19150 1365 19165 1385
rect 19185 1365 19200 1385
rect 19150 1335 19200 1365
rect 19150 1315 19165 1335
rect 19185 1315 19200 1335
rect 19150 1285 19200 1315
rect 19150 1265 19165 1285
rect 19185 1265 19200 1285
rect 19150 1235 19200 1265
rect 19150 1215 19165 1235
rect 19185 1215 19200 1235
rect 19150 1185 19200 1215
rect 19150 1165 19165 1185
rect 19185 1165 19200 1185
rect 19150 1135 19200 1165
rect 19150 1115 19165 1135
rect 19185 1115 19200 1135
rect 19150 1085 19200 1115
rect 19150 1065 19165 1085
rect 19185 1065 19200 1085
rect 19150 1035 19200 1065
rect 19150 1015 19165 1035
rect 19185 1015 19200 1035
rect 19150 985 19200 1015
rect 19150 965 19165 985
rect 19185 965 19200 985
rect 19150 935 19200 965
rect 19150 915 19165 935
rect 19185 915 19200 935
rect 19150 900 19200 915
rect 20350 1585 20400 1600
rect 20350 1565 20365 1585
rect 20385 1565 20400 1585
rect 20350 1535 20400 1565
rect 20350 1515 20365 1535
rect 20385 1515 20400 1535
rect 20350 1485 20400 1515
rect 20350 1465 20365 1485
rect 20385 1465 20400 1485
rect 20350 1435 20400 1465
rect 20350 1415 20365 1435
rect 20385 1415 20400 1435
rect 20350 1385 20400 1415
rect 20350 1365 20365 1385
rect 20385 1365 20400 1385
rect 20350 1335 20400 1365
rect 20350 1315 20365 1335
rect 20385 1315 20400 1335
rect 20350 1285 20400 1315
rect 20350 1265 20365 1285
rect 20385 1265 20400 1285
rect 20350 1235 20400 1265
rect 20350 1215 20365 1235
rect 20385 1215 20400 1235
rect 20350 1185 20400 1215
rect 20350 1165 20365 1185
rect 20385 1165 20400 1185
rect 20350 1135 20400 1165
rect 20350 1115 20365 1135
rect 20385 1115 20400 1135
rect 20350 1085 20400 1115
rect 20350 1065 20365 1085
rect 20385 1065 20400 1085
rect 20350 1035 20400 1065
rect 20350 1015 20365 1035
rect 20385 1015 20400 1035
rect 20350 985 20400 1015
rect 20350 965 20365 985
rect 20385 965 20400 985
rect 20350 935 20400 965
rect 20350 915 20365 935
rect 20385 915 20400 935
rect 20350 900 20400 915
rect 21550 1585 21600 1600
rect 21550 1565 21565 1585
rect 21585 1565 21600 1585
rect 21550 1535 21600 1565
rect 21550 1515 21565 1535
rect 21585 1515 21600 1535
rect 21550 1485 21600 1515
rect 21550 1465 21565 1485
rect 21585 1465 21600 1485
rect 21550 1435 21600 1465
rect 21550 1415 21565 1435
rect 21585 1415 21600 1435
rect 21550 1385 21600 1415
rect 21550 1365 21565 1385
rect 21585 1365 21600 1385
rect 21550 1335 21600 1365
rect 21550 1315 21565 1335
rect 21585 1315 21600 1335
rect 21550 1285 21600 1315
rect 21550 1265 21565 1285
rect 21585 1265 21600 1285
rect 21550 1235 21600 1265
rect 21550 1215 21565 1235
rect 21585 1215 21600 1235
rect 21550 1185 21600 1215
rect 21550 1165 21565 1185
rect 21585 1165 21600 1185
rect 21550 1135 21600 1165
rect 21550 1115 21565 1135
rect 21585 1115 21600 1135
rect 21550 1085 21600 1115
rect 21550 1065 21565 1085
rect 21585 1065 21600 1085
rect 21550 1035 21600 1065
rect 21550 1015 21565 1035
rect 21585 1015 21600 1035
rect 21550 985 21600 1015
rect 21550 965 21565 985
rect 21585 965 21600 985
rect 21550 935 21600 965
rect 21550 915 21565 935
rect 21585 915 21600 935
rect 21550 900 21600 915
rect 22450 1585 22500 1600
rect 22450 1565 22465 1585
rect 22485 1565 22500 1585
rect 22450 1535 22500 1565
rect 22450 1515 22465 1535
rect 22485 1515 22500 1535
rect 22450 1485 22500 1515
rect 22450 1465 22465 1485
rect 22485 1465 22500 1485
rect 22450 1435 22500 1465
rect 22450 1415 22465 1435
rect 22485 1415 22500 1435
rect 22450 1385 22500 1415
rect 22450 1365 22465 1385
rect 22485 1365 22500 1385
rect 22450 1335 22500 1365
rect 22450 1315 22465 1335
rect 22485 1315 22500 1335
rect 22450 1285 22500 1315
rect 22450 1265 22465 1285
rect 22485 1265 22500 1285
rect 22450 1235 22500 1265
rect 22450 1215 22465 1235
rect 22485 1215 22500 1235
rect 22450 1185 22500 1215
rect 22450 1165 22465 1185
rect 22485 1165 22500 1185
rect 22450 1135 22500 1165
rect 22450 1115 22465 1135
rect 22485 1115 22500 1135
rect 22450 1085 22500 1115
rect 22450 1065 22465 1085
rect 22485 1065 22500 1085
rect 22450 1035 22500 1065
rect 22450 1015 22465 1035
rect 22485 1015 22500 1035
rect 22450 985 22500 1015
rect 22450 965 22465 985
rect 22485 965 22500 985
rect 22450 935 22500 965
rect 22450 915 22465 935
rect 22485 915 22500 935
rect 22450 900 22500 915
rect 23350 1585 23400 1600
rect 23350 1565 23365 1585
rect 23385 1565 23400 1585
rect 23350 1535 23400 1565
rect 23350 1515 23365 1535
rect 23385 1515 23400 1535
rect 23350 1485 23400 1515
rect 23350 1465 23365 1485
rect 23385 1465 23400 1485
rect 23350 1435 23400 1465
rect 23350 1415 23365 1435
rect 23385 1415 23400 1435
rect 23350 1385 23400 1415
rect 23350 1365 23365 1385
rect 23385 1365 23400 1385
rect 23350 1335 23400 1365
rect 23350 1315 23365 1335
rect 23385 1315 23400 1335
rect 23350 1285 23400 1315
rect 23350 1265 23365 1285
rect 23385 1265 23400 1285
rect 23350 1235 23400 1265
rect 23350 1215 23365 1235
rect 23385 1215 23400 1235
rect 23350 1185 23400 1215
rect 23350 1165 23365 1185
rect 23385 1165 23400 1185
rect 23350 1135 23400 1165
rect 23350 1115 23365 1135
rect 23385 1115 23400 1135
rect 23350 1085 23400 1115
rect 23350 1065 23365 1085
rect 23385 1065 23400 1085
rect 23350 1035 23400 1065
rect 23350 1015 23365 1035
rect 23385 1015 23400 1035
rect 23350 985 23400 1015
rect 23350 965 23365 985
rect 23385 965 23400 985
rect 23350 935 23400 965
rect 23350 915 23365 935
rect 23385 915 23400 935
rect 23350 900 23400 915
rect 24550 1585 24600 1600
rect 24550 1565 24565 1585
rect 24585 1565 24600 1585
rect 24550 1535 24600 1565
rect 24550 1515 24565 1535
rect 24585 1515 24600 1535
rect 24550 1485 24600 1515
rect 24550 1465 24565 1485
rect 24585 1465 24600 1485
rect 24550 1435 24600 1465
rect 24550 1415 24565 1435
rect 24585 1415 24600 1435
rect 24550 1385 24600 1415
rect 24550 1365 24565 1385
rect 24585 1365 24600 1385
rect 24550 1335 24600 1365
rect 24550 1315 24565 1335
rect 24585 1315 24600 1335
rect 24550 1285 24600 1315
rect 24550 1265 24565 1285
rect 24585 1265 24600 1285
rect 24550 1235 24600 1265
rect 24550 1215 24565 1235
rect 24585 1215 24600 1235
rect 24550 1185 24600 1215
rect 24550 1165 24565 1185
rect 24585 1165 24600 1185
rect 24550 1135 24600 1165
rect 24550 1115 24565 1135
rect 24585 1115 24600 1135
rect 24550 1085 24600 1115
rect 24550 1065 24565 1085
rect 24585 1065 24600 1085
rect 24550 1035 24600 1065
rect 24550 1015 24565 1035
rect 24585 1015 24600 1035
rect 24550 985 24600 1015
rect 24550 965 24565 985
rect 24585 965 24600 985
rect 24550 935 24600 965
rect 24550 915 24565 935
rect 24585 915 24600 935
rect 24550 900 24600 915
rect 25750 1585 25800 1600
rect 25750 1565 25765 1585
rect 25785 1565 25800 1585
rect 25750 1535 25800 1565
rect 25750 1515 25765 1535
rect 25785 1515 25800 1535
rect 25750 1485 25800 1515
rect 25750 1465 25765 1485
rect 25785 1465 25800 1485
rect 25750 1435 25800 1465
rect 25750 1415 25765 1435
rect 25785 1415 25800 1435
rect 25750 1385 25800 1415
rect 25750 1365 25765 1385
rect 25785 1365 25800 1385
rect 25750 1335 25800 1365
rect 25750 1315 25765 1335
rect 25785 1315 25800 1335
rect 25750 1285 25800 1315
rect 25750 1265 25765 1285
rect 25785 1265 25800 1285
rect 25750 1235 25800 1265
rect 25750 1215 25765 1235
rect 25785 1215 25800 1235
rect 25750 1185 25800 1215
rect 25750 1165 25765 1185
rect 25785 1165 25800 1185
rect 25750 1135 25800 1165
rect 25750 1115 25765 1135
rect 25785 1115 25800 1135
rect 25750 1085 25800 1115
rect 25750 1065 25765 1085
rect 25785 1065 25800 1085
rect 25750 1035 25800 1065
rect 25750 1015 25765 1035
rect 25785 1015 25800 1035
rect 25750 985 25800 1015
rect 25750 965 25765 985
rect 25785 965 25800 985
rect 25750 935 25800 965
rect 25750 915 25765 935
rect 25785 915 25800 935
rect 25750 900 25800 915
rect 26650 1585 26700 1600
rect 26650 1565 26665 1585
rect 26685 1565 26700 1585
rect 26650 1535 26700 1565
rect 26650 1515 26665 1535
rect 26685 1515 26700 1535
rect 26650 1485 26700 1515
rect 26650 1465 26665 1485
rect 26685 1465 26700 1485
rect 26650 1435 26700 1465
rect 26650 1415 26665 1435
rect 26685 1415 26700 1435
rect 26650 1385 26700 1415
rect 26650 1365 26665 1385
rect 26685 1365 26700 1385
rect 26650 1335 26700 1365
rect 26650 1315 26665 1335
rect 26685 1315 26700 1335
rect 26650 1285 26700 1315
rect 26650 1265 26665 1285
rect 26685 1265 26700 1285
rect 26650 1235 26700 1265
rect 26650 1215 26665 1235
rect 26685 1215 26700 1235
rect 26650 1185 26700 1215
rect 26650 1165 26665 1185
rect 26685 1165 26700 1185
rect 26650 1135 26700 1165
rect 26650 1115 26665 1135
rect 26685 1115 26700 1135
rect 26650 1085 26700 1115
rect 26650 1065 26665 1085
rect 26685 1065 26700 1085
rect 26650 1035 26700 1065
rect 26650 1015 26665 1035
rect 26685 1015 26700 1035
rect 26650 985 26700 1015
rect 26650 965 26665 985
rect 26685 965 26700 985
rect 26650 935 26700 965
rect 26650 915 26665 935
rect 26685 915 26700 935
rect 26650 900 26700 915
rect 27550 1585 27600 1600
rect 27550 1565 27565 1585
rect 27585 1565 27600 1585
rect 27550 1535 27600 1565
rect 27550 1515 27565 1535
rect 27585 1515 27600 1535
rect 27550 1485 27600 1515
rect 27550 1465 27565 1485
rect 27585 1465 27600 1485
rect 27550 1435 27600 1465
rect 27550 1415 27565 1435
rect 27585 1415 27600 1435
rect 27550 1385 27600 1415
rect 27550 1365 27565 1385
rect 27585 1365 27600 1385
rect 27550 1335 27600 1365
rect 27550 1315 27565 1335
rect 27585 1315 27600 1335
rect 27550 1285 27600 1315
rect 27550 1265 27565 1285
rect 27585 1265 27600 1285
rect 27550 1235 27600 1265
rect 27550 1215 27565 1235
rect 27585 1215 27600 1235
rect 27550 1185 27600 1215
rect 27550 1165 27565 1185
rect 27585 1165 27600 1185
rect 27550 1135 27600 1165
rect 27550 1115 27565 1135
rect 27585 1115 27600 1135
rect 27550 1085 27600 1115
rect 27550 1065 27565 1085
rect 27585 1065 27600 1085
rect 27550 1035 27600 1065
rect 27550 1015 27565 1035
rect 27585 1015 27600 1035
rect 27550 985 27600 1015
rect 27550 965 27565 985
rect 27585 965 27600 985
rect 27550 935 27600 965
rect 27550 915 27565 935
rect 27585 915 27600 935
rect 27550 900 27600 915
rect 28750 1585 28800 1600
rect 28750 1565 28765 1585
rect 28785 1565 28800 1585
rect 28750 1535 28800 1565
rect 28750 1515 28765 1535
rect 28785 1515 28800 1535
rect 28750 1485 28800 1515
rect 28750 1465 28765 1485
rect 28785 1465 28800 1485
rect 28750 1435 28800 1465
rect 28750 1415 28765 1435
rect 28785 1415 28800 1435
rect 28750 1385 28800 1415
rect 28750 1365 28765 1385
rect 28785 1365 28800 1385
rect 28750 1335 28800 1365
rect 28750 1315 28765 1335
rect 28785 1315 28800 1335
rect 28750 1285 28800 1315
rect 28750 1265 28765 1285
rect 28785 1265 28800 1285
rect 28750 1235 28800 1265
rect 28750 1215 28765 1235
rect 28785 1215 28800 1235
rect 28750 1185 28800 1215
rect 28750 1165 28765 1185
rect 28785 1165 28800 1185
rect 28750 1135 28800 1165
rect 28750 1115 28765 1135
rect 28785 1115 28800 1135
rect 28750 1085 28800 1115
rect 28750 1065 28765 1085
rect 28785 1065 28800 1085
rect 28750 1035 28800 1065
rect 28750 1015 28765 1035
rect 28785 1015 28800 1035
rect 28750 985 28800 1015
rect 28750 965 28765 985
rect 28785 965 28800 985
rect 28750 935 28800 965
rect 28750 915 28765 935
rect 28785 915 28800 935
rect 28750 900 28800 915
rect -600 835 -350 850
rect -600 815 -585 835
rect -565 815 -535 835
rect -515 815 -485 835
rect -465 815 -435 835
rect -415 815 -385 835
rect -365 815 -350 835
rect -600 800 -350 815
rect -300 835 -50 850
rect -300 815 -285 835
rect -265 815 -235 835
rect -215 815 -185 835
rect -165 815 -135 835
rect -115 815 -85 835
rect -65 815 -50 835
rect -300 800 -50 815
rect 0 835 250 850
rect 0 815 15 835
rect 35 815 65 835
rect 85 815 115 835
rect 135 815 165 835
rect 185 815 215 835
rect 235 815 250 835
rect 0 800 250 815
rect 300 835 550 850
rect 300 815 315 835
rect 335 815 365 835
rect 385 815 415 835
rect 435 815 465 835
rect 485 815 515 835
rect 535 815 550 835
rect 300 800 550 815
rect 600 835 850 850
rect 600 815 615 835
rect 635 815 665 835
rect 685 815 715 835
rect 735 815 765 835
rect 785 815 815 835
rect 835 815 850 835
rect 600 800 850 815
rect 900 835 1150 850
rect 900 815 915 835
rect 935 815 965 835
rect 985 815 1015 835
rect 1035 815 1065 835
rect 1085 815 1115 835
rect 1135 815 1150 835
rect 900 800 1150 815
rect 1200 835 1450 850
rect 1200 815 1215 835
rect 1235 815 1265 835
rect 1285 815 1315 835
rect 1335 815 1365 835
rect 1385 815 1415 835
rect 1435 815 1450 835
rect 1200 800 1450 815
rect 1500 835 1750 850
rect 1500 815 1515 835
rect 1535 815 1565 835
rect 1585 815 1615 835
rect 1635 815 1665 835
rect 1685 815 1715 835
rect 1735 815 1750 835
rect 1500 800 1750 815
rect 1800 835 2050 850
rect 1800 815 1815 835
rect 1835 815 1865 835
rect 1885 815 1915 835
rect 1935 815 1965 835
rect 1985 815 2015 835
rect 2035 815 2050 835
rect 1800 800 2050 815
rect 2100 835 2350 850
rect 2100 815 2115 835
rect 2135 815 2165 835
rect 2185 815 2215 835
rect 2235 815 2265 835
rect 2285 815 2315 835
rect 2335 815 2350 835
rect 2100 800 2350 815
rect 2400 835 2650 850
rect 2400 815 2415 835
rect 2435 815 2465 835
rect 2485 815 2515 835
rect 2535 815 2565 835
rect 2585 815 2615 835
rect 2635 815 2650 835
rect 2400 800 2650 815
rect 2700 835 2950 850
rect 2700 815 2715 835
rect 2735 815 2765 835
rect 2785 815 2815 835
rect 2835 815 2865 835
rect 2885 815 2915 835
rect 2935 815 2950 835
rect 2700 800 2950 815
rect 3000 835 3250 850
rect 3000 815 3015 835
rect 3035 815 3065 835
rect 3085 815 3115 835
rect 3135 815 3165 835
rect 3185 815 3215 835
rect 3235 815 3250 835
rect 3000 800 3250 815
rect 3300 835 3550 850
rect 3300 815 3315 835
rect 3335 815 3365 835
rect 3385 815 3415 835
rect 3435 815 3465 835
rect 3485 815 3515 835
rect 3535 815 3550 835
rect 3300 800 3550 815
rect 3600 835 3850 850
rect 3600 815 3615 835
rect 3635 815 3665 835
rect 3685 815 3715 835
rect 3735 815 3765 835
rect 3785 815 3815 835
rect 3835 815 3850 835
rect 3600 800 3850 815
rect 3900 835 4150 850
rect 3900 815 3915 835
rect 3935 815 3965 835
rect 3985 815 4015 835
rect 4035 815 4065 835
rect 4085 815 4115 835
rect 4135 815 4150 835
rect 3900 800 4150 815
rect 4200 835 4450 850
rect 4200 815 4215 835
rect 4235 815 4265 835
rect 4285 815 4315 835
rect 4335 815 4365 835
rect 4385 815 4415 835
rect 4435 815 4450 835
rect 4200 800 4450 815
rect 4500 835 4750 850
rect 4500 815 4515 835
rect 4535 815 4565 835
rect 4585 815 4615 835
rect 4635 815 4665 835
rect 4685 815 4715 835
rect 4735 815 4750 835
rect 4500 800 4750 815
rect 4800 835 5050 850
rect 4800 815 4815 835
rect 4835 815 4865 835
rect 4885 815 4915 835
rect 4935 815 4965 835
rect 4985 815 5015 835
rect 5035 815 5050 835
rect 4800 800 5050 815
rect 5100 835 5350 850
rect 5100 815 5115 835
rect 5135 815 5165 835
rect 5185 815 5215 835
rect 5235 815 5265 835
rect 5285 815 5315 835
rect 5335 815 5350 835
rect 5100 800 5350 815
rect 5400 835 5650 850
rect 5400 815 5415 835
rect 5435 815 5465 835
rect 5485 815 5515 835
rect 5535 815 5565 835
rect 5585 815 5615 835
rect 5635 815 5650 835
rect 5400 800 5650 815
rect 5700 835 5950 850
rect 5700 815 5715 835
rect 5735 815 5765 835
rect 5785 815 5815 835
rect 5835 815 5865 835
rect 5885 815 5915 835
rect 5935 815 5950 835
rect 5700 800 5950 815
rect 6000 835 6250 850
rect 6000 815 6015 835
rect 6035 815 6065 835
rect 6085 815 6115 835
rect 6135 815 6165 835
rect 6185 815 6215 835
rect 6235 815 6250 835
rect 6000 800 6250 815
rect 6300 835 6550 850
rect 6300 815 6315 835
rect 6335 815 6365 835
rect 6385 815 6415 835
rect 6435 815 6465 835
rect 6485 815 6515 835
rect 6535 815 6550 835
rect 6300 800 6550 815
rect 6600 835 6850 850
rect 6600 815 6615 835
rect 6635 815 6665 835
rect 6685 815 6715 835
rect 6735 815 6765 835
rect 6785 815 6815 835
rect 6835 815 6850 835
rect 6600 800 6850 815
rect 6900 835 7150 850
rect 6900 815 6915 835
rect 6935 815 6965 835
rect 6985 815 7015 835
rect 7035 815 7065 835
rect 7085 815 7115 835
rect 7135 815 7150 835
rect 6900 800 7150 815
rect 7200 835 7450 850
rect 7200 815 7215 835
rect 7235 815 7265 835
rect 7285 815 7315 835
rect 7335 815 7365 835
rect 7385 815 7415 835
rect 7435 815 7450 835
rect 7200 800 7450 815
rect 7500 835 7750 850
rect 7500 815 7515 835
rect 7535 815 7565 835
rect 7585 815 7615 835
rect 7635 815 7665 835
rect 7685 815 7715 835
rect 7735 815 7750 835
rect 7500 800 7750 815
rect 7800 835 8050 850
rect 7800 815 7815 835
rect 7835 815 7865 835
rect 7885 815 7915 835
rect 7935 815 7965 835
rect 7985 815 8015 835
rect 8035 815 8050 835
rect 7800 800 8050 815
rect 8100 835 8350 850
rect 8100 815 8115 835
rect 8135 815 8165 835
rect 8185 815 8215 835
rect 8235 815 8265 835
rect 8285 815 8315 835
rect 8335 815 8350 835
rect 8100 800 8350 815
rect 8400 835 8650 850
rect 8400 815 8415 835
rect 8435 815 8465 835
rect 8485 815 8515 835
rect 8535 815 8565 835
rect 8585 815 8615 835
rect 8635 815 8650 835
rect 8400 800 8650 815
rect 8700 835 8950 850
rect 8700 815 8715 835
rect 8735 815 8765 835
rect 8785 815 8815 835
rect 8835 815 8865 835
rect 8885 815 8915 835
rect 8935 815 8950 835
rect 8700 800 8950 815
rect 9000 835 9250 850
rect 9000 815 9015 835
rect 9035 815 9065 835
rect 9085 815 9115 835
rect 9135 815 9165 835
rect 9185 815 9215 835
rect 9235 815 9250 835
rect 9000 800 9250 815
rect 9300 835 9550 850
rect 9300 815 9315 835
rect 9335 815 9365 835
rect 9385 815 9415 835
rect 9435 815 9465 835
rect 9485 815 9515 835
rect 9535 815 9550 835
rect 9300 800 9550 815
rect 9600 835 9850 850
rect 9600 815 9615 835
rect 9635 815 9665 835
rect 9685 815 9715 835
rect 9735 815 9765 835
rect 9785 815 9815 835
rect 9835 815 9850 835
rect 9600 800 9850 815
rect 9900 835 10150 850
rect 9900 815 9915 835
rect 9935 815 9965 835
rect 9985 815 10015 835
rect 10035 815 10065 835
rect 10085 815 10115 835
rect 10135 815 10150 835
rect 9900 800 10150 815
rect 10200 835 10450 850
rect 10200 815 10215 835
rect 10235 815 10265 835
rect 10285 815 10315 835
rect 10335 815 10365 835
rect 10385 815 10415 835
rect 10435 815 10450 835
rect 10200 800 10450 815
rect 10500 835 10750 850
rect 10500 815 10515 835
rect 10535 815 10565 835
rect 10585 815 10615 835
rect 10635 815 10665 835
rect 10685 815 10715 835
rect 10735 815 10750 835
rect 10500 800 10750 815
rect 10800 835 11050 850
rect 10800 815 10815 835
rect 10835 815 10865 835
rect 10885 815 10915 835
rect 10935 815 10965 835
rect 10985 815 11015 835
rect 11035 815 11050 835
rect 10800 800 11050 815
rect 11100 835 11350 850
rect 11100 815 11115 835
rect 11135 815 11165 835
rect 11185 815 11215 835
rect 11235 815 11265 835
rect 11285 815 11315 835
rect 11335 815 11350 835
rect 11100 800 11350 815
rect 11400 835 11650 850
rect 11400 815 11415 835
rect 11435 815 11465 835
rect 11485 815 11515 835
rect 11535 815 11565 835
rect 11585 815 11615 835
rect 11635 815 11650 835
rect 11400 800 11650 815
rect 11700 835 11950 850
rect 11700 815 11715 835
rect 11735 815 11765 835
rect 11785 815 11815 835
rect 11835 815 11865 835
rect 11885 815 11915 835
rect 11935 815 11950 835
rect 11700 800 11950 815
rect 12000 835 12250 850
rect 12000 815 12015 835
rect 12035 815 12065 835
rect 12085 815 12115 835
rect 12135 815 12165 835
rect 12185 815 12215 835
rect 12235 815 12250 835
rect 12000 800 12250 815
rect 12300 835 12550 850
rect 12300 815 12315 835
rect 12335 815 12365 835
rect 12385 815 12415 835
rect 12435 815 12465 835
rect 12485 815 12515 835
rect 12535 815 12550 835
rect 12300 800 12550 815
rect 12600 835 12850 850
rect 12600 815 12615 835
rect 12635 815 12665 835
rect 12685 815 12715 835
rect 12735 815 12765 835
rect 12785 815 12815 835
rect 12835 815 12850 835
rect 12600 800 12850 815
rect 12900 835 13150 850
rect 12900 815 12915 835
rect 12935 815 12965 835
rect 12985 815 13015 835
rect 13035 815 13065 835
rect 13085 815 13115 835
rect 13135 815 13150 835
rect 12900 800 13150 815
rect 13200 835 13450 850
rect 13200 815 13215 835
rect 13235 815 13265 835
rect 13285 815 13315 835
rect 13335 815 13365 835
rect 13385 815 13415 835
rect 13435 815 13450 835
rect 13200 800 13450 815
rect 13500 835 13750 850
rect 13500 815 13515 835
rect 13535 815 13565 835
rect 13585 815 13615 835
rect 13635 815 13665 835
rect 13685 815 13715 835
rect 13735 815 13750 835
rect 13500 800 13750 815
rect 13800 835 14050 850
rect 13800 815 13815 835
rect 13835 815 13865 835
rect 13885 815 13915 835
rect 13935 815 13965 835
rect 13985 815 14015 835
rect 14035 815 14050 835
rect 13800 800 14050 815
rect 14100 835 14350 850
rect 14100 815 14115 835
rect 14135 815 14165 835
rect 14185 815 14215 835
rect 14235 815 14265 835
rect 14285 815 14315 835
rect 14335 815 14350 835
rect 14100 800 14350 815
rect 14400 835 14650 850
rect 14400 815 14415 835
rect 14435 815 14465 835
rect 14485 815 14515 835
rect 14535 815 14565 835
rect 14585 815 14615 835
rect 14635 815 14650 835
rect 14400 800 14650 815
rect 14700 835 14950 850
rect 14700 815 14715 835
rect 14735 815 14765 835
rect 14785 815 14815 835
rect 14835 815 14865 835
rect 14885 815 14915 835
rect 14935 815 14950 835
rect 14700 800 14950 815
rect 15000 835 15250 850
rect 15000 815 15015 835
rect 15035 815 15065 835
rect 15085 815 15115 835
rect 15135 815 15165 835
rect 15185 815 15215 835
rect 15235 815 15250 835
rect 15000 800 15250 815
rect 15300 835 15550 850
rect 15300 815 15315 835
rect 15335 815 15365 835
rect 15385 815 15415 835
rect 15435 815 15465 835
rect 15485 815 15515 835
rect 15535 815 15550 835
rect 15300 800 15550 815
rect 15600 835 15850 850
rect 15600 815 15615 835
rect 15635 815 15665 835
rect 15685 815 15715 835
rect 15735 815 15765 835
rect 15785 815 15815 835
rect 15835 815 15850 835
rect 15600 800 15850 815
rect 15900 835 16150 850
rect 15900 815 15915 835
rect 15935 815 15965 835
rect 15985 815 16015 835
rect 16035 815 16065 835
rect 16085 815 16115 835
rect 16135 815 16150 835
rect 15900 800 16150 815
rect 16200 835 16450 850
rect 16200 815 16215 835
rect 16235 815 16265 835
rect 16285 815 16315 835
rect 16335 815 16365 835
rect 16385 815 16415 835
rect 16435 815 16450 835
rect 16200 800 16450 815
rect 16500 835 16750 850
rect 16500 815 16515 835
rect 16535 815 16565 835
rect 16585 815 16615 835
rect 16635 815 16665 835
rect 16685 815 16715 835
rect 16735 815 16750 835
rect 16500 800 16750 815
rect 16800 835 17050 850
rect 16800 815 16815 835
rect 16835 815 16865 835
rect 16885 815 16915 835
rect 16935 815 16965 835
rect 16985 815 17015 835
rect 17035 815 17050 835
rect 16800 800 17050 815
rect 17100 835 17350 850
rect 17100 815 17115 835
rect 17135 815 17165 835
rect 17185 815 17215 835
rect 17235 815 17265 835
rect 17285 815 17315 835
rect 17335 815 17350 835
rect 17100 800 17350 815
rect 17400 835 17650 850
rect 17400 815 17415 835
rect 17435 815 17465 835
rect 17485 815 17515 835
rect 17535 815 17565 835
rect 17585 815 17615 835
rect 17635 815 17650 835
rect 17400 800 17650 815
rect 17700 835 17950 850
rect 17700 815 17715 835
rect 17735 815 17765 835
rect 17785 815 17815 835
rect 17835 815 17865 835
rect 17885 815 17915 835
rect 17935 815 17950 835
rect 17700 800 17950 815
rect 18000 835 18250 850
rect 18000 815 18015 835
rect 18035 815 18065 835
rect 18085 815 18115 835
rect 18135 815 18165 835
rect 18185 815 18215 835
rect 18235 815 18250 835
rect 18000 800 18250 815
rect 18300 835 18550 850
rect 18300 815 18315 835
rect 18335 815 18365 835
rect 18385 815 18415 835
rect 18435 815 18465 835
rect 18485 815 18515 835
rect 18535 815 18550 835
rect 18300 800 18550 815
rect 18600 835 18850 850
rect 18600 815 18615 835
rect 18635 815 18665 835
rect 18685 815 18715 835
rect 18735 815 18765 835
rect 18785 815 18815 835
rect 18835 815 18850 835
rect 18600 800 18850 815
rect 18900 835 19150 850
rect 18900 815 18915 835
rect 18935 815 18965 835
rect 18985 815 19015 835
rect 19035 815 19065 835
rect 19085 815 19115 835
rect 19135 815 19150 835
rect 18900 800 19150 815
rect 19200 835 19450 850
rect 19200 815 19215 835
rect 19235 815 19265 835
rect 19285 815 19315 835
rect 19335 815 19365 835
rect 19385 815 19415 835
rect 19435 815 19450 835
rect 19200 800 19450 815
rect 19500 835 19750 850
rect 19500 815 19515 835
rect 19535 815 19565 835
rect 19585 815 19615 835
rect 19635 815 19665 835
rect 19685 815 19715 835
rect 19735 815 19750 835
rect 19500 800 19750 815
rect 19800 835 20050 850
rect 19800 815 19815 835
rect 19835 815 19865 835
rect 19885 815 19915 835
rect 19935 815 19965 835
rect 19985 815 20015 835
rect 20035 815 20050 835
rect 19800 800 20050 815
rect 20100 835 20350 850
rect 20100 815 20115 835
rect 20135 815 20165 835
rect 20185 815 20215 835
rect 20235 815 20265 835
rect 20285 815 20315 835
rect 20335 815 20350 835
rect 20100 800 20350 815
rect 20400 835 20650 850
rect 20400 815 20415 835
rect 20435 815 20465 835
rect 20485 815 20515 835
rect 20535 815 20565 835
rect 20585 815 20615 835
rect 20635 815 20650 835
rect 20400 800 20650 815
rect 20700 835 20950 850
rect 20700 815 20715 835
rect 20735 815 20765 835
rect 20785 815 20815 835
rect 20835 815 20865 835
rect 20885 815 20915 835
rect 20935 815 20950 835
rect 20700 800 20950 815
rect 21000 835 21250 850
rect 21000 815 21015 835
rect 21035 815 21065 835
rect 21085 815 21115 835
rect 21135 815 21165 835
rect 21185 815 21215 835
rect 21235 815 21250 835
rect 21000 800 21250 815
rect 21300 835 21550 850
rect 21300 815 21315 835
rect 21335 815 21365 835
rect 21385 815 21415 835
rect 21435 815 21465 835
rect 21485 815 21515 835
rect 21535 815 21550 835
rect 21300 800 21550 815
rect 21600 835 21850 850
rect 21600 815 21615 835
rect 21635 815 21665 835
rect 21685 815 21715 835
rect 21735 815 21765 835
rect 21785 815 21815 835
rect 21835 815 21850 835
rect 21600 800 21850 815
rect 21900 835 22150 850
rect 21900 815 21915 835
rect 21935 815 21965 835
rect 21985 815 22015 835
rect 22035 815 22065 835
rect 22085 815 22115 835
rect 22135 815 22150 835
rect 21900 800 22150 815
rect 22200 835 22450 850
rect 22200 815 22215 835
rect 22235 815 22265 835
rect 22285 815 22315 835
rect 22335 815 22365 835
rect 22385 815 22415 835
rect 22435 815 22450 835
rect 22200 800 22450 815
rect 22500 835 22750 850
rect 22500 815 22515 835
rect 22535 815 22565 835
rect 22585 815 22615 835
rect 22635 815 22665 835
rect 22685 815 22715 835
rect 22735 815 22750 835
rect 22500 800 22750 815
rect 22800 835 23050 850
rect 22800 815 22815 835
rect 22835 815 22865 835
rect 22885 815 22915 835
rect 22935 815 22965 835
rect 22985 815 23015 835
rect 23035 815 23050 835
rect 22800 800 23050 815
rect 23100 835 23350 850
rect 23100 815 23115 835
rect 23135 815 23165 835
rect 23185 815 23215 835
rect 23235 815 23265 835
rect 23285 815 23315 835
rect 23335 815 23350 835
rect 23100 800 23350 815
rect 23400 835 23650 850
rect 23400 815 23415 835
rect 23435 815 23465 835
rect 23485 815 23515 835
rect 23535 815 23565 835
rect 23585 815 23615 835
rect 23635 815 23650 835
rect 23400 800 23650 815
rect 23700 835 23950 850
rect 23700 815 23715 835
rect 23735 815 23765 835
rect 23785 815 23815 835
rect 23835 815 23865 835
rect 23885 815 23915 835
rect 23935 815 23950 835
rect 23700 800 23950 815
rect 24000 835 24250 850
rect 24000 815 24015 835
rect 24035 815 24065 835
rect 24085 815 24115 835
rect 24135 815 24165 835
rect 24185 815 24215 835
rect 24235 815 24250 835
rect 24000 800 24250 815
rect 24300 835 24550 850
rect 24300 815 24315 835
rect 24335 815 24365 835
rect 24385 815 24415 835
rect 24435 815 24465 835
rect 24485 815 24515 835
rect 24535 815 24550 835
rect 24300 800 24550 815
rect 24600 835 24850 850
rect 24600 815 24615 835
rect 24635 815 24665 835
rect 24685 815 24715 835
rect 24735 815 24765 835
rect 24785 815 24815 835
rect 24835 815 24850 835
rect 24600 800 24850 815
rect 24900 835 25150 850
rect 24900 815 24915 835
rect 24935 815 24965 835
rect 24985 815 25015 835
rect 25035 815 25065 835
rect 25085 815 25115 835
rect 25135 815 25150 835
rect 24900 800 25150 815
rect 25200 835 25450 850
rect 25200 815 25215 835
rect 25235 815 25265 835
rect 25285 815 25315 835
rect 25335 815 25365 835
rect 25385 815 25415 835
rect 25435 815 25450 835
rect 25200 800 25450 815
rect 25500 835 25750 850
rect 25500 815 25515 835
rect 25535 815 25565 835
rect 25585 815 25615 835
rect 25635 815 25665 835
rect 25685 815 25715 835
rect 25735 815 25750 835
rect 25500 800 25750 815
rect 25800 835 26050 850
rect 25800 815 25815 835
rect 25835 815 25865 835
rect 25885 815 25915 835
rect 25935 815 25965 835
rect 25985 815 26015 835
rect 26035 815 26050 835
rect 25800 800 26050 815
rect 26100 835 26350 850
rect 26100 815 26115 835
rect 26135 815 26165 835
rect 26185 815 26215 835
rect 26235 815 26265 835
rect 26285 815 26315 835
rect 26335 815 26350 835
rect 26100 800 26350 815
rect 26400 835 26650 850
rect 26400 815 26415 835
rect 26435 815 26465 835
rect 26485 815 26515 835
rect 26535 815 26565 835
rect 26585 815 26615 835
rect 26635 815 26650 835
rect 26400 800 26650 815
rect 26700 835 26950 850
rect 26700 815 26715 835
rect 26735 815 26765 835
rect 26785 815 26815 835
rect 26835 815 26865 835
rect 26885 815 26915 835
rect 26935 815 26950 835
rect 26700 800 26950 815
rect 27000 835 27250 850
rect 27000 815 27015 835
rect 27035 815 27065 835
rect 27085 815 27115 835
rect 27135 815 27165 835
rect 27185 815 27215 835
rect 27235 815 27250 835
rect 27000 800 27250 815
rect 27300 835 27550 850
rect 27300 815 27315 835
rect 27335 815 27365 835
rect 27385 815 27415 835
rect 27435 815 27465 835
rect 27485 815 27515 835
rect 27535 815 27550 835
rect 27300 800 27550 815
rect 27600 835 27850 850
rect 27600 815 27615 835
rect 27635 815 27665 835
rect 27685 815 27715 835
rect 27735 815 27765 835
rect 27785 815 27815 835
rect 27835 815 27850 835
rect 27600 800 27850 815
rect 27900 835 28150 850
rect 27900 815 27915 835
rect 27935 815 27965 835
rect 27985 815 28015 835
rect 28035 815 28065 835
rect 28085 815 28115 835
rect 28135 815 28150 835
rect 27900 800 28150 815
rect 28200 835 28450 850
rect 28200 815 28215 835
rect 28235 815 28265 835
rect 28285 815 28315 835
rect 28335 815 28365 835
rect 28385 815 28415 835
rect 28435 815 28450 835
rect 28200 800 28450 815
rect 28500 835 28750 850
rect 28500 815 28515 835
rect 28535 815 28565 835
rect 28585 815 28615 835
rect 28635 815 28665 835
rect 28685 815 28715 835
rect 28735 815 28750 835
rect 28500 800 28750 815
rect -650 735 -600 750
rect -650 715 -635 735
rect -615 715 -600 735
rect -650 685 -600 715
rect -650 665 -635 685
rect -615 665 -600 685
rect -650 635 -600 665
rect -650 615 -635 635
rect -615 615 -600 635
rect -650 585 -600 615
rect -650 565 -635 585
rect -615 565 -600 585
rect -650 535 -600 565
rect -650 515 -635 535
rect -615 515 -600 535
rect -650 485 -600 515
rect -650 465 -635 485
rect -615 465 -600 485
rect -650 435 -600 465
rect -650 415 -635 435
rect -615 415 -600 435
rect -650 385 -600 415
rect -650 365 -635 385
rect -615 365 -600 385
rect -650 335 -600 365
rect -650 315 -635 335
rect -615 315 -600 335
rect -650 285 -600 315
rect -650 265 -635 285
rect -615 265 -600 285
rect -650 235 -600 265
rect -650 215 -635 235
rect -615 215 -600 235
rect -650 185 -600 215
rect -650 165 -635 185
rect -615 165 -600 185
rect -650 135 -600 165
rect -650 115 -635 135
rect -615 115 -600 135
rect -650 85 -600 115
rect -650 65 -635 85
rect -615 65 -600 85
rect -650 50 -600 65
rect -500 735 -450 750
rect -500 715 -485 735
rect -465 715 -450 735
rect -500 685 -450 715
rect -500 665 -485 685
rect -465 665 -450 685
rect -500 635 -450 665
rect -500 615 -485 635
rect -465 615 -450 635
rect -500 585 -450 615
rect -500 565 -485 585
rect -465 565 -450 585
rect -500 535 -450 565
rect -500 515 -485 535
rect -465 515 -450 535
rect -500 485 -450 515
rect -500 465 -485 485
rect -465 465 -450 485
rect -500 435 -450 465
rect -500 415 -485 435
rect -465 415 -450 435
rect -500 385 -450 415
rect -500 365 -485 385
rect -465 365 -450 385
rect -500 335 -450 365
rect -500 315 -485 335
rect -465 315 -450 335
rect -500 285 -450 315
rect -500 265 -485 285
rect -465 265 -450 285
rect -500 235 -450 265
rect -500 215 -485 235
rect -465 215 -450 235
rect -500 185 -450 215
rect -500 165 -485 185
rect -465 165 -450 185
rect -500 135 -450 165
rect -500 115 -485 135
rect -465 115 -450 135
rect -500 85 -450 115
rect -500 65 -485 85
rect -465 65 -450 85
rect -500 50 -450 65
rect -350 735 -300 750
rect -350 715 -335 735
rect -315 715 -300 735
rect -350 685 -300 715
rect -350 665 -335 685
rect -315 665 -300 685
rect -350 635 -300 665
rect -350 615 -335 635
rect -315 615 -300 635
rect -350 585 -300 615
rect -350 565 -335 585
rect -315 565 -300 585
rect -350 535 -300 565
rect -350 515 -335 535
rect -315 515 -300 535
rect -350 485 -300 515
rect -350 465 -335 485
rect -315 465 -300 485
rect -350 435 -300 465
rect -350 415 -335 435
rect -315 415 -300 435
rect -350 385 -300 415
rect -350 365 -335 385
rect -315 365 -300 385
rect -350 335 -300 365
rect -350 315 -335 335
rect -315 315 -300 335
rect -350 285 -300 315
rect -350 265 -335 285
rect -315 265 -300 285
rect -350 235 -300 265
rect -350 215 -335 235
rect -315 215 -300 235
rect -350 185 -300 215
rect -350 165 -335 185
rect -315 165 -300 185
rect -350 135 -300 165
rect -350 115 -335 135
rect -315 115 -300 135
rect -350 85 -300 115
rect -350 65 -335 85
rect -315 65 -300 85
rect -350 50 -300 65
rect -200 735 -150 750
rect -200 715 -185 735
rect -165 715 -150 735
rect -200 685 -150 715
rect -200 665 -185 685
rect -165 665 -150 685
rect -200 635 -150 665
rect -200 615 -185 635
rect -165 615 -150 635
rect -200 585 -150 615
rect -200 565 -185 585
rect -165 565 -150 585
rect -200 535 -150 565
rect -200 515 -185 535
rect -165 515 -150 535
rect -200 485 -150 515
rect -200 465 -185 485
rect -165 465 -150 485
rect -200 435 -150 465
rect -200 415 -185 435
rect -165 415 -150 435
rect -200 385 -150 415
rect -200 365 -185 385
rect -165 365 -150 385
rect -200 335 -150 365
rect -200 315 -185 335
rect -165 315 -150 335
rect -200 285 -150 315
rect -200 265 -185 285
rect -165 265 -150 285
rect -200 235 -150 265
rect -200 215 -185 235
rect -165 215 -150 235
rect -200 185 -150 215
rect -200 165 -185 185
rect -165 165 -150 185
rect -200 135 -150 165
rect -200 115 -185 135
rect -165 115 -150 135
rect -200 85 -150 115
rect -200 65 -185 85
rect -165 65 -150 85
rect -200 50 -150 65
rect -50 735 0 750
rect -50 715 -35 735
rect -15 715 0 735
rect -50 685 0 715
rect -50 665 -35 685
rect -15 665 0 685
rect -50 635 0 665
rect -50 615 -35 635
rect -15 615 0 635
rect -50 585 0 615
rect -50 565 -35 585
rect -15 565 0 585
rect -50 535 0 565
rect -50 515 -35 535
rect -15 515 0 535
rect -50 485 0 515
rect -50 465 -35 485
rect -15 465 0 485
rect -50 435 0 465
rect -50 415 -35 435
rect -15 415 0 435
rect -50 385 0 415
rect -50 365 -35 385
rect -15 365 0 385
rect -50 335 0 365
rect -50 315 -35 335
rect -15 315 0 335
rect -50 285 0 315
rect -50 265 -35 285
rect -15 265 0 285
rect -50 235 0 265
rect -50 215 -35 235
rect -15 215 0 235
rect -50 185 0 215
rect -50 165 -35 185
rect -15 165 0 185
rect -50 135 0 165
rect -50 115 -35 135
rect -15 115 0 135
rect -50 85 0 115
rect -50 65 -35 85
rect -15 65 0 85
rect -50 50 0 65
rect 1150 735 1200 750
rect 1150 715 1165 735
rect 1185 715 1200 735
rect 1150 685 1200 715
rect 1150 665 1165 685
rect 1185 665 1200 685
rect 1150 635 1200 665
rect 1150 615 1165 635
rect 1185 615 1200 635
rect 1150 585 1200 615
rect 1150 565 1165 585
rect 1185 565 1200 585
rect 1150 535 1200 565
rect 1150 515 1165 535
rect 1185 515 1200 535
rect 1150 485 1200 515
rect 1150 465 1165 485
rect 1185 465 1200 485
rect 1150 435 1200 465
rect 1150 415 1165 435
rect 1185 415 1200 435
rect 1150 385 1200 415
rect 1150 365 1165 385
rect 1185 365 1200 385
rect 1150 335 1200 365
rect 1150 315 1165 335
rect 1185 315 1200 335
rect 1150 285 1200 315
rect 1150 265 1165 285
rect 1185 265 1200 285
rect 1150 235 1200 265
rect 1150 215 1165 235
rect 1185 215 1200 235
rect 1150 185 1200 215
rect 1150 165 1165 185
rect 1185 165 1200 185
rect 1150 135 1200 165
rect 1150 115 1165 135
rect 1185 115 1200 135
rect 1150 85 1200 115
rect 1150 65 1165 85
rect 1185 65 1200 85
rect 1150 50 1200 65
rect 1450 735 1500 750
rect 1450 715 1465 735
rect 1485 715 1500 735
rect 1450 685 1500 715
rect 1450 665 1465 685
rect 1485 665 1500 685
rect 1450 635 1500 665
rect 1450 615 1465 635
rect 1485 615 1500 635
rect 1450 585 1500 615
rect 1450 565 1465 585
rect 1485 565 1500 585
rect 1450 535 1500 565
rect 1450 515 1465 535
rect 1485 515 1500 535
rect 1450 485 1500 515
rect 1450 465 1465 485
rect 1485 465 1500 485
rect 1450 435 1500 465
rect 1450 415 1465 435
rect 1485 415 1500 435
rect 1450 385 1500 415
rect 1450 365 1465 385
rect 1485 365 1500 385
rect 1450 335 1500 365
rect 1450 315 1465 335
rect 1485 315 1500 335
rect 1450 285 1500 315
rect 1450 265 1465 285
rect 1485 265 1500 285
rect 1450 235 1500 265
rect 1450 215 1465 235
rect 1485 215 1500 235
rect 1450 185 1500 215
rect 1450 165 1465 185
rect 1485 165 1500 185
rect 1450 135 1500 165
rect 1450 115 1465 135
rect 1485 115 1500 135
rect 1450 85 1500 115
rect 1450 65 1465 85
rect 1485 65 1500 85
rect 1450 50 1500 65
rect 1750 735 1800 750
rect 1750 715 1765 735
rect 1785 715 1800 735
rect 1750 685 1800 715
rect 1750 665 1765 685
rect 1785 665 1800 685
rect 1750 635 1800 665
rect 1750 615 1765 635
rect 1785 615 1800 635
rect 1750 585 1800 615
rect 1750 565 1765 585
rect 1785 565 1800 585
rect 1750 535 1800 565
rect 1750 515 1765 535
rect 1785 515 1800 535
rect 1750 485 1800 515
rect 1750 465 1765 485
rect 1785 465 1800 485
rect 1750 435 1800 465
rect 1750 415 1765 435
rect 1785 415 1800 435
rect 1750 385 1800 415
rect 1750 365 1765 385
rect 1785 365 1800 385
rect 1750 335 1800 365
rect 1750 315 1765 335
rect 1785 315 1800 335
rect 1750 285 1800 315
rect 1750 265 1765 285
rect 1785 265 1800 285
rect 1750 235 1800 265
rect 1750 215 1765 235
rect 1785 215 1800 235
rect 1750 185 1800 215
rect 1750 165 1765 185
rect 1785 165 1800 185
rect 1750 135 1800 165
rect 1750 115 1765 135
rect 1785 115 1800 135
rect 1750 85 1800 115
rect 1750 65 1765 85
rect 1785 65 1800 85
rect 1750 50 1800 65
rect 2050 735 2100 750
rect 2050 715 2065 735
rect 2085 715 2100 735
rect 2050 685 2100 715
rect 2050 665 2065 685
rect 2085 665 2100 685
rect 2050 635 2100 665
rect 2050 615 2065 635
rect 2085 615 2100 635
rect 2050 585 2100 615
rect 2050 565 2065 585
rect 2085 565 2100 585
rect 2050 535 2100 565
rect 2050 515 2065 535
rect 2085 515 2100 535
rect 2050 485 2100 515
rect 2050 465 2065 485
rect 2085 465 2100 485
rect 2050 435 2100 465
rect 2050 415 2065 435
rect 2085 415 2100 435
rect 2050 385 2100 415
rect 2050 365 2065 385
rect 2085 365 2100 385
rect 2050 335 2100 365
rect 2050 315 2065 335
rect 2085 315 2100 335
rect 2050 285 2100 315
rect 2050 265 2065 285
rect 2085 265 2100 285
rect 2050 235 2100 265
rect 2050 215 2065 235
rect 2085 215 2100 235
rect 2050 185 2100 215
rect 2050 165 2065 185
rect 2085 165 2100 185
rect 2050 135 2100 165
rect 2050 115 2065 135
rect 2085 115 2100 135
rect 2050 85 2100 115
rect 2050 65 2065 85
rect 2085 65 2100 85
rect 2050 50 2100 65
rect 2350 735 2400 750
rect 2350 715 2365 735
rect 2385 715 2400 735
rect 2350 685 2400 715
rect 2350 665 2365 685
rect 2385 665 2400 685
rect 2350 635 2400 665
rect 2350 615 2365 635
rect 2385 615 2400 635
rect 2350 585 2400 615
rect 2350 565 2365 585
rect 2385 565 2400 585
rect 2350 535 2400 565
rect 2350 515 2365 535
rect 2385 515 2400 535
rect 2350 485 2400 515
rect 2350 465 2365 485
rect 2385 465 2400 485
rect 2350 435 2400 465
rect 2350 415 2365 435
rect 2385 415 2400 435
rect 2350 385 2400 415
rect 2350 365 2365 385
rect 2385 365 2400 385
rect 2350 335 2400 365
rect 2350 315 2365 335
rect 2385 315 2400 335
rect 2350 285 2400 315
rect 2350 265 2365 285
rect 2385 265 2400 285
rect 2350 235 2400 265
rect 2350 215 2365 235
rect 2385 215 2400 235
rect 2350 185 2400 215
rect 2350 165 2365 185
rect 2385 165 2400 185
rect 2350 135 2400 165
rect 2350 115 2365 135
rect 2385 115 2400 135
rect 2350 85 2400 115
rect 2350 65 2365 85
rect 2385 65 2400 85
rect 2350 50 2400 65
rect 2650 735 2700 750
rect 2650 715 2665 735
rect 2685 715 2700 735
rect 2650 685 2700 715
rect 2650 665 2665 685
rect 2685 665 2700 685
rect 2650 635 2700 665
rect 2650 615 2665 635
rect 2685 615 2700 635
rect 2650 585 2700 615
rect 2650 565 2665 585
rect 2685 565 2700 585
rect 2650 535 2700 565
rect 2650 515 2665 535
rect 2685 515 2700 535
rect 2650 485 2700 515
rect 2650 465 2665 485
rect 2685 465 2700 485
rect 2650 435 2700 465
rect 2650 415 2665 435
rect 2685 415 2700 435
rect 2650 385 2700 415
rect 2650 365 2665 385
rect 2685 365 2700 385
rect 2650 335 2700 365
rect 2650 315 2665 335
rect 2685 315 2700 335
rect 2650 285 2700 315
rect 2650 265 2665 285
rect 2685 265 2700 285
rect 2650 235 2700 265
rect 2650 215 2665 235
rect 2685 215 2700 235
rect 2650 185 2700 215
rect 2650 165 2665 185
rect 2685 165 2700 185
rect 2650 135 2700 165
rect 2650 115 2665 135
rect 2685 115 2700 135
rect 2650 85 2700 115
rect 2650 65 2665 85
rect 2685 65 2700 85
rect 2650 50 2700 65
rect 2950 735 3000 750
rect 2950 715 2965 735
rect 2985 715 3000 735
rect 2950 685 3000 715
rect 2950 665 2965 685
rect 2985 665 3000 685
rect 2950 635 3000 665
rect 2950 615 2965 635
rect 2985 615 3000 635
rect 2950 585 3000 615
rect 2950 565 2965 585
rect 2985 565 3000 585
rect 2950 535 3000 565
rect 2950 515 2965 535
rect 2985 515 3000 535
rect 2950 485 3000 515
rect 2950 465 2965 485
rect 2985 465 3000 485
rect 2950 435 3000 465
rect 2950 415 2965 435
rect 2985 415 3000 435
rect 2950 385 3000 415
rect 2950 365 2965 385
rect 2985 365 3000 385
rect 2950 335 3000 365
rect 2950 315 2965 335
rect 2985 315 3000 335
rect 2950 285 3000 315
rect 2950 265 2965 285
rect 2985 265 3000 285
rect 2950 235 3000 265
rect 2950 215 2965 235
rect 2985 215 3000 235
rect 2950 185 3000 215
rect 2950 165 2965 185
rect 2985 165 3000 185
rect 2950 135 3000 165
rect 2950 115 2965 135
rect 2985 115 3000 135
rect 2950 85 3000 115
rect 2950 65 2965 85
rect 2985 65 3000 85
rect 2950 50 3000 65
rect 3250 735 3300 750
rect 3250 715 3265 735
rect 3285 715 3300 735
rect 3250 685 3300 715
rect 3250 665 3265 685
rect 3285 665 3300 685
rect 3250 635 3300 665
rect 3250 615 3265 635
rect 3285 615 3300 635
rect 3250 585 3300 615
rect 3250 565 3265 585
rect 3285 565 3300 585
rect 3250 535 3300 565
rect 3250 515 3265 535
rect 3285 515 3300 535
rect 3250 485 3300 515
rect 3250 465 3265 485
rect 3285 465 3300 485
rect 3250 435 3300 465
rect 3250 415 3265 435
rect 3285 415 3300 435
rect 3250 385 3300 415
rect 3250 365 3265 385
rect 3285 365 3300 385
rect 3250 335 3300 365
rect 3250 315 3265 335
rect 3285 315 3300 335
rect 3250 285 3300 315
rect 3250 265 3265 285
rect 3285 265 3300 285
rect 3250 235 3300 265
rect 3250 215 3265 235
rect 3285 215 3300 235
rect 3250 185 3300 215
rect 3250 165 3265 185
rect 3285 165 3300 185
rect 3250 135 3300 165
rect 3250 115 3265 135
rect 3285 115 3300 135
rect 3250 85 3300 115
rect 3250 65 3265 85
rect 3285 65 3300 85
rect 3250 50 3300 65
rect 3550 735 3600 750
rect 3550 715 3565 735
rect 3585 715 3600 735
rect 3550 685 3600 715
rect 3550 665 3565 685
rect 3585 665 3600 685
rect 3550 635 3600 665
rect 3550 615 3565 635
rect 3585 615 3600 635
rect 3550 585 3600 615
rect 3550 565 3565 585
rect 3585 565 3600 585
rect 3550 535 3600 565
rect 3550 515 3565 535
rect 3585 515 3600 535
rect 3550 485 3600 515
rect 3550 465 3565 485
rect 3585 465 3600 485
rect 3550 435 3600 465
rect 3550 415 3565 435
rect 3585 415 3600 435
rect 3550 385 3600 415
rect 3550 365 3565 385
rect 3585 365 3600 385
rect 3550 335 3600 365
rect 3550 315 3565 335
rect 3585 315 3600 335
rect 3550 285 3600 315
rect 3550 265 3565 285
rect 3585 265 3600 285
rect 3550 235 3600 265
rect 3550 215 3565 235
rect 3585 215 3600 235
rect 3550 185 3600 215
rect 3550 165 3565 185
rect 3585 165 3600 185
rect 3550 135 3600 165
rect 3550 115 3565 135
rect 3585 115 3600 135
rect 3550 85 3600 115
rect 3550 65 3565 85
rect 3585 65 3600 85
rect 3550 50 3600 65
rect 3700 735 3750 750
rect 3700 715 3715 735
rect 3735 715 3750 735
rect 3700 685 3750 715
rect 3700 665 3715 685
rect 3735 665 3750 685
rect 3700 635 3750 665
rect 3700 615 3715 635
rect 3735 615 3750 635
rect 3700 585 3750 615
rect 3700 565 3715 585
rect 3735 565 3750 585
rect 3700 535 3750 565
rect 3700 515 3715 535
rect 3735 515 3750 535
rect 3700 485 3750 515
rect 3700 465 3715 485
rect 3735 465 3750 485
rect 3700 435 3750 465
rect 3700 415 3715 435
rect 3735 415 3750 435
rect 3700 385 3750 415
rect 3700 365 3715 385
rect 3735 365 3750 385
rect 3700 335 3750 365
rect 3700 315 3715 335
rect 3735 315 3750 335
rect 3700 285 3750 315
rect 3700 265 3715 285
rect 3735 265 3750 285
rect 3700 235 3750 265
rect 3700 215 3715 235
rect 3735 215 3750 235
rect 3700 185 3750 215
rect 3700 165 3715 185
rect 3735 165 3750 185
rect 3700 135 3750 165
rect 3700 115 3715 135
rect 3735 115 3750 135
rect 3700 85 3750 115
rect 3700 65 3715 85
rect 3735 65 3750 85
rect 3700 50 3750 65
rect 3850 735 3900 750
rect 3850 715 3865 735
rect 3885 715 3900 735
rect 3850 685 3900 715
rect 3850 665 3865 685
rect 3885 665 3900 685
rect 3850 635 3900 665
rect 3850 615 3865 635
rect 3885 615 3900 635
rect 3850 585 3900 615
rect 3850 565 3865 585
rect 3885 565 3900 585
rect 3850 535 3900 565
rect 3850 515 3865 535
rect 3885 515 3900 535
rect 3850 485 3900 515
rect 3850 465 3865 485
rect 3885 465 3900 485
rect 3850 435 3900 465
rect 3850 415 3865 435
rect 3885 415 3900 435
rect 3850 385 3900 415
rect 3850 365 3865 385
rect 3885 365 3900 385
rect 3850 335 3900 365
rect 3850 315 3865 335
rect 3885 315 3900 335
rect 3850 285 3900 315
rect 3850 265 3865 285
rect 3885 265 3900 285
rect 3850 235 3900 265
rect 3850 215 3865 235
rect 3885 215 3900 235
rect 3850 185 3900 215
rect 3850 165 3865 185
rect 3885 165 3900 185
rect 3850 135 3900 165
rect 3850 115 3865 135
rect 3885 115 3900 135
rect 3850 85 3900 115
rect 3850 65 3865 85
rect 3885 65 3900 85
rect 3850 50 3900 65
rect 4000 735 4050 750
rect 4000 715 4015 735
rect 4035 715 4050 735
rect 4000 685 4050 715
rect 4000 665 4015 685
rect 4035 665 4050 685
rect 4000 635 4050 665
rect 4000 615 4015 635
rect 4035 615 4050 635
rect 4000 585 4050 615
rect 4000 565 4015 585
rect 4035 565 4050 585
rect 4000 535 4050 565
rect 4000 515 4015 535
rect 4035 515 4050 535
rect 4000 485 4050 515
rect 4000 465 4015 485
rect 4035 465 4050 485
rect 4000 435 4050 465
rect 4000 415 4015 435
rect 4035 415 4050 435
rect 4000 385 4050 415
rect 4000 365 4015 385
rect 4035 365 4050 385
rect 4000 335 4050 365
rect 4000 315 4015 335
rect 4035 315 4050 335
rect 4000 285 4050 315
rect 4000 265 4015 285
rect 4035 265 4050 285
rect 4000 235 4050 265
rect 4000 215 4015 235
rect 4035 215 4050 235
rect 4000 185 4050 215
rect 4000 165 4015 185
rect 4035 165 4050 185
rect 4000 135 4050 165
rect 4000 115 4015 135
rect 4035 115 4050 135
rect 4000 85 4050 115
rect 4000 65 4015 85
rect 4035 65 4050 85
rect 4000 50 4050 65
rect 4150 735 4200 750
rect 4150 715 4165 735
rect 4185 715 4200 735
rect 4150 685 4200 715
rect 4150 665 4165 685
rect 4185 665 4200 685
rect 4150 635 4200 665
rect 4150 615 4165 635
rect 4185 615 4200 635
rect 4150 585 4200 615
rect 4150 565 4165 585
rect 4185 565 4200 585
rect 4150 535 4200 565
rect 4150 515 4165 535
rect 4185 515 4200 535
rect 4150 485 4200 515
rect 4150 465 4165 485
rect 4185 465 4200 485
rect 4150 435 4200 465
rect 4150 415 4165 435
rect 4185 415 4200 435
rect 4150 385 4200 415
rect 4150 365 4165 385
rect 4185 365 4200 385
rect 4150 335 4200 365
rect 4150 315 4165 335
rect 4185 315 4200 335
rect 4150 285 4200 315
rect 4150 265 4165 285
rect 4185 265 4200 285
rect 4150 235 4200 265
rect 4150 215 4165 235
rect 4185 215 4200 235
rect 4150 185 4200 215
rect 4150 165 4165 185
rect 4185 165 4200 185
rect 4150 135 4200 165
rect 4150 115 4165 135
rect 4185 115 4200 135
rect 4150 85 4200 115
rect 4150 65 4165 85
rect 4185 65 4200 85
rect 4150 50 4200 65
rect 4300 735 4350 750
rect 4300 715 4315 735
rect 4335 715 4350 735
rect 4300 685 4350 715
rect 4300 665 4315 685
rect 4335 665 4350 685
rect 4300 635 4350 665
rect 4300 615 4315 635
rect 4335 615 4350 635
rect 4300 585 4350 615
rect 4300 565 4315 585
rect 4335 565 4350 585
rect 4300 535 4350 565
rect 4300 515 4315 535
rect 4335 515 4350 535
rect 4300 485 4350 515
rect 4300 465 4315 485
rect 4335 465 4350 485
rect 4300 435 4350 465
rect 4300 415 4315 435
rect 4335 415 4350 435
rect 4300 385 4350 415
rect 4300 365 4315 385
rect 4335 365 4350 385
rect 4300 335 4350 365
rect 4300 315 4315 335
rect 4335 315 4350 335
rect 4300 285 4350 315
rect 4300 265 4315 285
rect 4335 265 4350 285
rect 4300 235 4350 265
rect 4300 215 4315 235
rect 4335 215 4350 235
rect 4300 185 4350 215
rect 4300 165 4315 185
rect 4335 165 4350 185
rect 4300 135 4350 165
rect 4300 115 4315 135
rect 4335 115 4350 135
rect 4300 85 4350 115
rect 4300 65 4315 85
rect 4335 65 4350 85
rect 4300 50 4350 65
rect 4450 735 4500 750
rect 4450 715 4465 735
rect 4485 715 4500 735
rect 4450 685 4500 715
rect 4450 665 4465 685
rect 4485 665 4500 685
rect 4450 635 4500 665
rect 4450 615 4465 635
rect 4485 615 4500 635
rect 4450 585 4500 615
rect 4450 565 4465 585
rect 4485 565 4500 585
rect 4450 535 4500 565
rect 4450 515 4465 535
rect 4485 515 4500 535
rect 4450 485 4500 515
rect 4450 465 4465 485
rect 4485 465 4500 485
rect 4450 435 4500 465
rect 4450 415 4465 435
rect 4485 415 4500 435
rect 4450 385 4500 415
rect 4450 365 4465 385
rect 4485 365 4500 385
rect 4450 335 4500 365
rect 4450 315 4465 335
rect 4485 315 4500 335
rect 4450 285 4500 315
rect 4450 265 4465 285
rect 4485 265 4500 285
rect 4450 235 4500 265
rect 4450 215 4465 235
rect 4485 215 4500 235
rect 4450 185 4500 215
rect 4450 165 4465 185
rect 4485 165 4500 185
rect 4450 135 4500 165
rect 4450 115 4465 135
rect 4485 115 4500 135
rect 4450 85 4500 115
rect 4450 65 4465 85
rect 4485 65 4500 85
rect 4450 50 4500 65
rect 4600 735 4650 750
rect 4600 715 4615 735
rect 4635 715 4650 735
rect 4600 685 4650 715
rect 4600 665 4615 685
rect 4635 665 4650 685
rect 4600 635 4650 665
rect 4600 615 4615 635
rect 4635 615 4650 635
rect 4600 585 4650 615
rect 4600 565 4615 585
rect 4635 565 4650 585
rect 4600 535 4650 565
rect 4600 515 4615 535
rect 4635 515 4650 535
rect 4600 485 4650 515
rect 4600 465 4615 485
rect 4635 465 4650 485
rect 4600 435 4650 465
rect 4600 415 4615 435
rect 4635 415 4650 435
rect 4600 385 4650 415
rect 4600 365 4615 385
rect 4635 365 4650 385
rect 4600 335 4650 365
rect 4600 315 4615 335
rect 4635 315 4650 335
rect 4600 285 4650 315
rect 4600 265 4615 285
rect 4635 265 4650 285
rect 4600 235 4650 265
rect 4600 215 4615 235
rect 4635 215 4650 235
rect 4600 185 4650 215
rect 4600 165 4615 185
rect 4635 165 4650 185
rect 4600 135 4650 165
rect 4600 115 4615 135
rect 4635 115 4650 135
rect 4600 85 4650 115
rect 4600 65 4615 85
rect 4635 65 4650 85
rect 4600 50 4650 65
rect 4750 735 4800 750
rect 4750 715 4765 735
rect 4785 715 4800 735
rect 4750 685 4800 715
rect 4750 665 4765 685
rect 4785 665 4800 685
rect 4750 635 4800 665
rect 4750 615 4765 635
rect 4785 615 4800 635
rect 4750 585 4800 615
rect 4750 565 4765 585
rect 4785 565 4800 585
rect 4750 535 4800 565
rect 4750 515 4765 535
rect 4785 515 4800 535
rect 4750 485 4800 515
rect 4750 465 4765 485
rect 4785 465 4800 485
rect 4750 435 4800 465
rect 4750 415 4765 435
rect 4785 415 4800 435
rect 4750 385 4800 415
rect 4750 365 4765 385
rect 4785 365 4800 385
rect 4750 335 4800 365
rect 4750 315 4765 335
rect 4785 315 4800 335
rect 4750 285 4800 315
rect 4750 265 4765 285
rect 4785 265 4800 285
rect 4750 235 4800 265
rect 4750 215 4765 235
rect 4785 215 4800 235
rect 4750 185 4800 215
rect 4750 165 4765 185
rect 4785 165 4800 185
rect 4750 135 4800 165
rect 4750 115 4765 135
rect 4785 115 4800 135
rect 4750 85 4800 115
rect 4750 65 4765 85
rect 4785 65 4800 85
rect 4750 50 4800 65
rect 5050 735 5100 750
rect 5050 715 5065 735
rect 5085 715 5100 735
rect 5050 685 5100 715
rect 5050 665 5065 685
rect 5085 665 5100 685
rect 5050 635 5100 665
rect 5050 615 5065 635
rect 5085 615 5100 635
rect 5050 585 5100 615
rect 5050 565 5065 585
rect 5085 565 5100 585
rect 5050 535 5100 565
rect 5050 515 5065 535
rect 5085 515 5100 535
rect 5050 485 5100 515
rect 5050 465 5065 485
rect 5085 465 5100 485
rect 5050 435 5100 465
rect 5050 415 5065 435
rect 5085 415 5100 435
rect 5050 385 5100 415
rect 5050 365 5065 385
rect 5085 365 5100 385
rect 5050 335 5100 365
rect 5050 315 5065 335
rect 5085 315 5100 335
rect 5050 285 5100 315
rect 5050 265 5065 285
rect 5085 265 5100 285
rect 5050 235 5100 265
rect 5050 215 5065 235
rect 5085 215 5100 235
rect 5050 185 5100 215
rect 5050 165 5065 185
rect 5085 165 5100 185
rect 5050 135 5100 165
rect 5050 115 5065 135
rect 5085 115 5100 135
rect 5050 85 5100 115
rect 5050 65 5065 85
rect 5085 65 5100 85
rect 5050 50 5100 65
rect 5350 735 5400 750
rect 5350 715 5365 735
rect 5385 715 5400 735
rect 5350 685 5400 715
rect 5350 665 5365 685
rect 5385 665 5400 685
rect 5350 635 5400 665
rect 5350 615 5365 635
rect 5385 615 5400 635
rect 5350 585 5400 615
rect 5350 565 5365 585
rect 5385 565 5400 585
rect 5350 535 5400 565
rect 5350 515 5365 535
rect 5385 515 5400 535
rect 5350 485 5400 515
rect 5350 465 5365 485
rect 5385 465 5400 485
rect 5350 435 5400 465
rect 5350 415 5365 435
rect 5385 415 5400 435
rect 5350 385 5400 415
rect 5350 365 5365 385
rect 5385 365 5400 385
rect 5350 335 5400 365
rect 5350 315 5365 335
rect 5385 315 5400 335
rect 5350 285 5400 315
rect 5350 265 5365 285
rect 5385 265 5400 285
rect 5350 235 5400 265
rect 5350 215 5365 235
rect 5385 215 5400 235
rect 5350 185 5400 215
rect 5350 165 5365 185
rect 5385 165 5400 185
rect 5350 135 5400 165
rect 5350 115 5365 135
rect 5385 115 5400 135
rect 5350 85 5400 115
rect 5350 65 5365 85
rect 5385 65 5400 85
rect 5350 50 5400 65
rect 5650 735 5700 750
rect 5650 715 5665 735
rect 5685 715 5700 735
rect 5650 685 5700 715
rect 5650 665 5665 685
rect 5685 665 5700 685
rect 5650 635 5700 665
rect 5650 615 5665 635
rect 5685 615 5700 635
rect 5650 585 5700 615
rect 5650 565 5665 585
rect 5685 565 5700 585
rect 5650 535 5700 565
rect 5650 515 5665 535
rect 5685 515 5700 535
rect 5650 485 5700 515
rect 5650 465 5665 485
rect 5685 465 5700 485
rect 5650 435 5700 465
rect 5650 415 5665 435
rect 5685 415 5700 435
rect 5650 385 5700 415
rect 5650 365 5665 385
rect 5685 365 5700 385
rect 5650 335 5700 365
rect 5650 315 5665 335
rect 5685 315 5700 335
rect 5650 285 5700 315
rect 5650 265 5665 285
rect 5685 265 5700 285
rect 5650 235 5700 265
rect 5650 215 5665 235
rect 5685 215 5700 235
rect 5650 185 5700 215
rect 5650 165 5665 185
rect 5685 165 5700 185
rect 5650 135 5700 165
rect 5650 115 5665 135
rect 5685 115 5700 135
rect 5650 85 5700 115
rect 5650 65 5665 85
rect 5685 65 5700 85
rect 5650 50 5700 65
rect 5950 735 6000 750
rect 5950 715 5965 735
rect 5985 715 6000 735
rect 5950 685 6000 715
rect 5950 665 5965 685
rect 5985 665 6000 685
rect 5950 635 6000 665
rect 5950 615 5965 635
rect 5985 615 6000 635
rect 5950 585 6000 615
rect 5950 565 5965 585
rect 5985 565 6000 585
rect 5950 535 6000 565
rect 5950 515 5965 535
rect 5985 515 6000 535
rect 5950 485 6000 515
rect 5950 465 5965 485
rect 5985 465 6000 485
rect 5950 435 6000 465
rect 5950 415 5965 435
rect 5985 415 6000 435
rect 5950 385 6000 415
rect 5950 365 5965 385
rect 5985 365 6000 385
rect 5950 335 6000 365
rect 5950 315 5965 335
rect 5985 315 6000 335
rect 5950 285 6000 315
rect 5950 265 5965 285
rect 5985 265 6000 285
rect 5950 235 6000 265
rect 5950 215 5965 235
rect 5985 215 6000 235
rect 5950 185 6000 215
rect 5950 165 5965 185
rect 5985 165 6000 185
rect 5950 135 6000 165
rect 5950 115 5965 135
rect 5985 115 6000 135
rect 5950 85 6000 115
rect 5950 65 5965 85
rect 5985 65 6000 85
rect 5950 50 6000 65
rect 6250 735 6300 750
rect 6250 715 6265 735
rect 6285 715 6300 735
rect 6250 685 6300 715
rect 6250 665 6265 685
rect 6285 665 6300 685
rect 6250 635 6300 665
rect 6250 615 6265 635
rect 6285 615 6300 635
rect 6250 585 6300 615
rect 6250 565 6265 585
rect 6285 565 6300 585
rect 6250 535 6300 565
rect 6250 515 6265 535
rect 6285 515 6300 535
rect 6250 485 6300 515
rect 6250 465 6265 485
rect 6285 465 6300 485
rect 6250 435 6300 465
rect 6250 415 6265 435
rect 6285 415 6300 435
rect 6250 385 6300 415
rect 6250 365 6265 385
rect 6285 365 6300 385
rect 6250 335 6300 365
rect 6250 315 6265 335
rect 6285 315 6300 335
rect 6250 285 6300 315
rect 6250 265 6265 285
rect 6285 265 6300 285
rect 6250 235 6300 265
rect 6250 215 6265 235
rect 6285 215 6300 235
rect 6250 185 6300 215
rect 6250 165 6265 185
rect 6285 165 6300 185
rect 6250 135 6300 165
rect 6250 115 6265 135
rect 6285 115 6300 135
rect 6250 85 6300 115
rect 6250 65 6265 85
rect 6285 65 6300 85
rect 6250 50 6300 65
rect 6550 735 6600 750
rect 6550 715 6565 735
rect 6585 715 6600 735
rect 6550 685 6600 715
rect 6550 665 6565 685
rect 6585 665 6600 685
rect 6550 635 6600 665
rect 6550 615 6565 635
rect 6585 615 6600 635
rect 6550 585 6600 615
rect 6550 565 6565 585
rect 6585 565 6600 585
rect 6550 535 6600 565
rect 6550 515 6565 535
rect 6585 515 6600 535
rect 6550 485 6600 515
rect 6550 465 6565 485
rect 6585 465 6600 485
rect 6550 435 6600 465
rect 6550 415 6565 435
rect 6585 415 6600 435
rect 6550 385 6600 415
rect 6550 365 6565 385
rect 6585 365 6600 385
rect 6550 335 6600 365
rect 6550 315 6565 335
rect 6585 315 6600 335
rect 6550 285 6600 315
rect 6550 265 6565 285
rect 6585 265 6600 285
rect 6550 235 6600 265
rect 6550 215 6565 235
rect 6585 215 6600 235
rect 6550 185 6600 215
rect 6550 165 6565 185
rect 6585 165 6600 185
rect 6550 135 6600 165
rect 6550 115 6565 135
rect 6585 115 6600 135
rect 6550 85 6600 115
rect 6550 65 6565 85
rect 6585 65 6600 85
rect 6550 50 6600 65
rect 6850 735 6900 750
rect 6850 715 6865 735
rect 6885 715 6900 735
rect 6850 685 6900 715
rect 6850 665 6865 685
rect 6885 665 6900 685
rect 6850 635 6900 665
rect 6850 615 6865 635
rect 6885 615 6900 635
rect 6850 585 6900 615
rect 6850 565 6865 585
rect 6885 565 6900 585
rect 6850 535 6900 565
rect 6850 515 6865 535
rect 6885 515 6900 535
rect 6850 485 6900 515
rect 6850 465 6865 485
rect 6885 465 6900 485
rect 6850 435 6900 465
rect 6850 415 6865 435
rect 6885 415 6900 435
rect 6850 385 6900 415
rect 6850 365 6865 385
rect 6885 365 6900 385
rect 6850 335 6900 365
rect 6850 315 6865 335
rect 6885 315 6900 335
rect 6850 285 6900 315
rect 6850 265 6865 285
rect 6885 265 6900 285
rect 6850 235 6900 265
rect 6850 215 6865 235
rect 6885 215 6900 235
rect 6850 185 6900 215
rect 6850 165 6865 185
rect 6885 165 6900 185
rect 6850 135 6900 165
rect 6850 115 6865 135
rect 6885 115 6900 135
rect 6850 85 6900 115
rect 6850 65 6865 85
rect 6885 65 6900 85
rect 6850 50 6900 65
rect 7150 735 7200 750
rect 7150 715 7165 735
rect 7185 715 7200 735
rect 7150 685 7200 715
rect 7150 665 7165 685
rect 7185 665 7200 685
rect 7150 635 7200 665
rect 7150 615 7165 635
rect 7185 615 7200 635
rect 7150 585 7200 615
rect 7150 565 7165 585
rect 7185 565 7200 585
rect 7150 535 7200 565
rect 7150 515 7165 535
rect 7185 515 7200 535
rect 7150 485 7200 515
rect 7150 465 7165 485
rect 7185 465 7200 485
rect 7150 435 7200 465
rect 7150 415 7165 435
rect 7185 415 7200 435
rect 7150 385 7200 415
rect 7150 365 7165 385
rect 7185 365 7200 385
rect 7150 335 7200 365
rect 7150 315 7165 335
rect 7185 315 7200 335
rect 7150 285 7200 315
rect 7150 265 7165 285
rect 7185 265 7200 285
rect 7150 235 7200 265
rect 7150 215 7165 235
rect 7185 215 7200 235
rect 7150 185 7200 215
rect 7150 165 7165 185
rect 7185 165 7200 185
rect 7150 135 7200 165
rect 7150 115 7165 135
rect 7185 115 7200 135
rect 7150 85 7200 115
rect 7150 65 7165 85
rect 7185 65 7200 85
rect 7150 50 7200 65
rect 8350 735 8400 750
rect 8350 715 8365 735
rect 8385 715 8400 735
rect 8350 685 8400 715
rect 8350 665 8365 685
rect 8385 665 8400 685
rect 8350 635 8400 665
rect 8350 615 8365 635
rect 8385 615 8400 635
rect 8350 585 8400 615
rect 8350 565 8365 585
rect 8385 565 8400 585
rect 8350 535 8400 565
rect 8350 515 8365 535
rect 8385 515 8400 535
rect 8350 485 8400 515
rect 8350 465 8365 485
rect 8385 465 8400 485
rect 8350 435 8400 465
rect 8350 415 8365 435
rect 8385 415 8400 435
rect 8350 385 8400 415
rect 8350 365 8365 385
rect 8385 365 8400 385
rect 8350 335 8400 365
rect 8350 315 8365 335
rect 8385 315 8400 335
rect 8350 285 8400 315
rect 8350 265 8365 285
rect 8385 265 8400 285
rect 8350 235 8400 265
rect 8350 215 8365 235
rect 8385 215 8400 235
rect 8350 185 8400 215
rect 8350 165 8365 185
rect 8385 165 8400 185
rect 8350 135 8400 165
rect 8350 115 8365 135
rect 8385 115 8400 135
rect 8350 85 8400 115
rect 8350 65 8365 85
rect 8385 65 8400 85
rect 8350 50 8400 65
rect 9550 735 9600 750
rect 9550 715 9565 735
rect 9585 715 9600 735
rect 9550 685 9600 715
rect 9550 665 9565 685
rect 9585 665 9600 685
rect 9550 635 9600 665
rect 9550 615 9565 635
rect 9585 615 9600 635
rect 9550 585 9600 615
rect 9550 565 9565 585
rect 9585 565 9600 585
rect 9550 535 9600 565
rect 9550 515 9565 535
rect 9585 515 9600 535
rect 9550 485 9600 515
rect 9550 465 9565 485
rect 9585 465 9600 485
rect 9550 435 9600 465
rect 9550 415 9565 435
rect 9585 415 9600 435
rect 9550 385 9600 415
rect 9550 365 9565 385
rect 9585 365 9600 385
rect 9550 335 9600 365
rect 9550 315 9565 335
rect 9585 315 9600 335
rect 9550 285 9600 315
rect 9550 265 9565 285
rect 9585 265 9600 285
rect 9550 235 9600 265
rect 9550 215 9565 235
rect 9585 215 9600 235
rect 9550 185 9600 215
rect 9550 165 9565 185
rect 9585 165 9600 185
rect 9550 135 9600 165
rect 9550 115 9565 135
rect 9585 115 9600 135
rect 9550 85 9600 115
rect 9550 65 9565 85
rect 9585 65 9600 85
rect 9550 50 9600 65
rect 10750 735 10800 750
rect 10750 715 10765 735
rect 10785 715 10800 735
rect 10750 685 10800 715
rect 10750 665 10765 685
rect 10785 665 10800 685
rect 10750 635 10800 665
rect 10750 615 10765 635
rect 10785 615 10800 635
rect 10750 585 10800 615
rect 10750 565 10765 585
rect 10785 565 10800 585
rect 10750 535 10800 565
rect 10750 515 10765 535
rect 10785 515 10800 535
rect 10750 485 10800 515
rect 10750 465 10765 485
rect 10785 465 10800 485
rect 10750 435 10800 465
rect 10750 415 10765 435
rect 10785 415 10800 435
rect 10750 385 10800 415
rect 10750 365 10765 385
rect 10785 365 10800 385
rect 10750 335 10800 365
rect 10750 315 10765 335
rect 10785 315 10800 335
rect 10750 285 10800 315
rect 10750 265 10765 285
rect 10785 265 10800 285
rect 10750 235 10800 265
rect 10750 215 10765 235
rect 10785 215 10800 235
rect 10750 185 10800 215
rect 10750 165 10765 185
rect 10785 165 10800 185
rect 10750 135 10800 165
rect 10750 115 10765 135
rect 10785 115 10800 135
rect 10750 85 10800 115
rect 10750 65 10765 85
rect 10785 65 10800 85
rect 10750 50 10800 65
rect 11950 735 12000 750
rect 11950 715 11965 735
rect 11985 715 12000 735
rect 11950 685 12000 715
rect 11950 665 11965 685
rect 11985 665 12000 685
rect 11950 635 12000 665
rect 11950 615 11965 635
rect 11985 615 12000 635
rect 11950 585 12000 615
rect 11950 565 11965 585
rect 11985 565 12000 585
rect 11950 535 12000 565
rect 11950 515 11965 535
rect 11985 515 12000 535
rect 11950 485 12000 515
rect 11950 465 11965 485
rect 11985 465 12000 485
rect 11950 435 12000 465
rect 11950 415 11965 435
rect 11985 415 12000 435
rect 11950 385 12000 415
rect 11950 365 11965 385
rect 11985 365 12000 385
rect 11950 335 12000 365
rect 11950 315 11965 335
rect 11985 315 12000 335
rect 11950 285 12000 315
rect 11950 265 11965 285
rect 11985 265 12000 285
rect 11950 235 12000 265
rect 11950 215 11965 235
rect 11985 215 12000 235
rect 11950 185 12000 215
rect 11950 165 11965 185
rect 11985 165 12000 185
rect 11950 135 12000 165
rect 11950 115 11965 135
rect 11985 115 12000 135
rect 11950 85 12000 115
rect 11950 65 11965 85
rect 11985 65 12000 85
rect 11950 50 12000 65
rect 12250 735 12300 750
rect 12250 715 12265 735
rect 12285 715 12300 735
rect 12250 685 12300 715
rect 12250 665 12265 685
rect 12285 665 12300 685
rect 12250 635 12300 665
rect 12250 615 12265 635
rect 12285 615 12300 635
rect 12250 585 12300 615
rect 12250 565 12265 585
rect 12285 565 12300 585
rect 12250 535 12300 565
rect 12250 515 12265 535
rect 12285 515 12300 535
rect 12250 485 12300 515
rect 12250 465 12265 485
rect 12285 465 12300 485
rect 12250 435 12300 465
rect 12250 415 12265 435
rect 12285 415 12300 435
rect 12250 385 12300 415
rect 12250 365 12265 385
rect 12285 365 12300 385
rect 12250 335 12300 365
rect 12250 315 12265 335
rect 12285 315 12300 335
rect 12250 285 12300 315
rect 12250 265 12265 285
rect 12285 265 12300 285
rect 12250 235 12300 265
rect 12250 215 12265 235
rect 12285 215 12300 235
rect 12250 185 12300 215
rect 12250 165 12265 185
rect 12285 165 12300 185
rect 12250 135 12300 165
rect 12250 115 12265 135
rect 12285 115 12300 135
rect 12250 85 12300 115
rect 12250 65 12265 85
rect 12285 65 12300 85
rect 12250 50 12300 65
rect 12550 735 12600 750
rect 12550 715 12565 735
rect 12585 715 12600 735
rect 12550 685 12600 715
rect 12550 665 12565 685
rect 12585 665 12600 685
rect 12550 635 12600 665
rect 12550 615 12565 635
rect 12585 615 12600 635
rect 12550 585 12600 615
rect 12550 565 12565 585
rect 12585 565 12600 585
rect 12550 535 12600 565
rect 12550 515 12565 535
rect 12585 515 12600 535
rect 12550 485 12600 515
rect 12550 465 12565 485
rect 12585 465 12600 485
rect 12550 435 12600 465
rect 12550 415 12565 435
rect 12585 415 12600 435
rect 12550 385 12600 415
rect 12550 365 12565 385
rect 12585 365 12600 385
rect 12550 335 12600 365
rect 12550 315 12565 335
rect 12585 315 12600 335
rect 12550 285 12600 315
rect 12550 265 12565 285
rect 12585 265 12600 285
rect 12550 235 12600 265
rect 12550 215 12565 235
rect 12585 215 12600 235
rect 12550 185 12600 215
rect 12550 165 12565 185
rect 12585 165 12600 185
rect 12550 135 12600 165
rect 12550 115 12565 135
rect 12585 115 12600 135
rect 12550 85 12600 115
rect 12550 65 12565 85
rect 12585 65 12600 85
rect 12550 50 12600 65
rect 12850 735 12900 750
rect 12850 715 12865 735
rect 12885 715 12900 735
rect 12850 685 12900 715
rect 12850 665 12865 685
rect 12885 665 12900 685
rect 12850 635 12900 665
rect 12850 615 12865 635
rect 12885 615 12900 635
rect 12850 585 12900 615
rect 12850 565 12865 585
rect 12885 565 12900 585
rect 12850 535 12900 565
rect 12850 515 12865 535
rect 12885 515 12900 535
rect 12850 485 12900 515
rect 12850 465 12865 485
rect 12885 465 12900 485
rect 12850 435 12900 465
rect 12850 415 12865 435
rect 12885 415 12900 435
rect 12850 385 12900 415
rect 12850 365 12865 385
rect 12885 365 12900 385
rect 12850 335 12900 365
rect 12850 315 12865 335
rect 12885 315 12900 335
rect 12850 285 12900 315
rect 12850 265 12865 285
rect 12885 265 12900 285
rect 12850 235 12900 265
rect 12850 215 12865 235
rect 12885 215 12900 235
rect 12850 185 12900 215
rect 12850 165 12865 185
rect 12885 165 12900 185
rect 12850 135 12900 165
rect 12850 115 12865 135
rect 12885 115 12900 135
rect 12850 85 12900 115
rect 12850 65 12865 85
rect 12885 65 12900 85
rect 12850 50 12900 65
rect 13150 735 13200 750
rect 13150 715 13165 735
rect 13185 715 13200 735
rect 13150 685 13200 715
rect 13150 665 13165 685
rect 13185 665 13200 685
rect 13150 635 13200 665
rect 13150 615 13165 635
rect 13185 615 13200 635
rect 13150 585 13200 615
rect 13150 565 13165 585
rect 13185 565 13200 585
rect 13150 535 13200 565
rect 13150 515 13165 535
rect 13185 515 13200 535
rect 13150 485 13200 515
rect 13150 465 13165 485
rect 13185 465 13200 485
rect 13150 435 13200 465
rect 13150 415 13165 435
rect 13185 415 13200 435
rect 13150 385 13200 415
rect 13150 365 13165 385
rect 13185 365 13200 385
rect 13150 335 13200 365
rect 13150 315 13165 335
rect 13185 315 13200 335
rect 13150 285 13200 315
rect 13150 265 13165 285
rect 13185 265 13200 285
rect 13150 235 13200 265
rect 13150 215 13165 235
rect 13185 215 13200 235
rect 13150 185 13200 215
rect 13150 165 13165 185
rect 13185 165 13200 185
rect 13150 135 13200 165
rect 13150 115 13165 135
rect 13185 115 13200 135
rect 13150 85 13200 115
rect 13150 65 13165 85
rect 13185 65 13200 85
rect 13150 50 13200 65
rect 13450 735 13500 750
rect 13450 715 13465 735
rect 13485 715 13500 735
rect 13450 685 13500 715
rect 13450 665 13465 685
rect 13485 665 13500 685
rect 13450 635 13500 665
rect 13450 615 13465 635
rect 13485 615 13500 635
rect 13450 585 13500 615
rect 13450 565 13465 585
rect 13485 565 13500 585
rect 13450 535 13500 565
rect 13450 515 13465 535
rect 13485 515 13500 535
rect 13450 485 13500 515
rect 13450 465 13465 485
rect 13485 465 13500 485
rect 13450 435 13500 465
rect 13450 415 13465 435
rect 13485 415 13500 435
rect 13450 385 13500 415
rect 13450 365 13465 385
rect 13485 365 13500 385
rect 13450 335 13500 365
rect 13450 315 13465 335
rect 13485 315 13500 335
rect 13450 285 13500 315
rect 13450 265 13465 285
rect 13485 265 13500 285
rect 13450 235 13500 265
rect 13450 215 13465 235
rect 13485 215 13500 235
rect 13450 185 13500 215
rect 13450 165 13465 185
rect 13485 165 13500 185
rect 13450 135 13500 165
rect 13450 115 13465 135
rect 13485 115 13500 135
rect 13450 85 13500 115
rect 13450 65 13465 85
rect 13485 65 13500 85
rect 13450 50 13500 65
rect 13750 735 13800 750
rect 13750 715 13765 735
rect 13785 715 13800 735
rect 13750 685 13800 715
rect 13750 665 13765 685
rect 13785 665 13800 685
rect 13750 635 13800 665
rect 13750 615 13765 635
rect 13785 615 13800 635
rect 13750 585 13800 615
rect 13750 565 13765 585
rect 13785 565 13800 585
rect 13750 535 13800 565
rect 13750 515 13765 535
rect 13785 515 13800 535
rect 13750 485 13800 515
rect 13750 465 13765 485
rect 13785 465 13800 485
rect 13750 435 13800 465
rect 13750 415 13765 435
rect 13785 415 13800 435
rect 13750 385 13800 415
rect 13750 365 13765 385
rect 13785 365 13800 385
rect 13750 335 13800 365
rect 13750 315 13765 335
rect 13785 315 13800 335
rect 13750 285 13800 315
rect 13750 265 13765 285
rect 13785 265 13800 285
rect 13750 235 13800 265
rect 13750 215 13765 235
rect 13785 215 13800 235
rect 13750 185 13800 215
rect 13750 165 13765 185
rect 13785 165 13800 185
rect 13750 135 13800 165
rect 13750 115 13765 135
rect 13785 115 13800 135
rect 13750 85 13800 115
rect 13750 65 13765 85
rect 13785 65 13800 85
rect 13750 50 13800 65
rect 14050 735 14100 750
rect 14050 715 14065 735
rect 14085 715 14100 735
rect 14050 685 14100 715
rect 14050 665 14065 685
rect 14085 665 14100 685
rect 14050 635 14100 665
rect 14050 615 14065 635
rect 14085 615 14100 635
rect 14050 585 14100 615
rect 14050 565 14065 585
rect 14085 565 14100 585
rect 14050 535 14100 565
rect 14050 515 14065 535
rect 14085 515 14100 535
rect 14050 485 14100 515
rect 14050 465 14065 485
rect 14085 465 14100 485
rect 14050 435 14100 465
rect 14050 415 14065 435
rect 14085 415 14100 435
rect 14050 385 14100 415
rect 14050 365 14065 385
rect 14085 365 14100 385
rect 14050 335 14100 365
rect 14050 315 14065 335
rect 14085 315 14100 335
rect 14050 285 14100 315
rect 14050 265 14065 285
rect 14085 265 14100 285
rect 14050 235 14100 265
rect 14050 215 14065 235
rect 14085 215 14100 235
rect 14050 185 14100 215
rect 14050 165 14065 185
rect 14085 165 14100 185
rect 14050 135 14100 165
rect 14050 115 14065 135
rect 14085 115 14100 135
rect 14050 85 14100 115
rect 14050 65 14065 85
rect 14085 65 14100 85
rect 14050 50 14100 65
rect 14350 735 14400 750
rect 14350 715 14365 735
rect 14385 715 14400 735
rect 14350 685 14400 715
rect 14350 665 14365 685
rect 14385 665 14400 685
rect 14350 635 14400 665
rect 14350 615 14365 635
rect 14385 615 14400 635
rect 14350 585 14400 615
rect 14350 565 14365 585
rect 14385 565 14400 585
rect 14350 535 14400 565
rect 14350 515 14365 535
rect 14385 515 14400 535
rect 14350 485 14400 515
rect 14350 465 14365 485
rect 14385 465 14400 485
rect 14350 435 14400 465
rect 14350 415 14365 435
rect 14385 415 14400 435
rect 14350 385 14400 415
rect 14350 365 14365 385
rect 14385 365 14400 385
rect 14350 335 14400 365
rect 14350 315 14365 335
rect 14385 315 14400 335
rect 14350 285 14400 315
rect 14350 265 14365 285
rect 14385 265 14400 285
rect 14350 235 14400 265
rect 14350 215 14365 235
rect 14385 215 14400 235
rect 14350 185 14400 215
rect 14350 165 14365 185
rect 14385 165 14400 185
rect 14350 135 14400 165
rect 14350 115 14365 135
rect 14385 115 14400 135
rect 14350 85 14400 115
rect 14350 65 14365 85
rect 14385 65 14400 85
rect 14350 50 14400 65
rect 15550 735 15600 750
rect 15550 715 15565 735
rect 15585 715 15600 735
rect 15550 685 15600 715
rect 15550 665 15565 685
rect 15585 665 15600 685
rect 15550 635 15600 665
rect 15550 615 15565 635
rect 15585 615 15600 635
rect 15550 585 15600 615
rect 15550 565 15565 585
rect 15585 565 15600 585
rect 15550 535 15600 565
rect 15550 515 15565 535
rect 15585 515 15600 535
rect 15550 485 15600 515
rect 15550 465 15565 485
rect 15585 465 15600 485
rect 15550 435 15600 465
rect 15550 415 15565 435
rect 15585 415 15600 435
rect 15550 385 15600 415
rect 15550 365 15565 385
rect 15585 365 15600 385
rect 15550 335 15600 365
rect 15550 315 15565 335
rect 15585 315 15600 335
rect 15550 285 15600 315
rect 15550 265 15565 285
rect 15585 265 15600 285
rect 15550 235 15600 265
rect 15550 215 15565 235
rect 15585 215 15600 235
rect 15550 185 15600 215
rect 15550 165 15565 185
rect 15585 165 15600 185
rect 15550 135 15600 165
rect 15550 115 15565 135
rect 15585 115 15600 135
rect 15550 85 15600 115
rect 15550 65 15565 85
rect 15585 65 15600 85
rect 15550 50 15600 65
rect 16750 735 16800 750
rect 16750 715 16765 735
rect 16785 715 16800 735
rect 16750 685 16800 715
rect 16750 665 16765 685
rect 16785 665 16800 685
rect 16750 635 16800 665
rect 16750 615 16765 635
rect 16785 615 16800 635
rect 16750 585 16800 615
rect 16750 565 16765 585
rect 16785 565 16800 585
rect 16750 535 16800 565
rect 16750 515 16765 535
rect 16785 515 16800 535
rect 16750 485 16800 515
rect 16750 465 16765 485
rect 16785 465 16800 485
rect 16750 435 16800 465
rect 16750 415 16765 435
rect 16785 415 16800 435
rect 16750 385 16800 415
rect 16750 365 16765 385
rect 16785 365 16800 385
rect 16750 335 16800 365
rect 16750 315 16765 335
rect 16785 315 16800 335
rect 16750 285 16800 315
rect 16750 265 16765 285
rect 16785 265 16800 285
rect 16750 235 16800 265
rect 16750 215 16765 235
rect 16785 215 16800 235
rect 16750 185 16800 215
rect 16750 165 16765 185
rect 16785 165 16800 185
rect 16750 135 16800 165
rect 16750 115 16765 135
rect 16785 115 16800 135
rect 16750 85 16800 115
rect 16750 65 16765 85
rect 16785 65 16800 85
rect 16750 50 16800 65
rect 17950 735 18000 750
rect 17950 715 17965 735
rect 17985 715 18000 735
rect 17950 685 18000 715
rect 17950 665 17965 685
rect 17985 665 18000 685
rect 17950 635 18000 665
rect 17950 615 17965 635
rect 17985 615 18000 635
rect 17950 585 18000 615
rect 17950 565 17965 585
rect 17985 565 18000 585
rect 17950 535 18000 565
rect 17950 515 17965 535
rect 17985 515 18000 535
rect 17950 485 18000 515
rect 17950 465 17965 485
rect 17985 465 18000 485
rect 17950 435 18000 465
rect 17950 415 17965 435
rect 17985 415 18000 435
rect 17950 385 18000 415
rect 17950 365 17965 385
rect 17985 365 18000 385
rect 17950 335 18000 365
rect 17950 315 17965 335
rect 17985 315 18000 335
rect 17950 285 18000 315
rect 17950 265 17965 285
rect 17985 265 18000 285
rect 17950 235 18000 265
rect 17950 215 17965 235
rect 17985 215 18000 235
rect 17950 185 18000 215
rect 17950 165 17965 185
rect 17985 165 18000 185
rect 17950 135 18000 165
rect 17950 115 17965 135
rect 17985 115 18000 135
rect 17950 85 18000 115
rect 17950 65 17965 85
rect 17985 65 18000 85
rect 17950 50 18000 65
rect 19150 735 19200 750
rect 19150 715 19165 735
rect 19185 715 19200 735
rect 19150 685 19200 715
rect 19150 665 19165 685
rect 19185 665 19200 685
rect 19150 635 19200 665
rect 19150 615 19165 635
rect 19185 615 19200 635
rect 19150 585 19200 615
rect 19150 565 19165 585
rect 19185 565 19200 585
rect 19150 535 19200 565
rect 19150 515 19165 535
rect 19185 515 19200 535
rect 19150 485 19200 515
rect 19150 465 19165 485
rect 19185 465 19200 485
rect 19150 435 19200 465
rect 19150 415 19165 435
rect 19185 415 19200 435
rect 19150 385 19200 415
rect 19150 365 19165 385
rect 19185 365 19200 385
rect 19150 335 19200 365
rect 19150 315 19165 335
rect 19185 315 19200 335
rect 19150 285 19200 315
rect 19150 265 19165 285
rect 19185 265 19200 285
rect 19150 235 19200 265
rect 19150 215 19165 235
rect 19185 215 19200 235
rect 19150 185 19200 215
rect 19150 165 19165 185
rect 19185 165 19200 185
rect 19150 135 19200 165
rect 19150 115 19165 135
rect 19185 115 19200 135
rect 19150 85 19200 115
rect 19150 65 19165 85
rect 19185 65 19200 85
rect 19150 50 19200 65
rect 20350 735 20400 750
rect 20350 715 20365 735
rect 20385 715 20400 735
rect 20350 685 20400 715
rect 20350 665 20365 685
rect 20385 665 20400 685
rect 20350 635 20400 665
rect 20350 615 20365 635
rect 20385 615 20400 635
rect 20350 585 20400 615
rect 20350 565 20365 585
rect 20385 565 20400 585
rect 20350 535 20400 565
rect 20350 515 20365 535
rect 20385 515 20400 535
rect 20350 485 20400 515
rect 20350 465 20365 485
rect 20385 465 20400 485
rect 20350 435 20400 465
rect 20350 415 20365 435
rect 20385 415 20400 435
rect 20350 385 20400 415
rect 20350 365 20365 385
rect 20385 365 20400 385
rect 20350 335 20400 365
rect 20350 315 20365 335
rect 20385 315 20400 335
rect 20350 285 20400 315
rect 20350 265 20365 285
rect 20385 265 20400 285
rect 20350 235 20400 265
rect 20350 215 20365 235
rect 20385 215 20400 235
rect 20350 185 20400 215
rect 20350 165 20365 185
rect 20385 165 20400 185
rect 20350 135 20400 165
rect 20350 115 20365 135
rect 20385 115 20400 135
rect 20350 85 20400 115
rect 20350 65 20365 85
rect 20385 65 20400 85
rect 20350 50 20400 65
rect 21550 735 21600 750
rect 21550 715 21565 735
rect 21585 715 21600 735
rect 21550 685 21600 715
rect 21550 665 21565 685
rect 21585 665 21600 685
rect 21550 635 21600 665
rect 21550 615 21565 635
rect 21585 615 21600 635
rect 21550 585 21600 615
rect 21550 565 21565 585
rect 21585 565 21600 585
rect 21550 535 21600 565
rect 21550 515 21565 535
rect 21585 515 21600 535
rect 21550 485 21600 515
rect 21550 465 21565 485
rect 21585 465 21600 485
rect 21550 435 21600 465
rect 21550 415 21565 435
rect 21585 415 21600 435
rect 21550 385 21600 415
rect 21550 365 21565 385
rect 21585 365 21600 385
rect 21550 335 21600 365
rect 21550 315 21565 335
rect 21585 315 21600 335
rect 21550 285 21600 315
rect 21550 265 21565 285
rect 21585 265 21600 285
rect 21550 235 21600 265
rect 21550 215 21565 235
rect 21585 215 21600 235
rect 21550 185 21600 215
rect 21550 165 21565 185
rect 21585 165 21600 185
rect 21550 135 21600 165
rect 21550 115 21565 135
rect 21585 115 21600 135
rect 21550 85 21600 115
rect 21550 65 21565 85
rect 21585 65 21600 85
rect 21550 50 21600 65
rect 22450 735 22500 750
rect 22450 715 22465 735
rect 22485 715 22500 735
rect 22450 685 22500 715
rect 22450 665 22465 685
rect 22485 665 22500 685
rect 22450 635 22500 665
rect 22450 615 22465 635
rect 22485 615 22500 635
rect 22450 585 22500 615
rect 22450 565 22465 585
rect 22485 565 22500 585
rect 22450 535 22500 565
rect 22450 515 22465 535
rect 22485 515 22500 535
rect 22450 485 22500 515
rect 22450 465 22465 485
rect 22485 465 22500 485
rect 22450 435 22500 465
rect 22450 415 22465 435
rect 22485 415 22500 435
rect 22450 385 22500 415
rect 22450 365 22465 385
rect 22485 365 22500 385
rect 22450 335 22500 365
rect 22450 315 22465 335
rect 22485 315 22500 335
rect 22450 285 22500 315
rect 22450 265 22465 285
rect 22485 265 22500 285
rect 22450 235 22500 265
rect 22450 215 22465 235
rect 22485 215 22500 235
rect 22450 185 22500 215
rect 22450 165 22465 185
rect 22485 165 22500 185
rect 22450 135 22500 165
rect 22450 115 22465 135
rect 22485 115 22500 135
rect 22450 85 22500 115
rect 22450 65 22465 85
rect 22485 65 22500 85
rect 22450 50 22500 65
rect 23350 735 23400 750
rect 23350 715 23365 735
rect 23385 715 23400 735
rect 23350 685 23400 715
rect 23350 665 23365 685
rect 23385 665 23400 685
rect 23350 635 23400 665
rect 23350 615 23365 635
rect 23385 615 23400 635
rect 23350 585 23400 615
rect 23350 565 23365 585
rect 23385 565 23400 585
rect 23350 535 23400 565
rect 23350 515 23365 535
rect 23385 515 23400 535
rect 23350 485 23400 515
rect 23350 465 23365 485
rect 23385 465 23400 485
rect 23350 435 23400 465
rect 23350 415 23365 435
rect 23385 415 23400 435
rect 23350 385 23400 415
rect 23350 365 23365 385
rect 23385 365 23400 385
rect 23350 335 23400 365
rect 23350 315 23365 335
rect 23385 315 23400 335
rect 23350 285 23400 315
rect 23350 265 23365 285
rect 23385 265 23400 285
rect 23350 235 23400 265
rect 23350 215 23365 235
rect 23385 215 23400 235
rect 23350 185 23400 215
rect 23350 165 23365 185
rect 23385 165 23400 185
rect 23350 135 23400 165
rect 23350 115 23365 135
rect 23385 115 23400 135
rect 23350 85 23400 115
rect 23350 65 23365 85
rect 23385 65 23400 85
rect 23350 50 23400 65
rect 24550 735 24600 750
rect 24550 715 24565 735
rect 24585 715 24600 735
rect 24550 685 24600 715
rect 24550 665 24565 685
rect 24585 665 24600 685
rect 24550 635 24600 665
rect 24550 615 24565 635
rect 24585 615 24600 635
rect 24550 585 24600 615
rect 24550 565 24565 585
rect 24585 565 24600 585
rect 24550 535 24600 565
rect 24550 515 24565 535
rect 24585 515 24600 535
rect 24550 485 24600 515
rect 24550 465 24565 485
rect 24585 465 24600 485
rect 24550 435 24600 465
rect 24550 415 24565 435
rect 24585 415 24600 435
rect 24550 385 24600 415
rect 24550 365 24565 385
rect 24585 365 24600 385
rect 24550 335 24600 365
rect 24550 315 24565 335
rect 24585 315 24600 335
rect 24550 285 24600 315
rect 24550 265 24565 285
rect 24585 265 24600 285
rect 24550 235 24600 265
rect 24550 215 24565 235
rect 24585 215 24600 235
rect 24550 185 24600 215
rect 24550 165 24565 185
rect 24585 165 24600 185
rect 24550 135 24600 165
rect 24550 115 24565 135
rect 24585 115 24600 135
rect 24550 85 24600 115
rect 24550 65 24565 85
rect 24585 65 24600 85
rect 24550 50 24600 65
rect 25750 735 25800 750
rect 25750 715 25765 735
rect 25785 715 25800 735
rect 25750 685 25800 715
rect 25750 665 25765 685
rect 25785 665 25800 685
rect 25750 635 25800 665
rect 25750 615 25765 635
rect 25785 615 25800 635
rect 25750 585 25800 615
rect 25750 565 25765 585
rect 25785 565 25800 585
rect 25750 535 25800 565
rect 25750 515 25765 535
rect 25785 515 25800 535
rect 25750 485 25800 515
rect 25750 465 25765 485
rect 25785 465 25800 485
rect 25750 435 25800 465
rect 25750 415 25765 435
rect 25785 415 25800 435
rect 25750 385 25800 415
rect 25750 365 25765 385
rect 25785 365 25800 385
rect 25750 335 25800 365
rect 25750 315 25765 335
rect 25785 315 25800 335
rect 25750 285 25800 315
rect 25750 265 25765 285
rect 25785 265 25800 285
rect 25750 235 25800 265
rect 25750 215 25765 235
rect 25785 215 25800 235
rect 25750 185 25800 215
rect 25750 165 25765 185
rect 25785 165 25800 185
rect 25750 135 25800 165
rect 25750 115 25765 135
rect 25785 115 25800 135
rect 25750 85 25800 115
rect 25750 65 25765 85
rect 25785 65 25800 85
rect 25750 50 25800 65
rect 26650 735 26700 750
rect 26650 715 26665 735
rect 26685 715 26700 735
rect 26650 685 26700 715
rect 26650 665 26665 685
rect 26685 665 26700 685
rect 26650 635 26700 665
rect 26650 615 26665 635
rect 26685 615 26700 635
rect 26650 585 26700 615
rect 26650 565 26665 585
rect 26685 565 26700 585
rect 26650 535 26700 565
rect 26650 515 26665 535
rect 26685 515 26700 535
rect 26650 485 26700 515
rect 26650 465 26665 485
rect 26685 465 26700 485
rect 26650 435 26700 465
rect 26650 415 26665 435
rect 26685 415 26700 435
rect 26650 385 26700 415
rect 26650 365 26665 385
rect 26685 365 26700 385
rect 26650 335 26700 365
rect 26650 315 26665 335
rect 26685 315 26700 335
rect 26650 285 26700 315
rect 26650 265 26665 285
rect 26685 265 26700 285
rect 26650 235 26700 265
rect 26650 215 26665 235
rect 26685 215 26700 235
rect 26650 185 26700 215
rect 26650 165 26665 185
rect 26685 165 26700 185
rect 26650 135 26700 165
rect 26650 115 26665 135
rect 26685 115 26700 135
rect 26650 85 26700 115
rect 26650 65 26665 85
rect 26685 65 26700 85
rect 26650 50 26700 65
rect 27550 735 27600 750
rect 27550 715 27565 735
rect 27585 715 27600 735
rect 27550 685 27600 715
rect 27550 665 27565 685
rect 27585 665 27600 685
rect 27550 635 27600 665
rect 27550 615 27565 635
rect 27585 615 27600 635
rect 27550 585 27600 615
rect 27550 565 27565 585
rect 27585 565 27600 585
rect 27550 535 27600 565
rect 27550 515 27565 535
rect 27585 515 27600 535
rect 27550 485 27600 515
rect 27550 465 27565 485
rect 27585 465 27600 485
rect 27550 435 27600 465
rect 27550 415 27565 435
rect 27585 415 27600 435
rect 27550 385 27600 415
rect 27550 365 27565 385
rect 27585 365 27600 385
rect 27550 335 27600 365
rect 27550 315 27565 335
rect 27585 315 27600 335
rect 27550 285 27600 315
rect 27550 265 27565 285
rect 27585 265 27600 285
rect 27550 235 27600 265
rect 27550 215 27565 235
rect 27585 215 27600 235
rect 27550 185 27600 215
rect 27550 165 27565 185
rect 27585 165 27600 185
rect 27550 135 27600 165
rect 27550 115 27565 135
rect 27585 115 27600 135
rect 27550 85 27600 115
rect 27550 65 27565 85
rect 27585 65 27600 85
rect 27550 50 27600 65
rect 28750 735 28800 750
rect 28750 715 28765 735
rect 28785 715 28800 735
rect 28750 685 28800 715
rect 28750 665 28765 685
rect 28785 665 28800 685
rect 28750 635 28800 665
rect 28750 615 28765 635
rect 28785 615 28800 635
rect 28750 585 28800 615
rect 28750 565 28765 585
rect 28785 565 28800 585
rect 28750 535 28800 565
rect 28750 515 28765 535
rect 28785 515 28800 535
rect 28750 485 28800 515
rect 28750 465 28765 485
rect 28785 465 28800 485
rect 28750 435 28800 465
rect 28750 415 28765 435
rect 28785 415 28800 435
rect 28750 385 28800 415
rect 28750 365 28765 385
rect 28785 365 28800 385
rect 28750 335 28800 365
rect 28750 315 28765 335
rect 28785 315 28800 335
rect 28750 285 28800 315
rect 28750 265 28765 285
rect 28785 265 28800 285
rect 28750 235 28800 265
rect 28750 215 28765 235
rect 28785 215 28800 235
rect 28750 185 28800 215
rect 28750 165 28765 185
rect 28785 165 28800 185
rect 28750 135 28800 165
rect 28750 115 28765 135
rect 28785 115 28800 135
rect 28750 85 28800 115
rect 28750 65 28765 85
rect 28785 65 28800 85
rect 28750 50 28800 65
rect -650 -15 28800 0
rect -650 -35 -635 -15
rect -615 -35 -585 -15
rect -565 -35 -535 -15
rect -515 -35 -485 -15
rect -465 -35 -435 -15
rect -415 -35 -385 -15
rect -365 -35 -335 -15
rect -315 -35 -285 -15
rect -265 -35 -235 -15
rect -215 -35 -185 -15
rect -165 -35 -135 -15
rect -115 -35 -85 -15
rect -65 -35 -35 -15
rect -15 -35 15 -15
rect 35 -35 65 -15
rect 85 -35 115 -15
rect 135 -35 165 -15
rect 185 -35 215 -15
rect 235 -35 265 -15
rect 285 -35 315 -15
rect 335 -35 365 -15
rect 385 -35 415 -15
rect 435 -35 465 -15
rect 485 -35 515 -15
rect 535 -35 565 -15
rect 585 -35 615 -15
rect 635 -35 665 -15
rect 685 -35 715 -15
rect 735 -35 765 -15
rect 785 -35 815 -15
rect 835 -35 865 -15
rect 885 -35 915 -15
rect 935 -35 965 -15
rect 985 -35 1015 -15
rect 1035 -35 1065 -15
rect 1085 -35 1115 -15
rect 1135 -35 1165 -15
rect 1185 -35 1215 -15
rect 1235 -35 1265 -15
rect 1285 -35 1315 -15
rect 1335 -35 1365 -15
rect 1385 -35 1415 -15
rect 1435 -35 1465 -15
rect 1485 -35 1515 -15
rect 1535 -35 1565 -15
rect 1585 -35 1615 -15
rect 1635 -35 1665 -15
rect 1685 -35 1715 -15
rect 1735 -35 1765 -15
rect 1785 -35 1815 -15
rect 1835 -35 1865 -15
rect 1885 -35 1915 -15
rect 1935 -35 1965 -15
rect 1985 -35 2015 -15
rect 2035 -35 2065 -15
rect 2085 -35 2115 -15
rect 2135 -35 2165 -15
rect 2185 -35 2215 -15
rect 2235 -35 2265 -15
rect 2285 -35 2315 -15
rect 2335 -35 2365 -15
rect 2385 -35 2415 -15
rect 2435 -35 2465 -15
rect 2485 -35 2515 -15
rect 2535 -35 2565 -15
rect 2585 -35 2615 -15
rect 2635 -35 2665 -15
rect 2685 -35 2715 -15
rect 2735 -35 2765 -15
rect 2785 -35 2815 -15
rect 2835 -35 2865 -15
rect 2885 -35 2915 -15
rect 2935 -35 2965 -15
rect 2985 -35 3015 -15
rect 3035 -35 3065 -15
rect 3085 -35 3115 -15
rect 3135 -35 3165 -15
rect 3185 -35 3215 -15
rect 3235 -35 3265 -15
rect 3285 -35 3315 -15
rect 3335 -35 3365 -15
rect 3385 -35 3415 -15
rect 3435 -35 3465 -15
rect 3485 -35 3515 -15
rect 3535 -35 3565 -15
rect 3585 -35 3615 -15
rect 3635 -35 3665 -15
rect 3685 -35 3715 -15
rect 3735 -35 3765 -15
rect 3785 -35 3815 -15
rect 3835 -35 3865 -15
rect 3885 -35 3915 -15
rect 3935 -35 3965 -15
rect 3985 -35 4015 -15
rect 4035 -35 4065 -15
rect 4085 -35 4115 -15
rect 4135 -35 4165 -15
rect 4185 -35 4215 -15
rect 4235 -35 4265 -15
rect 4285 -35 4315 -15
rect 4335 -35 4365 -15
rect 4385 -35 4415 -15
rect 4435 -35 4465 -15
rect 4485 -35 4515 -15
rect 4535 -35 4565 -15
rect 4585 -35 4615 -15
rect 4635 -35 4665 -15
rect 4685 -35 4715 -15
rect 4735 -35 4765 -15
rect 4785 -35 4815 -15
rect 4835 -35 4865 -15
rect 4885 -35 4915 -15
rect 4935 -35 4965 -15
rect 4985 -35 5015 -15
rect 5035 -35 5065 -15
rect 5085 -35 5115 -15
rect 5135 -35 5165 -15
rect 5185 -35 5215 -15
rect 5235 -35 5265 -15
rect 5285 -35 5315 -15
rect 5335 -35 5365 -15
rect 5385 -35 5415 -15
rect 5435 -35 5465 -15
rect 5485 -35 5515 -15
rect 5535 -35 5565 -15
rect 5585 -35 5615 -15
rect 5635 -35 5665 -15
rect 5685 -35 5715 -15
rect 5735 -35 5765 -15
rect 5785 -35 5815 -15
rect 5835 -35 5865 -15
rect 5885 -35 5915 -15
rect 5935 -35 5965 -15
rect 5985 -35 6015 -15
rect 6035 -35 6065 -15
rect 6085 -35 6115 -15
rect 6135 -35 6165 -15
rect 6185 -35 6215 -15
rect 6235 -35 6265 -15
rect 6285 -35 6315 -15
rect 6335 -35 6365 -15
rect 6385 -35 6415 -15
rect 6435 -35 6465 -15
rect 6485 -35 6515 -15
rect 6535 -35 6565 -15
rect 6585 -35 6615 -15
rect 6635 -35 6665 -15
rect 6685 -35 6715 -15
rect 6735 -35 6765 -15
rect 6785 -35 6815 -15
rect 6835 -35 6865 -15
rect 6885 -35 6915 -15
rect 6935 -35 6965 -15
rect 6985 -35 7015 -15
rect 7035 -35 7065 -15
rect 7085 -35 7115 -15
rect 7135 -35 7165 -15
rect 7185 -35 7215 -15
rect 7235 -35 7265 -15
rect 7285 -35 7315 -15
rect 7335 -35 7365 -15
rect 7385 -35 7415 -15
rect 7435 -35 7465 -15
rect 7485 -35 7515 -15
rect 7535 -35 7565 -15
rect 7585 -35 7615 -15
rect 7635 -35 7665 -15
rect 7685 -35 7715 -15
rect 7735 -35 7765 -15
rect 7785 -35 7815 -15
rect 7835 -35 7865 -15
rect 7885 -35 7915 -15
rect 7935 -35 7965 -15
rect 7985 -35 8015 -15
rect 8035 -35 8065 -15
rect 8085 -35 8115 -15
rect 8135 -35 8165 -15
rect 8185 -35 8215 -15
rect 8235 -35 8265 -15
rect 8285 -35 8315 -15
rect 8335 -35 8365 -15
rect 8385 -35 8415 -15
rect 8435 -35 8465 -15
rect 8485 -35 8515 -15
rect 8535 -35 8565 -15
rect 8585 -35 8615 -15
rect 8635 -35 8665 -15
rect 8685 -35 8715 -15
rect 8735 -35 8765 -15
rect 8785 -35 8815 -15
rect 8835 -35 8865 -15
rect 8885 -35 8915 -15
rect 8935 -35 8965 -15
rect 8985 -35 9015 -15
rect 9035 -35 9065 -15
rect 9085 -35 9115 -15
rect 9135 -35 9165 -15
rect 9185 -35 9215 -15
rect 9235 -35 9265 -15
rect 9285 -35 9315 -15
rect 9335 -35 9365 -15
rect 9385 -35 9415 -15
rect 9435 -35 9465 -15
rect 9485 -35 9515 -15
rect 9535 -35 9565 -15
rect 9585 -35 9615 -15
rect 9635 -35 9665 -15
rect 9685 -35 9715 -15
rect 9735 -35 9765 -15
rect 9785 -35 9815 -15
rect 9835 -35 9865 -15
rect 9885 -35 9915 -15
rect 9935 -35 9965 -15
rect 9985 -35 10015 -15
rect 10035 -35 10065 -15
rect 10085 -35 10115 -15
rect 10135 -35 10165 -15
rect 10185 -35 10215 -15
rect 10235 -35 10265 -15
rect 10285 -35 10315 -15
rect 10335 -35 10365 -15
rect 10385 -35 10415 -15
rect 10435 -35 10465 -15
rect 10485 -35 10515 -15
rect 10535 -35 10565 -15
rect 10585 -35 10615 -15
rect 10635 -35 10665 -15
rect 10685 -35 10715 -15
rect 10735 -35 10765 -15
rect 10785 -35 10815 -15
rect 10835 -35 10865 -15
rect 10885 -35 10915 -15
rect 10935 -35 10965 -15
rect 10985 -35 11015 -15
rect 11035 -35 11065 -15
rect 11085 -35 11115 -15
rect 11135 -35 11165 -15
rect 11185 -35 11215 -15
rect 11235 -35 11265 -15
rect 11285 -35 11315 -15
rect 11335 -35 11365 -15
rect 11385 -35 11415 -15
rect 11435 -35 11465 -15
rect 11485 -35 11515 -15
rect 11535 -35 11565 -15
rect 11585 -35 11615 -15
rect 11635 -35 11665 -15
rect 11685 -35 11715 -15
rect 11735 -35 11765 -15
rect 11785 -35 11815 -15
rect 11835 -35 11865 -15
rect 11885 -35 11915 -15
rect 11935 -35 11965 -15
rect 11985 -35 12015 -15
rect 12035 -35 12065 -15
rect 12085 -35 12115 -15
rect 12135 -35 12165 -15
rect 12185 -35 12215 -15
rect 12235 -35 12265 -15
rect 12285 -35 12315 -15
rect 12335 -35 12365 -15
rect 12385 -35 12415 -15
rect 12435 -35 12465 -15
rect 12485 -35 12515 -15
rect 12535 -35 12565 -15
rect 12585 -35 12615 -15
rect 12635 -35 12665 -15
rect 12685 -35 12715 -15
rect 12735 -35 12765 -15
rect 12785 -35 12815 -15
rect 12835 -35 12865 -15
rect 12885 -35 12915 -15
rect 12935 -35 12965 -15
rect 12985 -35 13015 -15
rect 13035 -35 13065 -15
rect 13085 -35 13115 -15
rect 13135 -35 13165 -15
rect 13185 -35 13215 -15
rect 13235 -35 13265 -15
rect 13285 -35 13315 -15
rect 13335 -35 13365 -15
rect 13385 -35 13415 -15
rect 13435 -35 13465 -15
rect 13485 -35 13515 -15
rect 13535 -35 13565 -15
rect 13585 -35 13615 -15
rect 13635 -35 13665 -15
rect 13685 -35 13715 -15
rect 13735 -35 13765 -15
rect 13785 -35 13815 -15
rect 13835 -35 13865 -15
rect 13885 -35 13915 -15
rect 13935 -35 13965 -15
rect 13985 -35 14015 -15
rect 14035 -35 14065 -15
rect 14085 -35 14115 -15
rect 14135 -35 14165 -15
rect 14185 -35 14215 -15
rect 14235 -35 14265 -15
rect 14285 -35 14315 -15
rect 14335 -35 14365 -15
rect 14385 -35 14415 -15
rect 14435 -35 14465 -15
rect 14485 -35 14515 -15
rect 14535 -35 14565 -15
rect 14585 -35 14615 -15
rect 14635 -35 14665 -15
rect 14685 -35 14715 -15
rect 14735 -35 14765 -15
rect 14785 -35 14815 -15
rect 14835 -35 14865 -15
rect 14885 -35 14915 -15
rect 14935 -35 14965 -15
rect 14985 -35 15015 -15
rect 15035 -35 15065 -15
rect 15085 -35 15115 -15
rect 15135 -35 15165 -15
rect 15185 -35 15215 -15
rect 15235 -35 15265 -15
rect 15285 -35 15315 -15
rect 15335 -35 15365 -15
rect 15385 -35 15415 -15
rect 15435 -35 15465 -15
rect 15485 -35 15515 -15
rect 15535 -35 15565 -15
rect 15585 -35 15615 -15
rect 15635 -35 15665 -15
rect 15685 -35 15715 -15
rect 15735 -35 15765 -15
rect 15785 -35 15815 -15
rect 15835 -35 15865 -15
rect 15885 -35 15915 -15
rect 15935 -35 15965 -15
rect 15985 -35 16015 -15
rect 16035 -35 16065 -15
rect 16085 -35 16115 -15
rect 16135 -35 16165 -15
rect 16185 -35 16215 -15
rect 16235 -35 16265 -15
rect 16285 -35 16315 -15
rect 16335 -35 16365 -15
rect 16385 -35 16415 -15
rect 16435 -35 16465 -15
rect 16485 -35 16515 -15
rect 16535 -35 16565 -15
rect 16585 -35 16615 -15
rect 16635 -35 16665 -15
rect 16685 -35 16715 -15
rect 16735 -35 16765 -15
rect 16785 -35 16815 -15
rect 16835 -35 16865 -15
rect 16885 -35 16915 -15
rect 16935 -35 16965 -15
rect 16985 -35 17015 -15
rect 17035 -35 17065 -15
rect 17085 -35 17115 -15
rect 17135 -35 17165 -15
rect 17185 -35 17215 -15
rect 17235 -35 17265 -15
rect 17285 -35 17315 -15
rect 17335 -35 17365 -15
rect 17385 -35 17415 -15
rect 17435 -35 17465 -15
rect 17485 -35 17515 -15
rect 17535 -35 17565 -15
rect 17585 -35 17615 -15
rect 17635 -35 17665 -15
rect 17685 -35 17715 -15
rect 17735 -35 17765 -15
rect 17785 -35 17815 -15
rect 17835 -35 17865 -15
rect 17885 -35 17915 -15
rect 17935 -35 17965 -15
rect 17985 -35 18015 -15
rect 18035 -35 18065 -15
rect 18085 -35 18115 -15
rect 18135 -35 18165 -15
rect 18185 -35 18215 -15
rect 18235 -35 18265 -15
rect 18285 -35 18315 -15
rect 18335 -35 18365 -15
rect 18385 -35 18415 -15
rect 18435 -35 18465 -15
rect 18485 -35 18515 -15
rect 18535 -35 18565 -15
rect 18585 -35 18615 -15
rect 18635 -35 18665 -15
rect 18685 -35 18715 -15
rect 18735 -35 18765 -15
rect 18785 -35 18815 -15
rect 18835 -35 18865 -15
rect 18885 -35 18915 -15
rect 18935 -35 18965 -15
rect 18985 -35 19015 -15
rect 19035 -35 19065 -15
rect 19085 -35 19115 -15
rect 19135 -35 19165 -15
rect 19185 -35 19215 -15
rect 19235 -35 19265 -15
rect 19285 -35 19315 -15
rect 19335 -35 19365 -15
rect 19385 -35 19415 -15
rect 19435 -35 19465 -15
rect 19485 -35 19515 -15
rect 19535 -35 19565 -15
rect 19585 -35 19615 -15
rect 19635 -35 19665 -15
rect 19685 -35 19715 -15
rect 19735 -35 19765 -15
rect 19785 -35 19815 -15
rect 19835 -35 19865 -15
rect 19885 -35 19915 -15
rect 19935 -35 19965 -15
rect 19985 -35 20015 -15
rect 20035 -35 20065 -15
rect 20085 -35 20115 -15
rect 20135 -35 20165 -15
rect 20185 -35 20215 -15
rect 20235 -35 20265 -15
rect 20285 -35 20315 -15
rect 20335 -35 20365 -15
rect 20385 -35 20415 -15
rect 20435 -35 20465 -15
rect 20485 -35 20515 -15
rect 20535 -35 20565 -15
rect 20585 -35 20615 -15
rect 20635 -35 20665 -15
rect 20685 -35 20715 -15
rect 20735 -35 20765 -15
rect 20785 -35 20815 -15
rect 20835 -35 20865 -15
rect 20885 -35 20915 -15
rect 20935 -35 20965 -15
rect 20985 -35 21015 -15
rect 21035 -35 21065 -15
rect 21085 -35 21115 -15
rect 21135 -35 21165 -15
rect 21185 -35 21215 -15
rect 21235 -35 21265 -15
rect 21285 -35 21315 -15
rect 21335 -35 21365 -15
rect 21385 -35 21415 -15
rect 21435 -35 21465 -15
rect 21485 -35 21515 -15
rect 21535 -35 21565 -15
rect 21585 -35 21615 -15
rect 21635 -35 21665 -15
rect 21685 -35 21715 -15
rect 21735 -35 21765 -15
rect 21785 -35 21815 -15
rect 21835 -35 21865 -15
rect 21885 -35 21915 -15
rect 21935 -35 21965 -15
rect 21985 -35 22015 -15
rect 22035 -35 22065 -15
rect 22085 -35 22115 -15
rect 22135 -35 22165 -15
rect 22185 -35 22215 -15
rect 22235 -35 22265 -15
rect 22285 -35 22315 -15
rect 22335 -35 22365 -15
rect 22385 -35 22415 -15
rect 22435 -35 22465 -15
rect 22485 -35 22515 -15
rect 22535 -35 22565 -15
rect 22585 -35 22615 -15
rect 22635 -35 22665 -15
rect 22685 -35 22715 -15
rect 22735 -35 22765 -15
rect 22785 -35 22815 -15
rect 22835 -35 22865 -15
rect 22885 -35 22915 -15
rect 22935 -35 22965 -15
rect 22985 -35 23015 -15
rect 23035 -35 23065 -15
rect 23085 -35 23115 -15
rect 23135 -35 23165 -15
rect 23185 -35 23215 -15
rect 23235 -35 23265 -15
rect 23285 -35 23315 -15
rect 23335 -35 23365 -15
rect 23385 -35 23415 -15
rect 23435 -35 23465 -15
rect 23485 -35 23515 -15
rect 23535 -35 23565 -15
rect 23585 -35 23615 -15
rect 23635 -35 23665 -15
rect 23685 -35 23715 -15
rect 23735 -35 23765 -15
rect 23785 -35 23815 -15
rect 23835 -35 23865 -15
rect 23885 -35 23915 -15
rect 23935 -35 23965 -15
rect 23985 -35 24015 -15
rect 24035 -35 24065 -15
rect 24085 -35 24115 -15
rect 24135 -35 24165 -15
rect 24185 -35 24215 -15
rect 24235 -35 24265 -15
rect 24285 -35 24315 -15
rect 24335 -35 24365 -15
rect 24385 -35 24415 -15
rect 24435 -35 24465 -15
rect 24485 -35 24515 -15
rect 24535 -35 24565 -15
rect 24585 -35 24615 -15
rect 24635 -35 24665 -15
rect 24685 -35 24715 -15
rect 24735 -35 24765 -15
rect 24785 -35 24815 -15
rect 24835 -35 24865 -15
rect 24885 -35 24915 -15
rect 24935 -35 24965 -15
rect 24985 -35 25015 -15
rect 25035 -35 25065 -15
rect 25085 -35 25115 -15
rect 25135 -35 25165 -15
rect 25185 -35 25215 -15
rect 25235 -35 25265 -15
rect 25285 -35 25315 -15
rect 25335 -35 25365 -15
rect 25385 -35 25415 -15
rect 25435 -35 25465 -15
rect 25485 -35 25515 -15
rect 25535 -35 25565 -15
rect 25585 -35 25615 -15
rect 25635 -35 25665 -15
rect 25685 -35 25715 -15
rect 25735 -35 25765 -15
rect 25785 -35 25815 -15
rect 25835 -35 25865 -15
rect 25885 -35 25915 -15
rect 25935 -35 25965 -15
rect 25985 -35 26015 -15
rect 26035 -35 26065 -15
rect 26085 -35 26115 -15
rect 26135 -35 26165 -15
rect 26185 -35 26215 -15
rect 26235 -35 26265 -15
rect 26285 -35 26315 -15
rect 26335 -35 26365 -15
rect 26385 -35 26415 -15
rect 26435 -35 26465 -15
rect 26485 -35 26515 -15
rect 26535 -35 26565 -15
rect 26585 -35 26615 -15
rect 26635 -35 26665 -15
rect 26685 -35 26715 -15
rect 26735 -35 26765 -15
rect 26785 -35 26815 -15
rect 26835 -35 26865 -15
rect 26885 -35 26915 -15
rect 26935 -35 26965 -15
rect 26985 -35 27015 -15
rect 27035 -35 27065 -15
rect 27085 -35 27115 -15
rect 27135 -35 27165 -15
rect 27185 -35 27215 -15
rect 27235 -35 27265 -15
rect 27285 -35 27315 -15
rect 27335 -35 27365 -15
rect 27385 -35 27415 -15
rect 27435 -35 27465 -15
rect 27485 -35 27515 -15
rect 27535 -35 27565 -15
rect 27585 -35 27615 -15
rect 27635 -35 27665 -15
rect 27685 -35 27715 -15
rect 27735 -35 27765 -15
rect 27785 -35 27815 -15
rect 27835 -35 27865 -15
rect 27885 -35 27915 -15
rect 27935 -35 27965 -15
rect 27985 -35 28015 -15
rect 28035 -35 28065 -15
rect 28085 -35 28115 -15
rect 28135 -35 28165 -15
rect 28185 -35 28215 -15
rect 28235 -35 28265 -15
rect 28285 -35 28315 -15
rect 28335 -35 28365 -15
rect 28385 -35 28415 -15
rect 28435 -35 28465 -15
rect 28485 -35 28515 -15
rect 28535 -35 28565 -15
rect 28585 -35 28615 -15
rect 28635 -35 28665 -15
rect 28685 -35 28715 -15
rect 28735 -35 28765 -15
rect 28785 -35 28800 -15
rect -650 -50 28800 -35
rect -650 -115 -600 -100
rect -650 -135 -635 -115
rect -615 -135 -600 -115
rect -650 -165 -600 -135
rect -650 -185 -635 -165
rect -615 -185 -600 -165
rect -650 -215 -600 -185
rect -650 -235 -635 -215
rect -615 -235 -600 -215
rect -650 -265 -600 -235
rect -650 -285 -635 -265
rect -615 -285 -600 -265
rect -650 -315 -600 -285
rect -650 -335 -635 -315
rect -615 -335 -600 -315
rect -650 -365 -600 -335
rect -650 -385 -635 -365
rect -615 -385 -600 -365
rect -650 -415 -600 -385
rect -650 -435 -635 -415
rect -615 -435 -600 -415
rect -650 -465 -600 -435
rect -650 -485 -635 -465
rect -615 -485 -600 -465
rect -650 -515 -600 -485
rect -650 -535 -635 -515
rect -615 -535 -600 -515
rect -650 -565 -600 -535
rect -650 -585 -635 -565
rect -615 -585 -600 -565
rect -650 -615 -600 -585
rect -650 -635 -635 -615
rect -615 -635 -600 -615
rect -650 -665 -600 -635
rect -650 -685 -635 -665
rect -615 -685 -600 -665
rect -650 -715 -600 -685
rect -650 -735 -635 -715
rect -615 -735 -600 -715
rect -650 -765 -600 -735
rect -650 -785 -635 -765
rect -615 -785 -600 -765
rect -650 -800 -600 -785
rect -500 -115 -450 -100
rect -500 -135 -485 -115
rect -465 -135 -450 -115
rect -500 -165 -450 -135
rect -500 -185 -485 -165
rect -465 -185 -450 -165
rect -500 -215 -450 -185
rect -500 -235 -485 -215
rect -465 -235 -450 -215
rect -500 -265 -450 -235
rect -500 -285 -485 -265
rect -465 -285 -450 -265
rect -500 -315 -450 -285
rect -500 -335 -485 -315
rect -465 -335 -450 -315
rect -500 -365 -450 -335
rect -500 -385 -485 -365
rect -465 -385 -450 -365
rect -500 -415 -450 -385
rect -500 -435 -485 -415
rect -465 -435 -450 -415
rect -500 -465 -450 -435
rect -500 -485 -485 -465
rect -465 -485 -450 -465
rect -500 -515 -450 -485
rect -500 -535 -485 -515
rect -465 -535 -450 -515
rect -500 -565 -450 -535
rect -500 -585 -485 -565
rect -465 -585 -450 -565
rect -500 -615 -450 -585
rect -500 -635 -485 -615
rect -465 -635 -450 -615
rect -500 -665 -450 -635
rect -500 -685 -485 -665
rect -465 -685 -450 -665
rect -500 -715 -450 -685
rect -500 -735 -485 -715
rect -465 -735 -450 -715
rect -500 -765 -450 -735
rect -500 -785 -485 -765
rect -465 -785 -450 -765
rect -500 -800 -450 -785
rect -350 -115 -300 -100
rect -350 -135 -335 -115
rect -315 -135 -300 -115
rect -350 -165 -300 -135
rect -350 -185 -335 -165
rect -315 -185 -300 -165
rect -350 -215 -300 -185
rect -350 -235 -335 -215
rect -315 -235 -300 -215
rect -350 -265 -300 -235
rect -350 -285 -335 -265
rect -315 -285 -300 -265
rect -350 -315 -300 -285
rect -350 -335 -335 -315
rect -315 -335 -300 -315
rect -350 -365 -300 -335
rect -350 -385 -335 -365
rect -315 -385 -300 -365
rect -350 -415 -300 -385
rect -350 -435 -335 -415
rect -315 -435 -300 -415
rect -350 -465 -300 -435
rect -350 -485 -335 -465
rect -315 -485 -300 -465
rect -350 -515 -300 -485
rect -350 -535 -335 -515
rect -315 -535 -300 -515
rect -350 -565 -300 -535
rect -350 -585 -335 -565
rect -315 -585 -300 -565
rect -350 -615 -300 -585
rect -350 -635 -335 -615
rect -315 -635 -300 -615
rect -350 -665 -300 -635
rect -350 -685 -335 -665
rect -315 -685 -300 -665
rect -350 -715 -300 -685
rect -350 -735 -335 -715
rect -315 -735 -300 -715
rect -350 -765 -300 -735
rect -350 -785 -335 -765
rect -315 -785 -300 -765
rect -350 -800 -300 -785
rect -200 -115 -150 -100
rect -200 -135 -185 -115
rect -165 -135 -150 -115
rect -200 -165 -150 -135
rect -200 -185 -185 -165
rect -165 -185 -150 -165
rect -200 -215 -150 -185
rect -200 -235 -185 -215
rect -165 -235 -150 -215
rect -200 -265 -150 -235
rect -200 -285 -185 -265
rect -165 -285 -150 -265
rect -200 -315 -150 -285
rect -200 -335 -185 -315
rect -165 -335 -150 -315
rect -200 -365 -150 -335
rect -200 -385 -185 -365
rect -165 -385 -150 -365
rect -200 -415 -150 -385
rect -200 -435 -185 -415
rect -165 -435 -150 -415
rect -200 -465 -150 -435
rect -200 -485 -185 -465
rect -165 -485 -150 -465
rect -200 -515 -150 -485
rect -200 -535 -185 -515
rect -165 -535 -150 -515
rect -200 -565 -150 -535
rect -200 -585 -185 -565
rect -165 -585 -150 -565
rect -200 -615 -150 -585
rect -200 -635 -185 -615
rect -165 -635 -150 -615
rect -200 -665 -150 -635
rect -200 -685 -185 -665
rect -165 -685 -150 -665
rect -200 -715 -150 -685
rect -200 -735 -185 -715
rect -165 -735 -150 -715
rect -200 -765 -150 -735
rect -200 -785 -185 -765
rect -165 -785 -150 -765
rect -200 -800 -150 -785
rect -50 -115 0 -100
rect -50 -135 -35 -115
rect -15 -135 0 -115
rect -50 -165 0 -135
rect -50 -185 -35 -165
rect -15 -185 0 -165
rect -50 -215 0 -185
rect -50 -235 -35 -215
rect -15 -235 0 -215
rect -50 -265 0 -235
rect -50 -285 -35 -265
rect -15 -285 0 -265
rect -50 -315 0 -285
rect -50 -335 -35 -315
rect -15 -335 0 -315
rect -50 -365 0 -335
rect -50 -385 -35 -365
rect -15 -385 0 -365
rect -50 -415 0 -385
rect -50 -435 -35 -415
rect -15 -435 0 -415
rect -50 -465 0 -435
rect -50 -485 -35 -465
rect -15 -485 0 -465
rect -50 -515 0 -485
rect -50 -535 -35 -515
rect -15 -535 0 -515
rect -50 -565 0 -535
rect -50 -585 -35 -565
rect -15 -585 0 -565
rect -50 -615 0 -585
rect -50 -635 -35 -615
rect -15 -635 0 -615
rect -50 -665 0 -635
rect -50 -685 -35 -665
rect -15 -685 0 -665
rect -50 -715 0 -685
rect -50 -735 -35 -715
rect -15 -735 0 -715
rect -50 -765 0 -735
rect -50 -785 -35 -765
rect -15 -785 0 -765
rect -50 -800 0 -785
rect 1150 -115 1200 -100
rect 1150 -135 1165 -115
rect 1185 -135 1200 -115
rect 1150 -165 1200 -135
rect 1150 -185 1165 -165
rect 1185 -185 1200 -165
rect 1150 -215 1200 -185
rect 1150 -235 1165 -215
rect 1185 -235 1200 -215
rect 1150 -265 1200 -235
rect 1150 -285 1165 -265
rect 1185 -285 1200 -265
rect 1150 -315 1200 -285
rect 1150 -335 1165 -315
rect 1185 -335 1200 -315
rect 1150 -365 1200 -335
rect 1150 -385 1165 -365
rect 1185 -385 1200 -365
rect 1150 -415 1200 -385
rect 1150 -435 1165 -415
rect 1185 -435 1200 -415
rect 1150 -465 1200 -435
rect 1150 -485 1165 -465
rect 1185 -485 1200 -465
rect 1150 -515 1200 -485
rect 1150 -535 1165 -515
rect 1185 -535 1200 -515
rect 1150 -565 1200 -535
rect 1150 -585 1165 -565
rect 1185 -585 1200 -565
rect 1150 -615 1200 -585
rect 1150 -635 1165 -615
rect 1185 -635 1200 -615
rect 1150 -665 1200 -635
rect 1150 -685 1165 -665
rect 1185 -685 1200 -665
rect 1150 -715 1200 -685
rect 1150 -735 1165 -715
rect 1185 -735 1200 -715
rect 1150 -765 1200 -735
rect 1150 -785 1165 -765
rect 1185 -785 1200 -765
rect 1150 -800 1200 -785
rect 1450 -115 1500 -100
rect 1450 -135 1465 -115
rect 1485 -135 1500 -115
rect 1450 -165 1500 -135
rect 1450 -185 1465 -165
rect 1485 -185 1500 -165
rect 1450 -215 1500 -185
rect 1450 -235 1465 -215
rect 1485 -235 1500 -215
rect 1450 -265 1500 -235
rect 1450 -285 1465 -265
rect 1485 -285 1500 -265
rect 1450 -315 1500 -285
rect 1450 -335 1465 -315
rect 1485 -335 1500 -315
rect 1450 -365 1500 -335
rect 1450 -385 1465 -365
rect 1485 -385 1500 -365
rect 1450 -415 1500 -385
rect 1450 -435 1465 -415
rect 1485 -435 1500 -415
rect 1450 -465 1500 -435
rect 1450 -485 1465 -465
rect 1485 -485 1500 -465
rect 1450 -515 1500 -485
rect 1450 -535 1465 -515
rect 1485 -535 1500 -515
rect 1450 -565 1500 -535
rect 1450 -585 1465 -565
rect 1485 -585 1500 -565
rect 1450 -615 1500 -585
rect 1450 -635 1465 -615
rect 1485 -635 1500 -615
rect 1450 -665 1500 -635
rect 1450 -685 1465 -665
rect 1485 -685 1500 -665
rect 1450 -715 1500 -685
rect 1450 -735 1465 -715
rect 1485 -735 1500 -715
rect 1450 -765 1500 -735
rect 1450 -785 1465 -765
rect 1485 -785 1500 -765
rect 1450 -800 1500 -785
rect 1750 -115 1800 -100
rect 1750 -135 1765 -115
rect 1785 -135 1800 -115
rect 1750 -165 1800 -135
rect 1750 -185 1765 -165
rect 1785 -185 1800 -165
rect 1750 -215 1800 -185
rect 1750 -235 1765 -215
rect 1785 -235 1800 -215
rect 1750 -265 1800 -235
rect 1750 -285 1765 -265
rect 1785 -285 1800 -265
rect 1750 -315 1800 -285
rect 1750 -335 1765 -315
rect 1785 -335 1800 -315
rect 1750 -365 1800 -335
rect 1750 -385 1765 -365
rect 1785 -385 1800 -365
rect 1750 -415 1800 -385
rect 1750 -435 1765 -415
rect 1785 -435 1800 -415
rect 1750 -465 1800 -435
rect 1750 -485 1765 -465
rect 1785 -485 1800 -465
rect 1750 -515 1800 -485
rect 1750 -535 1765 -515
rect 1785 -535 1800 -515
rect 1750 -565 1800 -535
rect 1750 -585 1765 -565
rect 1785 -585 1800 -565
rect 1750 -615 1800 -585
rect 1750 -635 1765 -615
rect 1785 -635 1800 -615
rect 1750 -665 1800 -635
rect 1750 -685 1765 -665
rect 1785 -685 1800 -665
rect 1750 -715 1800 -685
rect 1750 -735 1765 -715
rect 1785 -735 1800 -715
rect 1750 -765 1800 -735
rect 1750 -785 1765 -765
rect 1785 -785 1800 -765
rect 1750 -800 1800 -785
rect 2050 -115 2100 -100
rect 2050 -135 2065 -115
rect 2085 -135 2100 -115
rect 2050 -165 2100 -135
rect 2050 -185 2065 -165
rect 2085 -185 2100 -165
rect 2050 -215 2100 -185
rect 2050 -235 2065 -215
rect 2085 -235 2100 -215
rect 2050 -265 2100 -235
rect 2050 -285 2065 -265
rect 2085 -285 2100 -265
rect 2050 -315 2100 -285
rect 2050 -335 2065 -315
rect 2085 -335 2100 -315
rect 2050 -365 2100 -335
rect 2050 -385 2065 -365
rect 2085 -385 2100 -365
rect 2050 -415 2100 -385
rect 2050 -435 2065 -415
rect 2085 -435 2100 -415
rect 2050 -465 2100 -435
rect 2050 -485 2065 -465
rect 2085 -485 2100 -465
rect 2050 -515 2100 -485
rect 2050 -535 2065 -515
rect 2085 -535 2100 -515
rect 2050 -565 2100 -535
rect 2050 -585 2065 -565
rect 2085 -585 2100 -565
rect 2050 -615 2100 -585
rect 2050 -635 2065 -615
rect 2085 -635 2100 -615
rect 2050 -665 2100 -635
rect 2050 -685 2065 -665
rect 2085 -685 2100 -665
rect 2050 -715 2100 -685
rect 2050 -735 2065 -715
rect 2085 -735 2100 -715
rect 2050 -765 2100 -735
rect 2050 -785 2065 -765
rect 2085 -785 2100 -765
rect 2050 -800 2100 -785
rect 2350 -115 2400 -100
rect 2350 -135 2365 -115
rect 2385 -135 2400 -115
rect 2350 -165 2400 -135
rect 2350 -185 2365 -165
rect 2385 -185 2400 -165
rect 2350 -215 2400 -185
rect 2350 -235 2365 -215
rect 2385 -235 2400 -215
rect 2350 -265 2400 -235
rect 2350 -285 2365 -265
rect 2385 -285 2400 -265
rect 2350 -315 2400 -285
rect 2350 -335 2365 -315
rect 2385 -335 2400 -315
rect 2350 -365 2400 -335
rect 2350 -385 2365 -365
rect 2385 -385 2400 -365
rect 2350 -415 2400 -385
rect 2350 -435 2365 -415
rect 2385 -435 2400 -415
rect 2350 -465 2400 -435
rect 2350 -485 2365 -465
rect 2385 -485 2400 -465
rect 2350 -515 2400 -485
rect 2350 -535 2365 -515
rect 2385 -535 2400 -515
rect 2350 -565 2400 -535
rect 2350 -585 2365 -565
rect 2385 -585 2400 -565
rect 2350 -615 2400 -585
rect 2350 -635 2365 -615
rect 2385 -635 2400 -615
rect 2350 -665 2400 -635
rect 2350 -685 2365 -665
rect 2385 -685 2400 -665
rect 2350 -715 2400 -685
rect 2350 -735 2365 -715
rect 2385 -735 2400 -715
rect 2350 -765 2400 -735
rect 2350 -785 2365 -765
rect 2385 -785 2400 -765
rect 2350 -800 2400 -785
rect 2650 -115 2700 -100
rect 2650 -135 2665 -115
rect 2685 -135 2700 -115
rect 2650 -165 2700 -135
rect 2650 -185 2665 -165
rect 2685 -185 2700 -165
rect 2650 -215 2700 -185
rect 2650 -235 2665 -215
rect 2685 -235 2700 -215
rect 2650 -265 2700 -235
rect 2650 -285 2665 -265
rect 2685 -285 2700 -265
rect 2650 -315 2700 -285
rect 2650 -335 2665 -315
rect 2685 -335 2700 -315
rect 2650 -365 2700 -335
rect 2650 -385 2665 -365
rect 2685 -385 2700 -365
rect 2650 -415 2700 -385
rect 2650 -435 2665 -415
rect 2685 -435 2700 -415
rect 2650 -465 2700 -435
rect 2650 -485 2665 -465
rect 2685 -485 2700 -465
rect 2650 -515 2700 -485
rect 2650 -535 2665 -515
rect 2685 -535 2700 -515
rect 2650 -565 2700 -535
rect 2650 -585 2665 -565
rect 2685 -585 2700 -565
rect 2650 -615 2700 -585
rect 2650 -635 2665 -615
rect 2685 -635 2700 -615
rect 2650 -665 2700 -635
rect 2650 -685 2665 -665
rect 2685 -685 2700 -665
rect 2650 -715 2700 -685
rect 2650 -735 2665 -715
rect 2685 -735 2700 -715
rect 2650 -765 2700 -735
rect 2650 -785 2665 -765
rect 2685 -785 2700 -765
rect 2650 -800 2700 -785
rect 2950 -115 3000 -100
rect 2950 -135 2965 -115
rect 2985 -135 3000 -115
rect 2950 -165 3000 -135
rect 2950 -185 2965 -165
rect 2985 -185 3000 -165
rect 2950 -215 3000 -185
rect 2950 -235 2965 -215
rect 2985 -235 3000 -215
rect 2950 -265 3000 -235
rect 2950 -285 2965 -265
rect 2985 -285 3000 -265
rect 2950 -315 3000 -285
rect 2950 -335 2965 -315
rect 2985 -335 3000 -315
rect 2950 -365 3000 -335
rect 2950 -385 2965 -365
rect 2985 -385 3000 -365
rect 2950 -415 3000 -385
rect 2950 -435 2965 -415
rect 2985 -435 3000 -415
rect 2950 -465 3000 -435
rect 2950 -485 2965 -465
rect 2985 -485 3000 -465
rect 2950 -515 3000 -485
rect 2950 -535 2965 -515
rect 2985 -535 3000 -515
rect 2950 -565 3000 -535
rect 2950 -585 2965 -565
rect 2985 -585 3000 -565
rect 2950 -615 3000 -585
rect 2950 -635 2965 -615
rect 2985 -635 3000 -615
rect 2950 -665 3000 -635
rect 2950 -685 2965 -665
rect 2985 -685 3000 -665
rect 2950 -715 3000 -685
rect 2950 -735 2965 -715
rect 2985 -735 3000 -715
rect 2950 -765 3000 -735
rect 2950 -785 2965 -765
rect 2985 -785 3000 -765
rect 2950 -800 3000 -785
rect 3250 -115 3300 -100
rect 3250 -135 3265 -115
rect 3285 -135 3300 -115
rect 3250 -165 3300 -135
rect 3250 -185 3265 -165
rect 3285 -185 3300 -165
rect 3250 -215 3300 -185
rect 3250 -235 3265 -215
rect 3285 -235 3300 -215
rect 3250 -265 3300 -235
rect 3250 -285 3265 -265
rect 3285 -285 3300 -265
rect 3250 -315 3300 -285
rect 3250 -335 3265 -315
rect 3285 -335 3300 -315
rect 3250 -365 3300 -335
rect 3250 -385 3265 -365
rect 3285 -385 3300 -365
rect 3250 -415 3300 -385
rect 3250 -435 3265 -415
rect 3285 -435 3300 -415
rect 3250 -465 3300 -435
rect 3250 -485 3265 -465
rect 3285 -485 3300 -465
rect 3250 -515 3300 -485
rect 3250 -535 3265 -515
rect 3285 -535 3300 -515
rect 3250 -565 3300 -535
rect 3250 -585 3265 -565
rect 3285 -585 3300 -565
rect 3250 -615 3300 -585
rect 3250 -635 3265 -615
rect 3285 -635 3300 -615
rect 3250 -665 3300 -635
rect 3250 -685 3265 -665
rect 3285 -685 3300 -665
rect 3250 -715 3300 -685
rect 3250 -735 3265 -715
rect 3285 -735 3300 -715
rect 3250 -765 3300 -735
rect 3250 -785 3265 -765
rect 3285 -785 3300 -765
rect 3250 -800 3300 -785
rect 3550 -115 3600 -100
rect 3550 -135 3565 -115
rect 3585 -135 3600 -115
rect 3550 -165 3600 -135
rect 3550 -185 3565 -165
rect 3585 -185 3600 -165
rect 3550 -215 3600 -185
rect 3550 -235 3565 -215
rect 3585 -235 3600 -215
rect 3550 -265 3600 -235
rect 3550 -285 3565 -265
rect 3585 -285 3600 -265
rect 3550 -315 3600 -285
rect 3550 -335 3565 -315
rect 3585 -335 3600 -315
rect 3550 -365 3600 -335
rect 3550 -385 3565 -365
rect 3585 -385 3600 -365
rect 3550 -415 3600 -385
rect 3550 -435 3565 -415
rect 3585 -435 3600 -415
rect 3550 -465 3600 -435
rect 3550 -485 3565 -465
rect 3585 -485 3600 -465
rect 3550 -515 3600 -485
rect 3550 -535 3565 -515
rect 3585 -535 3600 -515
rect 3550 -565 3600 -535
rect 3550 -585 3565 -565
rect 3585 -585 3600 -565
rect 3550 -615 3600 -585
rect 3550 -635 3565 -615
rect 3585 -635 3600 -615
rect 3550 -665 3600 -635
rect 3550 -685 3565 -665
rect 3585 -685 3600 -665
rect 3550 -715 3600 -685
rect 3550 -735 3565 -715
rect 3585 -735 3600 -715
rect 3550 -765 3600 -735
rect 3550 -785 3565 -765
rect 3585 -785 3600 -765
rect 3550 -800 3600 -785
rect 3700 -115 3750 -100
rect 3700 -135 3715 -115
rect 3735 -135 3750 -115
rect 3700 -165 3750 -135
rect 3700 -185 3715 -165
rect 3735 -185 3750 -165
rect 3700 -215 3750 -185
rect 3700 -235 3715 -215
rect 3735 -235 3750 -215
rect 3700 -265 3750 -235
rect 3700 -285 3715 -265
rect 3735 -285 3750 -265
rect 3700 -315 3750 -285
rect 3700 -335 3715 -315
rect 3735 -335 3750 -315
rect 3700 -365 3750 -335
rect 3700 -385 3715 -365
rect 3735 -385 3750 -365
rect 3700 -415 3750 -385
rect 3700 -435 3715 -415
rect 3735 -435 3750 -415
rect 3700 -465 3750 -435
rect 3700 -485 3715 -465
rect 3735 -485 3750 -465
rect 3700 -515 3750 -485
rect 3700 -535 3715 -515
rect 3735 -535 3750 -515
rect 3700 -565 3750 -535
rect 3700 -585 3715 -565
rect 3735 -585 3750 -565
rect 3700 -615 3750 -585
rect 3700 -635 3715 -615
rect 3735 -635 3750 -615
rect 3700 -665 3750 -635
rect 3700 -685 3715 -665
rect 3735 -685 3750 -665
rect 3700 -715 3750 -685
rect 3700 -735 3715 -715
rect 3735 -735 3750 -715
rect 3700 -765 3750 -735
rect 3700 -785 3715 -765
rect 3735 -785 3750 -765
rect 3700 -800 3750 -785
rect 3850 -115 3900 -100
rect 3850 -135 3865 -115
rect 3885 -135 3900 -115
rect 3850 -165 3900 -135
rect 3850 -185 3865 -165
rect 3885 -185 3900 -165
rect 3850 -215 3900 -185
rect 3850 -235 3865 -215
rect 3885 -235 3900 -215
rect 3850 -265 3900 -235
rect 3850 -285 3865 -265
rect 3885 -285 3900 -265
rect 3850 -315 3900 -285
rect 3850 -335 3865 -315
rect 3885 -335 3900 -315
rect 3850 -365 3900 -335
rect 3850 -385 3865 -365
rect 3885 -385 3900 -365
rect 3850 -415 3900 -385
rect 3850 -435 3865 -415
rect 3885 -435 3900 -415
rect 3850 -465 3900 -435
rect 3850 -485 3865 -465
rect 3885 -485 3900 -465
rect 3850 -515 3900 -485
rect 3850 -535 3865 -515
rect 3885 -535 3900 -515
rect 3850 -565 3900 -535
rect 3850 -585 3865 -565
rect 3885 -585 3900 -565
rect 3850 -615 3900 -585
rect 3850 -635 3865 -615
rect 3885 -635 3900 -615
rect 3850 -665 3900 -635
rect 3850 -685 3865 -665
rect 3885 -685 3900 -665
rect 3850 -715 3900 -685
rect 3850 -735 3865 -715
rect 3885 -735 3900 -715
rect 3850 -765 3900 -735
rect 3850 -785 3865 -765
rect 3885 -785 3900 -765
rect 3850 -800 3900 -785
rect 4000 -115 4050 -100
rect 4000 -135 4015 -115
rect 4035 -135 4050 -115
rect 4000 -165 4050 -135
rect 4000 -185 4015 -165
rect 4035 -185 4050 -165
rect 4000 -215 4050 -185
rect 4000 -235 4015 -215
rect 4035 -235 4050 -215
rect 4000 -265 4050 -235
rect 4000 -285 4015 -265
rect 4035 -285 4050 -265
rect 4000 -315 4050 -285
rect 4000 -335 4015 -315
rect 4035 -335 4050 -315
rect 4000 -365 4050 -335
rect 4000 -385 4015 -365
rect 4035 -385 4050 -365
rect 4000 -415 4050 -385
rect 4000 -435 4015 -415
rect 4035 -435 4050 -415
rect 4000 -465 4050 -435
rect 4000 -485 4015 -465
rect 4035 -485 4050 -465
rect 4000 -515 4050 -485
rect 4000 -535 4015 -515
rect 4035 -535 4050 -515
rect 4000 -565 4050 -535
rect 4000 -585 4015 -565
rect 4035 -585 4050 -565
rect 4000 -615 4050 -585
rect 4000 -635 4015 -615
rect 4035 -635 4050 -615
rect 4000 -665 4050 -635
rect 4000 -685 4015 -665
rect 4035 -685 4050 -665
rect 4000 -715 4050 -685
rect 4000 -735 4015 -715
rect 4035 -735 4050 -715
rect 4000 -765 4050 -735
rect 4000 -785 4015 -765
rect 4035 -785 4050 -765
rect 4000 -800 4050 -785
rect 4150 -115 4200 -100
rect 4150 -135 4165 -115
rect 4185 -135 4200 -115
rect 4150 -165 4200 -135
rect 4150 -185 4165 -165
rect 4185 -185 4200 -165
rect 4150 -215 4200 -185
rect 4150 -235 4165 -215
rect 4185 -235 4200 -215
rect 4150 -265 4200 -235
rect 4150 -285 4165 -265
rect 4185 -285 4200 -265
rect 4150 -315 4200 -285
rect 4150 -335 4165 -315
rect 4185 -335 4200 -315
rect 4150 -365 4200 -335
rect 4150 -385 4165 -365
rect 4185 -385 4200 -365
rect 4150 -415 4200 -385
rect 4150 -435 4165 -415
rect 4185 -435 4200 -415
rect 4150 -465 4200 -435
rect 4150 -485 4165 -465
rect 4185 -485 4200 -465
rect 4150 -515 4200 -485
rect 4150 -535 4165 -515
rect 4185 -535 4200 -515
rect 4150 -565 4200 -535
rect 4150 -585 4165 -565
rect 4185 -585 4200 -565
rect 4150 -615 4200 -585
rect 4150 -635 4165 -615
rect 4185 -635 4200 -615
rect 4150 -665 4200 -635
rect 4150 -685 4165 -665
rect 4185 -685 4200 -665
rect 4150 -715 4200 -685
rect 4150 -735 4165 -715
rect 4185 -735 4200 -715
rect 4150 -765 4200 -735
rect 4150 -785 4165 -765
rect 4185 -785 4200 -765
rect 4150 -800 4200 -785
rect 4300 -115 4350 -100
rect 4300 -135 4315 -115
rect 4335 -135 4350 -115
rect 4300 -165 4350 -135
rect 4300 -185 4315 -165
rect 4335 -185 4350 -165
rect 4300 -215 4350 -185
rect 4300 -235 4315 -215
rect 4335 -235 4350 -215
rect 4300 -265 4350 -235
rect 4300 -285 4315 -265
rect 4335 -285 4350 -265
rect 4300 -315 4350 -285
rect 4300 -335 4315 -315
rect 4335 -335 4350 -315
rect 4300 -365 4350 -335
rect 4300 -385 4315 -365
rect 4335 -385 4350 -365
rect 4300 -415 4350 -385
rect 4300 -435 4315 -415
rect 4335 -435 4350 -415
rect 4300 -465 4350 -435
rect 4300 -485 4315 -465
rect 4335 -485 4350 -465
rect 4300 -515 4350 -485
rect 4300 -535 4315 -515
rect 4335 -535 4350 -515
rect 4300 -565 4350 -535
rect 4300 -585 4315 -565
rect 4335 -585 4350 -565
rect 4300 -615 4350 -585
rect 4300 -635 4315 -615
rect 4335 -635 4350 -615
rect 4300 -665 4350 -635
rect 4300 -685 4315 -665
rect 4335 -685 4350 -665
rect 4300 -715 4350 -685
rect 4300 -735 4315 -715
rect 4335 -735 4350 -715
rect 4300 -765 4350 -735
rect 4300 -785 4315 -765
rect 4335 -785 4350 -765
rect 4300 -800 4350 -785
rect 4450 -115 4500 -100
rect 4450 -135 4465 -115
rect 4485 -135 4500 -115
rect 4450 -165 4500 -135
rect 4450 -185 4465 -165
rect 4485 -185 4500 -165
rect 4450 -215 4500 -185
rect 4450 -235 4465 -215
rect 4485 -235 4500 -215
rect 4450 -265 4500 -235
rect 4450 -285 4465 -265
rect 4485 -285 4500 -265
rect 4450 -315 4500 -285
rect 4450 -335 4465 -315
rect 4485 -335 4500 -315
rect 4450 -365 4500 -335
rect 4450 -385 4465 -365
rect 4485 -385 4500 -365
rect 4450 -415 4500 -385
rect 4450 -435 4465 -415
rect 4485 -435 4500 -415
rect 4450 -465 4500 -435
rect 4450 -485 4465 -465
rect 4485 -485 4500 -465
rect 4450 -515 4500 -485
rect 4450 -535 4465 -515
rect 4485 -535 4500 -515
rect 4450 -565 4500 -535
rect 4450 -585 4465 -565
rect 4485 -585 4500 -565
rect 4450 -615 4500 -585
rect 4450 -635 4465 -615
rect 4485 -635 4500 -615
rect 4450 -665 4500 -635
rect 4450 -685 4465 -665
rect 4485 -685 4500 -665
rect 4450 -715 4500 -685
rect 4450 -735 4465 -715
rect 4485 -735 4500 -715
rect 4450 -765 4500 -735
rect 4450 -785 4465 -765
rect 4485 -785 4500 -765
rect 4450 -800 4500 -785
rect 4600 -115 4650 -100
rect 4600 -135 4615 -115
rect 4635 -135 4650 -115
rect 4600 -165 4650 -135
rect 4600 -185 4615 -165
rect 4635 -185 4650 -165
rect 4600 -215 4650 -185
rect 4600 -235 4615 -215
rect 4635 -235 4650 -215
rect 4600 -265 4650 -235
rect 4600 -285 4615 -265
rect 4635 -285 4650 -265
rect 4600 -315 4650 -285
rect 4600 -335 4615 -315
rect 4635 -335 4650 -315
rect 4600 -365 4650 -335
rect 4600 -385 4615 -365
rect 4635 -385 4650 -365
rect 4600 -415 4650 -385
rect 4600 -435 4615 -415
rect 4635 -435 4650 -415
rect 4600 -465 4650 -435
rect 4600 -485 4615 -465
rect 4635 -485 4650 -465
rect 4600 -515 4650 -485
rect 4600 -535 4615 -515
rect 4635 -535 4650 -515
rect 4600 -565 4650 -535
rect 4600 -585 4615 -565
rect 4635 -585 4650 -565
rect 4600 -615 4650 -585
rect 4600 -635 4615 -615
rect 4635 -635 4650 -615
rect 4600 -665 4650 -635
rect 4600 -685 4615 -665
rect 4635 -685 4650 -665
rect 4600 -715 4650 -685
rect 4600 -735 4615 -715
rect 4635 -735 4650 -715
rect 4600 -765 4650 -735
rect 4600 -785 4615 -765
rect 4635 -785 4650 -765
rect 4600 -800 4650 -785
rect 4750 -115 4800 -100
rect 4750 -135 4765 -115
rect 4785 -135 4800 -115
rect 4750 -165 4800 -135
rect 4750 -185 4765 -165
rect 4785 -185 4800 -165
rect 4750 -215 4800 -185
rect 4750 -235 4765 -215
rect 4785 -235 4800 -215
rect 4750 -265 4800 -235
rect 4750 -285 4765 -265
rect 4785 -285 4800 -265
rect 4750 -315 4800 -285
rect 4750 -335 4765 -315
rect 4785 -335 4800 -315
rect 4750 -365 4800 -335
rect 4750 -385 4765 -365
rect 4785 -385 4800 -365
rect 4750 -415 4800 -385
rect 4750 -435 4765 -415
rect 4785 -435 4800 -415
rect 4750 -465 4800 -435
rect 4750 -485 4765 -465
rect 4785 -485 4800 -465
rect 4750 -515 4800 -485
rect 4750 -535 4765 -515
rect 4785 -535 4800 -515
rect 4750 -565 4800 -535
rect 4750 -585 4765 -565
rect 4785 -585 4800 -565
rect 4750 -615 4800 -585
rect 4750 -635 4765 -615
rect 4785 -635 4800 -615
rect 4750 -665 4800 -635
rect 4750 -685 4765 -665
rect 4785 -685 4800 -665
rect 4750 -715 4800 -685
rect 4750 -735 4765 -715
rect 4785 -735 4800 -715
rect 4750 -765 4800 -735
rect 4750 -785 4765 -765
rect 4785 -785 4800 -765
rect 4750 -800 4800 -785
rect 5050 -115 5100 -100
rect 5050 -135 5065 -115
rect 5085 -135 5100 -115
rect 5050 -165 5100 -135
rect 5050 -185 5065 -165
rect 5085 -185 5100 -165
rect 5050 -215 5100 -185
rect 5050 -235 5065 -215
rect 5085 -235 5100 -215
rect 5050 -265 5100 -235
rect 5050 -285 5065 -265
rect 5085 -285 5100 -265
rect 5050 -315 5100 -285
rect 5050 -335 5065 -315
rect 5085 -335 5100 -315
rect 5050 -365 5100 -335
rect 5050 -385 5065 -365
rect 5085 -385 5100 -365
rect 5050 -415 5100 -385
rect 5050 -435 5065 -415
rect 5085 -435 5100 -415
rect 5050 -465 5100 -435
rect 5050 -485 5065 -465
rect 5085 -485 5100 -465
rect 5050 -515 5100 -485
rect 5050 -535 5065 -515
rect 5085 -535 5100 -515
rect 5050 -565 5100 -535
rect 5050 -585 5065 -565
rect 5085 -585 5100 -565
rect 5050 -615 5100 -585
rect 5050 -635 5065 -615
rect 5085 -635 5100 -615
rect 5050 -665 5100 -635
rect 5050 -685 5065 -665
rect 5085 -685 5100 -665
rect 5050 -715 5100 -685
rect 5050 -735 5065 -715
rect 5085 -735 5100 -715
rect 5050 -765 5100 -735
rect 5050 -785 5065 -765
rect 5085 -785 5100 -765
rect 5050 -800 5100 -785
rect 5350 -115 5400 -100
rect 5350 -135 5365 -115
rect 5385 -135 5400 -115
rect 5350 -165 5400 -135
rect 5350 -185 5365 -165
rect 5385 -185 5400 -165
rect 5350 -215 5400 -185
rect 5350 -235 5365 -215
rect 5385 -235 5400 -215
rect 5350 -265 5400 -235
rect 5350 -285 5365 -265
rect 5385 -285 5400 -265
rect 5350 -315 5400 -285
rect 5350 -335 5365 -315
rect 5385 -335 5400 -315
rect 5350 -365 5400 -335
rect 5350 -385 5365 -365
rect 5385 -385 5400 -365
rect 5350 -415 5400 -385
rect 5350 -435 5365 -415
rect 5385 -435 5400 -415
rect 5350 -465 5400 -435
rect 5350 -485 5365 -465
rect 5385 -485 5400 -465
rect 5350 -515 5400 -485
rect 5350 -535 5365 -515
rect 5385 -535 5400 -515
rect 5350 -565 5400 -535
rect 5350 -585 5365 -565
rect 5385 -585 5400 -565
rect 5350 -615 5400 -585
rect 5350 -635 5365 -615
rect 5385 -635 5400 -615
rect 5350 -665 5400 -635
rect 5350 -685 5365 -665
rect 5385 -685 5400 -665
rect 5350 -715 5400 -685
rect 5350 -735 5365 -715
rect 5385 -735 5400 -715
rect 5350 -765 5400 -735
rect 5350 -785 5365 -765
rect 5385 -785 5400 -765
rect 5350 -800 5400 -785
rect 5650 -115 5700 -100
rect 5650 -135 5665 -115
rect 5685 -135 5700 -115
rect 5650 -165 5700 -135
rect 5650 -185 5665 -165
rect 5685 -185 5700 -165
rect 5650 -215 5700 -185
rect 5650 -235 5665 -215
rect 5685 -235 5700 -215
rect 5650 -265 5700 -235
rect 5650 -285 5665 -265
rect 5685 -285 5700 -265
rect 5650 -315 5700 -285
rect 5650 -335 5665 -315
rect 5685 -335 5700 -315
rect 5650 -365 5700 -335
rect 5650 -385 5665 -365
rect 5685 -385 5700 -365
rect 5650 -415 5700 -385
rect 5650 -435 5665 -415
rect 5685 -435 5700 -415
rect 5650 -465 5700 -435
rect 5650 -485 5665 -465
rect 5685 -485 5700 -465
rect 5650 -515 5700 -485
rect 5650 -535 5665 -515
rect 5685 -535 5700 -515
rect 5650 -565 5700 -535
rect 5650 -585 5665 -565
rect 5685 -585 5700 -565
rect 5650 -615 5700 -585
rect 5650 -635 5665 -615
rect 5685 -635 5700 -615
rect 5650 -665 5700 -635
rect 5650 -685 5665 -665
rect 5685 -685 5700 -665
rect 5650 -715 5700 -685
rect 5650 -735 5665 -715
rect 5685 -735 5700 -715
rect 5650 -765 5700 -735
rect 5650 -785 5665 -765
rect 5685 -785 5700 -765
rect 5650 -800 5700 -785
rect 5950 -115 6000 -100
rect 5950 -135 5965 -115
rect 5985 -135 6000 -115
rect 5950 -165 6000 -135
rect 5950 -185 5965 -165
rect 5985 -185 6000 -165
rect 5950 -215 6000 -185
rect 5950 -235 5965 -215
rect 5985 -235 6000 -215
rect 5950 -265 6000 -235
rect 5950 -285 5965 -265
rect 5985 -285 6000 -265
rect 5950 -315 6000 -285
rect 5950 -335 5965 -315
rect 5985 -335 6000 -315
rect 5950 -365 6000 -335
rect 5950 -385 5965 -365
rect 5985 -385 6000 -365
rect 5950 -415 6000 -385
rect 5950 -435 5965 -415
rect 5985 -435 6000 -415
rect 5950 -465 6000 -435
rect 5950 -485 5965 -465
rect 5985 -485 6000 -465
rect 5950 -515 6000 -485
rect 5950 -535 5965 -515
rect 5985 -535 6000 -515
rect 5950 -565 6000 -535
rect 5950 -585 5965 -565
rect 5985 -585 6000 -565
rect 5950 -615 6000 -585
rect 5950 -635 5965 -615
rect 5985 -635 6000 -615
rect 5950 -665 6000 -635
rect 5950 -685 5965 -665
rect 5985 -685 6000 -665
rect 5950 -715 6000 -685
rect 5950 -735 5965 -715
rect 5985 -735 6000 -715
rect 5950 -765 6000 -735
rect 5950 -785 5965 -765
rect 5985 -785 6000 -765
rect 5950 -800 6000 -785
rect 6250 -115 6300 -100
rect 6250 -135 6265 -115
rect 6285 -135 6300 -115
rect 6250 -165 6300 -135
rect 6250 -185 6265 -165
rect 6285 -185 6300 -165
rect 6250 -215 6300 -185
rect 6250 -235 6265 -215
rect 6285 -235 6300 -215
rect 6250 -265 6300 -235
rect 6250 -285 6265 -265
rect 6285 -285 6300 -265
rect 6250 -315 6300 -285
rect 6250 -335 6265 -315
rect 6285 -335 6300 -315
rect 6250 -365 6300 -335
rect 6250 -385 6265 -365
rect 6285 -385 6300 -365
rect 6250 -415 6300 -385
rect 6250 -435 6265 -415
rect 6285 -435 6300 -415
rect 6250 -465 6300 -435
rect 6250 -485 6265 -465
rect 6285 -485 6300 -465
rect 6250 -515 6300 -485
rect 6250 -535 6265 -515
rect 6285 -535 6300 -515
rect 6250 -565 6300 -535
rect 6250 -585 6265 -565
rect 6285 -585 6300 -565
rect 6250 -615 6300 -585
rect 6250 -635 6265 -615
rect 6285 -635 6300 -615
rect 6250 -665 6300 -635
rect 6250 -685 6265 -665
rect 6285 -685 6300 -665
rect 6250 -715 6300 -685
rect 6250 -735 6265 -715
rect 6285 -735 6300 -715
rect 6250 -765 6300 -735
rect 6250 -785 6265 -765
rect 6285 -785 6300 -765
rect 6250 -800 6300 -785
rect 6550 -115 6600 -100
rect 6550 -135 6565 -115
rect 6585 -135 6600 -115
rect 6550 -165 6600 -135
rect 6550 -185 6565 -165
rect 6585 -185 6600 -165
rect 6550 -215 6600 -185
rect 6550 -235 6565 -215
rect 6585 -235 6600 -215
rect 6550 -265 6600 -235
rect 6550 -285 6565 -265
rect 6585 -285 6600 -265
rect 6550 -315 6600 -285
rect 6550 -335 6565 -315
rect 6585 -335 6600 -315
rect 6550 -365 6600 -335
rect 6550 -385 6565 -365
rect 6585 -385 6600 -365
rect 6550 -415 6600 -385
rect 6550 -435 6565 -415
rect 6585 -435 6600 -415
rect 6550 -465 6600 -435
rect 6550 -485 6565 -465
rect 6585 -485 6600 -465
rect 6550 -515 6600 -485
rect 6550 -535 6565 -515
rect 6585 -535 6600 -515
rect 6550 -565 6600 -535
rect 6550 -585 6565 -565
rect 6585 -585 6600 -565
rect 6550 -615 6600 -585
rect 6550 -635 6565 -615
rect 6585 -635 6600 -615
rect 6550 -665 6600 -635
rect 6550 -685 6565 -665
rect 6585 -685 6600 -665
rect 6550 -715 6600 -685
rect 6550 -735 6565 -715
rect 6585 -735 6600 -715
rect 6550 -765 6600 -735
rect 6550 -785 6565 -765
rect 6585 -785 6600 -765
rect 6550 -800 6600 -785
rect 6850 -115 6900 -100
rect 6850 -135 6865 -115
rect 6885 -135 6900 -115
rect 6850 -165 6900 -135
rect 6850 -185 6865 -165
rect 6885 -185 6900 -165
rect 6850 -215 6900 -185
rect 6850 -235 6865 -215
rect 6885 -235 6900 -215
rect 6850 -265 6900 -235
rect 6850 -285 6865 -265
rect 6885 -285 6900 -265
rect 6850 -315 6900 -285
rect 6850 -335 6865 -315
rect 6885 -335 6900 -315
rect 6850 -365 6900 -335
rect 6850 -385 6865 -365
rect 6885 -385 6900 -365
rect 6850 -415 6900 -385
rect 6850 -435 6865 -415
rect 6885 -435 6900 -415
rect 6850 -465 6900 -435
rect 6850 -485 6865 -465
rect 6885 -485 6900 -465
rect 6850 -515 6900 -485
rect 6850 -535 6865 -515
rect 6885 -535 6900 -515
rect 6850 -565 6900 -535
rect 6850 -585 6865 -565
rect 6885 -585 6900 -565
rect 6850 -615 6900 -585
rect 6850 -635 6865 -615
rect 6885 -635 6900 -615
rect 6850 -665 6900 -635
rect 6850 -685 6865 -665
rect 6885 -685 6900 -665
rect 6850 -715 6900 -685
rect 6850 -735 6865 -715
rect 6885 -735 6900 -715
rect 6850 -765 6900 -735
rect 6850 -785 6865 -765
rect 6885 -785 6900 -765
rect 6850 -800 6900 -785
rect 7150 -115 7200 -100
rect 7150 -135 7165 -115
rect 7185 -135 7200 -115
rect 7150 -165 7200 -135
rect 7150 -185 7165 -165
rect 7185 -185 7200 -165
rect 7150 -215 7200 -185
rect 7150 -235 7165 -215
rect 7185 -235 7200 -215
rect 7150 -265 7200 -235
rect 7150 -285 7165 -265
rect 7185 -285 7200 -265
rect 7150 -315 7200 -285
rect 7150 -335 7165 -315
rect 7185 -335 7200 -315
rect 7150 -365 7200 -335
rect 7150 -385 7165 -365
rect 7185 -385 7200 -365
rect 7150 -415 7200 -385
rect 7150 -435 7165 -415
rect 7185 -435 7200 -415
rect 7150 -465 7200 -435
rect 7150 -485 7165 -465
rect 7185 -485 7200 -465
rect 7150 -515 7200 -485
rect 7150 -535 7165 -515
rect 7185 -535 7200 -515
rect 7150 -565 7200 -535
rect 7150 -585 7165 -565
rect 7185 -585 7200 -565
rect 7150 -615 7200 -585
rect 7150 -635 7165 -615
rect 7185 -635 7200 -615
rect 7150 -665 7200 -635
rect 7150 -685 7165 -665
rect 7185 -685 7200 -665
rect 7150 -715 7200 -685
rect 7150 -735 7165 -715
rect 7185 -735 7200 -715
rect 7150 -765 7200 -735
rect 7150 -785 7165 -765
rect 7185 -785 7200 -765
rect 7150 -800 7200 -785
rect 8350 -115 8400 -100
rect 8350 -135 8365 -115
rect 8385 -135 8400 -115
rect 8350 -165 8400 -135
rect 8350 -185 8365 -165
rect 8385 -185 8400 -165
rect 8350 -215 8400 -185
rect 8350 -235 8365 -215
rect 8385 -235 8400 -215
rect 8350 -265 8400 -235
rect 8350 -285 8365 -265
rect 8385 -285 8400 -265
rect 8350 -315 8400 -285
rect 8350 -335 8365 -315
rect 8385 -335 8400 -315
rect 8350 -365 8400 -335
rect 8350 -385 8365 -365
rect 8385 -385 8400 -365
rect 8350 -415 8400 -385
rect 8350 -435 8365 -415
rect 8385 -435 8400 -415
rect 8350 -465 8400 -435
rect 8350 -485 8365 -465
rect 8385 -485 8400 -465
rect 8350 -515 8400 -485
rect 8350 -535 8365 -515
rect 8385 -535 8400 -515
rect 8350 -565 8400 -535
rect 8350 -585 8365 -565
rect 8385 -585 8400 -565
rect 8350 -615 8400 -585
rect 8350 -635 8365 -615
rect 8385 -635 8400 -615
rect 8350 -665 8400 -635
rect 8350 -685 8365 -665
rect 8385 -685 8400 -665
rect 8350 -715 8400 -685
rect 8350 -735 8365 -715
rect 8385 -735 8400 -715
rect 8350 -765 8400 -735
rect 8350 -785 8365 -765
rect 8385 -785 8400 -765
rect 8350 -800 8400 -785
rect 9550 -115 9600 -100
rect 9550 -135 9565 -115
rect 9585 -135 9600 -115
rect 9550 -165 9600 -135
rect 9550 -185 9565 -165
rect 9585 -185 9600 -165
rect 9550 -215 9600 -185
rect 9550 -235 9565 -215
rect 9585 -235 9600 -215
rect 9550 -265 9600 -235
rect 9550 -285 9565 -265
rect 9585 -285 9600 -265
rect 9550 -315 9600 -285
rect 9550 -335 9565 -315
rect 9585 -335 9600 -315
rect 9550 -365 9600 -335
rect 9550 -385 9565 -365
rect 9585 -385 9600 -365
rect 9550 -415 9600 -385
rect 9550 -435 9565 -415
rect 9585 -435 9600 -415
rect 9550 -465 9600 -435
rect 9550 -485 9565 -465
rect 9585 -485 9600 -465
rect 9550 -515 9600 -485
rect 9550 -535 9565 -515
rect 9585 -535 9600 -515
rect 9550 -565 9600 -535
rect 9550 -585 9565 -565
rect 9585 -585 9600 -565
rect 9550 -615 9600 -585
rect 9550 -635 9565 -615
rect 9585 -635 9600 -615
rect 9550 -665 9600 -635
rect 9550 -685 9565 -665
rect 9585 -685 9600 -665
rect 9550 -715 9600 -685
rect 9550 -735 9565 -715
rect 9585 -735 9600 -715
rect 9550 -765 9600 -735
rect 9550 -785 9565 -765
rect 9585 -785 9600 -765
rect 9550 -800 9600 -785
rect 10750 -115 10800 -100
rect 10750 -135 10765 -115
rect 10785 -135 10800 -115
rect 10750 -165 10800 -135
rect 10750 -185 10765 -165
rect 10785 -185 10800 -165
rect 10750 -215 10800 -185
rect 10750 -235 10765 -215
rect 10785 -235 10800 -215
rect 10750 -265 10800 -235
rect 10750 -285 10765 -265
rect 10785 -285 10800 -265
rect 10750 -315 10800 -285
rect 10750 -335 10765 -315
rect 10785 -335 10800 -315
rect 10750 -365 10800 -335
rect 10750 -385 10765 -365
rect 10785 -385 10800 -365
rect 10750 -415 10800 -385
rect 10750 -435 10765 -415
rect 10785 -435 10800 -415
rect 10750 -465 10800 -435
rect 10750 -485 10765 -465
rect 10785 -485 10800 -465
rect 10750 -515 10800 -485
rect 10750 -535 10765 -515
rect 10785 -535 10800 -515
rect 10750 -565 10800 -535
rect 10750 -585 10765 -565
rect 10785 -585 10800 -565
rect 10750 -615 10800 -585
rect 10750 -635 10765 -615
rect 10785 -635 10800 -615
rect 10750 -665 10800 -635
rect 10750 -685 10765 -665
rect 10785 -685 10800 -665
rect 10750 -715 10800 -685
rect 10750 -735 10765 -715
rect 10785 -735 10800 -715
rect 10750 -765 10800 -735
rect 10750 -785 10765 -765
rect 10785 -785 10800 -765
rect 10750 -800 10800 -785
rect 11950 -115 12000 -100
rect 11950 -135 11965 -115
rect 11985 -135 12000 -115
rect 11950 -165 12000 -135
rect 11950 -185 11965 -165
rect 11985 -185 12000 -165
rect 11950 -215 12000 -185
rect 11950 -235 11965 -215
rect 11985 -235 12000 -215
rect 11950 -265 12000 -235
rect 11950 -285 11965 -265
rect 11985 -285 12000 -265
rect 11950 -315 12000 -285
rect 11950 -335 11965 -315
rect 11985 -335 12000 -315
rect 11950 -365 12000 -335
rect 11950 -385 11965 -365
rect 11985 -385 12000 -365
rect 11950 -415 12000 -385
rect 11950 -435 11965 -415
rect 11985 -435 12000 -415
rect 11950 -465 12000 -435
rect 11950 -485 11965 -465
rect 11985 -485 12000 -465
rect 11950 -515 12000 -485
rect 11950 -535 11965 -515
rect 11985 -535 12000 -515
rect 11950 -565 12000 -535
rect 11950 -585 11965 -565
rect 11985 -585 12000 -565
rect 11950 -615 12000 -585
rect 11950 -635 11965 -615
rect 11985 -635 12000 -615
rect 11950 -665 12000 -635
rect 11950 -685 11965 -665
rect 11985 -685 12000 -665
rect 11950 -715 12000 -685
rect 11950 -735 11965 -715
rect 11985 -735 12000 -715
rect 11950 -765 12000 -735
rect 11950 -785 11965 -765
rect 11985 -785 12000 -765
rect 11950 -800 12000 -785
rect 12250 -115 12300 -100
rect 12250 -135 12265 -115
rect 12285 -135 12300 -115
rect 12250 -165 12300 -135
rect 12250 -185 12265 -165
rect 12285 -185 12300 -165
rect 12250 -215 12300 -185
rect 12250 -235 12265 -215
rect 12285 -235 12300 -215
rect 12250 -265 12300 -235
rect 12250 -285 12265 -265
rect 12285 -285 12300 -265
rect 12250 -315 12300 -285
rect 12250 -335 12265 -315
rect 12285 -335 12300 -315
rect 12250 -365 12300 -335
rect 12250 -385 12265 -365
rect 12285 -385 12300 -365
rect 12250 -415 12300 -385
rect 12250 -435 12265 -415
rect 12285 -435 12300 -415
rect 12250 -465 12300 -435
rect 12250 -485 12265 -465
rect 12285 -485 12300 -465
rect 12250 -515 12300 -485
rect 12250 -535 12265 -515
rect 12285 -535 12300 -515
rect 12250 -565 12300 -535
rect 12250 -585 12265 -565
rect 12285 -585 12300 -565
rect 12250 -615 12300 -585
rect 12250 -635 12265 -615
rect 12285 -635 12300 -615
rect 12250 -665 12300 -635
rect 12250 -685 12265 -665
rect 12285 -685 12300 -665
rect 12250 -715 12300 -685
rect 12250 -735 12265 -715
rect 12285 -735 12300 -715
rect 12250 -765 12300 -735
rect 12250 -785 12265 -765
rect 12285 -785 12300 -765
rect 12250 -800 12300 -785
rect 12550 -115 12600 -100
rect 12550 -135 12565 -115
rect 12585 -135 12600 -115
rect 12550 -165 12600 -135
rect 12550 -185 12565 -165
rect 12585 -185 12600 -165
rect 12550 -215 12600 -185
rect 12550 -235 12565 -215
rect 12585 -235 12600 -215
rect 12550 -265 12600 -235
rect 12550 -285 12565 -265
rect 12585 -285 12600 -265
rect 12550 -315 12600 -285
rect 12550 -335 12565 -315
rect 12585 -335 12600 -315
rect 12550 -365 12600 -335
rect 12550 -385 12565 -365
rect 12585 -385 12600 -365
rect 12550 -415 12600 -385
rect 12550 -435 12565 -415
rect 12585 -435 12600 -415
rect 12550 -465 12600 -435
rect 12550 -485 12565 -465
rect 12585 -485 12600 -465
rect 12550 -515 12600 -485
rect 12550 -535 12565 -515
rect 12585 -535 12600 -515
rect 12550 -565 12600 -535
rect 12550 -585 12565 -565
rect 12585 -585 12600 -565
rect 12550 -615 12600 -585
rect 12550 -635 12565 -615
rect 12585 -635 12600 -615
rect 12550 -665 12600 -635
rect 12550 -685 12565 -665
rect 12585 -685 12600 -665
rect 12550 -715 12600 -685
rect 12550 -735 12565 -715
rect 12585 -735 12600 -715
rect 12550 -765 12600 -735
rect 12550 -785 12565 -765
rect 12585 -785 12600 -765
rect 12550 -800 12600 -785
rect 12850 -115 12900 -100
rect 12850 -135 12865 -115
rect 12885 -135 12900 -115
rect 12850 -165 12900 -135
rect 12850 -185 12865 -165
rect 12885 -185 12900 -165
rect 12850 -215 12900 -185
rect 12850 -235 12865 -215
rect 12885 -235 12900 -215
rect 12850 -265 12900 -235
rect 12850 -285 12865 -265
rect 12885 -285 12900 -265
rect 12850 -315 12900 -285
rect 12850 -335 12865 -315
rect 12885 -335 12900 -315
rect 12850 -365 12900 -335
rect 12850 -385 12865 -365
rect 12885 -385 12900 -365
rect 12850 -415 12900 -385
rect 12850 -435 12865 -415
rect 12885 -435 12900 -415
rect 12850 -465 12900 -435
rect 12850 -485 12865 -465
rect 12885 -485 12900 -465
rect 12850 -515 12900 -485
rect 12850 -535 12865 -515
rect 12885 -535 12900 -515
rect 12850 -565 12900 -535
rect 12850 -585 12865 -565
rect 12885 -585 12900 -565
rect 12850 -615 12900 -585
rect 12850 -635 12865 -615
rect 12885 -635 12900 -615
rect 12850 -665 12900 -635
rect 12850 -685 12865 -665
rect 12885 -685 12900 -665
rect 12850 -715 12900 -685
rect 12850 -735 12865 -715
rect 12885 -735 12900 -715
rect 12850 -765 12900 -735
rect 12850 -785 12865 -765
rect 12885 -785 12900 -765
rect 12850 -800 12900 -785
rect 13150 -115 13200 -100
rect 13150 -135 13165 -115
rect 13185 -135 13200 -115
rect 13150 -165 13200 -135
rect 13150 -185 13165 -165
rect 13185 -185 13200 -165
rect 13150 -215 13200 -185
rect 13150 -235 13165 -215
rect 13185 -235 13200 -215
rect 13150 -265 13200 -235
rect 13150 -285 13165 -265
rect 13185 -285 13200 -265
rect 13150 -315 13200 -285
rect 13150 -335 13165 -315
rect 13185 -335 13200 -315
rect 13150 -365 13200 -335
rect 13150 -385 13165 -365
rect 13185 -385 13200 -365
rect 13150 -415 13200 -385
rect 13150 -435 13165 -415
rect 13185 -435 13200 -415
rect 13150 -465 13200 -435
rect 13150 -485 13165 -465
rect 13185 -485 13200 -465
rect 13150 -515 13200 -485
rect 13150 -535 13165 -515
rect 13185 -535 13200 -515
rect 13150 -565 13200 -535
rect 13150 -585 13165 -565
rect 13185 -585 13200 -565
rect 13150 -615 13200 -585
rect 13150 -635 13165 -615
rect 13185 -635 13200 -615
rect 13150 -665 13200 -635
rect 13150 -685 13165 -665
rect 13185 -685 13200 -665
rect 13150 -715 13200 -685
rect 13150 -735 13165 -715
rect 13185 -735 13200 -715
rect 13150 -765 13200 -735
rect 13150 -785 13165 -765
rect 13185 -785 13200 -765
rect 13150 -800 13200 -785
rect 13450 -115 13500 -100
rect 13450 -135 13465 -115
rect 13485 -135 13500 -115
rect 13450 -165 13500 -135
rect 13450 -185 13465 -165
rect 13485 -185 13500 -165
rect 13450 -215 13500 -185
rect 13450 -235 13465 -215
rect 13485 -235 13500 -215
rect 13450 -265 13500 -235
rect 13450 -285 13465 -265
rect 13485 -285 13500 -265
rect 13450 -315 13500 -285
rect 13450 -335 13465 -315
rect 13485 -335 13500 -315
rect 13450 -365 13500 -335
rect 13450 -385 13465 -365
rect 13485 -385 13500 -365
rect 13450 -415 13500 -385
rect 13450 -435 13465 -415
rect 13485 -435 13500 -415
rect 13450 -465 13500 -435
rect 13450 -485 13465 -465
rect 13485 -485 13500 -465
rect 13450 -515 13500 -485
rect 13450 -535 13465 -515
rect 13485 -535 13500 -515
rect 13450 -565 13500 -535
rect 13450 -585 13465 -565
rect 13485 -585 13500 -565
rect 13450 -615 13500 -585
rect 13450 -635 13465 -615
rect 13485 -635 13500 -615
rect 13450 -665 13500 -635
rect 13450 -685 13465 -665
rect 13485 -685 13500 -665
rect 13450 -715 13500 -685
rect 13450 -735 13465 -715
rect 13485 -735 13500 -715
rect 13450 -765 13500 -735
rect 13450 -785 13465 -765
rect 13485 -785 13500 -765
rect 13450 -800 13500 -785
rect 13750 -115 13800 -100
rect 13750 -135 13765 -115
rect 13785 -135 13800 -115
rect 13750 -165 13800 -135
rect 13750 -185 13765 -165
rect 13785 -185 13800 -165
rect 13750 -215 13800 -185
rect 13750 -235 13765 -215
rect 13785 -235 13800 -215
rect 13750 -265 13800 -235
rect 13750 -285 13765 -265
rect 13785 -285 13800 -265
rect 13750 -315 13800 -285
rect 13750 -335 13765 -315
rect 13785 -335 13800 -315
rect 13750 -365 13800 -335
rect 13750 -385 13765 -365
rect 13785 -385 13800 -365
rect 13750 -415 13800 -385
rect 13750 -435 13765 -415
rect 13785 -435 13800 -415
rect 13750 -465 13800 -435
rect 13750 -485 13765 -465
rect 13785 -485 13800 -465
rect 13750 -515 13800 -485
rect 13750 -535 13765 -515
rect 13785 -535 13800 -515
rect 13750 -565 13800 -535
rect 13750 -585 13765 -565
rect 13785 -585 13800 -565
rect 13750 -615 13800 -585
rect 13750 -635 13765 -615
rect 13785 -635 13800 -615
rect 13750 -665 13800 -635
rect 13750 -685 13765 -665
rect 13785 -685 13800 -665
rect 13750 -715 13800 -685
rect 13750 -735 13765 -715
rect 13785 -735 13800 -715
rect 13750 -765 13800 -735
rect 13750 -785 13765 -765
rect 13785 -785 13800 -765
rect 13750 -800 13800 -785
rect 14050 -115 14100 -100
rect 14050 -135 14065 -115
rect 14085 -135 14100 -115
rect 14050 -165 14100 -135
rect 14050 -185 14065 -165
rect 14085 -185 14100 -165
rect 14050 -215 14100 -185
rect 14050 -235 14065 -215
rect 14085 -235 14100 -215
rect 14050 -265 14100 -235
rect 14050 -285 14065 -265
rect 14085 -285 14100 -265
rect 14050 -315 14100 -285
rect 14050 -335 14065 -315
rect 14085 -335 14100 -315
rect 14050 -365 14100 -335
rect 14050 -385 14065 -365
rect 14085 -385 14100 -365
rect 14050 -415 14100 -385
rect 14050 -435 14065 -415
rect 14085 -435 14100 -415
rect 14050 -465 14100 -435
rect 14050 -485 14065 -465
rect 14085 -485 14100 -465
rect 14050 -515 14100 -485
rect 14050 -535 14065 -515
rect 14085 -535 14100 -515
rect 14050 -565 14100 -535
rect 14050 -585 14065 -565
rect 14085 -585 14100 -565
rect 14050 -615 14100 -585
rect 14050 -635 14065 -615
rect 14085 -635 14100 -615
rect 14050 -665 14100 -635
rect 14050 -685 14065 -665
rect 14085 -685 14100 -665
rect 14050 -715 14100 -685
rect 14050 -735 14065 -715
rect 14085 -735 14100 -715
rect 14050 -765 14100 -735
rect 14050 -785 14065 -765
rect 14085 -785 14100 -765
rect 14050 -800 14100 -785
rect 14350 -115 14400 -100
rect 14350 -135 14365 -115
rect 14385 -135 14400 -115
rect 14350 -165 14400 -135
rect 14350 -185 14365 -165
rect 14385 -185 14400 -165
rect 14350 -215 14400 -185
rect 14350 -235 14365 -215
rect 14385 -235 14400 -215
rect 14350 -265 14400 -235
rect 14350 -285 14365 -265
rect 14385 -285 14400 -265
rect 14350 -315 14400 -285
rect 14350 -335 14365 -315
rect 14385 -335 14400 -315
rect 14350 -365 14400 -335
rect 14350 -385 14365 -365
rect 14385 -385 14400 -365
rect 14350 -415 14400 -385
rect 14350 -435 14365 -415
rect 14385 -435 14400 -415
rect 14350 -465 14400 -435
rect 14350 -485 14365 -465
rect 14385 -485 14400 -465
rect 14350 -515 14400 -485
rect 14350 -535 14365 -515
rect 14385 -535 14400 -515
rect 14350 -565 14400 -535
rect 14350 -585 14365 -565
rect 14385 -585 14400 -565
rect 14350 -615 14400 -585
rect 14350 -635 14365 -615
rect 14385 -635 14400 -615
rect 14350 -665 14400 -635
rect 14350 -685 14365 -665
rect 14385 -685 14400 -665
rect 14350 -715 14400 -685
rect 14350 -735 14365 -715
rect 14385 -735 14400 -715
rect 14350 -765 14400 -735
rect 14350 -785 14365 -765
rect 14385 -785 14400 -765
rect 14350 -800 14400 -785
rect 15550 -115 15600 -100
rect 15550 -135 15565 -115
rect 15585 -135 15600 -115
rect 15550 -165 15600 -135
rect 15550 -185 15565 -165
rect 15585 -185 15600 -165
rect 15550 -215 15600 -185
rect 15550 -235 15565 -215
rect 15585 -235 15600 -215
rect 15550 -265 15600 -235
rect 15550 -285 15565 -265
rect 15585 -285 15600 -265
rect 15550 -315 15600 -285
rect 15550 -335 15565 -315
rect 15585 -335 15600 -315
rect 15550 -365 15600 -335
rect 15550 -385 15565 -365
rect 15585 -385 15600 -365
rect 15550 -415 15600 -385
rect 15550 -435 15565 -415
rect 15585 -435 15600 -415
rect 15550 -465 15600 -435
rect 15550 -485 15565 -465
rect 15585 -485 15600 -465
rect 15550 -515 15600 -485
rect 15550 -535 15565 -515
rect 15585 -535 15600 -515
rect 15550 -565 15600 -535
rect 15550 -585 15565 -565
rect 15585 -585 15600 -565
rect 15550 -615 15600 -585
rect 15550 -635 15565 -615
rect 15585 -635 15600 -615
rect 15550 -665 15600 -635
rect 15550 -685 15565 -665
rect 15585 -685 15600 -665
rect 15550 -715 15600 -685
rect 15550 -735 15565 -715
rect 15585 -735 15600 -715
rect 15550 -765 15600 -735
rect 15550 -785 15565 -765
rect 15585 -785 15600 -765
rect 15550 -800 15600 -785
rect 16750 -115 16800 -100
rect 16750 -135 16765 -115
rect 16785 -135 16800 -115
rect 16750 -165 16800 -135
rect 16750 -185 16765 -165
rect 16785 -185 16800 -165
rect 16750 -215 16800 -185
rect 16750 -235 16765 -215
rect 16785 -235 16800 -215
rect 16750 -265 16800 -235
rect 16750 -285 16765 -265
rect 16785 -285 16800 -265
rect 16750 -315 16800 -285
rect 16750 -335 16765 -315
rect 16785 -335 16800 -315
rect 16750 -365 16800 -335
rect 16750 -385 16765 -365
rect 16785 -385 16800 -365
rect 16750 -415 16800 -385
rect 16750 -435 16765 -415
rect 16785 -435 16800 -415
rect 16750 -465 16800 -435
rect 16750 -485 16765 -465
rect 16785 -485 16800 -465
rect 16750 -515 16800 -485
rect 16750 -535 16765 -515
rect 16785 -535 16800 -515
rect 16750 -565 16800 -535
rect 16750 -585 16765 -565
rect 16785 -585 16800 -565
rect 16750 -615 16800 -585
rect 16750 -635 16765 -615
rect 16785 -635 16800 -615
rect 16750 -665 16800 -635
rect 16750 -685 16765 -665
rect 16785 -685 16800 -665
rect 16750 -715 16800 -685
rect 16750 -735 16765 -715
rect 16785 -735 16800 -715
rect 16750 -765 16800 -735
rect 16750 -785 16765 -765
rect 16785 -785 16800 -765
rect 16750 -800 16800 -785
rect 17950 -115 18000 -100
rect 17950 -135 17965 -115
rect 17985 -135 18000 -115
rect 17950 -165 18000 -135
rect 17950 -185 17965 -165
rect 17985 -185 18000 -165
rect 17950 -215 18000 -185
rect 17950 -235 17965 -215
rect 17985 -235 18000 -215
rect 17950 -265 18000 -235
rect 17950 -285 17965 -265
rect 17985 -285 18000 -265
rect 17950 -315 18000 -285
rect 17950 -335 17965 -315
rect 17985 -335 18000 -315
rect 17950 -365 18000 -335
rect 17950 -385 17965 -365
rect 17985 -385 18000 -365
rect 17950 -415 18000 -385
rect 17950 -435 17965 -415
rect 17985 -435 18000 -415
rect 17950 -465 18000 -435
rect 17950 -485 17965 -465
rect 17985 -485 18000 -465
rect 17950 -515 18000 -485
rect 17950 -535 17965 -515
rect 17985 -535 18000 -515
rect 17950 -565 18000 -535
rect 17950 -585 17965 -565
rect 17985 -585 18000 -565
rect 17950 -615 18000 -585
rect 17950 -635 17965 -615
rect 17985 -635 18000 -615
rect 17950 -665 18000 -635
rect 17950 -685 17965 -665
rect 17985 -685 18000 -665
rect 17950 -715 18000 -685
rect 17950 -735 17965 -715
rect 17985 -735 18000 -715
rect 17950 -765 18000 -735
rect 17950 -785 17965 -765
rect 17985 -785 18000 -765
rect 17950 -800 18000 -785
rect 19150 -115 19200 -100
rect 19150 -135 19165 -115
rect 19185 -135 19200 -115
rect 19150 -165 19200 -135
rect 19150 -185 19165 -165
rect 19185 -185 19200 -165
rect 19150 -215 19200 -185
rect 19150 -235 19165 -215
rect 19185 -235 19200 -215
rect 19150 -265 19200 -235
rect 19150 -285 19165 -265
rect 19185 -285 19200 -265
rect 19150 -315 19200 -285
rect 19150 -335 19165 -315
rect 19185 -335 19200 -315
rect 19150 -365 19200 -335
rect 19150 -385 19165 -365
rect 19185 -385 19200 -365
rect 19150 -415 19200 -385
rect 19150 -435 19165 -415
rect 19185 -435 19200 -415
rect 19150 -465 19200 -435
rect 19150 -485 19165 -465
rect 19185 -485 19200 -465
rect 19150 -515 19200 -485
rect 19150 -535 19165 -515
rect 19185 -535 19200 -515
rect 19150 -565 19200 -535
rect 19150 -585 19165 -565
rect 19185 -585 19200 -565
rect 19150 -615 19200 -585
rect 19150 -635 19165 -615
rect 19185 -635 19200 -615
rect 19150 -665 19200 -635
rect 19150 -685 19165 -665
rect 19185 -685 19200 -665
rect 19150 -715 19200 -685
rect 19150 -735 19165 -715
rect 19185 -735 19200 -715
rect 19150 -765 19200 -735
rect 19150 -785 19165 -765
rect 19185 -785 19200 -765
rect 19150 -800 19200 -785
rect 20350 -115 20400 -100
rect 20350 -135 20365 -115
rect 20385 -135 20400 -115
rect 20350 -165 20400 -135
rect 20350 -185 20365 -165
rect 20385 -185 20400 -165
rect 20350 -215 20400 -185
rect 20350 -235 20365 -215
rect 20385 -235 20400 -215
rect 20350 -265 20400 -235
rect 20350 -285 20365 -265
rect 20385 -285 20400 -265
rect 20350 -315 20400 -285
rect 20350 -335 20365 -315
rect 20385 -335 20400 -315
rect 20350 -365 20400 -335
rect 20350 -385 20365 -365
rect 20385 -385 20400 -365
rect 20350 -415 20400 -385
rect 20350 -435 20365 -415
rect 20385 -435 20400 -415
rect 20350 -465 20400 -435
rect 20350 -485 20365 -465
rect 20385 -485 20400 -465
rect 20350 -515 20400 -485
rect 20350 -535 20365 -515
rect 20385 -535 20400 -515
rect 20350 -565 20400 -535
rect 20350 -585 20365 -565
rect 20385 -585 20400 -565
rect 20350 -615 20400 -585
rect 20350 -635 20365 -615
rect 20385 -635 20400 -615
rect 20350 -665 20400 -635
rect 20350 -685 20365 -665
rect 20385 -685 20400 -665
rect 20350 -715 20400 -685
rect 20350 -735 20365 -715
rect 20385 -735 20400 -715
rect 20350 -765 20400 -735
rect 20350 -785 20365 -765
rect 20385 -785 20400 -765
rect 20350 -800 20400 -785
rect 21550 -115 21600 -100
rect 21550 -135 21565 -115
rect 21585 -135 21600 -115
rect 21550 -165 21600 -135
rect 21550 -185 21565 -165
rect 21585 -185 21600 -165
rect 21550 -215 21600 -185
rect 21550 -235 21565 -215
rect 21585 -235 21600 -215
rect 21550 -265 21600 -235
rect 21550 -285 21565 -265
rect 21585 -285 21600 -265
rect 21550 -315 21600 -285
rect 21550 -335 21565 -315
rect 21585 -335 21600 -315
rect 21550 -365 21600 -335
rect 21550 -385 21565 -365
rect 21585 -385 21600 -365
rect 21550 -415 21600 -385
rect 21550 -435 21565 -415
rect 21585 -435 21600 -415
rect 21550 -465 21600 -435
rect 21550 -485 21565 -465
rect 21585 -485 21600 -465
rect 21550 -515 21600 -485
rect 21550 -535 21565 -515
rect 21585 -535 21600 -515
rect 21550 -565 21600 -535
rect 21550 -585 21565 -565
rect 21585 -585 21600 -565
rect 21550 -615 21600 -585
rect 21550 -635 21565 -615
rect 21585 -635 21600 -615
rect 21550 -665 21600 -635
rect 21550 -685 21565 -665
rect 21585 -685 21600 -665
rect 21550 -715 21600 -685
rect 21550 -735 21565 -715
rect 21585 -735 21600 -715
rect 21550 -765 21600 -735
rect 21550 -785 21565 -765
rect 21585 -785 21600 -765
rect 21550 -800 21600 -785
rect 22450 -115 22500 -100
rect 22450 -135 22465 -115
rect 22485 -135 22500 -115
rect 22450 -165 22500 -135
rect 22450 -185 22465 -165
rect 22485 -185 22500 -165
rect 22450 -215 22500 -185
rect 22450 -235 22465 -215
rect 22485 -235 22500 -215
rect 22450 -265 22500 -235
rect 22450 -285 22465 -265
rect 22485 -285 22500 -265
rect 22450 -315 22500 -285
rect 22450 -335 22465 -315
rect 22485 -335 22500 -315
rect 22450 -365 22500 -335
rect 22450 -385 22465 -365
rect 22485 -385 22500 -365
rect 22450 -415 22500 -385
rect 22450 -435 22465 -415
rect 22485 -435 22500 -415
rect 22450 -465 22500 -435
rect 22450 -485 22465 -465
rect 22485 -485 22500 -465
rect 22450 -515 22500 -485
rect 22450 -535 22465 -515
rect 22485 -535 22500 -515
rect 22450 -565 22500 -535
rect 22450 -585 22465 -565
rect 22485 -585 22500 -565
rect 22450 -615 22500 -585
rect 22450 -635 22465 -615
rect 22485 -635 22500 -615
rect 22450 -665 22500 -635
rect 22450 -685 22465 -665
rect 22485 -685 22500 -665
rect 22450 -715 22500 -685
rect 22450 -735 22465 -715
rect 22485 -735 22500 -715
rect 22450 -765 22500 -735
rect 22450 -785 22465 -765
rect 22485 -785 22500 -765
rect 22450 -800 22500 -785
rect 23350 -115 23400 -100
rect 23350 -135 23365 -115
rect 23385 -135 23400 -115
rect 23350 -165 23400 -135
rect 23350 -185 23365 -165
rect 23385 -185 23400 -165
rect 23350 -215 23400 -185
rect 23350 -235 23365 -215
rect 23385 -235 23400 -215
rect 23350 -265 23400 -235
rect 23350 -285 23365 -265
rect 23385 -285 23400 -265
rect 23350 -315 23400 -285
rect 23350 -335 23365 -315
rect 23385 -335 23400 -315
rect 23350 -365 23400 -335
rect 23350 -385 23365 -365
rect 23385 -385 23400 -365
rect 23350 -415 23400 -385
rect 23350 -435 23365 -415
rect 23385 -435 23400 -415
rect 23350 -465 23400 -435
rect 23350 -485 23365 -465
rect 23385 -485 23400 -465
rect 23350 -515 23400 -485
rect 23350 -535 23365 -515
rect 23385 -535 23400 -515
rect 23350 -565 23400 -535
rect 23350 -585 23365 -565
rect 23385 -585 23400 -565
rect 23350 -615 23400 -585
rect 23350 -635 23365 -615
rect 23385 -635 23400 -615
rect 23350 -665 23400 -635
rect 23350 -685 23365 -665
rect 23385 -685 23400 -665
rect 23350 -715 23400 -685
rect 23350 -735 23365 -715
rect 23385 -735 23400 -715
rect 23350 -765 23400 -735
rect 23350 -785 23365 -765
rect 23385 -785 23400 -765
rect 23350 -800 23400 -785
rect 24550 -115 24600 -100
rect 24550 -135 24565 -115
rect 24585 -135 24600 -115
rect 24550 -165 24600 -135
rect 24550 -185 24565 -165
rect 24585 -185 24600 -165
rect 24550 -215 24600 -185
rect 24550 -235 24565 -215
rect 24585 -235 24600 -215
rect 24550 -265 24600 -235
rect 24550 -285 24565 -265
rect 24585 -285 24600 -265
rect 24550 -315 24600 -285
rect 24550 -335 24565 -315
rect 24585 -335 24600 -315
rect 24550 -365 24600 -335
rect 24550 -385 24565 -365
rect 24585 -385 24600 -365
rect 24550 -415 24600 -385
rect 24550 -435 24565 -415
rect 24585 -435 24600 -415
rect 24550 -465 24600 -435
rect 24550 -485 24565 -465
rect 24585 -485 24600 -465
rect 24550 -515 24600 -485
rect 24550 -535 24565 -515
rect 24585 -535 24600 -515
rect 24550 -565 24600 -535
rect 24550 -585 24565 -565
rect 24585 -585 24600 -565
rect 24550 -615 24600 -585
rect 24550 -635 24565 -615
rect 24585 -635 24600 -615
rect 24550 -665 24600 -635
rect 24550 -685 24565 -665
rect 24585 -685 24600 -665
rect 24550 -715 24600 -685
rect 24550 -735 24565 -715
rect 24585 -735 24600 -715
rect 24550 -765 24600 -735
rect 24550 -785 24565 -765
rect 24585 -785 24600 -765
rect 24550 -800 24600 -785
rect 25750 -115 25800 -100
rect 25750 -135 25765 -115
rect 25785 -135 25800 -115
rect 25750 -165 25800 -135
rect 25750 -185 25765 -165
rect 25785 -185 25800 -165
rect 25750 -215 25800 -185
rect 25750 -235 25765 -215
rect 25785 -235 25800 -215
rect 25750 -265 25800 -235
rect 25750 -285 25765 -265
rect 25785 -285 25800 -265
rect 25750 -315 25800 -285
rect 25750 -335 25765 -315
rect 25785 -335 25800 -315
rect 25750 -365 25800 -335
rect 25750 -385 25765 -365
rect 25785 -385 25800 -365
rect 25750 -415 25800 -385
rect 25750 -435 25765 -415
rect 25785 -435 25800 -415
rect 25750 -465 25800 -435
rect 25750 -485 25765 -465
rect 25785 -485 25800 -465
rect 25750 -515 25800 -485
rect 25750 -535 25765 -515
rect 25785 -535 25800 -515
rect 25750 -565 25800 -535
rect 25750 -585 25765 -565
rect 25785 -585 25800 -565
rect 25750 -615 25800 -585
rect 25750 -635 25765 -615
rect 25785 -635 25800 -615
rect 25750 -665 25800 -635
rect 25750 -685 25765 -665
rect 25785 -685 25800 -665
rect 25750 -715 25800 -685
rect 25750 -735 25765 -715
rect 25785 -735 25800 -715
rect 25750 -765 25800 -735
rect 25750 -785 25765 -765
rect 25785 -785 25800 -765
rect 25750 -800 25800 -785
rect 26650 -115 26700 -100
rect 26650 -135 26665 -115
rect 26685 -135 26700 -115
rect 26650 -165 26700 -135
rect 26650 -185 26665 -165
rect 26685 -185 26700 -165
rect 26650 -215 26700 -185
rect 26650 -235 26665 -215
rect 26685 -235 26700 -215
rect 26650 -265 26700 -235
rect 26650 -285 26665 -265
rect 26685 -285 26700 -265
rect 26650 -315 26700 -285
rect 26650 -335 26665 -315
rect 26685 -335 26700 -315
rect 26650 -365 26700 -335
rect 26650 -385 26665 -365
rect 26685 -385 26700 -365
rect 26650 -415 26700 -385
rect 26650 -435 26665 -415
rect 26685 -435 26700 -415
rect 26650 -465 26700 -435
rect 26650 -485 26665 -465
rect 26685 -485 26700 -465
rect 26650 -515 26700 -485
rect 26650 -535 26665 -515
rect 26685 -535 26700 -515
rect 26650 -565 26700 -535
rect 26650 -585 26665 -565
rect 26685 -585 26700 -565
rect 26650 -615 26700 -585
rect 26650 -635 26665 -615
rect 26685 -635 26700 -615
rect 26650 -665 26700 -635
rect 26650 -685 26665 -665
rect 26685 -685 26700 -665
rect 26650 -715 26700 -685
rect 26650 -735 26665 -715
rect 26685 -735 26700 -715
rect 26650 -765 26700 -735
rect 26650 -785 26665 -765
rect 26685 -785 26700 -765
rect 26650 -800 26700 -785
rect 27550 -115 27600 -100
rect 27550 -135 27565 -115
rect 27585 -135 27600 -115
rect 27550 -165 27600 -135
rect 27550 -185 27565 -165
rect 27585 -185 27600 -165
rect 27550 -215 27600 -185
rect 27550 -235 27565 -215
rect 27585 -235 27600 -215
rect 27550 -265 27600 -235
rect 27550 -285 27565 -265
rect 27585 -285 27600 -265
rect 27550 -315 27600 -285
rect 27550 -335 27565 -315
rect 27585 -335 27600 -315
rect 27550 -365 27600 -335
rect 27550 -385 27565 -365
rect 27585 -385 27600 -365
rect 27550 -415 27600 -385
rect 27550 -435 27565 -415
rect 27585 -435 27600 -415
rect 27550 -465 27600 -435
rect 27550 -485 27565 -465
rect 27585 -485 27600 -465
rect 27550 -515 27600 -485
rect 27550 -535 27565 -515
rect 27585 -535 27600 -515
rect 27550 -565 27600 -535
rect 27550 -585 27565 -565
rect 27585 -585 27600 -565
rect 27550 -615 27600 -585
rect 27550 -635 27565 -615
rect 27585 -635 27600 -615
rect 27550 -665 27600 -635
rect 27550 -685 27565 -665
rect 27585 -685 27600 -665
rect 27550 -715 27600 -685
rect 27550 -735 27565 -715
rect 27585 -735 27600 -715
rect 27550 -765 27600 -735
rect 27550 -785 27565 -765
rect 27585 -785 27600 -765
rect 27550 -800 27600 -785
rect 28750 -115 28800 -100
rect 28750 -135 28765 -115
rect 28785 -135 28800 -115
rect 28750 -165 28800 -135
rect 28750 -185 28765 -165
rect 28785 -185 28800 -165
rect 28750 -215 28800 -185
rect 28750 -235 28765 -215
rect 28785 -235 28800 -215
rect 28750 -265 28800 -235
rect 28750 -285 28765 -265
rect 28785 -285 28800 -265
rect 28750 -315 28800 -285
rect 28750 -335 28765 -315
rect 28785 -335 28800 -315
rect 28750 -365 28800 -335
rect 28750 -385 28765 -365
rect 28785 -385 28800 -365
rect 28750 -415 28800 -385
rect 28750 -435 28765 -415
rect 28785 -435 28800 -415
rect 28750 -465 28800 -435
rect 28750 -485 28765 -465
rect 28785 -485 28800 -465
rect 28750 -515 28800 -485
rect 28750 -535 28765 -515
rect 28785 -535 28800 -515
rect 28750 -565 28800 -535
rect 28750 -585 28765 -565
rect 28785 -585 28800 -565
rect 28750 -615 28800 -585
rect 28750 -635 28765 -615
rect 28785 -635 28800 -615
rect 28750 -665 28800 -635
rect 28750 -685 28765 -665
rect 28785 -685 28800 -665
rect 28750 -715 28800 -685
rect 28750 -735 28765 -715
rect 28785 -735 28800 -715
rect 28750 -765 28800 -735
rect 28750 -785 28765 -765
rect 28785 -785 28800 -765
rect 28750 -800 28800 -785
rect -600 -865 -350 -850
rect -600 -885 -585 -865
rect -565 -885 -535 -865
rect -515 -885 -485 -865
rect -465 -885 -435 -865
rect -415 -885 -385 -865
rect -365 -885 -350 -865
rect -600 -900 -350 -885
rect -300 -865 -50 -850
rect -300 -885 -285 -865
rect -265 -885 -235 -865
rect -215 -885 -185 -865
rect -165 -885 -135 -865
rect -115 -885 -85 -865
rect -65 -885 -50 -865
rect -300 -900 -50 -885
rect 0 -865 250 -850
rect 0 -885 15 -865
rect 35 -885 65 -865
rect 85 -885 115 -865
rect 135 -885 165 -865
rect 185 -885 215 -865
rect 235 -885 250 -865
rect 0 -900 250 -885
rect 300 -865 550 -850
rect 300 -885 315 -865
rect 335 -885 365 -865
rect 385 -885 415 -865
rect 435 -885 465 -865
rect 485 -885 515 -865
rect 535 -885 550 -865
rect 300 -900 550 -885
rect 600 -865 850 -850
rect 600 -885 615 -865
rect 635 -885 665 -865
rect 685 -885 715 -865
rect 735 -885 765 -865
rect 785 -885 815 -865
rect 835 -885 850 -865
rect 600 -900 850 -885
rect 900 -865 1150 -850
rect 900 -885 915 -865
rect 935 -885 965 -865
rect 985 -885 1015 -865
rect 1035 -885 1065 -865
rect 1085 -885 1115 -865
rect 1135 -885 1150 -865
rect 900 -900 1150 -885
rect 1200 -865 1450 -850
rect 1200 -885 1215 -865
rect 1235 -885 1265 -865
rect 1285 -885 1315 -865
rect 1335 -885 1365 -865
rect 1385 -885 1415 -865
rect 1435 -885 1450 -865
rect 1200 -900 1450 -885
rect 1500 -865 1750 -850
rect 1500 -885 1515 -865
rect 1535 -885 1565 -865
rect 1585 -885 1615 -865
rect 1635 -885 1665 -865
rect 1685 -885 1715 -865
rect 1735 -885 1750 -865
rect 1500 -900 1750 -885
rect 1800 -865 2050 -850
rect 1800 -885 1815 -865
rect 1835 -885 1865 -865
rect 1885 -885 1915 -865
rect 1935 -885 1965 -865
rect 1985 -885 2015 -865
rect 2035 -885 2050 -865
rect 1800 -900 2050 -885
rect 2100 -865 2350 -850
rect 2100 -885 2115 -865
rect 2135 -885 2165 -865
rect 2185 -885 2215 -865
rect 2235 -885 2265 -865
rect 2285 -885 2315 -865
rect 2335 -885 2350 -865
rect 2100 -900 2350 -885
rect 2400 -865 2650 -850
rect 2400 -885 2415 -865
rect 2435 -885 2465 -865
rect 2485 -885 2515 -865
rect 2535 -885 2565 -865
rect 2585 -885 2615 -865
rect 2635 -885 2650 -865
rect 2400 -900 2650 -885
rect 2700 -865 2950 -850
rect 2700 -885 2715 -865
rect 2735 -885 2765 -865
rect 2785 -885 2815 -865
rect 2835 -885 2865 -865
rect 2885 -885 2915 -865
rect 2935 -885 2950 -865
rect 2700 -900 2950 -885
rect 3000 -865 3250 -850
rect 3000 -885 3015 -865
rect 3035 -885 3065 -865
rect 3085 -885 3115 -865
rect 3135 -885 3165 -865
rect 3185 -885 3215 -865
rect 3235 -885 3250 -865
rect 3000 -900 3250 -885
rect 3300 -865 3550 -850
rect 3300 -885 3315 -865
rect 3335 -885 3365 -865
rect 3385 -885 3415 -865
rect 3435 -885 3465 -865
rect 3485 -885 3515 -865
rect 3535 -885 3550 -865
rect 3300 -900 3550 -885
rect 3600 -865 3850 -850
rect 3600 -885 3615 -865
rect 3635 -885 3665 -865
rect 3685 -885 3715 -865
rect 3735 -885 3765 -865
rect 3785 -885 3815 -865
rect 3835 -885 3850 -865
rect 3600 -900 3850 -885
rect 3900 -865 4150 -850
rect 3900 -885 3915 -865
rect 3935 -885 3965 -865
rect 3985 -885 4015 -865
rect 4035 -885 4065 -865
rect 4085 -885 4115 -865
rect 4135 -885 4150 -865
rect 3900 -900 4150 -885
rect 4200 -865 4450 -850
rect 4200 -885 4215 -865
rect 4235 -885 4265 -865
rect 4285 -885 4315 -865
rect 4335 -885 4365 -865
rect 4385 -885 4415 -865
rect 4435 -885 4450 -865
rect 4200 -900 4450 -885
rect 4500 -865 4750 -850
rect 4500 -885 4515 -865
rect 4535 -885 4565 -865
rect 4585 -885 4615 -865
rect 4635 -885 4665 -865
rect 4685 -885 4715 -865
rect 4735 -885 4750 -865
rect 4500 -900 4750 -885
rect 4800 -865 5050 -850
rect 4800 -885 4815 -865
rect 4835 -885 4865 -865
rect 4885 -885 4915 -865
rect 4935 -885 4965 -865
rect 4985 -885 5015 -865
rect 5035 -885 5050 -865
rect 4800 -900 5050 -885
rect 5100 -865 5350 -850
rect 5100 -885 5115 -865
rect 5135 -885 5165 -865
rect 5185 -885 5215 -865
rect 5235 -885 5265 -865
rect 5285 -885 5315 -865
rect 5335 -885 5350 -865
rect 5100 -900 5350 -885
rect 5400 -865 5650 -850
rect 5400 -885 5415 -865
rect 5435 -885 5465 -865
rect 5485 -885 5515 -865
rect 5535 -885 5565 -865
rect 5585 -885 5615 -865
rect 5635 -885 5650 -865
rect 5400 -900 5650 -885
rect 5700 -865 5950 -850
rect 5700 -885 5715 -865
rect 5735 -885 5765 -865
rect 5785 -885 5815 -865
rect 5835 -885 5865 -865
rect 5885 -885 5915 -865
rect 5935 -885 5950 -865
rect 5700 -900 5950 -885
rect 6000 -865 6250 -850
rect 6000 -885 6015 -865
rect 6035 -885 6065 -865
rect 6085 -885 6115 -865
rect 6135 -885 6165 -865
rect 6185 -885 6215 -865
rect 6235 -885 6250 -865
rect 6000 -900 6250 -885
rect 6300 -865 6550 -850
rect 6300 -885 6315 -865
rect 6335 -885 6365 -865
rect 6385 -885 6415 -865
rect 6435 -885 6465 -865
rect 6485 -885 6515 -865
rect 6535 -885 6550 -865
rect 6300 -900 6550 -885
rect 6600 -865 6850 -850
rect 6600 -885 6615 -865
rect 6635 -885 6665 -865
rect 6685 -885 6715 -865
rect 6735 -885 6765 -865
rect 6785 -885 6815 -865
rect 6835 -885 6850 -865
rect 6600 -900 6850 -885
rect 6900 -865 7150 -850
rect 6900 -885 6915 -865
rect 6935 -885 6965 -865
rect 6985 -885 7015 -865
rect 7035 -885 7065 -865
rect 7085 -885 7115 -865
rect 7135 -885 7150 -865
rect 6900 -900 7150 -885
rect 7200 -865 7450 -850
rect 7200 -885 7215 -865
rect 7235 -885 7265 -865
rect 7285 -885 7315 -865
rect 7335 -885 7365 -865
rect 7385 -885 7415 -865
rect 7435 -885 7450 -865
rect 7200 -900 7450 -885
rect 7500 -865 7750 -850
rect 7500 -885 7515 -865
rect 7535 -885 7565 -865
rect 7585 -885 7615 -865
rect 7635 -885 7665 -865
rect 7685 -885 7715 -865
rect 7735 -885 7750 -865
rect 7500 -900 7750 -885
rect 7800 -865 8050 -850
rect 7800 -885 7815 -865
rect 7835 -885 7865 -865
rect 7885 -885 7915 -865
rect 7935 -885 7965 -865
rect 7985 -885 8015 -865
rect 8035 -885 8050 -865
rect 7800 -900 8050 -885
rect 8100 -865 8350 -850
rect 8100 -885 8115 -865
rect 8135 -885 8165 -865
rect 8185 -885 8215 -865
rect 8235 -885 8265 -865
rect 8285 -885 8315 -865
rect 8335 -885 8350 -865
rect 8100 -900 8350 -885
rect 8400 -865 8650 -850
rect 8400 -885 8415 -865
rect 8435 -885 8465 -865
rect 8485 -885 8515 -865
rect 8535 -885 8565 -865
rect 8585 -885 8615 -865
rect 8635 -885 8650 -865
rect 8400 -900 8650 -885
rect 8700 -865 8950 -850
rect 8700 -885 8715 -865
rect 8735 -885 8765 -865
rect 8785 -885 8815 -865
rect 8835 -885 8865 -865
rect 8885 -885 8915 -865
rect 8935 -885 8950 -865
rect 8700 -900 8950 -885
rect 9000 -865 9250 -850
rect 9000 -885 9015 -865
rect 9035 -885 9065 -865
rect 9085 -885 9115 -865
rect 9135 -885 9165 -865
rect 9185 -885 9215 -865
rect 9235 -885 9250 -865
rect 9000 -900 9250 -885
rect 9300 -865 9550 -850
rect 9300 -885 9315 -865
rect 9335 -885 9365 -865
rect 9385 -885 9415 -865
rect 9435 -885 9465 -865
rect 9485 -885 9515 -865
rect 9535 -885 9550 -865
rect 9300 -900 9550 -885
rect 9600 -865 9850 -850
rect 9600 -885 9615 -865
rect 9635 -885 9665 -865
rect 9685 -885 9715 -865
rect 9735 -885 9765 -865
rect 9785 -885 9815 -865
rect 9835 -885 9850 -865
rect 9600 -900 9850 -885
rect 9900 -865 10150 -850
rect 9900 -885 9915 -865
rect 9935 -885 9965 -865
rect 9985 -885 10015 -865
rect 10035 -885 10065 -865
rect 10085 -885 10115 -865
rect 10135 -885 10150 -865
rect 9900 -900 10150 -885
rect 10200 -865 10450 -850
rect 10200 -885 10215 -865
rect 10235 -885 10265 -865
rect 10285 -885 10315 -865
rect 10335 -885 10365 -865
rect 10385 -885 10415 -865
rect 10435 -885 10450 -865
rect 10200 -900 10450 -885
rect 10500 -865 10750 -850
rect 10500 -885 10515 -865
rect 10535 -885 10565 -865
rect 10585 -885 10615 -865
rect 10635 -885 10665 -865
rect 10685 -885 10715 -865
rect 10735 -885 10750 -865
rect 10500 -900 10750 -885
rect 10800 -865 11050 -850
rect 10800 -885 10815 -865
rect 10835 -885 10865 -865
rect 10885 -885 10915 -865
rect 10935 -885 10965 -865
rect 10985 -885 11015 -865
rect 11035 -885 11050 -865
rect 10800 -900 11050 -885
rect 11100 -865 11350 -850
rect 11100 -885 11115 -865
rect 11135 -885 11165 -865
rect 11185 -885 11215 -865
rect 11235 -885 11265 -865
rect 11285 -885 11315 -865
rect 11335 -885 11350 -865
rect 11100 -900 11350 -885
rect 11400 -865 11650 -850
rect 11400 -885 11415 -865
rect 11435 -885 11465 -865
rect 11485 -885 11515 -865
rect 11535 -885 11565 -865
rect 11585 -885 11615 -865
rect 11635 -885 11650 -865
rect 11400 -900 11650 -885
rect 11700 -865 11950 -850
rect 11700 -885 11715 -865
rect 11735 -885 11765 -865
rect 11785 -885 11815 -865
rect 11835 -885 11865 -865
rect 11885 -885 11915 -865
rect 11935 -885 11950 -865
rect 11700 -900 11950 -885
rect 12000 -865 12250 -850
rect 12000 -885 12015 -865
rect 12035 -885 12065 -865
rect 12085 -885 12115 -865
rect 12135 -885 12165 -865
rect 12185 -885 12215 -865
rect 12235 -885 12250 -865
rect 12000 -900 12250 -885
rect 12300 -865 12550 -850
rect 12300 -885 12315 -865
rect 12335 -885 12365 -865
rect 12385 -885 12415 -865
rect 12435 -885 12465 -865
rect 12485 -885 12515 -865
rect 12535 -885 12550 -865
rect 12300 -900 12550 -885
rect 12600 -865 12850 -850
rect 12600 -885 12615 -865
rect 12635 -885 12665 -865
rect 12685 -885 12715 -865
rect 12735 -885 12765 -865
rect 12785 -885 12815 -865
rect 12835 -885 12850 -865
rect 12600 -900 12850 -885
rect 12900 -865 13150 -850
rect 12900 -885 12915 -865
rect 12935 -885 12965 -865
rect 12985 -885 13015 -865
rect 13035 -885 13065 -865
rect 13085 -885 13115 -865
rect 13135 -885 13150 -865
rect 12900 -900 13150 -885
rect 13200 -865 13450 -850
rect 13200 -885 13215 -865
rect 13235 -885 13265 -865
rect 13285 -885 13315 -865
rect 13335 -885 13365 -865
rect 13385 -885 13415 -865
rect 13435 -885 13450 -865
rect 13200 -900 13450 -885
rect 13500 -865 13750 -850
rect 13500 -885 13515 -865
rect 13535 -885 13565 -865
rect 13585 -885 13615 -865
rect 13635 -885 13665 -865
rect 13685 -885 13715 -865
rect 13735 -885 13750 -865
rect 13500 -900 13750 -885
rect 13800 -865 14050 -850
rect 13800 -885 13815 -865
rect 13835 -885 13865 -865
rect 13885 -885 13915 -865
rect 13935 -885 13965 -865
rect 13985 -885 14015 -865
rect 14035 -885 14050 -865
rect 13800 -900 14050 -885
rect 14100 -865 14350 -850
rect 14100 -885 14115 -865
rect 14135 -885 14165 -865
rect 14185 -885 14215 -865
rect 14235 -885 14265 -865
rect 14285 -885 14315 -865
rect 14335 -885 14350 -865
rect 14100 -900 14350 -885
rect 14400 -865 14650 -850
rect 14400 -885 14415 -865
rect 14435 -885 14465 -865
rect 14485 -885 14515 -865
rect 14535 -885 14565 -865
rect 14585 -885 14615 -865
rect 14635 -885 14650 -865
rect 14400 -900 14650 -885
rect 14700 -865 14950 -850
rect 14700 -885 14715 -865
rect 14735 -885 14765 -865
rect 14785 -885 14815 -865
rect 14835 -885 14865 -865
rect 14885 -885 14915 -865
rect 14935 -885 14950 -865
rect 14700 -900 14950 -885
rect 15000 -865 15250 -850
rect 15000 -885 15015 -865
rect 15035 -885 15065 -865
rect 15085 -885 15115 -865
rect 15135 -885 15165 -865
rect 15185 -885 15215 -865
rect 15235 -885 15250 -865
rect 15000 -900 15250 -885
rect 15300 -865 15550 -850
rect 15300 -885 15315 -865
rect 15335 -885 15365 -865
rect 15385 -885 15415 -865
rect 15435 -885 15465 -865
rect 15485 -885 15515 -865
rect 15535 -885 15550 -865
rect 15300 -900 15550 -885
rect 15600 -865 15850 -850
rect 15600 -885 15615 -865
rect 15635 -885 15665 -865
rect 15685 -885 15715 -865
rect 15735 -885 15765 -865
rect 15785 -885 15815 -865
rect 15835 -885 15850 -865
rect 15600 -900 15850 -885
rect 15900 -865 16150 -850
rect 15900 -885 15915 -865
rect 15935 -885 15965 -865
rect 15985 -885 16015 -865
rect 16035 -885 16065 -865
rect 16085 -885 16115 -865
rect 16135 -885 16150 -865
rect 15900 -900 16150 -885
rect 16200 -865 16450 -850
rect 16200 -885 16215 -865
rect 16235 -885 16265 -865
rect 16285 -885 16315 -865
rect 16335 -885 16365 -865
rect 16385 -885 16415 -865
rect 16435 -885 16450 -865
rect 16200 -900 16450 -885
rect 16500 -865 16750 -850
rect 16500 -885 16515 -865
rect 16535 -885 16565 -865
rect 16585 -885 16615 -865
rect 16635 -885 16665 -865
rect 16685 -885 16715 -865
rect 16735 -885 16750 -865
rect 16500 -900 16750 -885
rect 16800 -865 17050 -850
rect 16800 -885 16815 -865
rect 16835 -885 16865 -865
rect 16885 -885 16915 -865
rect 16935 -885 16965 -865
rect 16985 -885 17015 -865
rect 17035 -885 17050 -865
rect 16800 -900 17050 -885
rect 17100 -865 17350 -850
rect 17100 -885 17115 -865
rect 17135 -885 17165 -865
rect 17185 -885 17215 -865
rect 17235 -885 17265 -865
rect 17285 -885 17315 -865
rect 17335 -885 17350 -865
rect 17100 -900 17350 -885
rect 17400 -865 17650 -850
rect 17400 -885 17415 -865
rect 17435 -885 17465 -865
rect 17485 -885 17515 -865
rect 17535 -885 17565 -865
rect 17585 -885 17615 -865
rect 17635 -885 17650 -865
rect 17400 -900 17650 -885
rect 17700 -865 17950 -850
rect 17700 -885 17715 -865
rect 17735 -885 17765 -865
rect 17785 -885 17815 -865
rect 17835 -885 17865 -865
rect 17885 -885 17915 -865
rect 17935 -885 17950 -865
rect 17700 -900 17950 -885
rect 18000 -865 18250 -850
rect 18000 -885 18015 -865
rect 18035 -885 18065 -865
rect 18085 -885 18115 -865
rect 18135 -885 18165 -865
rect 18185 -885 18215 -865
rect 18235 -885 18250 -865
rect 18000 -900 18250 -885
rect 18300 -865 18550 -850
rect 18300 -885 18315 -865
rect 18335 -885 18365 -865
rect 18385 -885 18415 -865
rect 18435 -885 18465 -865
rect 18485 -885 18515 -865
rect 18535 -885 18550 -865
rect 18300 -900 18550 -885
rect 18600 -865 18850 -850
rect 18600 -885 18615 -865
rect 18635 -885 18665 -865
rect 18685 -885 18715 -865
rect 18735 -885 18765 -865
rect 18785 -885 18815 -865
rect 18835 -885 18850 -865
rect 18600 -900 18850 -885
rect 18900 -865 19150 -850
rect 18900 -885 18915 -865
rect 18935 -885 18965 -865
rect 18985 -885 19015 -865
rect 19035 -885 19065 -865
rect 19085 -885 19115 -865
rect 19135 -885 19150 -865
rect 18900 -900 19150 -885
rect 19200 -865 19450 -850
rect 19200 -885 19215 -865
rect 19235 -885 19265 -865
rect 19285 -885 19315 -865
rect 19335 -885 19365 -865
rect 19385 -885 19415 -865
rect 19435 -885 19450 -865
rect 19200 -900 19450 -885
rect 19500 -865 19750 -850
rect 19500 -885 19515 -865
rect 19535 -885 19565 -865
rect 19585 -885 19615 -865
rect 19635 -885 19665 -865
rect 19685 -885 19715 -865
rect 19735 -885 19750 -865
rect 19500 -900 19750 -885
rect 19800 -865 20050 -850
rect 19800 -885 19815 -865
rect 19835 -885 19865 -865
rect 19885 -885 19915 -865
rect 19935 -885 19965 -865
rect 19985 -885 20015 -865
rect 20035 -885 20050 -865
rect 19800 -900 20050 -885
rect 20100 -865 20350 -850
rect 20100 -885 20115 -865
rect 20135 -885 20165 -865
rect 20185 -885 20215 -865
rect 20235 -885 20265 -865
rect 20285 -885 20315 -865
rect 20335 -885 20350 -865
rect 20100 -900 20350 -885
rect 20400 -865 20650 -850
rect 20400 -885 20415 -865
rect 20435 -885 20465 -865
rect 20485 -885 20515 -865
rect 20535 -885 20565 -865
rect 20585 -885 20615 -865
rect 20635 -885 20650 -865
rect 20400 -900 20650 -885
rect 20700 -865 20950 -850
rect 20700 -885 20715 -865
rect 20735 -885 20765 -865
rect 20785 -885 20815 -865
rect 20835 -885 20865 -865
rect 20885 -885 20915 -865
rect 20935 -885 20950 -865
rect 20700 -900 20950 -885
rect 21000 -865 21250 -850
rect 21000 -885 21015 -865
rect 21035 -885 21065 -865
rect 21085 -885 21115 -865
rect 21135 -885 21165 -865
rect 21185 -885 21215 -865
rect 21235 -885 21250 -865
rect 21000 -900 21250 -885
rect 21300 -865 21550 -850
rect 21300 -885 21315 -865
rect 21335 -885 21365 -865
rect 21385 -885 21415 -865
rect 21435 -885 21465 -865
rect 21485 -885 21515 -865
rect 21535 -885 21550 -865
rect 21300 -900 21550 -885
rect 21600 -865 21850 -850
rect 21600 -885 21615 -865
rect 21635 -885 21665 -865
rect 21685 -885 21715 -865
rect 21735 -885 21765 -865
rect 21785 -885 21815 -865
rect 21835 -885 21850 -865
rect 21600 -900 21850 -885
rect 21900 -865 22150 -850
rect 21900 -885 21915 -865
rect 21935 -885 21965 -865
rect 21985 -885 22015 -865
rect 22035 -885 22065 -865
rect 22085 -885 22115 -865
rect 22135 -885 22150 -865
rect 21900 -900 22150 -885
rect 22200 -865 22450 -850
rect 22200 -885 22215 -865
rect 22235 -885 22265 -865
rect 22285 -885 22315 -865
rect 22335 -885 22365 -865
rect 22385 -885 22415 -865
rect 22435 -885 22450 -865
rect 22200 -900 22450 -885
rect 22500 -865 22750 -850
rect 22500 -885 22515 -865
rect 22535 -885 22565 -865
rect 22585 -885 22615 -865
rect 22635 -885 22665 -865
rect 22685 -885 22715 -865
rect 22735 -885 22750 -865
rect 22500 -900 22750 -885
rect 22800 -865 23050 -850
rect 22800 -885 22815 -865
rect 22835 -885 22865 -865
rect 22885 -885 22915 -865
rect 22935 -885 22965 -865
rect 22985 -885 23015 -865
rect 23035 -885 23050 -865
rect 22800 -900 23050 -885
rect 23100 -865 23350 -850
rect 23100 -885 23115 -865
rect 23135 -885 23165 -865
rect 23185 -885 23215 -865
rect 23235 -885 23265 -865
rect 23285 -885 23315 -865
rect 23335 -885 23350 -865
rect 23100 -900 23350 -885
rect 23400 -865 23650 -850
rect 23400 -885 23415 -865
rect 23435 -885 23465 -865
rect 23485 -885 23515 -865
rect 23535 -885 23565 -865
rect 23585 -885 23615 -865
rect 23635 -885 23650 -865
rect 23400 -900 23650 -885
rect 23700 -865 23950 -850
rect 23700 -885 23715 -865
rect 23735 -885 23765 -865
rect 23785 -885 23815 -865
rect 23835 -885 23865 -865
rect 23885 -885 23915 -865
rect 23935 -885 23950 -865
rect 23700 -900 23950 -885
rect 24000 -865 24250 -850
rect 24000 -885 24015 -865
rect 24035 -885 24065 -865
rect 24085 -885 24115 -865
rect 24135 -885 24165 -865
rect 24185 -885 24215 -865
rect 24235 -885 24250 -865
rect 24000 -900 24250 -885
rect 24300 -865 24550 -850
rect 24300 -885 24315 -865
rect 24335 -885 24365 -865
rect 24385 -885 24415 -865
rect 24435 -885 24465 -865
rect 24485 -885 24515 -865
rect 24535 -885 24550 -865
rect 24300 -900 24550 -885
rect 24600 -865 24850 -850
rect 24600 -885 24615 -865
rect 24635 -885 24665 -865
rect 24685 -885 24715 -865
rect 24735 -885 24765 -865
rect 24785 -885 24815 -865
rect 24835 -885 24850 -865
rect 24600 -900 24850 -885
rect 24900 -865 25150 -850
rect 24900 -885 24915 -865
rect 24935 -885 24965 -865
rect 24985 -885 25015 -865
rect 25035 -885 25065 -865
rect 25085 -885 25115 -865
rect 25135 -885 25150 -865
rect 24900 -900 25150 -885
rect 25200 -865 25450 -850
rect 25200 -885 25215 -865
rect 25235 -885 25265 -865
rect 25285 -885 25315 -865
rect 25335 -885 25365 -865
rect 25385 -885 25415 -865
rect 25435 -885 25450 -865
rect 25200 -900 25450 -885
rect 25500 -865 25750 -850
rect 25500 -885 25515 -865
rect 25535 -885 25565 -865
rect 25585 -885 25615 -865
rect 25635 -885 25665 -865
rect 25685 -885 25715 -865
rect 25735 -885 25750 -865
rect 25500 -900 25750 -885
rect 25800 -865 26050 -850
rect 25800 -885 25815 -865
rect 25835 -885 25865 -865
rect 25885 -885 25915 -865
rect 25935 -885 25965 -865
rect 25985 -885 26015 -865
rect 26035 -885 26050 -865
rect 25800 -900 26050 -885
rect 26100 -865 26350 -850
rect 26100 -885 26115 -865
rect 26135 -885 26165 -865
rect 26185 -885 26215 -865
rect 26235 -885 26265 -865
rect 26285 -885 26315 -865
rect 26335 -885 26350 -865
rect 26100 -900 26350 -885
rect 26400 -865 26650 -850
rect 26400 -885 26415 -865
rect 26435 -885 26465 -865
rect 26485 -885 26515 -865
rect 26535 -885 26565 -865
rect 26585 -885 26615 -865
rect 26635 -885 26650 -865
rect 26400 -900 26650 -885
rect 26700 -865 26950 -850
rect 26700 -885 26715 -865
rect 26735 -885 26765 -865
rect 26785 -885 26815 -865
rect 26835 -885 26865 -865
rect 26885 -885 26915 -865
rect 26935 -885 26950 -865
rect 26700 -900 26950 -885
rect 27000 -865 27250 -850
rect 27000 -885 27015 -865
rect 27035 -885 27065 -865
rect 27085 -885 27115 -865
rect 27135 -885 27165 -865
rect 27185 -885 27215 -865
rect 27235 -885 27250 -865
rect 27000 -900 27250 -885
rect 27300 -865 27550 -850
rect 27300 -885 27315 -865
rect 27335 -885 27365 -865
rect 27385 -885 27415 -865
rect 27435 -885 27465 -865
rect 27485 -885 27515 -865
rect 27535 -885 27550 -865
rect 27300 -900 27550 -885
rect 27600 -865 27850 -850
rect 27600 -885 27615 -865
rect 27635 -885 27665 -865
rect 27685 -885 27715 -865
rect 27735 -885 27765 -865
rect 27785 -885 27815 -865
rect 27835 -885 27850 -865
rect 27600 -900 27850 -885
rect 27900 -865 28150 -850
rect 27900 -885 27915 -865
rect 27935 -885 27965 -865
rect 27985 -885 28015 -865
rect 28035 -885 28065 -865
rect 28085 -885 28115 -865
rect 28135 -885 28150 -865
rect 27900 -900 28150 -885
rect 28200 -865 28450 -850
rect 28200 -885 28215 -865
rect 28235 -885 28265 -865
rect 28285 -885 28315 -865
rect 28335 -885 28365 -865
rect 28385 -885 28415 -865
rect 28435 -885 28450 -865
rect 28200 -900 28450 -885
rect 28500 -865 28750 -850
rect 28500 -885 28515 -865
rect 28535 -885 28565 -865
rect 28585 -885 28615 -865
rect 28635 -885 28665 -865
rect 28685 -885 28715 -865
rect 28735 -885 28750 -865
rect 28500 -900 28750 -885
rect -650 -965 -600 -950
rect -650 -985 -635 -965
rect -615 -985 -600 -965
rect -650 -1015 -600 -985
rect -650 -1035 -635 -1015
rect -615 -1035 -600 -1015
rect -650 -1065 -600 -1035
rect -650 -1085 -635 -1065
rect -615 -1085 -600 -1065
rect -650 -1115 -600 -1085
rect -650 -1135 -635 -1115
rect -615 -1135 -600 -1115
rect -650 -1165 -600 -1135
rect -650 -1185 -635 -1165
rect -615 -1185 -600 -1165
rect -650 -1215 -600 -1185
rect -650 -1235 -635 -1215
rect -615 -1235 -600 -1215
rect -650 -1265 -600 -1235
rect -650 -1285 -635 -1265
rect -615 -1285 -600 -1265
rect -650 -1315 -600 -1285
rect -650 -1335 -635 -1315
rect -615 -1335 -600 -1315
rect -650 -1365 -600 -1335
rect -650 -1385 -635 -1365
rect -615 -1385 -600 -1365
rect -650 -1415 -600 -1385
rect -650 -1435 -635 -1415
rect -615 -1435 -600 -1415
rect -650 -1465 -600 -1435
rect -650 -1485 -635 -1465
rect -615 -1485 -600 -1465
rect -650 -1515 -600 -1485
rect -650 -1535 -635 -1515
rect -615 -1535 -600 -1515
rect -650 -1565 -600 -1535
rect -650 -1585 -635 -1565
rect -615 -1585 -600 -1565
rect -650 -1615 -600 -1585
rect -650 -1635 -635 -1615
rect -615 -1635 -600 -1615
rect -650 -1650 -600 -1635
rect -500 -965 -450 -950
rect -500 -985 -485 -965
rect -465 -985 -450 -965
rect -500 -1015 -450 -985
rect -500 -1035 -485 -1015
rect -465 -1035 -450 -1015
rect -500 -1065 -450 -1035
rect -500 -1085 -485 -1065
rect -465 -1085 -450 -1065
rect -500 -1115 -450 -1085
rect -500 -1135 -485 -1115
rect -465 -1135 -450 -1115
rect -500 -1165 -450 -1135
rect -500 -1185 -485 -1165
rect -465 -1185 -450 -1165
rect -500 -1215 -450 -1185
rect -500 -1235 -485 -1215
rect -465 -1235 -450 -1215
rect -500 -1265 -450 -1235
rect -500 -1285 -485 -1265
rect -465 -1285 -450 -1265
rect -500 -1315 -450 -1285
rect -500 -1335 -485 -1315
rect -465 -1335 -450 -1315
rect -500 -1365 -450 -1335
rect -500 -1385 -485 -1365
rect -465 -1385 -450 -1365
rect -500 -1415 -450 -1385
rect -500 -1435 -485 -1415
rect -465 -1435 -450 -1415
rect -500 -1465 -450 -1435
rect -500 -1485 -485 -1465
rect -465 -1485 -450 -1465
rect -500 -1515 -450 -1485
rect -500 -1535 -485 -1515
rect -465 -1535 -450 -1515
rect -500 -1565 -450 -1535
rect -500 -1585 -485 -1565
rect -465 -1585 -450 -1565
rect -500 -1615 -450 -1585
rect -500 -1635 -485 -1615
rect -465 -1635 -450 -1615
rect -500 -1650 -450 -1635
rect -350 -965 -300 -950
rect -350 -985 -335 -965
rect -315 -985 -300 -965
rect -350 -1015 -300 -985
rect -350 -1035 -335 -1015
rect -315 -1035 -300 -1015
rect -350 -1065 -300 -1035
rect -350 -1085 -335 -1065
rect -315 -1085 -300 -1065
rect -350 -1115 -300 -1085
rect -350 -1135 -335 -1115
rect -315 -1135 -300 -1115
rect -350 -1165 -300 -1135
rect -350 -1185 -335 -1165
rect -315 -1185 -300 -1165
rect -350 -1215 -300 -1185
rect -350 -1235 -335 -1215
rect -315 -1235 -300 -1215
rect -350 -1265 -300 -1235
rect -350 -1285 -335 -1265
rect -315 -1285 -300 -1265
rect -350 -1315 -300 -1285
rect -350 -1335 -335 -1315
rect -315 -1335 -300 -1315
rect -350 -1365 -300 -1335
rect -350 -1385 -335 -1365
rect -315 -1385 -300 -1365
rect -350 -1415 -300 -1385
rect -350 -1435 -335 -1415
rect -315 -1435 -300 -1415
rect -350 -1465 -300 -1435
rect -350 -1485 -335 -1465
rect -315 -1485 -300 -1465
rect -350 -1515 -300 -1485
rect -350 -1535 -335 -1515
rect -315 -1535 -300 -1515
rect -350 -1565 -300 -1535
rect -350 -1585 -335 -1565
rect -315 -1585 -300 -1565
rect -350 -1615 -300 -1585
rect -350 -1635 -335 -1615
rect -315 -1635 -300 -1615
rect -350 -1650 -300 -1635
rect -200 -965 -150 -950
rect -200 -985 -185 -965
rect -165 -985 -150 -965
rect -200 -1015 -150 -985
rect -200 -1035 -185 -1015
rect -165 -1035 -150 -1015
rect -200 -1065 -150 -1035
rect -200 -1085 -185 -1065
rect -165 -1085 -150 -1065
rect -200 -1115 -150 -1085
rect -200 -1135 -185 -1115
rect -165 -1135 -150 -1115
rect -200 -1165 -150 -1135
rect -200 -1185 -185 -1165
rect -165 -1185 -150 -1165
rect -200 -1215 -150 -1185
rect -200 -1235 -185 -1215
rect -165 -1235 -150 -1215
rect -200 -1265 -150 -1235
rect -200 -1285 -185 -1265
rect -165 -1285 -150 -1265
rect -200 -1315 -150 -1285
rect -200 -1335 -185 -1315
rect -165 -1335 -150 -1315
rect -200 -1365 -150 -1335
rect -200 -1385 -185 -1365
rect -165 -1385 -150 -1365
rect -200 -1415 -150 -1385
rect -200 -1435 -185 -1415
rect -165 -1435 -150 -1415
rect -200 -1465 -150 -1435
rect -200 -1485 -185 -1465
rect -165 -1485 -150 -1465
rect -200 -1515 -150 -1485
rect -200 -1535 -185 -1515
rect -165 -1535 -150 -1515
rect -200 -1565 -150 -1535
rect -200 -1585 -185 -1565
rect -165 -1585 -150 -1565
rect -200 -1615 -150 -1585
rect -200 -1635 -185 -1615
rect -165 -1635 -150 -1615
rect -200 -1650 -150 -1635
rect -50 -965 0 -950
rect -50 -985 -35 -965
rect -15 -985 0 -965
rect -50 -1015 0 -985
rect -50 -1035 -35 -1015
rect -15 -1035 0 -1015
rect -50 -1065 0 -1035
rect -50 -1085 -35 -1065
rect -15 -1085 0 -1065
rect -50 -1115 0 -1085
rect -50 -1135 -35 -1115
rect -15 -1135 0 -1115
rect -50 -1165 0 -1135
rect -50 -1185 -35 -1165
rect -15 -1185 0 -1165
rect -50 -1215 0 -1185
rect -50 -1235 -35 -1215
rect -15 -1235 0 -1215
rect -50 -1265 0 -1235
rect -50 -1285 -35 -1265
rect -15 -1285 0 -1265
rect -50 -1315 0 -1285
rect -50 -1335 -35 -1315
rect -15 -1335 0 -1315
rect -50 -1365 0 -1335
rect -50 -1385 -35 -1365
rect -15 -1385 0 -1365
rect -50 -1415 0 -1385
rect -50 -1435 -35 -1415
rect -15 -1435 0 -1415
rect -50 -1465 0 -1435
rect -50 -1485 -35 -1465
rect -15 -1485 0 -1465
rect -50 -1515 0 -1485
rect -50 -1535 -35 -1515
rect -15 -1535 0 -1515
rect -50 -1565 0 -1535
rect -50 -1585 -35 -1565
rect -15 -1585 0 -1565
rect -50 -1615 0 -1585
rect -50 -1635 -35 -1615
rect -15 -1635 0 -1615
rect -50 -1650 0 -1635
rect 1150 -965 1200 -950
rect 1150 -985 1165 -965
rect 1185 -985 1200 -965
rect 1150 -1015 1200 -985
rect 1150 -1035 1165 -1015
rect 1185 -1035 1200 -1015
rect 1150 -1065 1200 -1035
rect 1150 -1085 1165 -1065
rect 1185 -1085 1200 -1065
rect 1150 -1115 1200 -1085
rect 1150 -1135 1165 -1115
rect 1185 -1135 1200 -1115
rect 1150 -1165 1200 -1135
rect 1150 -1185 1165 -1165
rect 1185 -1185 1200 -1165
rect 1150 -1215 1200 -1185
rect 1150 -1235 1165 -1215
rect 1185 -1235 1200 -1215
rect 1150 -1265 1200 -1235
rect 1150 -1285 1165 -1265
rect 1185 -1285 1200 -1265
rect 1150 -1315 1200 -1285
rect 1150 -1335 1165 -1315
rect 1185 -1335 1200 -1315
rect 1150 -1365 1200 -1335
rect 1150 -1385 1165 -1365
rect 1185 -1385 1200 -1365
rect 1150 -1415 1200 -1385
rect 1150 -1435 1165 -1415
rect 1185 -1435 1200 -1415
rect 1150 -1465 1200 -1435
rect 1150 -1485 1165 -1465
rect 1185 -1485 1200 -1465
rect 1150 -1515 1200 -1485
rect 1150 -1535 1165 -1515
rect 1185 -1535 1200 -1515
rect 1150 -1565 1200 -1535
rect 1150 -1585 1165 -1565
rect 1185 -1585 1200 -1565
rect 1150 -1615 1200 -1585
rect 1150 -1635 1165 -1615
rect 1185 -1635 1200 -1615
rect 1150 -1650 1200 -1635
rect 1450 -965 1500 -950
rect 1450 -985 1465 -965
rect 1485 -985 1500 -965
rect 1450 -1015 1500 -985
rect 1450 -1035 1465 -1015
rect 1485 -1035 1500 -1015
rect 1450 -1065 1500 -1035
rect 1450 -1085 1465 -1065
rect 1485 -1085 1500 -1065
rect 1450 -1115 1500 -1085
rect 1450 -1135 1465 -1115
rect 1485 -1135 1500 -1115
rect 1450 -1165 1500 -1135
rect 1450 -1185 1465 -1165
rect 1485 -1185 1500 -1165
rect 1450 -1215 1500 -1185
rect 1450 -1235 1465 -1215
rect 1485 -1235 1500 -1215
rect 1450 -1265 1500 -1235
rect 1450 -1285 1465 -1265
rect 1485 -1285 1500 -1265
rect 1450 -1315 1500 -1285
rect 1450 -1335 1465 -1315
rect 1485 -1335 1500 -1315
rect 1450 -1365 1500 -1335
rect 1450 -1385 1465 -1365
rect 1485 -1385 1500 -1365
rect 1450 -1415 1500 -1385
rect 1450 -1435 1465 -1415
rect 1485 -1435 1500 -1415
rect 1450 -1465 1500 -1435
rect 1450 -1485 1465 -1465
rect 1485 -1485 1500 -1465
rect 1450 -1515 1500 -1485
rect 1450 -1535 1465 -1515
rect 1485 -1535 1500 -1515
rect 1450 -1565 1500 -1535
rect 1450 -1585 1465 -1565
rect 1485 -1585 1500 -1565
rect 1450 -1615 1500 -1585
rect 1450 -1635 1465 -1615
rect 1485 -1635 1500 -1615
rect 1450 -1650 1500 -1635
rect 1750 -965 1800 -950
rect 1750 -985 1765 -965
rect 1785 -985 1800 -965
rect 1750 -1015 1800 -985
rect 1750 -1035 1765 -1015
rect 1785 -1035 1800 -1015
rect 1750 -1065 1800 -1035
rect 1750 -1085 1765 -1065
rect 1785 -1085 1800 -1065
rect 1750 -1115 1800 -1085
rect 1750 -1135 1765 -1115
rect 1785 -1135 1800 -1115
rect 1750 -1165 1800 -1135
rect 1750 -1185 1765 -1165
rect 1785 -1185 1800 -1165
rect 1750 -1215 1800 -1185
rect 1750 -1235 1765 -1215
rect 1785 -1235 1800 -1215
rect 1750 -1265 1800 -1235
rect 1750 -1285 1765 -1265
rect 1785 -1285 1800 -1265
rect 1750 -1315 1800 -1285
rect 1750 -1335 1765 -1315
rect 1785 -1335 1800 -1315
rect 1750 -1365 1800 -1335
rect 1750 -1385 1765 -1365
rect 1785 -1385 1800 -1365
rect 1750 -1415 1800 -1385
rect 1750 -1435 1765 -1415
rect 1785 -1435 1800 -1415
rect 1750 -1465 1800 -1435
rect 1750 -1485 1765 -1465
rect 1785 -1485 1800 -1465
rect 1750 -1515 1800 -1485
rect 1750 -1535 1765 -1515
rect 1785 -1535 1800 -1515
rect 1750 -1565 1800 -1535
rect 1750 -1585 1765 -1565
rect 1785 -1585 1800 -1565
rect 1750 -1615 1800 -1585
rect 1750 -1635 1765 -1615
rect 1785 -1635 1800 -1615
rect 1750 -1650 1800 -1635
rect 2050 -965 2100 -950
rect 2050 -985 2065 -965
rect 2085 -985 2100 -965
rect 2050 -1015 2100 -985
rect 2050 -1035 2065 -1015
rect 2085 -1035 2100 -1015
rect 2050 -1065 2100 -1035
rect 2050 -1085 2065 -1065
rect 2085 -1085 2100 -1065
rect 2050 -1115 2100 -1085
rect 2050 -1135 2065 -1115
rect 2085 -1135 2100 -1115
rect 2050 -1165 2100 -1135
rect 2050 -1185 2065 -1165
rect 2085 -1185 2100 -1165
rect 2050 -1215 2100 -1185
rect 2050 -1235 2065 -1215
rect 2085 -1235 2100 -1215
rect 2050 -1265 2100 -1235
rect 2050 -1285 2065 -1265
rect 2085 -1285 2100 -1265
rect 2050 -1315 2100 -1285
rect 2050 -1335 2065 -1315
rect 2085 -1335 2100 -1315
rect 2050 -1365 2100 -1335
rect 2050 -1385 2065 -1365
rect 2085 -1385 2100 -1365
rect 2050 -1415 2100 -1385
rect 2050 -1435 2065 -1415
rect 2085 -1435 2100 -1415
rect 2050 -1465 2100 -1435
rect 2050 -1485 2065 -1465
rect 2085 -1485 2100 -1465
rect 2050 -1515 2100 -1485
rect 2050 -1535 2065 -1515
rect 2085 -1535 2100 -1515
rect 2050 -1565 2100 -1535
rect 2050 -1585 2065 -1565
rect 2085 -1585 2100 -1565
rect 2050 -1615 2100 -1585
rect 2050 -1635 2065 -1615
rect 2085 -1635 2100 -1615
rect 2050 -1650 2100 -1635
rect 2350 -965 2400 -950
rect 2350 -985 2365 -965
rect 2385 -985 2400 -965
rect 2350 -1015 2400 -985
rect 2350 -1035 2365 -1015
rect 2385 -1035 2400 -1015
rect 2350 -1065 2400 -1035
rect 2350 -1085 2365 -1065
rect 2385 -1085 2400 -1065
rect 2350 -1115 2400 -1085
rect 2350 -1135 2365 -1115
rect 2385 -1135 2400 -1115
rect 2350 -1165 2400 -1135
rect 2350 -1185 2365 -1165
rect 2385 -1185 2400 -1165
rect 2350 -1215 2400 -1185
rect 2350 -1235 2365 -1215
rect 2385 -1235 2400 -1215
rect 2350 -1265 2400 -1235
rect 2350 -1285 2365 -1265
rect 2385 -1285 2400 -1265
rect 2350 -1315 2400 -1285
rect 2350 -1335 2365 -1315
rect 2385 -1335 2400 -1315
rect 2350 -1365 2400 -1335
rect 2350 -1385 2365 -1365
rect 2385 -1385 2400 -1365
rect 2350 -1415 2400 -1385
rect 2350 -1435 2365 -1415
rect 2385 -1435 2400 -1415
rect 2350 -1465 2400 -1435
rect 2350 -1485 2365 -1465
rect 2385 -1485 2400 -1465
rect 2350 -1515 2400 -1485
rect 2350 -1535 2365 -1515
rect 2385 -1535 2400 -1515
rect 2350 -1565 2400 -1535
rect 2350 -1585 2365 -1565
rect 2385 -1585 2400 -1565
rect 2350 -1615 2400 -1585
rect 2350 -1635 2365 -1615
rect 2385 -1635 2400 -1615
rect 2350 -1650 2400 -1635
rect 2650 -965 2700 -950
rect 2650 -985 2665 -965
rect 2685 -985 2700 -965
rect 2650 -1015 2700 -985
rect 2650 -1035 2665 -1015
rect 2685 -1035 2700 -1015
rect 2650 -1065 2700 -1035
rect 2650 -1085 2665 -1065
rect 2685 -1085 2700 -1065
rect 2650 -1115 2700 -1085
rect 2650 -1135 2665 -1115
rect 2685 -1135 2700 -1115
rect 2650 -1165 2700 -1135
rect 2650 -1185 2665 -1165
rect 2685 -1185 2700 -1165
rect 2650 -1215 2700 -1185
rect 2650 -1235 2665 -1215
rect 2685 -1235 2700 -1215
rect 2650 -1265 2700 -1235
rect 2650 -1285 2665 -1265
rect 2685 -1285 2700 -1265
rect 2650 -1315 2700 -1285
rect 2650 -1335 2665 -1315
rect 2685 -1335 2700 -1315
rect 2650 -1365 2700 -1335
rect 2650 -1385 2665 -1365
rect 2685 -1385 2700 -1365
rect 2650 -1415 2700 -1385
rect 2650 -1435 2665 -1415
rect 2685 -1435 2700 -1415
rect 2650 -1465 2700 -1435
rect 2650 -1485 2665 -1465
rect 2685 -1485 2700 -1465
rect 2650 -1515 2700 -1485
rect 2650 -1535 2665 -1515
rect 2685 -1535 2700 -1515
rect 2650 -1565 2700 -1535
rect 2650 -1585 2665 -1565
rect 2685 -1585 2700 -1565
rect 2650 -1615 2700 -1585
rect 2650 -1635 2665 -1615
rect 2685 -1635 2700 -1615
rect 2650 -1650 2700 -1635
rect 2950 -965 3000 -950
rect 2950 -985 2965 -965
rect 2985 -985 3000 -965
rect 2950 -1015 3000 -985
rect 2950 -1035 2965 -1015
rect 2985 -1035 3000 -1015
rect 2950 -1065 3000 -1035
rect 2950 -1085 2965 -1065
rect 2985 -1085 3000 -1065
rect 2950 -1115 3000 -1085
rect 2950 -1135 2965 -1115
rect 2985 -1135 3000 -1115
rect 2950 -1165 3000 -1135
rect 2950 -1185 2965 -1165
rect 2985 -1185 3000 -1165
rect 2950 -1215 3000 -1185
rect 2950 -1235 2965 -1215
rect 2985 -1235 3000 -1215
rect 2950 -1265 3000 -1235
rect 2950 -1285 2965 -1265
rect 2985 -1285 3000 -1265
rect 2950 -1315 3000 -1285
rect 2950 -1335 2965 -1315
rect 2985 -1335 3000 -1315
rect 2950 -1365 3000 -1335
rect 2950 -1385 2965 -1365
rect 2985 -1385 3000 -1365
rect 2950 -1415 3000 -1385
rect 2950 -1435 2965 -1415
rect 2985 -1435 3000 -1415
rect 2950 -1465 3000 -1435
rect 2950 -1485 2965 -1465
rect 2985 -1485 3000 -1465
rect 2950 -1515 3000 -1485
rect 2950 -1535 2965 -1515
rect 2985 -1535 3000 -1515
rect 2950 -1565 3000 -1535
rect 2950 -1585 2965 -1565
rect 2985 -1585 3000 -1565
rect 2950 -1615 3000 -1585
rect 2950 -1635 2965 -1615
rect 2985 -1635 3000 -1615
rect 2950 -1650 3000 -1635
rect 3250 -965 3300 -950
rect 3250 -985 3265 -965
rect 3285 -985 3300 -965
rect 3250 -1015 3300 -985
rect 3250 -1035 3265 -1015
rect 3285 -1035 3300 -1015
rect 3250 -1065 3300 -1035
rect 3250 -1085 3265 -1065
rect 3285 -1085 3300 -1065
rect 3250 -1115 3300 -1085
rect 3250 -1135 3265 -1115
rect 3285 -1135 3300 -1115
rect 3250 -1165 3300 -1135
rect 3250 -1185 3265 -1165
rect 3285 -1185 3300 -1165
rect 3250 -1215 3300 -1185
rect 3250 -1235 3265 -1215
rect 3285 -1235 3300 -1215
rect 3250 -1265 3300 -1235
rect 3250 -1285 3265 -1265
rect 3285 -1285 3300 -1265
rect 3250 -1315 3300 -1285
rect 3250 -1335 3265 -1315
rect 3285 -1335 3300 -1315
rect 3250 -1365 3300 -1335
rect 3250 -1385 3265 -1365
rect 3285 -1385 3300 -1365
rect 3250 -1415 3300 -1385
rect 3250 -1435 3265 -1415
rect 3285 -1435 3300 -1415
rect 3250 -1465 3300 -1435
rect 3250 -1485 3265 -1465
rect 3285 -1485 3300 -1465
rect 3250 -1515 3300 -1485
rect 3250 -1535 3265 -1515
rect 3285 -1535 3300 -1515
rect 3250 -1565 3300 -1535
rect 3250 -1585 3265 -1565
rect 3285 -1585 3300 -1565
rect 3250 -1615 3300 -1585
rect 3250 -1635 3265 -1615
rect 3285 -1635 3300 -1615
rect 3250 -1650 3300 -1635
rect 3550 -965 3600 -950
rect 3550 -985 3565 -965
rect 3585 -985 3600 -965
rect 3550 -1015 3600 -985
rect 3550 -1035 3565 -1015
rect 3585 -1035 3600 -1015
rect 3550 -1065 3600 -1035
rect 3550 -1085 3565 -1065
rect 3585 -1085 3600 -1065
rect 3550 -1115 3600 -1085
rect 3550 -1135 3565 -1115
rect 3585 -1135 3600 -1115
rect 3550 -1165 3600 -1135
rect 3550 -1185 3565 -1165
rect 3585 -1185 3600 -1165
rect 3550 -1215 3600 -1185
rect 3550 -1235 3565 -1215
rect 3585 -1235 3600 -1215
rect 3550 -1265 3600 -1235
rect 3550 -1285 3565 -1265
rect 3585 -1285 3600 -1265
rect 3550 -1315 3600 -1285
rect 3550 -1335 3565 -1315
rect 3585 -1335 3600 -1315
rect 3550 -1365 3600 -1335
rect 3550 -1385 3565 -1365
rect 3585 -1385 3600 -1365
rect 3550 -1415 3600 -1385
rect 3550 -1435 3565 -1415
rect 3585 -1435 3600 -1415
rect 3550 -1465 3600 -1435
rect 3550 -1485 3565 -1465
rect 3585 -1485 3600 -1465
rect 3550 -1515 3600 -1485
rect 3550 -1535 3565 -1515
rect 3585 -1535 3600 -1515
rect 3550 -1565 3600 -1535
rect 3550 -1585 3565 -1565
rect 3585 -1585 3600 -1565
rect 3550 -1615 3600 -1585
rect 3550 -1635 3565 -1615
rect 3585 -1635 3600 -1615
rect 3550 -1650 3600 -1635
rect 3700 -965 3750 -950
rect 3700 -985 3715 -965
rect 3735 -985 3750 -965
rect 3700 -1015 3750 -985
rect 3700 -1035 3715 -1015
rect 3735 -1035 3750 -1015
rect 3700 -1065 3750 -1035
rect 3700 -1085 3715 -1065
rect 3735 -1085 3750 -1065
rect 3700 -1115 3750 -1085
rect 3700 -1135 3715 -1115
rect 3735 -1135 3750 -1115
rect 3700 -1165 3750 -1135
rect 3700 -1185 3715 -1165
rect 3735 -1185 3750 -1165
rect 3700 -1215 3750 -1185
rect 3700 -1235 3715 -1215
rect 3735 -1235 3750 -1215
rect 3700 -1265 3750 -1235
rect 3700 -1285 3715 -1265
rect 3735 -1285 3750 -1265
rect 3700 -1315 3750 -1285
rect 3700 -1335 3715 -1315
rect 3735 -1335 3750 -1315
rect 3700 -1365 3750 -1335
rect 3700 -1385 3715 -1365
rect 3735 -1385 3750 -1365
rect 3700 -1415 3750 -1385
rect 3700 -1435 3715 -1415
rect 3735 -1435 3750 -1415
rect 3700 -1465 3750 -1435
rect 3700 -1485 3715 -1465
rect 3735 -1485 3750 -1465
rect 3700 -1515 3750 -1485
rect 3700 -1535 3715 -1515
rect 3735 -1535 3750 -1515
rect 3700 -1565 3750 -1535
rect 3700 -1585 3715 -1565
rect 3735 -1585 3750 -1565
rect 3700 -1615 3750 -1585
rect 3700 -1635 3715 -1615
rect 3735 -1635 3750 -1615
rect 3700 -1650 3750 -1635
rect 3850 -965 3900 -950
rect 3850 -985 3865 -965
rect 3885 -985 3900 -965
rect 3850 -1015 3900 -985
rect 3850 -1035 3865 -1015
rect 3885 -1035 3900 -1015
rect 3850 -1065 3900 -1035
rect 3850 -1085 3865 -1065
rect 3885 -1085 3900 -1065
rect 3850 -1115 3900 -1085
rect 3850 -1135 3865 -1115
rect 3885 -1135 3900 -1115
rect 3850 -1165 3900 -1135
rect 3850 -1185 3865 -1165
rect 3885 -1185 3900 -1165
rect 3850 -1215 3900 -1185
rect 3850 -1235 3865 -1215
rect 3885 -1235 3900 -1215
rect 3850 -1265 3900 -1235
rect 3850 -1285 3865 -1265
rect 3885 -1285 3900 -1265
rect 3850 -1315 3900 -1285
rect 3850 -1335 3865 -1315
rect 3885 -1335 3900 -1315
rect 3850 -1365 3900 -1335
rect 3850 -1385 3865 -1365
rect 3885 -1385 3900 -1365
rect 3850 -1415 3900 -1385
rect 3850 -1435 3865 -1415
rect 3885 -1435 3900 -1415
rect 3850 -1465 3900 -1435
rect 3850 -1485 3865 -1465
rect 3885 -1485 3900 -1465
rect 3850 -1515 3900 -1485
rect 3850 -1535 3865 -1515
rect 3885 -1535 3900 -1515
rect 3850 -1565 3900 -1535
rect 3850 -1585 3865 -1565
rect 3885 -1585 3900 -1565
rect 3850 -1615 3900 -1585
rect 3850 -1635 3865 -1615
rect 3885 -1635 3900 -1615
rect 3850 -1650 3900 -1635
rect 4000 -965 4050 -950
rect 4000 -985 4015 -965
rect 4035 -985 4050 -965
rect 4000 -1015 4050 -985
rect 4000 -1035 4015 -1015
rect 4035 -1035 4050 -1015
rect 4000 -1065 4050 -1035
rect 4000 -1085 4015 -1065
rect 4035 -1085 4050 -1065
rect 4000 -1115 4050 -1085
rect 4000 -1135 4015 -1115
rect 4035 -1135 4050 -1115
rect 4000 -1165 4050 -1135
rect 4000 -1185 4015 -1165
rect 4035 -1185 4050 -1165
rect 4000 -1215 4050 -1185
rect 4000 -1235 4015 -1215
rect 4035 -1235 4050 -1215
rect 4000 -1265 4050 -1235
rect 4000 -1285 4015 -1265
rect 4035 -1285 4050 -1265
rect 4000 -1315 4050 -1285
rect 4000 -1335 4015 -1315
rect 4035 -1335 4050 -1315
rect 4000 -1365 4050 -1335
rect 4000 -1385 4015 -1365
rect 4035 -1385 4050 -1365
rect 4000 -1415 4050 -1385
rect 4000 -1435 4015 -1415
rect 4035 -1435 4050 -1415
rect 4000 -1465 4050 -1435
rect 4000 -1485 4015 -1465
rect 4035 -1485 4050 -1465
rect 4000 -1515 4050 -1485
rect 4000 -1535 4015 -1515
rect 4035 -1535 4050 -1515
rect 4000 -1565 4050 -1535
rect 4000 -1585 4015 -1565
rect 4035 -1585 4050 -1565
rect 4000 -1615 4050 -1585
rect 4000 -1635 4015 -1615
rect 4035 -1635 4050 -1615
rect 4000 -1650 4050 -1635
rect 4150 -965 4200 -950
rect 4150 -985 4165 -965
rect 4185 -985 4200 -965
rect 4150 -1015 4200 -985
rect 4150 -1035 4165 -1015
rect 4185 -1035 4200 -1015
rect 4150 -1065 4200 -1035
rect 4150 -1085 4165 -1065
rect 4185 -1085 4200 -1065
rect 4150 -1115 4200 -1085
rect 4150 -1135 4165 -1115
rect 4185 -1135 4200 -1115
rect 4150 -1165 4200 -1135
rect 4150 -1185 4165 -1165
rect 4185 -1185 4200 -1165
rect 4150 -1215 4200 -1185
rect 4150 -1235 4165 -1215
rect 4185 -1235 4200 -1215
rect 4150 -1265 4200 -1235
rect 4150 -1285 4165 -1265
rect 4185 -1285 4200 -1265
rect 4150 -1315 4200 -1285
rect 4150 -1335 4165 -1315
rect 4185 -1335 4200 -1315
rect 4150 -1365 4200 -1335
rect 4150 -1385 4165 -1365
rect 4185 -1385 4200 -1365
rect 4150 -1415 4200 -1385
rect 4150 -1435 4165 -1415
rect 4185 -1435 4200 -1415
rect 4150 -1465 4200 -1435
rect 4150 -1485 4165 -1465
rect 4185 -1485 4200 -1465
rect 4150 -1515 4200 -1485
rect 4150 -1535 4165 -1515
rect 4185 -1535 4200 -1515
rect 4150 -1565 4200 -1535
rect 4150 -1585 4165 -1565
rect 4185 -1585 4200 -1565
rect 4150 -1615 4200 -1585
rect 4150 -1635 4165 -1615
rect 4185 -1635 4200 -1615
rect 4150 -1650 4200 -1635
rect 4300 -965 4350 -950
rect 4300 -985 4315 -965
rect 4335 -985 4350 -965
rect 4300 -1015 4350 -985
rect 4300 -1035 4315 -1015
rect 4335 -1035 4350 -1015
rect 4300 -1065 4350 -1035
rect 4300 -1085 4315 -1065
rect 4335 -1085 4350 -1065
rect 4300 -1115 4350 -1085
rect 4300 -1135 4315 -1115
rect 4335 -1135 4350 -1115
rect 4300 -1165 4350 -1135
rect 4300 -1185 4315 -1165
rect 4335 -1185 4350 -1165
rect 4300 -1215 4350 -1185
rect 4300 -1235 4315 -1215
rect 4335 -1235 4350 -1215
rect 4300 -1265 4350 -1235
rect 4300 -1285 4315 -1265
rect 4335 -1285 4350 -1265
rect 4300 -1315 4350 -1285
rect 4300 -1335 4315 -1315
rect 4335 -1335 4350 -1315
rect 4300 -1365 4350 -1335
rect 4300 -1385 4315 -1365
rect 4335 -1385 4350 -1365
rect 4300 -1415 4350 -1385
rect 4300 -1435 4315 -1415
rect 4335 -1435 4350 -1415
rect 4300 -1465 4350 -1435
rect 4300 -1485 4315 -1465
rect 4335 -1485 4350 -1465
rect 4300 -1515 4350 -1485
rect 4300 -1535 4315 -1515
rect 4335 -1535 4350 -1515
rect 4300 -1565 4350 -1535
rect 4300 -1585 4315 -1565
rect 4335 -1585 4350 -1565
rect 4300 -1615 4350 -1585
rect 4300 -1635 4315 -1615
rect 4335 -1635 4350 -1615
rect 4300 -1650 4350 -1635
rect 4450 -965 4500 -950
rect 4450 -985 4465 -965
rect 4485 -985 4500 -965
rect 4450 -1015 4500 -985
rect 4450 -1035 4465 -1015
rect 4485 -1035 4500 -1015
rect 4450 -1065 4500 -1035
rect 4450 -1085 4465 -1065
rect 4485 -1085 4500 -1065
rect 4450 -1115 4500 -1085
rect 4450 -1135 4465 -1115
rect 4485 -1135 4500 -1115
rect 4450 -1165 4500 -1135
rect 4450 -1185 4465 -1165
rect 4485 -1185 4500 -1165
rect 4450 -1215 4500 -1185
rect 4450 -1235 4465 -1215
rect 4485 -1235 4500 -1215
rect 4450 -1265 4500 -1235
rect 4450 -1285 4465 -1265
rect 4485 -1285 4500 -1265
rect 4450 -1315 4500 -1285
rect 4450 -1335 4465 -1315
rect 4485 -1335 4500 -1315
rect 4450 -1365 4500 -1335
rect 4450 -1385 4465 -1365
rect 4485 -1385 4500 -1365
rect 4450 -1415 4500 -1385
rect 4450 -1435 4465 -1415
rect 4485 -1435 4500 -1415
rect 4450 -1465 4500 -1435
rect 4450 -1485 4465 -1465
rect 4485 -1485 4500 -1465
rect 4450 -1515 4500 -1485
rect 4450 -1535 4465 -1515
rect 4485 -1535 4500 -1515
rect 4450 -1565 4500 -1535
rect 4450 -1585 4465 -1565
rect 4485 -1585 4500 -1565
rect 4450 -1615 4500 -1585
rect 4450 -1635 4465 -1615
rect 4485 -1635 4500 -1615
rect 4450 -1650 4500 -1635
rect 4600 -965 4650 -950
rect 4600 -985 4615 -965
rect 4635 -985 4650 -965
rect 4600 -1015 4650 -985
rect 4600 -1035 4615 -1015
rect 4635 -1035 4650 -1015
rect 4600 -1065 4650 -1035
rect 4600 -1085 4615 -1065
rect 4635 -1085 4650 -1065
rect 4600 -1115 4650 -1085
rect 4600 -1135 4615 -1115
rect 4635 -1135 4650 -1115
rect 4600 -1165 4650 -1135
rect 4600 -1185 4615 -1165
rect 4635 -1185 4650 -1165
rect 4600 -1215 4650 -1185
rect 4600 -1235 4615 -1215
rect 4635 -1235 4650 -1215
rect 4600 -1265 4650 -1235
rect 4600 -1285 4615 -1265
rect 4635 -1285 4650 -1265
rect 4600 -1315 4650 -1285
rect 4600 -1335 4615 -1315
rect 4635 -1335 4650 -1315
rect 4600 -1365 4650 -1335
rect 4600 -1385 4615 -1365
rect 4635 -1385 4650 -1365
rect 4600 -1415 4650 -1385
rect 4600 -1435 4615 -1415
rect 4635 -1435 4650 -1415
rect 4600 -1465 4650 -1435
rect 4600 -1485 4615 -1465
rect 4635 -1485 4650 -1465
rect 4600 -1515 4650 -1485
rect 4600 -1535 4615 -1515
rect 4635 -1535 4650 -1515
rect 4600 -1565 4650 -1535
rect 4600 -1585 4615 -1565
rect 4635 -1585 4650 -1565
rect 4600 -1615 4650 -1585
rect 4600 -1635 4615 -1615
rect 4635 -1635 4650 -1615
rect 4600 -1650 4650 -1635
rect 4750 -965 4800 -950
rect 4750 -985 4765 -965
rect 4785 -985 4800 -965
rect 4750 -1015 4800 -985
rect 4750 -1035 4765 -1015
rect 4785 -1035 4800 -1015
rect 4750 -1065 4800 -1035
rect 4750 -1085 4765 -1065
rect 4785 -1085 4800 -1065
rect 4750 -1115 4800 -1085
rect 4750 -1135 4765 -1115
rect 4785 -1135 4800 -1115
rect 4750 -1165 4800 -1135
rect 4750 -1185 4765 -1165
rect 4785 -1185 4800 -1165
rect 4750 -1215 4800 -1185
rect 4750 -1235 4765 -1215
rect 4785 -1235 4800 -1215
rect 4750 -1265 4800 -1235
rect 4750 -1285 4765 -1265
rect 4785 -1285 4800 -1265
rect 4750 -1315 4800 -1285
rect 4750 -1335 4765 -1315
rect 4785 -1335 4800 -1315
rect 4750 -1365 4800 -1335
rect 4750 -1385 4765 -1365
rect 4785 -1385 4800 -1365
rect 4750 -1415 4800 -1385
rect 4750 -1435 4765 -1415
rect 4785 -1435 4800 -1415
rect 4750 -1465 4800 -1435
rect 4750 -1485 4765 -1465
rect 4785 -1485 4800 -1465
rect 4750 -1515 4800 -1485
rect 4750 -1535 4765 -1515
rect 4785 -1535 4800 -1515
rect 4750 -1565 4800 -1535
rect 4750 -1585 4765 -1565
rect 4785 -1585 4800 -1565
rect 4750 -1615 4800 -1585
rect 4750 -1635 4765 -1615
rect 4785 -1635 4800 -1615
rect 4750 -1650 4800 -1635
rect 5050 -965 5100 -950
rect 5050 -985 5065 -965
rect 5085 -985 5100 -965
rect 5050 -1015 5100 -985
rect 5050 -1035 5065 -1015
rect 5085 -1035 5100 -1015
rect 5050 -1065 5100 -1035
rect 5050 -1085 5065 -1065
rect 5085 -1085 5100 -1065
rect 5050 -1115 5100 -1085
rect 5050 -1135 5065 -1115
rect 5085 -1135 5100 -1115
rect 5050 -1165 5100 -1135
rect 5050 -1185 5065 -1165
rect 5085 -1185 5100 -1165
rect 5050 -1215 5100 -1185
rect 5050 -1235 5065 -1215
rect 5085 -1235 5100 -1215
rect 5050 -1265 5100 -1235
rect 5050 -1285 5065 -1265
rect 5085 -1285 5100 -1265
rect 5050 -1315 5100 -1285
rect 5050 -1335 5065 -1315
rect 5085 -1335 5100 -1315
rect 5050 -1365 5100 -1335
rect 5050 -1385 5065 -1365
rect 5085 -1385 5100 -1365
rect 5050 -1415 5100 -1385
rect 5050 -1435 5065 -1415
rect 5085 -1435 5100 -1415
rect 5050 -1465 5100 -1435
rect 5050 -1485 5065 -1465
rect 5085 -1485 5100 -1465
rect 5050 -1515 5100 -1485
rect 5050 -1535 5065 -1515
rect 5085 -1535 5100 -1515
rect 5050 -1565 5100 -1535
rect 5050 -1585 5065 -1565
rect 5085 -1585 5100 -1565
rect 5050 -1615 5100 -1585
rect 5050 -1635 5065 -1615
rect 5085 -1635 5100 -1615
rect 5050 -1650 5100 -1635
rect 5350 -965 5400 -950
rect 5350 -985 5365 -965
rect 5385 -985 5400 -965
rect 5350 -1015 5400 -985
rect 5350 -1035 5365 -1015
rect 5385 -1035 5400 -1015
rect 5350 -1065 5400 -1035
rect 5350 -1085 5365 -1065
rect 5385 -1085 5400 -1065
rect 5350 -1115 5400 -1085
rect 5350 -1135 5365 -1115
rect 5385 -1135 5400 -1115
rect 5350 -1165 5400 -1135
rect 5350 -1185 5365 -1165
rect 5385 -1185 5400 -1165
rect 5350 -1215 5400 -1185
rect 5350 -1235 5365 -1215
rect 5385 -1235 5400 -1215
rect 5350 -1265 5400 -1235
rect 5350 -1285 5365 -1265
rect 5385 -1285 5400 -1265
rect 5350 -1315 5400 -1285
rect 5350 -1335 5365 -1315
rect 5385 -1335 5400 -1315
rect 5350 -1365 5400 -1335
rect 5350 -1385 5365 -1365
rect 5385 -1385 5400 -1365
rect 5350 -1415 5400 -1385
rect 5350 -1435 5365 -1415
rect 5385 -1435 5400 -1415
rect 5350 -1465 5400 -1435
rect 5350 -1485 5365 -1465
rect 5385 -1485 5400 -1465
rect 5350 -1515 5400 -1485
rect 5350 -1535 5365 -1515
rect 5385 -1535 5400 -1515
rect 5350 -1565 5400 -1535
rect 5350 -1585 5365 -1565
rect 5385 -1585 5400 -1565
rect 5350 -1615 5400 -1585
rect 5350 -1635 5365 -1615
rect 5385 -1635 5400 -1615
rect 5350 -1650 5400 -1635
rect 5650 -965 5700 -950
rect 5650 -985 5665 -965
rect 5685 -985 5700 -965
rect 5650 -1015 5700 -985
rect 5650 -1035 5665 -1015
rect 5685 -1035 5700 -1015
rect 5650 -1065 5700 -1035
rect 5650 -1085 5665 -1065
rect 5685 -1085 5700 -1065
rect 5650 -1115 5700 -1085
rect 5650 -1135 5665 -1115
rect 5685 -1135 5700 -1115
rect 5650 -1165 5700 -1135
rect 5650 -1185 5665 -1165
rect 5685 -1185 5700 -1165
rect 5650 -1215 5700 -1185
rect 5650 -1235 5665 -1215
rect 5685 -1235 5700 -1215
rect 5650 -1265 5700 -1235
rect 5650 -1285 5665 -1265
rect 5685 -1285 5700 -1265
rect 5650 -1315 5700 -1285
rect 5650 -1335 5665 -1315
rect 5685 -1335 5700 -1315
rect 5650 -1365 5700 -1335
rect 5650 -1385 5665 -1365
rect 5685 -1385 5700 -1365
rect 5650 -1415 5700 -1385
rect 5650 -1435 5665 -1415
rect 5685 -1435 5700 -1415
rect 5650 -1465 5700 -1435
rect 5650 -1485 5665 -1465
rect 5685 -1485 5700 -1465
rect 5650 -1515 5700 -1485
rect 5650 -1535 5665 -1515
rect 5685 -1535 5700 -1515
rect 5650 -1565 5700 -1535
rect 5650 -1585 5665 -1565
rect 5685 -1585 5700 -1565
rect 5650 -1615 5700 -1585
rect 5650 -1635 5665 -1615
rect 5685 -1635 5700 -1615
rect 5650 -1650 5700 -1635
rect 5950 -965 6000 -950
rect 5950 -985 5965 -965
rect 5985 -985 6000 -965
rect 5950 -1015 6000 -985
rect 5950 -1035 5965 -1015
rect 5985 -1035 6000 -1015
rect 5950 -1065 6000 -1035
rect 5950 -1085 5965 -1065
rect 5985 -1085 6000 -1065
rect 5950 -1115 6000 -1085
rect 5950 -1135 5965 -1115
rect 5985 -1135 6000 -1115
rect 5950 -1165 6000 -1135
rect 5950 -1185 5965 -1165
rect 5985 -1185 6000 -1165
rect 5950 -1215 6000 -1185
rect 5950 -1235 5965 -1215
rect 5985 -1235 6000 -1215
rect 5950 -1265 6000 -1235
rect 5950 -1285 5965 -1265
rect 5985 -1285 6000 -1265
rect 5950 -1315 6000 -1285
rect 5950 -1335 5965 -1315
rect 5985 -1335 6000 -1315
rect 5950 -1365 6000 -1335
rect 5950 -1385 5965 -1365
rect 5985 -1385 6000 -1365
rect 5950 -1415 6000 -1385
rect 5950 -1435 5965 -1415
rect 5985 -1435 6000 -1415
rect 5950 -1465 6000 -1435
rect 5950 -1485 5965 -1465
rect 5985 -1485 6000 -1465
rect 5950 -1515 6000 -1485
rect 5950 -1535 5965 -1515
rect 5985 -1535 6000 -1515
rect 5950 -1565 6000 -1535
rect 5950 -1585 5965 -1565
rect 5985 -1585 6000 -1565
rect 5950 -1615 6000 -1585
rect 5950 -1635 5965 -1615
rect 5985 -1635 6000 -1615
rect 5950 -1650 6000 -1635
rect 6250 -965 6300 -950
rect 6250 -985 6265 -965
rect 6285 -985 6300 -965
rect 6250 -1015 6300 -985
rect 6250 -1035 6265 -1015
rect 6285 -1035 6300 -1015
rect 6250 -1065 6300 -1035
rect 6250 -1085 6265 -1065
rect 6285 -1085 6300 -1065
rect 6250 -1115 6300 -1085
rect 6250 -1135 6265 -1115
rect 6285 -1135 6300 -1115
rect 6250 -1165 6300 -1135
rect 6250 -1185 6265 -1165
rect 6285 -1185 6300 -1165
rect 6250 -1215 6300 -1185
rect 6250 -1235 6265 -1215
rect 6285 -1235 6300 -1215
rect 6250 -1265 6300 -1235
rect 6250 -1285 6265 -1265
rect 6285 -1285 6300 -1265
rect 6250 -1315 6300 -1285
rect 6250 -1335 6265 -1315
rect 6285 -1335 6300 -1315
rect 6250 -1365 6300 -1335
rect 6250 -1385 6265 -1365
rect 6285 -1385 6300 -1365
rect 6250 -1415 6300 -1385
rect 6250 -1435 6265 -1415
rect 6285 -1435 6300 -1415
rect 6250 -1465 6300 -1435
rect 6250 -1485 6265 -1465
rect 6285 -1485 6300 -1465
rect 6250 -1515 6300 -1485
rect 6250 -1535 6265 -1515
rect 6285 -1535 6300 -1515
rect 6250 -1565 6300 -1535
rect 6250 -1585 6265 -1565
rect 6285 -1585 6300 -1565
rect 6250 -1615 6300 -1585
rect 6250 -1635 6265 -1615
rect 6285 -1635 6300 -1615
rect 6250 -1650 6300 -1635
rect 6550 -965 6600 -950
rect 6550 -985 6565 -965
rect 6585 -985 6600 -965
rect 6550 -1015 6600 -985
rect 6550 -1035 6565 -1015
rect 6585 -1035 6600 -1015
rect 6550 -1065 6600 -1035
rect 6550 -1085 6565 -1065
rect 6585 -1085 6600 -1065
rect 6550 -1115 6600 -1085
rect 6550 -1135 6565 -1115
rect 6585 -1135 6600 -1115
rect 6550 -1165 6600 -1135
rect 6550 -1185 6565 -1165
rect 6585 -1185 6600 -1165
rect 6550 -1215 6600 -1185
rect 6550 -1235 6565 -1215
rect 6585 -1235 6600 -1215
rect 6550 -1265 6600 -1235
rect 6550 -1285 6565 -1265
rect 6585 -1285 6600 -1265
rect 6550 -1315 6600 -1285
rect 6550 -1335 6565 -1315
rect 6585 -1335 6600 -1315
rect 6550 -1365 6600 -1335
rect 6550 -1385 6565 -1365
rect 6585 -1385 6600 -1365
rect 6550 -1415 6600 -1385
rect 6550 -1435 6565 -1415
rect 6585 -1435 6600 -1415
rect 6550 -1465 6600 -1435
rect 6550 -1485 6565 -1465
rect 6585 -1485 6600 -1465
rect 6550 -1515 6600 -1485
rect 6550 -1535 6565 -1515
rect 6585 -1535 6600 -1515
rect 6550 -1565 6600 -1535
rect 6550 -1585 6565 -1565
rect 6585 -1585 6600 -1565
rect 6550 -1615 6600 -1585
rect 6550 -1635 6565 -1615
rect 6585 -1635 6600 -1615
rect 6550 -1650 6600 -1635
rect 6850 -965 6900 -950
rect 6850 -985 6865 -965
rect 6885 -985 6900 -965
rect 6850 -1015 6900 -985
rect 6850 -1035 6865 -1015
rect 6885 -1035 6900 -1015
rect 6850 -1065 6900 -1035
rect 6850 -1085 6865 -1065
rect 6885 -1085 6900 -1065
rect 6850 -1115 6900 -1085
rect 6850 -1135 6865 -1115
rect 6885 -1135 6900 -1115
rect 6850 -1165 6900 -1135
rect 6850 -1185 6865 -1165
rect 6885 -1185 6900 -1165
rect 6850 -1215 6900 -1185
rect 6850 -1235 6865 -1215
rect 6885 -1235 6900 -1215
rect 6850 -1265 6900 -1235
rect 6850 -1285 6865 -1265
rect 6885 -1285 6900 -1265
rect 6850 -1315 6900 -1285
rect 6850 -1335 6865 -1315
rect 6885 -1335 6900 -1315
rect 6850 -1365 6900 -1335
rect 6850 -1385 6865 -1365
rect 6885 -1385 6900 -1365
rect 6850 -1415 6900 -1385
rect 6850 -1435 6865 -1415
rect 6885 -1435 6900 -1415
rect 6850 -1465 6900 -1435
rect 6850 -1485 6865 -1465
rect 6885 -1485 6900 -1465
rect 6850 -1515 6900 -1485
rect 6850 -1535 6865 -1515
rect 6885 -1535 6900 -1515
rect 6850 -1565 6900 -1535
rect 6850 -1585 6865 -1565
rect 6885 -1585 6900 -1565
rect 6850 -1615 6900 -1585
rect 6850 -1635 6865 -1615
rect 6885 -1635 6900 -1615
rect 6850 -1650 6900 -1635
rect 7150 -965 7200 -950
rect 7150 -985 7165 -965
rect 7185 -985 7200 -965
rect 7150 -1015 7200 -985
rect 7150 -1035 7165 -1015
rect 7185 -1035 7200 -1015
rect 7150 -1065 7200 -1035
rect 7150 -1085 7165 -1065
rect 7185 -1085 7200 -1065
rect 7150 -1115 7200 -1085
rect 7150 -1135 7165 -1115
rect 7185 -1135 7200 -1115
rect 7150 -1165 7200 -1135
rect 7150 -1185 7165 -1165
rect 7185 -1185 7200 -1165
rect 7150 -1215 7200 -1185
rect 7150 -1235 7165 -1215
rect 7185 -1235 7200 -1215
rect 7150 -1265 7200 -1235
rect 7150 -1285 7165 -1265
rect 7185 -1285 7200 -1265
rect 7150 -1315 7200 -1285
rect 7150 -1335 7165 -1315
rect 7185 -1335 7200 -1315
rect 7150 -1365 7200 -1335
rect 7150 -1385 7165 -1365
rect 7185 -1385 7200 -1365
rect 7150 -1415 7200 -1385
rect 7150 -1435 7165 -1415
rect 7185 -1435 7200 -1415
rect 7150 -1465 7200 -1435
rect 7150 -1485 7165 -1465
rect 7185 -1485 7200 -1465
rect 7150 -1515 7200 -1485
rect 7150 -1535 7165 -1515
rect 7185 -1535 7200 -1515
rect 7150 -1565 7200 -1535
rect 7150 -1585 7165 -1565
rect 7185 -1585 7200 -1565
rect 7150 -1615 7200 -1585
rect 7150 -1635 7165 -1615
rect 7185 -1635 7200 -1615
rect 7150 -1650 7200 -1635
rect 8350 -965 8400 -950
rect 8350 -985 8365 -965
rect 8385 -985 8400 -965
rect 8350 -1015 8400 -985
rect 8350 -1035 8365 -1015
rect 8385 -1035 8400 -1015
rect 8350 -1065 8400 -1035
rect 8350 -1085 8365 -1065
rect 8385 -1085 8400 -1065
rect 8350 -1115 8400 -1085
rect 8350 -1135 8365 -1115
rect 8385 -1135 8400 -1115
rect 8350 -1165 8400 -1135
rect 8350 -1185 8365 -1165
rect 8385 -1185 8400 -1165
rect 8350 -1215 8400 -1185
rect 8350 -1235 8365 -1215
rect 8385 -1235 8400 -1215
rect 8350 -1265 8400 -1235
rect 8350 -1285 8365 -1265
rect 8385 -1285 8400 -1265
rect 8350 -1315 8400 -1285
rect 8350 -1335 8365 -1315
rect 8385 -1335 8400 -1315
rect 8350 -1365 8400 -1335
rect 8350 -1385 8365 -1365
rect 8385 -1385 8400 -1365
rect 8350 -1415 8400 -1385
rect 8350 -1435 8365 -1415
rect 8385 -1435 8400 -1415
rect 8350 -1465 8400 -1435
rect 8350 -1485 8365 -1465
rect 8385 -1485 8400 -1465
rect 8350 -1515 8400 -1485
rect 8350 -1535 8365 -1515
rect 8385 -1535 8400 -1515
rect 8350 -1565 8400 -1535
rect 8350 -1585 8365 -1565
rect 8385 -1585 8400 -1565
rect 8350 -1615 8400 -1585
rect 8350 -1635 8365 -1615
rect 8385 -1635 8400 -1615
rect 8350 -1650 8400 -1635
rect 9550 -965 9600 -950
rect 9550 -985 9565 -965
rect 9585 -985 9600 -965
rect 9550 -1015 9600 -985
rect 9550 -1035 9565 -1015
rect 9585 -1035 9600 -1015
rect 9550 -1065 9600 -1035
rect 9550 -1085 9565 -1065
rect 9585 -1085 9600 -1065
rect 9550 -1115 9600 -1085
rect 9550 -1135 9565 -1115
rect 9585 -1135 9600 -1115
rect 9550 -1165 9600 -1135
rect 9550 -1185 9565 -1165
rect 9585 -1185 9600 -1165
rect 9550 -1215 9600 -1185
rect 9550 -1235 9565 -1215
rect 9585 -1235 9600 -1215
rect 9550 -1265 9600 -1235
rect 9550 -1285 9565 -1265
rect 9585 -1285 9600 -1265
rect 9550 -1315 9600 -1285
rect 9550 -1335 9565 -1315
rect 9585 -1335 9600 -1315
rect 9550 -1365 9600 -1335
rect 9550 -1385 9565 -1365
rect 9585 -1385 9600 -1365
rect 9550 -1415 9600 -1385
rect 9550 -1435 9565 -1415
rect 9585 -1435 9600 -1415
rect 9550 -1465 9600 -1435
rect 9550 -1485 9565 -1465
rect 9585 -1485 9600 -1465
rect 9550 -1515 9600 -1485
rect 9550 -1535 9565 -1515
rect 9585 -1535 9600 -1515
rect 9550 -1565 9600 -1535
rect 9550 -1585 9565 -1565
rect 9585 -1585 9600 -1565
rect 9550 -1615 9600 -1585
rect 9550 -1635 9565 -1615
rect 9585 -1635 9600 -1615
rect 9550 -1650 9600 -1635
rect 10750 -965 10800 -950
rect 10750 -985 10765 -965
rect 10785 -985 10800 -965
rect 10750 -1015 10800 -985
rect 10750 -1035 10765 -1015
rect 10785 -1035 10800 -1015
rect 10750 -1065 10800 -1035
rect 10750 -1085 10765 -1065
rect 10785 -1085 10800 -1065
rect 10750 -1115 10800 -1085
rect 10750 -1135 10765 -1115
rect 10785 -1135 10800 -1115
rect 10750 -1165 10800 -1135
rect 10750 -1185 10765 -1165
rect 10785 -1185 10800 -1165
rect 10750 -1215 10800 -1185
rect 10750 -1235 10765 -1215
rect 10785 -1235 10800 -1215
rect 10750 -1265 10800 -1235
rect 10750 -1285 10765 -1265
rect 10785 -1285 10800 -1265
rect 10750 -1315 10800 -1285
rect 10750 -1335 10765 -1315
rect 10785 -1335 10800 -1315
rect 10750 -1365 10800 -1335
rect 10750 -1385 10765 -1365
rect 10785 -1385 10800 -1365
rect 10750 -1415 10800 -1385
rect 10750 -1435 10765 -1415
rect 10785 -1435 10800 -1415
rect 10750 -1465 10800 -1435
rect 10750 -1485 10765 -1465
rect 10785 -1485 10800 -1465
rect 10750 -1515 10800 -1485
rect 10750 -1535 10765 -1515
rect 10785 -1535 10800 -1515
rect 10750 -1565 10800 -1535
rect 10750 -1585 10765 -1565
rect 10785 -1585 10800 -1565
rect 10750 -1615 10800 -1585
rect 10750 -1635 10765 -1615
rect 10785 -1635 10800 -1615
rect 10750 -1650 10800 -1635
rect 11950 -965 12000 -950
rect 11950 -985 11965 -965
rect 11985 -985 12000 -965
rect 11950 -1015 12000 -985
rect 11950 -1035 11965 -1015
rect 11985 -1035 12000 -1015
rect 11950 -1065 12000 -1035
rect 11950 -1085 11965 -1065
rect 11985 -1085 12000 -1065
rect 11950 -1115 12000 -1085
rect 11950 -1135 11965 -1115
rect 11985 -1135 12000 -1115
rect 11950 -1165 12000 -1135
rect 11950 -1185 11965 -1165
rect 11985 -1185 12000 -1165
rect 11950 -1215 12000 -1185
rect 11950 -1235 11965 -1215
rect 11985 -1235 12000 -1215
rect 11950 -1265 12000 -1235
rect 11950 -1285 11965 -1265
rect 11985 -1285 12000 -1265
rect 11950 -1315 12000 -1285
rect 11950 -1335 11965 -1315
rect 11985 -1335 12000 -1315
rect 11950 -1365 12000 -1335
rect 11950 -1385 11965 -1365
rect 11985 -1385 12000 -1365
rect 11950 -1415 12000 -1385
rect 11950 -1435 11965 -1415
rect 11985 -1435 12000 -1415
rect 11950 -1465 12000 -1435
rect 11950 -1485 11965 -1465
rect 11985 -1485 12000 -1465
rect 11950 -1515 12000 -1485
rect 11950 -1535 11965 -1515
rect 11985 -1535 12000 -1515
rect 11950 -1565 12000 -1535
rect 11950 -1585 11965 -1565
rect 11985 -1585 12000 -1565
rect 11950 -1615 12000 -1585
rect 11950 -1635 11965 -1615
rect 11985 -1635 12000 -1615
rect 11950 -1650 12000 -1635
rect 12250 -965 12300 -950
rect 12250 -985 12265 -965
rect 12285 -985 12300 -965
rect 12250 -1015 12300 -985
rect 12250 -1035 12265 -1015
rect 12285 -1035 12300 -1015
rect 12250 -1065 12300 -1035
rect 12250 -1085 12265 -1065
rect 12285 -1085 12300 -1065
rect 12250 -1115 12300 -1085
rect 12250 -1135 12265 -1115
rect 12285 -1135 12300 -1115
rect 12250 -1165 12300 -1135
rect 12250 -1185 12265 -1165
rect 12285 -1185 12300 -1165
rect 12250 -1215 12300 -1185
rect 12250 -1235 12265 -1215
rect 12285 -1235 12300 -1215
rect 12250 -1265 12300 -1235
rect 12250 -1285 12265 -1265
rect 12285 -1285 12300 -1265
rect 12250 -1315 12300 -1285
rect 12250 -1335 12265 -1315
rect 12285 -1335 12300 -1315
rect 12250 -1365 12300 -1335
rect 12250 -1385 12265 -1365
rect 12285 -1385 12300 -1365
rect 12250 -1415 12300 -1385
rect 12250 -1435 12265 -1415
rect 12285 -1435 12300 -1415
rect 12250 -1465 12300 -1435
rect 12250 -1485 12265 -1465
rect 12285 -1485 12300 -1465
rect 12250 -1515 12300 -1485
rect 12250 -1535 12265 -1515
rect 12285 -1535 12300 -1515
rect 12250 -1565 12300 -1535
rect 12250 -1585 12265 -1565
rect 12285 -1585 12300 -1565
rect 12250 -1615 12300 -1585
rect 12250 -1635 12265 -1615
rect 12285 -1635 12300 -1615
rect 12250 -1650 12300 -1635
rect 12550 -965 12600 -950
rect 12550 -985 12565 -965
rect 12585 -985 12600 -965
rect 12550 -1015 12600 -985
rect 12550 -1035 12565 -1015
rect 12585 -1035 12600 -1015
rect 12550 -1065 12600 -1035
rect 12550 -1085 12565 -1065
rect 12585 -1085 12600 -1065
rect 12550 -1115 12600 -1085
rect 12550 -1135 12565 -1115
rect 12585 -1135 12600 -1115
rect 12550 -1165 12600 -1135
rect 12550 -1185 12565 -1165
rect 12585 -1185 12600 -1165
rect 12550 -1215 12600 -1185
rect 12550 -1235 12565 -1215
rect 12585 -1235 12600 -1215
rect 12550 -1265 12600 -1235
rect 12550 -1285 12565 -1265
rect 12585 -1285 12600 -1265
rect 12550 -1315 12600 -1285
rect 12550 -1335 12565 -1315
rect 12585 -1335 12600 -1315
rect 12550 -1365 12600 -1335
rect 12550 -1385 12565 -1365
rect 12585 -1385 12600 -1365
rect 12550 -1415 12600 -1385
rect 12550 -1435 12565 -1415
rect 12585 -1435 12600 -1415
rect 12550 -1465 12600 -1435
rect 12550 -1485 12565 -1465
rect 12585 -1485 12600 -1465
rect 12550 -1515 12600 -1485
rect 12550 -1535 12565 -1515
rect 12585 -1535 12600 -1515
rect 12550 -1565 12600 -1535
rect 12550 -1585 12565 -1565
rect 12585 -1585 12600 -1565
rect 12550 -1615 12600 -1585
rect 12550 -1635 12565 -1615
rect 12585 -1635 12600 -1615
rect 12550 -1650 12600 -1635
rect 12850 -965 12900 -950
rect 12850 -985 12865 -965
rect 12885 -985 12900 -965
rect 12850 -1015 12900 -985
rect 12850 -1035 12865 -1015
rect 12885 -1035 12900 -1015
rect 12850 -1065 12900 -1035
rect 12850 -1085 12865 -1065
rect 12885 -1085 12900 -1065
rect 12850 -1115 12900 -1085
rect 12850 -1135 12865 -1115
rect 12885 -1135 12900 -1115
rect 12850 -1165 12900 -1135
rect 12850 -1185 12865 -1165
rect 12885 -1185 12900 -1165
rect 12850 -1215 12900 -1185
rect 12850 -1235 12865 -1215
rect 12885 -1235 12900 -1215
rect 12850 -1265 12900 -1235
rect 12850 -1285 12865 -1265
rect 12885 -1285 12900 -1265
rect 12850 -1315 12900 -1285
rect 12850 -1335 12865 -1315
rect 12885 -1335 12900 -1315
rect 12850 -1365 12900 -1335
rect 12850 -1385 12865 -1365
rect 12885 -1385 12900 -1365
rect 12850 -1415 12900 -1385
rect 12850 -1435 12865 -1415
rect 12885 -1435 12900 -1415
rect 12850 -1465 12900 -1435
rect 12850 -1485 12865 -1465
rect 12885 -1485 12900 -1465
rect 12850 -1515 12900 -1485
rect 12850 -1535 12865 -1515
rect 12885 -1535 12900 -1515
rect 12850 -1565 12900 -1535
rect 12850 -1585 12865 -1565
rect 12885 -1585 12900 -1565
rect 12850 -1615 12900 -1585
rect 12850 -1635 12865 -1615
rect 12885 -1635 12900 -1615
rect 12850 -1650 12900 -1635
rect 13150 -965 13200 -950
rect 13150 -985 13165 -965
rect 13185 -985 13200 -965
rect 13150 -1015 13200 -985
rect 13150 -1035 13165 -1015
rect 13185 -1035 13200 -1015
rect 13150 -1065 13200 -1035
rect 13150 -1085 13165 -1065
rect 13185 -1085 13200 -1065
rect 13150 -1115 13200 -1085
rect 13150 -1135 13165 -1115
rect 13185 -1135 13200 -1115
rect 13150 -1165 13200 -1135
rect 13150 -1185 13165 -1165
rect 13185 -1185 13200 -1165
rect 13150 -1215 13200 -1185
rect 13150 -1235 13165 -1215
rect 13185 -1235 13200 -1215
rect 13150 -1265 13200 -1235
rect 13150 -1285 13165 -1265
rect 13185 -1285 13200 -1265
rect 13150 -1315 13200 -1285
rect 13150 -1335 13165 -1315
rect 13185 -1335 13200 -1315
rect 13150 -1365 13200 -1335
rect 13150 -1385 13165 -1365
rect 13185 -1385 13200 -1365
rect 13150 -1415 13200 -1385
rect 13150 -1435 13165 -1415
rect 13185 -1435 13200 -1415
rect 13150 -1465 13200 -1435
rect 13150 -1485 13165 -1465
rect 13185 -1485 13200 -1465
rect 13150 -1515 13200 -1485
rect 13150 -1535 13165 -1515
rect 13185 -1535 13200 -1515
rect 13150 -1565 13200 -1535
rect 13150 -1585 13165 -1565
rect 13185 -1585 13200 -1565
rect 13150 -1615 13200 -1585
rect 13150 -1635 13165 -1615
rect 13185 -1635 13200 -1615
rect 13150 -1650 13200 -1635
rect 13450 -965 13500 -950
rect 13450 -985 13465 -965
rect 13485 -985 13500 -965
rect 13450 -1015 13500 -985
rect 13450 -1035 13465 -1015
rect 13485 -1035 13500 -1015
rect 13450 -1065 13500 -1035
rect 13450 -1085 13465 -1065
rect 13485 -1085 13500 -1065
rect 13450 -1115 13500 -1085
rect 13450 -1135 13465 -1115
rect 13485 -1135 13500 -1115
rect 13450 -1165 13500 -1135
rect 13450 -1185 13465 -1165
rect 13485 -1185 13500 -1165
rect 13450 -1215 13500 -1185
rect 13450 -1235 13465 -1215
rect 13485 -1235 13500 -1215
rect 13450 -1265 13500 -1235
rect 13450 -1285 13465 -1265
rect 13485 -1285 13500 -1265
rect 13450 -1315 13500 -1285
rect 13450 -1335 13465 -1315
rect 13485 -1335 13500 -1315
rect 13450 -1365 13500 -1335
rect 13450 -1385 13465 -1365
rect 13485 -1385 13500 -1365
rect 13450 -1415 13500 -1385
rect 13450 -1435 13465 -1415
rect 13485 -1435 13500 -1415
rect 13450 -1465 13500 -1435
rect 13450 -1485 13465 -1465
rect 13485 -1485 13500 -1465
rect 13450 -1515 13500 -1485
rect 13450 -1535 13465 -1515
rect 13485 -1535 13500 -1515
rect 13450 -1565 13500 -1535
rect 13450 -1585 13465 -1565
rect 13485 -1585 13500 -1565
rect 13450 -1615 13500 -1585
rect 13450 -1635 13465 -1615
rect 13485 -1635 13500 -1615
rect 13450 -1650 13500 -1635
rect 13750 -965 13800 -950
rect 13750 -985 13765 -965
rect 13785 -985 13800 -965
rect 13750 -1015 13800 -985
rect 13750 -1035 13765 -1015
rect 13785 -1035 13800 -1015
rect 13750 -1065 13800 -1035
rect 13750 -1085 13765 -1065
rect 13785 -1085 13800 -1065
rect 13750 -1115 13800 -1085
rect 13750 -1135 13765 -1115
rect 13785 -1135 13800 -1115
rect 13750 -1165 13800 -1135
rect 13750 -1185 13765 -1165
rect 13785 -1185 13800 -1165
rect 13750 -1215 13800 -1185
rect 13750 -1235 13765 -1215
rect 13785 -1235 13800 -1215
rect 13750 -1265 13800 -1235
rect 13750 -1285 13765 -1265
rect 13785 -1285 13800 -1265
rect 13750 -1315 13800 -1285
rect 13750 -1335 13765 -1315
rect 13785 -1335 13800 -1315
rect 13750 -1365 13800 -1335
rect 13750 -1385 13765 -1365
rect 13785 -1385 13800 -1365
rect 13750 -1415 13800 -1385
rect 13750 -1435 13765 -1415
rect 13785 -1435 13800 -1415
rect 13750 -1465 13800 -1435
rect 13750 -1485 13765 -1465
rect 13785 -1485 13800 -1465
rect 13750 -1515 13800 -1485
rect 13750 -1535 13765 -1515
rect 13785 -1535 13800 -1515
rect 13750 -1565 13800 -1535
rect 13750 -1585 13765 -1565
rect 13785 -1585 13800 -1565
rect 13750 -1615 13800 -1585
rect 13750 -1635 13765 -1615
rect 13785 -1635 13800 -1615
rect 13750 -1650 13800 -1635
rect 14050 -965 14100 -950
rect 14050 -985 14065 -965
rect 14085 -985 14100 -965
rect 14050 -1015 14100 -985
rect 14050 -1035 14065 -1015
rect 14085 -1035 14100 -1015
rect 14050 -1065 14100 -1035
rect 14050 -1085 14065 -1065
rect 14085 -1085 14100 -1065
rect 14050 -1115 14100 -1085
rect 14050 -1135 14065 -1115
rect 14085 -1135 14100 -1115
rect 14050 -1165 14100 -1135
rect 14050 -1185 14065 -1165
rect 14085 -1185 14100 -1165
rect 14050 -1215 14100 -1185
rect 14050 -1235 14065 -1215
rect 14085 -1235 14100 -1215
rect 14050 -1265 14100 -1235
rect 14050 -1285 14065 -1265
rect 14085 -1285 14100 -1265
rect 14050 -1315 14100 -1285
rect 14050 -1335 14065 -1315
rect 14085 -1335 14100 -1315
rect 14050 -1365 14100 -1335
rect 14050 -1385 14065 -1365
rect 14085 -1385 14100 -1365
rect 14050 -1415 14100 -1385
rect 14050 -1435 14065 -1415
rect 14085 -1435 14100 -1415
rect 14050 -1465 14100 -1435
rect 14050 -1485 14065 -1465
rect 14085 -1485 14100 -1465
rect 14050 -1515 14100 -1485
rect 14050 -1535 14065 -1515
rect 14085 -1535 14100 -1515
rect 14050 -1565 14100 -1535
rect 14050 -1585 14065 -1565
rect 14085 -1585 14100 -1565
rect 14050 -1615 14100 -1585
rect 14050 -1635 14065 -1615
rect 14085 -1635 14100 -1615
rect 14050 -1650 14100 -1635
rect 14350 -965 14400 -950
rect 14350 -985 14365 -965
rect 14385 -985 14400 -965
rect 14350 -1015 14400 -985
rect 14350 -1035 14365 -1015
rect 14385 -1035 14400 -1015
rect 14350 -1065 14400 -1035
rect 14350 -1085 14365 -1065
rect 14385 -1085 14400 -1065
rect 14350 -1115 14400 -1085
rect 14350 -1135 14365 -1115
rect 14385 -1135 14400 -1115
rect 14350 -1165 14400 -1135
rect 14350 -1185 14365 -1165
rect 14385 -1185 14400 -1165
rect 14350 -1215 14400 -1185
rect 14350 -1235 14365 -1215
rect 14385 -1235 14400 -1215
rect 14350 -1265 14400 -1235
rect 14350 -1285 14365 -1265
rect 14385 -1285 14400 -1265
rect 14350 -1315 14400 -1285
rect 14350 -1335 14365 -1315
rect 14385 -1335 14400 -1315
rect 14350 -1365 14400 -1335
rect 14350 -1385 14365 -1365
rect 14385 -1385 14400 -1365
rect 14350 -1415 14400 -1385
rect 14350 -1435 14365 -1415
rect 14385 -1435 14400 -1415
rect 14350 -1465 14400 -1435
rect 14350 -1485 14365 -1465
rect 14385 -1485 14400 -1465
rect 14350 -1515 14400 -1485
rect 14350 -1535 14365 -1515
rect 14385 -1535 14400 -1515
rect 14350 -1565 14400 -1535
rect 14350 -1585 14365 -1565
rect 14385 -1585 14400 -1565
rect 14350 -1615 14400 -1585
rect 14350 -1635 14365 -1615
rect 14385 -1635 14400 -1615
rect 14350 -1650 14400 -1635
rect 15550 -965 15600 -950
rect 15550 -985 15565 -965
rect 15585 -985 15600 -965
rect 15550 -1015 15600 -985
rect 15550 -1035 15565 -1015
rect 15585 -1035 15600 -1015
rect 15550 -1065 15600 -1035
rect 15550 -1085 15565 -1065
rect 15585 -1085 15600 -1065
rect 15550 -1115 15600 -1085
rect 15550 -1135 15565 -1115
rect 15585 -1135 15600 -1115
rect 15550 -1165 15600 -1135
rect 15550 -1185 15565 -1165
rect 15585 -1185 15600 -1165
rect 15550 -1215 15600 -1185
rect 15550 -1235 15565 -1215
rect 15585 -1235 15600 -1215
rect 15550 -1265 15600 -1235
rect 15550 -1285 15565 -1265
rect 15585 -1285 15600 -1265
rect 15550 -1315 15600 -1285
rect 15550 -1335 15565 -1315
rect 15585 -1335 15600 -1315
rect 15550 -1365 15600 -1335
rect 15550 -1385 15565 -1365
rect 15585 -1385 15600 -1365
rect 15550 -1415 15600 -1385
rect 15550 -1435 15565 -1415
rect 15585 -1435 15600 -1415
rect 15550 -1465 15600 -1435
rect 15550 -1485 15565 -1465
rect 15585 -1485 15600 -1465
rect 15550 -1515 15600 -1485
rect 15550 -1535 15565 -1515
rect 15585 -1535 15600 -1515
rect 15550 -1565 15600 -1535
rect 15550 -1585 15565 -1565
rect 15585 -1585 15600 -1565
rect 15550 -1615 15600 -1585
rect 15550 -1635 15565 -1615
rect 15585 -1635 15600 -1615
rect 15550 -1650 15600 -1635
rect 16750 -965 16800 -950
rect 16750 -985 16765 -965
rect 16785 -985 16800 -965
rect 16750 -1015 16800 -985
rect 16750 -1035 16765 -1015
rect 16785 -1035 16800 -1015
rect 16750 -1065 16800 -1035
rect 16750 -1085 16765 -1065
rect 16785 -1085 16800 -1065
rect 16750 -1115 16800 -1085
rect 16750 -1135 16765 -1115
rect 16785 -1135 16800 -1115
rect 16750 -1165 16800 -1135
rect 16750 -1185 16765 -1165
rect 16785 -1185 16800 -1165
rect 16750 -1215 16800 -1185
rect 16750 -1235 16765 -1215
rect 16785 -1235 16800 -1215
rect 16750 -1265 16800 -1235
rect 16750 -1285 16765 -1265
rect 16785 -1285 16800 -1265
rect 16750 -1315 16800 -1285
rect 16750 -1335 16765 -1315
rect 16785 -1335 16800 -1315
rect 16750 -1365 16800 -1335
rect 16750 -1385 16765 -1365
rect 16785 -1385 16800 -1365
rect 16750 -1415 16800 -1385
rect 16750 -1435 16765 -1415
rect 16785 -1435 16800 -1415
rect 16750 -1465 16800 -1435
rect 16750 -1485 16765 -1465
rect 16785 -1485 16800 -1465
rect 16750 -1515 16800 -1485
rect 16750 -1535 16765 -1515
rect 16785 -1535 16800 -1515
rect 16750 -1565 16800 -1535
rect 16750 -1585 16765 -1565
rect 16785 -1585 16800 -1565
rect 16750 -1615 16800 -1585
rect 16750 -1635 16765 -1615
rect 16785 -1635 16800 -1615
rect 16750 -1650 16800 -1635
rect 17950 -965 18000 -950
rect 17950 -985 17965 -965
rect 17985 -985 18000 -965
rect 17950 -1015 18000 -985
rect 17950 -1035 17965 -1015
rect 17985 -1035 18000 -1015
rect 17950 -1065 18000 -1035
rect 17950 -1085 17965 -1065
rect 17985 -1085 18000 -1065
rect 17950 -1115 18000 -1085
rect 17950 -1135 17965 -1115
rect 17985 -1135 18000 -1115
rect 17950 -1165 18000 -1135
rect 17950 -1185 17965 -1165
rect 17985 -1185 18000 -1165
rect 17950 -1215 18000 -1185
rect 17950 -1235 17965 -1215
rect 17985 -1235 18000 -1215
rect 17950 -1265 18000 -1235
rect 17950 -1285 17965 -1265
rect 17985 -1285 18000 -1265
rect 17950 -1315 18000 -1285
rect 17950 -1335 17965 -1315
rect 17985 -1335 18000 -1315
rect 17950 -1365 18000 -1335
rect 17950 -1385 17965 -1365
rect 17985 -1385 18000 -1365
rect 17950 -1415 18000 -1385
rect 17950 -1435 17965 -1415
rect 17985 -1435 18000 -1415
rect 17950 -1465 18000 -1435
rect 17950 -1485 17965 -1465
rect 17985 -1485 18000 -1465
rect 17950 -1515 18000 -1485
rect 17950 -1535 17965 -1515
rect 17985 -1535 18000 -1515
rect 17950 -1565 18000 -1535
rect 17950 -1585 17965 -1565
rect 17985 -1585 18000 -1565
rect 17950 -1615 18000 -1585
rect 17950 -1635 17965 -1615
rect 17985 -1635 18000 -1615
rect 17950 -1650 18000 -1635
rect 19150 -965 19200 -950
rect 19150 -985 19165 -965
rect 19185 -985 19200 -965
rect 19150 -1015 19200 -985
rect 19150 -1035 19165 -1015
rect 19185 -1035 19200 -1015
rect 19150 -1065 19200 -1035
rect 19150 -1085 19165 -1065
rect 19185 -1085 19200 -1065
rect 19150 -1115 19200 -1085
rect 19150 -1135 19165 -1115
rect 19185 -1135 19200 -1115
rect 19150 -1165 19200 -1135
rect 19150 -1185 19165 -1165
rect 19185 -1185 19200 -1165
rect 19150 -1215 19200 -1185
rect 19150 -1235 19165 -1215
rect 19185 -1235 19200 -1215
rect 19150 -1265 19200 -1235
rect 19150 -1285 19165 -1265
rect 19185 -1285 19200 -1265
rect 19150 -1315 19200 -1285
rect 19150 -1335 19165 -1315
rect 19185 -1335 19200 -1315
rect 19150 -1365 19200 -1335
rect 19150 -1385 19165 -1365
rect 19185 -1385 19200 -1365
rect 19150 -1415 19200 -1385
rect 19150 -1435 19165 -1415
rect 19185 -1435 19200 -1415
rect 19150 -1465 19200 -1435
rect 19150 -1485 19165 -1465
rect 19185 -1485 19200 -1465
rect 19150 -1515 19200 -1485
rect 19150 -1535 19165 -1515
rect 19185 -1535 19200 -1515
rect 19150 -1565 19200 -1535
rect 19150 -1585 19165 -1565
rect 19185 -1585 19200 -1565
rect 19150 -1615 19200 -1585
rect 19150 -1635 19165 -1615
rect 19185 -1635 19200 -1615
rect 19150 -1650 19200 -1635
rect 20350 -965 20400 -950
rect 20350 -985 20365 -965
rect 20385 -985 20400 -965
rect 20350 -1015 20400 -985
rect 20350 -1035 20365 -1015
rect 20385 -1035 20400 -1015
rect 20350 -1065 20400 -1035
rect 20350 -1085 20365 -1065
rect 20385 -1085 20400 -1065
rect 20350 -1115 20400 -1085
rect 20350 -1135 20365 -1115
rect 20385 -1135 20400 -1115
rect 20350 -1165 20400 -1135
rect 20350 -1185 20365 -1165
rect 20385 -1185 20400 -1165
rect 20350 -1215 20400 -1185
rect 20350 -1235 20365 -1215
rect 20385 -1235 20400 -1215
rect 20350 -1265 20400 -1235
rect 20350 -1285 20365 -1265
rect 20385 -1285 20400 -1265
rect 20350 -1315 20400 -1285
rect 20350 -1335 20365 -1315
rect 20385 -1335 20400 -1315
rect 20350 -1365 20400 -1335
rect 20350 -1385 20365 -1365
rect 20385 -1385 20400 -1365
rect 20350 -1415 20400 -1385
rect 20350 -1435 20365 -1415
rect 20385 -1435 20400 -1415
rect 20350 -1465 20400 -1435
rect 20350 -1485 20365 -1465
rect 20385 -1485 20400 -1465
rect 20350 -1515 20400 -1485
rect 20350 -1535 20365 -1515
rect 20385 -1535 20400 -1515
rect 20350 -1565 20400 -1535
rect 20350 -1585 20365 -1565
rect 20385 -1585 20400 -1565
rect 20350 -1615 20400 -1585
rect 20350 -1635 20365 -1615
rect 20385 -1635 20400 -1615
rect 20350 -1650 20400 -1635
rect 21550 -965 21600 -950
rect 21550 -985 21565 -965
rect 21585 -985 21600 -965
rect 21550 -1015 21600 -985
rect 21550 -1035 21565 -1015
rect 21585 -1035 21600 -1015
rect 21550 -1065 21600 -1035
rect 21550 -1085 21565 -1065
rect 21585 -1085 21600 -1065
rect 21550 -1115 21600 -1085
rect 21550 -1135 21565 -1115
rect 21585 -1135 21600 -1115
rect 21550 -1165 21600 -1135
rect 21550 -1185 21565 -1165
rect 21585 -1185 21600 -1165
rect 21550 -1215 21600 -1185
rect 21550 -1235 21565 -1215
rect 21585 -1235 21600 -1215
rect 21550 -1265 21600 -1235
rect 21550 -1285 21565 -1265
rect 21585 -1285 21600 -1265
rect 21550 -1315 21600 -1285
rect 21550 -1335 21565 -1315
rect 21585 -1335 21600 -1315
rect 21550 -1365 21600 -1335
rect 21550 -1385 21565 -1365
rect 21585 -1385 21600 -1365
rect 21550 -1415 21600 -1385
rect 21550 -1435 21565 -1415
rect 21585 -1435 21600 -1415
rect 21550 -1465 21600 -1435
rect 21550 -1485 21565 -1465
rect 21585 -1485 21600 -1465
rect 21550 -1515 21600 -1485
rect 21550 -1535 21565 -1515
rect 21585 -1535 21600 -1515
rect 21550 -1565 21600 -1535
rect 21550 -1585 21565 -1565
rect 21585 -1585 21600 -1565
rect 21550 -1615 21600 -1585
rect 21550 -1635 21565 -1615
rect 21585 -1635 21600 -1615
rect 21550 -1650 21600 -1635
rect 22450 -965 22500 -950
rect 22450 -985 22465 -965
rect 22485 -985 22500 -965
rect 22450 -1015 22500 -985
rect 22450 -1035 22465 -1015
rect 22485 -1035 22500 -1015
rect 22450 -1065 22500 -1035
rect 22450 -1085 22465 -1065
rect 22485 -1085 22500 -1065
rect 22450 -1115 22500 -1085
rect 22450 -1135 22465 -1115
rect 22485 -1135 22500 -1115
rect 22450 -1165 22500 -1135
rect 22450 -1185 22465 -1165
rect 22485 -1185 22500 -1165
rect 22450 -1215 22500 -1185
rect 22450 -1235 22465 -1215
rect 22485 -1235 22500 -1215
rect 22450 -1265 22500 -1235
rect 22450 -1285 22465 -1265
rect 22485 -1285 22500 -1265
rect 22450 -1315 22500 -1285
rect 22450 -1335 22465 -1315
rect 22485 -1335 22500 -1315
rect 22450 -1365 22500 -1335
rect 22450 -1385 22465 -1365
rect 22485 -1385 22500 -1365
rect 22450 -1415 22500 -1385
rect 22450 -1435 22465 -1415
rect 22485 -1435 22500 -1415
rect 22450 -1465 22500 -1435
rect 22450 -1485 22465 -1465
rect 22485 -1485 22500 -1465
rect 22450 -1515 22500 -1485
rect 22450 -1535 22465 -1515
rect 22485 -1535 22500 -1515
rect 22450 -1565 22500 -1535
rect 22450 -1585 22465 -1565
rect 22485 -1585 22500 -1565
rect 22450 -1615 22500 -1585
rect 22450 -1635 22465 -1615
rect 22485 -1635 22500 -1615
rect 22450 -1650 22500 -1635
rect 23350 -965 23400 -950
rect 23350 -985 23365 -965
rect 23385 -985 23400 -965
rect 23350 -1015 23400 -985
rect 23350 -1035 23365 -1015
rect 23385 -1035 23400 -1015
rect 23350 -1065 23400 -1035
rect 23350 -1085 23365 -1065
rect 23385 -1085 23400 -1065
rect 23350 -1115 23400 -1085
rect 23350 -1135 23365 -1115
rect 23385 -1135 23400 -1115
rect 23350 -1165 23400 -1135
rect 23350 -1185 23365 -1165
rect 23385 -1185 23400 -1165
rect 23350 -1215 23400 -1185
rect 23350 -1235 23365 -1215
rect 23385 -1235 23400 -1215
rect 23350 -1265 23400 -1235
rect 23350 -1285 23365 -1265
rect 23385 -1285 23400 -1265
rect 23350 -1315 23400 -1285
rect 23350 -1335 23365 -1315
rect 23385 -1335 23400 -1315
rect 23350 -1365 23400 -1335
rect 23350 -1385 23365 -1365
rect 23385 -1385 23400 -1365
rect 23350 -1415 23400 -1385
rect 23350 -1435 23365 -1415
rect 23385 -1435 23400 -1415
rect 23350 -1465 23400 -1435
rect 23350 -1485 23365 -1465
rect 23385 -1485 23400 -1465
rect 23350 -1515 23400 -1485
rect 23350 -1535 23365 -1515
rect 23385 -1535 23400 -1515
rect 23350 -1565 23400 -1535
rect 23350 -1585 23365 -1565
rect 23385 -1585 23400 -1565
rect 23350 -1615 23400 -1585
rect 23350 -1635 23365 -1615
rect 23385 -1635 23400 -1615
rect 23350 -1650 23400 -1635
rect 24550 -965 24600 -950
rect 24550 -985 24565 -965
rect 24585 -985 24600 -965
rect 24550 -1015 24600 -985
rect 24550 -1035 24565 -1015
rect 24585 -1035 24600 -1015
rect 24550 -1065 24600 -1035
rect 24550 -1085 24565 -1065
rect 24585 -1085 24600 -1065
rect 24550 -1115 24600 -1085
rect 24550 -1135 24565 -1115
rect 24585 -1135 24600 -1115
rect 24550 -1165 24600 -1135
rect 24550 -1185 24565 -1165
rect 24585 -1185 24600 -1165
rect 24550 -1215 24600 -1185
rect 24550 -1235 24565 -1215
rect 24585 -1235 24600 -1215
rect 24550 -1265 24600 -1235
rect 24550 -1285 24565 -1265
rect 24585 -1285 24600 -1265
rect 24550 -1315 24600 -1285
rect 24550 -1335 24565 -1315
rect 24585 -1335 24600 -1315
rect 24550 -1365 24600 -1335
rect 24550 -1385 24565 -1365
rect 24585 -1385 24600 -1365
rect 24550 -1415 24600 -1385
rect 24550 -1435 24565 -1415
rect 24585 -1435 24600 -1415
rect 24550 -1465 24600 -1435
rect 24550 -1485 24565 -1465
rect 24585 -1485 24600 -1465
rect 24550 -1515 24600 -1485
rect 24550 -1535 24565 -1515
rect 24585 -1535 24600 -1515
rect 24550 -1565 24600 -1535
rect 24550 -1585 24565 -1565
rect 24585 -1585 24600 -1565
rect 24550 -1615 24600 -1585
rect 24550 -1635 24565 -1615
rect 24585 -1635 24600 -1615
rect 24550 -1650 24600 -1635
rect 25750 -965 25800 -950
rect 25750 -985 25765 -965
rect 25785 -985 25800 -965
rect 25750 -1015 25800 -985
rect 25750 -1035 25765 -1015
rect 25785 -1035 25800 -1015
rect 25750 -1065 25800 -1035
rect 25750 -1085 25765 -1065
rect 25785 -1085 25800 -1065
rect 25750 -1115 25800 -1085
rect 25750 -1135 25765 -1115
rect 25785 -1135 25800 -1115
rect 25750 -1165 25800 -1135
rect 25750 -1185 25765 -1165
rect 25785 -1185 25800 -1165
rect 25750 -1215 25800 -1185
rect 25750 -1235 25765 -1215
rect 25785 -1235 25800 -1215
rect 25750 -1265 25800 -1235
rect 25750 -1285 25765 -1265
rect 25785 -1285 25800 -1265
rect 25750 -1315 25800 -1285
rect 25750 -1335 25765 -1315
rect 25785 -1335 25800 -1315
rect 25750 -1365 25800 -1335
rect 25750 -1385 25765 -1365
rect 25785 -1385 25800 -1365
rect 25750 -1415 25800 -1385
rect 25750 -1435 25765 -1415
rect 25785 -1435 25800 -1415
rect 25750 -1465 25800 -1435
rect 25750 -1485 25765 -1465
rect 25785 -1485 25800 -1465
rect 25750 -1515 25800 -1485
rect 25750 -1535 25765 -1515
rect 25785 -1535 25800 -1515
rect 25750 -1565 25800 -1535
rect 25750 -1585 25765 -1565
rect 25785 -1585 25800 -1565
rect 25750 -1615 25800 -1585
rect 25750 -1635 25765 -1615
rect 25785 -1635 25800 -1615
rect 25750 -1650 25800 -1635
rect 26650 -965 26700 -950
rect 26650 -985 26665 -965
rect 26685 -985 26700 -965
rect 26650 -1015 26700 -985
rect 26650 -1035 26665 -1015
rect 26685 -1035 26700 -1015
rect 26650 -1065 26700 -1035
rect 26650 -1085 26665 -1065
rect 26685 -1085 26700 -1065
rect 26650 -1115 26700 -1085
rect 26650 -1135 26665 -1115
rect 26685 -1135 26700 -1115
rect 26650 -1165 26700 -1135
rect 26650 -1185 26665 -1165
rect 26685 -1185 26700 -1165
rect 26650 -1215 26700 -1185
rect 26650 -1235 26665 -1215
rect 26685 -1235 26700 -1215
rect 26650 -1265 26700 -1235
rect 26650 -1285 26665 -1265
rect 26685 -1285 26700 -1265
rect 26650 -1315 26700 -1285
rect 26650 -1335 26665 -1315
rect 26685 -1335 26700 -1315
rect 26650 -1365 26700 -1335
rect 26650 -1385 26665 -1365
rect 26685 -1385 26700 -1365
rect 26650 -1415 26700 -1385
rect 26650 -1435 26665 -1415
rect 26685 -1435 26700 -1415
rect 26650 -1465 26700 -1435
rect 26650 -1485 26665 -1465
rect 26685 -1485 26700 -1465
rect 26650 -1515 26700 -1485
rect 26650 -1535 26665 -1515
rect 26685 -1535 26700 -1515
rect 26650 -1565 26700 -1535
rect 26650 -1585 26665 -1565
rect 26685 -1585 26700 -1565
rect 26650 -1615 26700 -1585
rect 26650 -1635 26665 -1615
rect 26685 -1635 26700 -1615
rect 26650 -1650 26700 -1635
rect 27550 -965 27600 -950
rect 27550 -985 27565 -965
rect 27585 -985 27600 -965
rect 27550 -1015 27600 -985
rect 27550 -1035 27565 -1015
rect 27585 -1035 27600 -1015
rect 27550 -1065 27600 -1035
rect 27550 -1085 27565 -1065
rect 27585 -1085 27600 -1065
rect 27550 -1115 27600 -1085
rect 27550 -1135 27565 -1115
rect 27585 -1135 27600 -1115
rect 27550 -1165 27600 -1135
rect 27550 -1185 27565 -1165
rect 27585 -1185 27600 -1165
rect 27550 -1215 27600 -1185
rect 27550 -1235 27565 -1215
rect 27585 -1235 27600 -1215
rect 27550 -1265 27600 -1235
rect 27550 -1285 27565 -1265
rect 27585 -1285 27600 -1265
rect 27550 -1315 27600 -1285
rect 27550 -1335 27565 -1315
rect 27585 -1335 27600 -1315
rect 27550 -1365 27600 -1335
rect 27550 -1385 27565 -1365
rect 27585 -1385 27600 -1365
rect 27550 -1415 27600 -1385
rect 27550 -1435 27565 -1415
rect 27585 -1435 27600 -1415
rect 27550 -1465 27600 -1435
rect 27550 -1485 27565 -1465
rect 27585 -1485 27600 -1465
rect 27550 -1515 27600 -1485
rect 27550 -1535 27565 -1515
rect 27585 -1535 27600 -1515
rect 27550 -1565 27600 -1535
rect 27550 -1585 27565 -1565
rect 27585 -1585 27600 -1565
rect 27550 -1615 27600 -1585
rect 27550 -1635 27565 -1615
rect 27585 -1635 27600 -1615
rect 27550 -1650 27600 -1635
rect 28750 -965 28800 -950
rect 28750 -985 28765 -965
rect 28785 -985 28800 -965
rect 28750 -1015 28800 -985
rect 28750 -1035 28765 -1015
rect 28785 -1035 28800 -1015
rect 28750 -1065 28800 -1035
rect 28750 -1085 28765 -1065
rect 28785 -1085 28800 -1065
rect 28750 -1115 28800 -1085
rect 28750 -1135 28765 -1115
rect 28785 -1135 28800 -1115
rect 28750 -1165 28800 -1135
rect 28750 -1185 28765 -1165
rect 28785 -1185 28800 -1165
rect 28750 -1215 28800 -1185
rect 28750 -1235 28765 -1215
rect 28785 -1235 28800 -1215
rect 28750 -1265 28800 -1235
rect 28750 -1285 28765 -1265
rect 28785 -1285 28800 -1265
rect 28750 -1315 28800 -1285
rect 28750 -1335 28765 -1315
rect 28785 -1335 28800 -1315
rect 28750 -1365 28800 -1335
rect 28750 -1385 28765 -1365
rect 28785 -1385 28800 -1365
rect 28750 -1415 28800 -1385
rect 28750 -1435 28765 -1415
rect 28785 -1435 28800 -1415
rect 28750 -1465 28800 -1435
rect 28750 -1485 28765 -1465
rect 28785 -1485 28800 -1465
rect 28750 -1515 28800 -1485
rect 28750 -1535 28765 -1515
rect 28785 -1535 28800 -1515
rect 28750 -1565 28800 -1535
rect 28750 -1585 28765 -1565
rect 28785 -1585 28800 -1565
rect 28750 -1615 28800 -1585
rect 28750 -1635 28765 -1615
rect 28785 -1635 28800 -1615
rect 28750 -1650 28800 -1635
rect -650 -1715 28800 -1700
rect -650 -1735 -635 -1715
rect -615 -1735 -585 -1715
rect -565 -1735 -535 -1715
rect -515 -1735 -485 -1715
rect -465 -1735 -435 -1715
rect -415 -1735 -385 -1715
rect -365 -1735 -335 -1715
rect -315 -1735 -285 -1715
rect -265 -1735 -235 -1715
rect -215 -1735 -185 -1715
rect -165 -1735 -135 -1715
rect -115 -1735 -85 -1715
rect -65 -1735 -35 -1715
rect -15 -1735 15 -1715
rect 35 -1735 65 -1715
rect 85 -1735 115 -1715
rect 135 -1735 165 -1715
rect 185 -1735 215 -1715
rect 235 -1735 265 -1715
rect 285 -1735 315 -1715
rect 335 -1735 365 -1715
rect 385 -1735 415 -1715
rect 435 -1735 465 -1715
rect 485 -1735 515 -1715
rect 535 -1735 565 -1715
rect 585 -1735 615 -1715
rect 635 -1735 665 -1715
rect 685 -1735 715 -1715
rect 735 -1735 765 -1715
rect 785 -1735 815 -1715
rect 835 -1735 865 -1715
rect 885 -1735 915 -1715
rect 935 -1735 965 -1715
rect 985 -1735 1015 -1715
rect 1035 -1735 1065 -1715
rect 1085 -1735 1115 -1715
rect 1135 -1735 1165 -1715
rect 1185 -1735 1215 -1715
rect 1235 -1735 1265 -1715
rect 1285 -1735 1315 -1715
rect 1335 -1735 1365 -1715
rect 1385 -1735 1415 -1715
rect 1435 -1735 1465 -1715
rect 1485 -1735 1515 -1715
rect 1535 -1735 1565 -1715
rect 1585 -1735 1615 -1715
rect 1635 -1735 1665 -1715
rect 1685 -1735 1715 -1715
rect 1735 -1735 1765 -1715
rect 1785 -1735 1815 -1715
rect 1835 -1735 1865 -1715
rect 1885 -1735 1915 -1715
rect 1935 -1735 1965 -1715
rect 1985 -1735 2015 -1715
rect 2035 -1735 2065 -1715
rect 2085 -1735 2115 -1715
rect 2135 -1735 2165 -1715
rect 2185 -1735 2215 -1715
rect 2235 -1735 2265 -1715
rect 2285 -1735 2315 -1715
rect 2335 -1735 2365 -1715
rect 2385 -1735 2415 -1715
rect 2435 -1735 2465 -1715
rect 2485 -1735 2515 -1715
rect 2535 -1735 2565 -1715
rect 2585 -1735 2615 -1715
rect 2635 -1735 2665 -1715
rect 2685 -1735 2715 -1715
rect 2735 -1735 2765 -1715
rect 2785 -1735 2815 -1715
rect 2835 -1735 2865 -1715
rect 2885 -1735 2915 -1715
rect 2935 -1735 2965 -1715
rect 2985 -1735 3015 -1715
rect 3035 -1735 3065 -1715
rect 3085 -1735 3115 -1715
rect 3135 -1735 3165 -1715
rect 3185 -1735 3215 -1715
rect 3235 -1735 3265 -1715
rect 3285 -1735 3315 -1715
rect 3335 -1735 3365 -1715
rect 3385 -1735 3415 -1715
rect 3435 -1735 3465 -1715
rect 3485 -1735 3515 -1715
rect 3535 -1735 3565 -1715
rect 3585 -1735 3615 -1715
rect 3635 -1735 3665 -1715
rect 3685 -1735 3715 -1715
rect 3735 -1735 3765 -1715
rect 3785 -1735 3815 -1715
rect 3835 -1735 3865 -1715
rect 3885 -1735 3915 -1715
rect 3935 -1735 3965 -1715
rect 3985 -1735 4015 -1715
rect 4035 -1735 4065 -1715
rect 4085 -1735 4115 -1715
rect 4135 -1735 4165 -1715
rect 4185 -1735 4215 -1715
rect 4235 -1735 4265 -1715
rect 4285 -1735 4315 -1715
rect 4335 -1735 4365 -1715
rect 4385 -1735 4415 -1715
rect 4435 -1735 4465 -1715
rect 4485 -1735 4515 -1715
rect 4535 -1735 4565 -1715
rect 4585 -1735 4615 -1715
rect 4635 -1735 4665 -1715
rect 4685 -1735 4715 -1715
rect 4735 -1735 4765 -1715
rect 4785 -1735 4815 -1715
rect 4835 -1735 4865 -1715
rect 4885 -1735 4915 -1715
rect 4935 -1735 4965 -1715
rect 4985 -1735 5015 -1715
rect 5035 -1735 5065 -1715
rect 5085 -1735 5115 -1715
rect 5135 -1735 5165 -1715
rect 5185 -1735 5215 -1715
rect 5235 -1735 5265 -1715
rect 5285 -1735 5315 -1715
rect 5335 -1735 5365 -1715
rect 5385 -1735 5415 -1715
rect 5435 -1735 5465 -1715
rect 5485 -1735 5515 -1715
rect 5535 -1735 5565 -1715
rect 5585 -1735 5615 -1715
rect 5635 -1735 5665 -1715
rect 5685 -1735 5715 -1715
rect 5735 -1735 5765 -1715
rect 5785 -1735 5815 -1715
rect 5835 -1735 5865 -1715
rect 5885 -1735 5915 -1715
rect 5935 -1735 5965 -1715
rect 5985 -1735 6015 -1715
rect 6035 -1735 6065 -1715
rect 6085 -1735 6115 -1715
rect 6135 -1735 6165 -1715
rect 6185 -1735 6215 -1715
rect 6235 -1735 6265 -1715
rect 6285 -1735 6315 -1715
rect 6335 -1735 6365 -1715
rect 6385 -1735 6415 -1715
rect 6435 -1735 6465 -1715
rect 6485 -1735 6515 -1715
rect 6535 -1735 6565 -1715
rect 6585 -1735 6615 -1715
rect 6635 -1735 6665 -1715
rect 6685 -1735 6715 -1715
rect 6735 -1735 6765 -1715
rect 6785 -1735 6815 -1715
rect 6835 -1735 6865 -1715
rect 6885 -1735 6915 -1715
rect 6935 -1735 6965 -1715
rect 6985 -1735 7015 -1715
rect 7035 -1735 7065 -1715
rect 7085 -1735 7115 -1715
rect 7135 -1735 7165 -1715
rect 7185 -1735 7215 -1715
rect 7235 -1735 7265 -1715
rect 7285 -1735 7315 -1715
rect 7335 -1735 7365 -1715
rect 7385 -1735 7415 -1715
rect 7435 -1735 7465 -1715
rect 7485 -1735 7515 -1715
rect 7535 -1735 7565 -1715
rect 7585 -1735 7615 -1715
rect 7635 -1735 7665 -1715
rect 7685 -1735 7715 -1715
rect 7735 -1735 7765 -1715
rect 7785 -1735 7815 -1715
rect 7835 -1735 7865 -1715
rect 7885 -1735 7915 -1715
rect 7935 -1735 7965 -1715
rect 7985 -1735 8015 -1715
rect 8035 -1735 8065 -1715
rect 8085 -1735 8115 -1715
rect 8135 -1735 8165 -1715
rect 8185 -1735 8215 -1715
rect 8235 -1735 8265 -1715
rect 8285 -1735 8315 -1715
rect 8335 -1735 8365 -1715
rect 8385 -1735 8415 -1715
rect 8435 -1735 8465 -1715
rect 8485 -1735 8515 -1715
rect 8535 -1735 8565 -1715
rect 8585 -1735 8615 -1715
rect 8635 -1735 8665 -1715
rect 8685 -1735 8715 -1715
rect 8735 -1735 8765 -1715
rect 8785 -1735 8815 -1715
rect 8835 -1735 8865 -1715
rect 8885 -1735 8915 -1715
rect 8935 -1735 8965 -1715
rect 8985 -1735 9015 -1715
rect 9035 -1735 9065 -1715
rect 9085 -1735 9115 -1715
rect 9135 -1735 9165 -1715
rect 9185 -1735 9215 -1715
rect 9235 -1735 9265 -1715
rect 9285 -1735 9315 -1715
rect 9335 -1735 9365 -1715
rect 9385 -1735 9415 -1715
rect 9435 -1735 9465 -1715
rect 9485 -1735 9515 -1715
rect 9535 -1735 9565 -1715
rect 9585 -1735 9615 -1715
rect 9635 -1735 9665 -1715
rect 9685 -1735 9715 -1715
rect 9735 -1735 9765 -1715
rect 9785 -1735 9815 -1715
rect 9835 -1735 9865 -1715
rect 9885 -1735 9915 -1715
rect 9935 -1735 9965 -1715
rect 9985 -1735 10015 -1715
rect 10035 -1735 10065 -1715
rect 10085 -1735 10115 -1715
rect 10135 -1735 10165 -1715
rect 10185 -1735 10215 -1715
rect 10235 -1735 10265 -1715
rect 10285 -1735 10315 -1715
rect 10335 -1735 10365 -1715
rect 10385 -1735 10415 -1715
rect 10435 -1735 10465 -1715
rect 10485 -1735 10515 -1715
rect 10535 -1735 10565 -1715
rect 10585 -1735 10615 -1715
rect 10635 -1735 10665 -1715
rect 10685 -1735 10715 -1715
rect 10735 -1735 10765 -1715
rect 10785 -1735 10815 -1715
rect 10835 -1735 10865 -1715
rect 10885 -1735 10915 -1715
rect 10935 -1735 10965 -1715
rect 10985 -1735 11015 -1715
rect 11035 -1735 11065 -1715
rect 11085 -1735 11115 -1715
rect 11135 -1735 11165 -1715
rect 11185 -1735 11215 -1715
rect 11235 -1735 11265 -1715
rect 11285 -1735 11315 -1715
rect 11335 -1735 11365 -1715
rect 11385 -1735 11415 -1715
rect 11435 -1735 11465 -1715
rect 11485 -1735 11515 -1715
rect 11535 -1735 11565 -1715
rect 11585 -1735 11615 -1715
rect 11635 -1735 11665 -1715
rect 11685 -1735 11715 -1715
rect 11735 -1735 11765 -1715
rect 11785 -1735 11815 -1715
rect 11835 -1735 11865 -1715
rect 11885 -1735 11915 -1715
rect 11935 -1735 11965 -1715
rect 11985 -1735 12015 -1715
rect 12035 -1735 12065 -1715
rect 12085 -1735 12115 -1715
rect 12135 -1735 12165 -1715
rect 12185 -1735 12215 -1715
rect 12235 -1735 12265 -1715
rect 12285 -1735 12315 -1715
rect 12335 -1735 12365 -1715
rect 12385 -1735 12415 -1715
rect 12435 -1735 12465 -1715
rect 12485 -1735 12515 -1715
rect 12535 -1735 12565 -1715
rect 12585 -1735 12615 -1715
rect 12635 -1735 12665 -1715
rect 12685 -1735 12715 -1715
rect 12735 -1735 12765 -1715
rect 12785 -1735 12815 -1715
rect 12835 -1735 12865 -1715
rect 12885 -1735 12915 -1715
rect 12935 -1735 12965 -1715
rect 12985 -1735 13015 -1715
rect 13035 -1735 13065 -1715
rect 13085 -1735 13115 -1715
rect 13135 -1735 13165 -1715
rect 13185 -1735 13215 -1715
rect 13235 -1735 13265 -1715
rect 13285 -1735 13315 -1715
rect 13335 -1735 13365 -1715
rect 13385 -1735 13415 -1715
rect 13435 -1735 13465 -1715
rect 13485 -1735 13515 -1715
rect 13535 -1735 13565 -1715
rect 13585 -1735 13615 -1715
rect 13635 -1735 13665 -1715
rect 13685 -1735 13715 -1715
rect 13735 -1735 13765 -1715
rect 13785 -1735 13815 -1715
rect 13835 -1735 13865 -1715
rect 13885 -1735 13915 -1715
rect 13935 -1735 13965 -1715
rect 13985 -1735 14015 -1715
rect 14035 -1735 14065 -1715
rect 14085 -1735 14115 -1715
rect 14135 -1735 14165 -1715
rect 14185 -1735 14215 -1715
rect 14235 -1735 14265 -1715
rect 14285 -1735 14315 -1715
rect 14335 -1735 14365 -1715
rect 14385 -1735 14415 -1715
rect 14435 -1735 14465 -1715
rect 14485 -1735 14515 -1715
rect 14535 -1735 14565 -1715
rect 14585 -1735 14615 -1715
rect 14635 -1735 14665 -1715
rect 14685 -1735 14715 -1715
rect 14735 -1735 14765 -1715
rect 14785 -1735 14815 -1715
rect 14835 -1735 14865 -1715
rect 14885 -1735 14915 -1715
rect 14935 -1735 14965 -1715
rect 14985 -1735 15015 -1715
rect 15035 -1735 15065 -1715
rect 15085 -1735 15115 -1715
rect 15135 -1735 15165 -1715
rect 15185 -1735 15215 -1715
rect 15235 -1735 15265 -1715
rect 15285 -1735 15315 -1715
rect 15335 -1735 15365 -1715
rect 15385 -1735 15415 -1715
rect 15435 -1735 15465 -1715
rect 15485 -1735 15515 -1715
rect 15535 -1735 15565 -1715
rect 15585 -1735 15615 -1715
rect 15635 -1735 15665 -1715
rect 15685 -1735 15715 -1715
rect 15735 -1735 15765 -1715
rect 15785 -1735 15815 -1715
rect 15835 -1735 15865 -1715
rect 15885 -1735 15915 -1715
rect 15935 -1735 15965 -1715
rect 15985 -1735 16015 -1715
rect 16035 -1735 16065 -1715
rect 16085 -1735 16115 -1715
rect 16135 -1735 16165 -1715
rect 16185 -1735 16215 -1715
rect 16235 -1735 16265 -1715
rect 16285 -1735 16315 -1715
rect 16335 -1735 16365 -1715
rect 16385 -1735 16415 -1715
rect 16435 -1735 16465 -1715
rect 16485 -1735 16515 -1715
rect 16535 -1735 16565 -1715
rect 16585 -1735 16615 -1715
rect 16635 -1735 16665 -1715
rect 16685 -1735 16715 -1715
rect 16735 -1735 16765 -1715
rect 16785 -1735 16815 -1715
rect 16835 -1735 16865 -1715
rect 16885 -1735 16915 -1715
rect 16935 -1735 16965 -1715
rect 16985 -1735 17015 -1715
rect 17035 -1735 17065 -1715
rect 17085 -1735 17115 -1715
rect 17135 -1735 17165 -1715
rect 17185 -1735 17215 -1715
rect 17235 -1735 17265 -1715
rect 17285 -1735 17315 -1715
rect 17335 -1735 17365 -1715
rect 17385 -1735 17415 -1715
rect 17435 -1735 17465 -1715
rect 17485 -1735 17515 -1715
rect 17535 -1735 17565 -1715
rect 17585 -1735 17615 -1715
rect 17635 -1735 17665 -1715
rect 17685 -1735 17715 -1715
rect 17735 -1735 17765 -1715
rect 17785 -1735 17815 -1715
rect 17835 -1735 17865 -1715
rect 17885 -1735 17915 -1715
rect 17935 -1735 17965 -1715
rect 17985 -1735 18015 -1715
rect 18035 -1735 18065 -1715
rect 18085 -1735 18115 -1715
rect 18135 -1735 18165 -1715
rect 18185 -1735 18215 -1715
rect 18235 -1735 18265 -1715
rect 18285 -1735 18315 -1715
rect 18335 -1735 18365 -1715
rect 18385 -1735 18415 -1715
rect 18435 -1735 18465 -1715
rect 18485 -1735 18515 -1715
rect 18535 -1735 18565 -1715
rect 18585 -1735 18615 -1715
rect 18635 -1735 18665 -1715
rect 18685 -1735 18715 -1715
rect 18735 -1735 18765 -1715
rect 18785 -1735 18815 -1715
rect 18835 -1735 18865 -1715
rect 18885 -1735 18915 -1715
rect 18935 -1735 18965 -1715
rect 18985 -1735 19015 -1715
rect 19035 -1735 19065 -1715
rect 19085 -1735 19115 -1715
rect 19135 -1735 19165 -1715
rect 19185 -1735 19215 -1715
rect 19235 -1735 19265 -1715
rect 19285 -1735 19315 -1715
rect 19335 -1735 19365 -1715
rect 19385 -1735 19415 -1715
rect 19435 -1735 19465 -1715
rect 19485 -1735 19515 -1715
rect 19535 -1735 19565 -1715
rect 19585 -1735 19615 -1715
rect 19635 -1735 19665 -1715
rect 19685 -1735 19715 -1715
rect 19735 -1735 19765 -1715
rect 19785 -1735 19815 -1715
rect 19835 -1735 19865 -1715
rect 19885 -1735 19915 -1715
rect 19935 -1735 19965 -1715
rect 19985 -1735 20015 -1715
rect 20035 -1735 20065 -1715
rect 20085 -1735 20115 -1715
rect 20135 -1735 20165 -1715
rect 20185 -1735 20215 -1715
rect 20235 -1735 20265 -1715
rect 20285 -1735 20315 -1715
rect 20335 -1735 20365 -1715
rect 20385 -1735 20415 -1715
rect 20435 -1735 20465 -1715
rect 20485 -1735 20515 -1715
rect 20535 -1735 20565 -1715
rect 20585 -1735 20615 -1715
rect 20635 -1735 20665 -1715
rect 20685 -1735 20715 -1715
rect 20735 -1735 20765 -1715
rect 20785 -1735 20815 -1715
rect 20835 -1735 20865 -1715
rect 20885 -1735 20915 -1715
rect 20935 -1735 20965 -1715
rect 20985 -1735 21015 -1715
rect 21035 -1735 21065 -1715
rect 21085 -1735 21115 -1715
rect 21135 -1735 21165 -1715
rect 21185 -1735 21215 -1715
rect 21235 -1735 21265 -1715
rect 21285 -1735 21315 -1715
rect 21335 -1735 21365 -1715
rect 21385 -1735 21415 -1715
rect 21435 -1735 21465 -1715
rect 21485 -1735 21515 -1715
rect 21535 -1735 21565 -1715
rect 21585 -1735 21615 -1715
rect 21635 -1735 21665 -1715
rect 21685 -1735 21715 -1715
rect 21735 -1735 21765 -1715
rect 21785 -1735 21815 -1715
rect 21835 -1735 21865 -1715
rect 21885 -1735 21915 -1715
rect 21935 -1735 21965 -1715
rect 21985 -1735 22015 -1715
rect 22035 -1735 22065 -1715
rect 22085 -1735 22115 -1715
rect 22135 -1735 22165 -1715
rect 22185 -1735 22215 -1715
rect 22235 -1735 22265 -1715
rect 22285 -1735 22315 -1715
rect 22335 -1735 22365 -1715
rect 22385 -1735 22415 -1715
rect 22435 -1735 22465 -1715
rect 22485 -1735 22515 -1715
rect 22535 -1735 22565 -1715
rect 22585 -1735 22615 -1715
rect 22635 -1735 22665 -1715
rect 22685 -1735 22715 -1715
rect 22735 -1735 22765 -1715
rect 22785 -1735 22815 -1715
rect 22835 -1735 22865 -1715
rect 22885 -1735 22915 -1715
rect 22935 -1735 22965 -1715
rect 22985 -1735 23015 -1715
rect 23035 -1735 23065 -1715
rect 23085 -1735 23115 -1715
rect 23135 -1735 23165 -1715
rect 23185 -1735 23215 -1715
rect 23235 -1735 23265 -1715
rect 23285 -1735 23315 -1715
rect 23335 -1735 23365 -1715
rect 23385 -1735 23415 -1715
rect 23435 -1735 23465 -1715
rect 23485 -1735 23515 -1715
rect 23535 -1735 23565 -1715
rect 23585 -1735 23615 -1715
rect 23635 -1735 23665 -1715
rect 23685 -1735 23715 -1715
rect 23735 -1735 23765 -1715
rect 23785 -1735 23815 -1715
rect 23835 -1735 23865 -1715
rect 23885 -1735 23915 -1715
rect 23935 -1735 23965 -1715
rect 23985 -1735 24015 -1715
rect 24035 -1735 24065 -1715
rect 24085 -1735 24115 -1715
rect 24135 -1735 24165 -1715
rect 24185 -1735 24215 -1715
rect 24235 -1735 24265 -1715
rect 24285 -1735 24315 -1715
rect 24335 -1735 24365 -1715
rect 24385 -1735 24415 -1715
rect 24435 -1735 24465 -1715
rect 24485 -1735 24515 -1715
rect 24535 -1735 24565 -1715
rect 24585 -1735 24615 -1715
rect 24635 -1735 24665 -1715
rect 24685 -1735 24715 -1715
rect 24735 -1735 24765 -1715
rect 24785 -1735 24815 -1715
rect 24835 -1735 24865 -1715
rect 24885 -1735 24915 -1715
rect 24935 -1735 24965 -1715
rect 24985 -1735 25015 -1715
rect 25035 -1735 25065 -1715
rect 25085 -1735 25115 -1715
rect 25135 -1735 25165 -1715
rect 25185 -1735 25215 -1715
rect 25235 -1735 25265 -1715
rect 25285 -1735 25315 -1715
rect 25335 -1735 25365 -1715
rect 25385 -1735 25415 -1715
rect 25435 -1735 25465 -1715
rect 25485 -1735 25515 -1715
rect 25535 -1735 25565 -1715
rect 25585 -1735 25615 -1715
rect 25635 -1735 25665 -1715
rect 25685 -1735 25715 -1715
rect 25735 -1735 25765 -1715
rect 25785 -1735 25815 -1715
rect 25835 -1735 25865 -1715
rect 25885 -1735 25915 -1715
rect 25935 -1735 25965 -1715
rect 25985 -1735 26015 -1715
rect 26035 -1735 26065 -1715
rect 26085 -1735 26115 -1715
rect 26135 -1735 26165 -1715
rect 26185 -1735 26215 -1715
rect 26235 -1735 26265 -1715
rect 26285 -1735 26315 -1715
rect 26335 -1735 26365 -1715
rect 26385 -1735 26415 -1715
rect 26435 -1735 26465 -1715
rect 26485 -1735 26515 -1715
rect 26535 -1735 26565 -1715
rect 26585 -1735 26615 -1715
rect 26635 -1735 26665 -1715
rect 26685 -1735 26715 -1715
rect 26735 -1735 26765 -1715
rect 26785 -1735 26815 -1715
rect 26835 -1735 26865 -1715
rect 26885 -1735 26915 -1715
rect 26935 -1735 26965 -1715
rect 26985 -1735 27015 -1715
rect 27035 -1735 27065 -1715
rect 27085 -1735 27115 -1715
rect 27135 -1735 27165 -1715
rect 27185 -1735 27215 -1715
rect 27235 -1735 27265 -1715
rect 27285 -1735 27315 -1715
rect 27335 -1735 27365 -1715
rect 27385 -1735 27415 -1715
rect 27435 -1735 27465 -1715
rect 27485 -1735 27515 -1715
rect 27535 -1735 27565 -1715
rect 27585 -1735 27615 -1715
rect 27635 -1735 27665 -1715
rect 27685 -1735 27715 -1715
rect 27735 -1735 27765 -1715
rect 27785 -1735 27815 -1715
rect 27835 -1735 27865 -1715
rect 27885 -1735 27915 -1715
rect 27935 -1735 27965 -1715
rect 27985 -1735 28015 -1715
rect 28035 -1735 28065 -1715
rect 28085 -1735 28115 -1715
rect 28135 -1735 28165 -1715
rect 28185 -1735 28215 -1715
rect 28235 -1735 28265 -1715
rect 28285 -1735 28315 -1715
rect 28335 -1735 28365 -1715
rect 28385 -1735 28415 -1715
rect 28435 -1735 28465 -1715
rect 28485 -1735 28515 -1715
rect 28535 -1735 28565 -1715
rect 28585 -1735 28615 -1715
rect 28635 -1735 28665 -1715
rect 28685 -1735 28715 -1715
rect 28735 -1735 28765 -1715
rect 28785 -1735 28800 -1715
rect -650 -1750 28800 -1735
rect -650 -1865 28800 -1850
rect -650 -1885 -635 -1865
rect -615 -1885 -585 -1865
rect -565 -1885 -535 -1865
rect -515 -1885 -485 -1865
rect -465 -1885 -435 -1865
rect -415 -1885 -385 -1865
rect -365 -1885 -335 -1865
rect -315 -1885 -285 -1865
rect -265 -1885 -235 -1865
rect -215 -1885 -185 -1865
rect -165 -1885 -135 -1865
rect -115 -1885 -85 -1865
rect -65 -1885 -35 -1865
rect -15 -1885 15 -1865
rect 35 -1885 65 -1865
rect 85 -1885 115 -1865
rect 135 -1885 165 -1865
rect 185 -1885 215 -1865
rect 235 -1885 265 -1865
rect 285 -1885 315 -1865
rect 335 -1885 365 -1865
rect 385 -1885 415 -1865
rect 435 -1885 465 -1865
rect 485 -1885 515 -1865
rect 535 -1885 565 -1865
rect 585 -1885 615 -1865
rect 635 -1885 665 -1865
rect 685 -1885 715 -1865
rect 735 -1885 765 -1865
rect 785 -1885 815 -1865
rect 835 -1885 865 -1865
rect 885 -1885 915 -1865
rect 935 -1885 965 -1865
rect 985 -1885 1015 -1865
rect 1035 -1885 1065 -1865
rect 1085 -1885 1115 -1865
rect 1135 -1885 1165 -1865
rect 1185 -1885 1215 -1865
rect 1235 -1885 1265 -1865
rect 1285 -1885 1315 -1865
rect 1335 -1885 1365 -1865
rect 1385 -1885 1415 -1865
rect 1435 -1885 1465 -1865
rect 1485 -1885 1515 -1865
rect 1535 -1885 1565 -1865
rect 1585 -1885 1615 -1865
rect 1635 -1885 1665 -1865
rect 1685 -1885 1715 -1865
rect 1735 -1885 1765 -1865
rect 1785 -1885 1815 -1865
rect 1835 -1885 1865 -1865
rect 1885 -1885 1915 -1865
rect 1935 -1885 1965 -1865
rect 1985 -1885 2015 -1865
rect 2035 -1885 2065 -1865
rect 2085 -1885 2115 -1865
rect 2135 -1885 2165 -1865
rect 2185 -1885 2215 -1865
rect 2235 -1885 2265 -1865
rect 2285 -1885 2315 -1865
rect 2335 -1885 2365 -1865
rect 2385 -1885 2415 -1865
rect 2435 -1885 2465 -1865
rect 2485 -1885 2515 -1865
rect 2535 -1885 2565 -1865
rect 2585 -1885 2615 -1865
rect 2635 -1885 2665 -1865
rect 2685 -1885 2715 -1865
rect 2735 -1885 2765 -1865
rect 2785 -1885 2815 -1865
rect 2835 -1885 2865 -1865
rect 2885 -1885 2915 -1865
rect 2935 -1885 2965 -1865
rect 2985 -1885 3015 -1865
rect 3035 -1885 3065 -1865
rect 3085 -1885 3115 -1865
rect 3135 -1885 3165 -1865
rect 3185 -1885 3215 -1865
rect 3235 -1885 3265 -1865
rect 3285 -1885 3315 -1865
rect 3335 -1885 3365 -1865
rect 3385 -1885 3415 -1865
rect 3435 -1885 3465 -1865
rect 3485 -1885 3515 -1865
rect 3535 -1885 3565 -1865
rect 3585 -1885 3615 -1865
rect 3635 -1885 3665 -1865
rect 3685 -1885 3715 -1865
rect 3735 -1885 3765 -1865
rect 3785 -1885 3815 -1865
rect 3835 -1885 3865 -1865
rect 3885 -1885 3915 -1865
rect 3935 -1885 3965 -1865
rect 3985 -1885 4015 -1865
rect 4035 -1885 4065 -1865
rect 4085 -1885 4115 -1865
rect 4135 -1885 4165 -1865
rect 4185 -1885 4215 -1865
rect 4235 -1885 4265 -1865
rect 4285 -1885 4315 -1865
rect 4335 -1885 4365 -1865
rect 4385 -1885 4415 -1865
rect 4435 -1885 4465 -1865
rect 4485 -1885 4515 -1865
rect 4535 -1885 4565 -1865
rect 4585 -1885 4615 -1865
rect 4635 -1885 4665 -1865
rect 4685 -1885 4715 -1865
rect 4735 -1885 4765 -1865
rect 4785 -1885 4815 -1865
rect 4835 -1885 4865 -1865
rect 4885 -1885 4915 -1865
rect 4935 -1885 4965 -1865
rect 4985 -1885 5015 -1865
rect 5035 -1885 5065 -1865
rect 5085 -1885 5115 -1865
rect 5135 -1885 5165 -1865
rect 5185 -1885 5215 -1865
rect 5235 -1885 5265 -1865
rect 5285 -1885 5315 -1865
rect 5335 -1885 5365 -1865
rect 5385 -1885 5415 -1865
rect 5435 -1885 5465 -1865
rect 5485 -1885 5515 -1865
rect 5535 -1885 5565 -1865
rect 5585 -1885 5615 -1865
rect 5635 -1885 5665 -1865
rect 5685 -1885 5715 -1865
rect 5735 -1885 5765 -1865
rect 5785 -1885 5815 -1865
rect 5835 -1885 5865 -1865
rect 5885 -1885 5915 -1865
rect 5935 -1885 5965 -1865
rect 5985 -1885 6015 -1865
rect 6035 -1885 6065 -1865
rect 6085 -1885 6115 -1865
rect 6135 -1885 6165 -1865
rect 6185 -1885 6215 -1865
rect 6235 -1885 6265 -1865
rect 6285 -1885 6315 -1865
rect 6335 -1885 6365 -1865
rect 6385 -1885 6415 -1865
rect 6435 -1885 6465 -1865
rect 6485 -1885 6515 -1865
rect 6535 -1885 6565 -1865
rect 6585 -1885 6615 -1865
rect 6635 -1885 6665 -1865
rect 6685 -1885 6715 -1865
rect 6735 -1885 6765 -1865
rect 6785 -1885 6815 -1865
rect 6835 -1885 6865 -1865
rect 6885 -1885 6915 -1865
rect 6935 -1885 6965 -1865
rect 6985 -1885 7015 -1865
rect 7035 -1885 7065 -1865
rect 7085 -1885 7115 -1865
rect 7135 -1885 7165 -1865
rect 7185 -1885 7215 -1865
rect 7235 -1885 7265 -1865
rect 7285 -1885 7315 -1865
rect 7335 -1885 7365 -1865
rect 7385 -1885 7415 -1865
rect 7435 -1885 7465 -1865
rect 7485 -1885 7515 -1865
rect 7535 -1885 7565 -1865
rect 7585 -1885 7615 -1865
rect 7635 -1885 7665 -1865
rect 7685 -1885 7715 -1865
rect 7735 -1885 7765 -1865
rect 7785 -1885 7815 -1865
rect 7835 -1885 7865 -1865
rect 7885 -1885 7915 -1865
rect 7935 -1885 7965 -1865
rect 7985 -1885 8015 -1865
rect 8035 -1885 8065 -1865
rect 8085 -1885 8115 -1865
rect 8135 -1885 8165 -1865
rect 8185 -1885 8215 -1865
rect 8235 -1885 8265 -1865
rect 8285 -1885 8315 -1865
rect 8335 -1885 8365 -1865
rect 8385 -1885 8415 -1865
rect 8435 -1885 8465 -1865
rect 8485 -1885 8515 -1865
rect 8535 -1885 8565 -1865
rect 8585 -1885 8615 -1865
rect 8635 -1885 8665 -1865
rect 8685 -1885 8715 -1865
rect 8735 -1885 8765 -1865
rect 8785 -1885 8815 -1865
rect 8835 -1885 8865 -1865
rect 8885 -1885 8915 -1865
rect 8935 -1885 8965 -1865
rect 8985 -1885 9015 -1865
rect 9035 -1885 9065 -1865
rect 9085 -1885 9115 -1865
rect 9135 -1885 9165 -1865
rect 9185 -1885 9215 -1865
rect 9235 -1885 9265 -1865
rect 9285 -1885 9315 -1865
rect 9335 -1885 9365 -1865
rect 9385 -1885 9415 -1865
rect 9435 -1885 9465 -1865
rect 9485 -1885 9515 -1865
rect 9535 -1885 9565 -1865
rect 9585 -1885 9615 -1865
rect 9635 -1885 9665 -1865
rect 9685 -1885 9715 -1865
rect 9735 -1885 9765 -1865
rect 9785 -1885 9815 -1865
rect 9835 -1885 9865 -1865
rect 9885 -1885 9915 -1865
rect 9935 -1885 9965 -1865
rect 9985 -1885 10015 -1865
rect 10035 -1885 10065 -1865
rect 10085 -1885 10115 -1865
rect 10135 -1885 10165 -1865
rect 10185 -1885 10215 -1865
rect 10235 -1885 10265 -1865
rect 10285 -1885 10315 -1865
rect 10335 -1885 10365 -1865
rect 10385 -1885 10415 -1865
rect 10435 -1885 10465 -1865
rect 10485 -1885 10515 -1865
rect 10535 -1885 10565 -1865
rect 10585 -1885 10615 -1865
rect 10635 -1885 10665 -1865
rect 10685 -1885 10715 -1865
rect 10735 -1885 10765 -1865
rect 10785 -1885 10815 -1865
rect 10835 -1885 10865 -1865
rect 10885 -1885 10915 -1865
rect 10935 -1885 10965 -1865
rect 10985 -1885 11015 -1865
rect 11035 -1885 11065 -1865
rect 11085 -1885 11115 -1865
rect 11135 -1885 11165 -1865
rect 11185 -1885 11215 -1865
rect 11235 -1885 11265 -1865
rect 11285 -1885 11315 -1865
rect 11335 -1885 11365 -1865
rect 11385 -1885 11415 -1865
rect 11435 -1885 11465 -1865
rect 11485 -1885 11515 -1865
rect 11535 -1885 11565 -1865
rect 11585 -1885 11615 -1865
rect 11635 -1885 11665 -1865
rect 11685 -1885 11715 -1865
rect 11735 -1885 11765 -1865
rect 11785 -1885 11815 -1865
rect 11835 -1885 11865 -1865
rect 11885 -1885 11915 -1865
rect 11935 -1885 11965 -1865
rect 11985 -1885 12015 -1865
rect 12035 -1885 12065 -1865
rect 12085 -1885 12115 -1865
rect 12135 -1885 12165 -1865
rect 12185 -1885 12215 -1865
rect 12235 -1885 12265 -1865
rect 12285 -1885 12315 -1865
rect 12335 -1885 12365 -1865
rect 12385 -1885 12415 -1865
rect 12435 -1885 12465 -1865
rect 12485 -1885 12515 -1865
rect 12535 -1885 12565 -1865
rect 12585 -1885 12615 -1865
rect 12635 -1885 12665 -1865
rect 12685 -1885 12715 -1865
rect 12735 -1885 12765 -1865
rect 12785 -1885 12815 -1865
rect 12835 -1885 12865 -1865
rect 12885 -1885 12915 -1865
rect 12935 -1885 12965 -1865
rect 12985 -1885 13015 -1865
rect 13035 -1885 13065 -1865
rect 13085 -1885 13115 -1865
rect 13135 -1885 13165 -1865
rect 13185 -1885 13215 -1865
rect 13235 -1885 13265 -1865
rect 13285 -1885 13315 -1865
rect 13335 -1885 13365 -1865
rect 13385 -1885 13415 -1865
rect 13435 -1885 13465 -1865
rect 13485 -1885 13515 -1865
rect 13535 -1885 13565 -1865
rect 13585 -1885 13615 -1865
rect 13635 -1885 13665 -1865
rect 13685 -1885 13715 -1865
rect 13735 -1885 13765 -1865
rect 13785 -1885 13815 -1865
rect 13835 -1885 13865 -1865
rect 13885 -1885 13915 -1865
rect 13935 -1885 13965 -1865
rect 13985 -1885 14015 -1865
rect 14035 -1885 14065 -1865
rect 14085 -1885 14115 -1865
rect 14135 -1885 14165 -1865
rect 14185 -1885 14215 -1865
rect 14235 -1885 14265 -1865
rect 14285 -1885 14315 -1865
rect 14335 -1885 14365 -1865
rect 14385 -1885 14415 -1865
rect 14435 -1885 14465 -1865
rect 14485 -1885 14515 -1865
rect 14535 -1885 14565 -1865
rect 14585 -1885 14615 -1865
rect 14635 -1885 14665 -1865
rect 14685 -1885 14715 -1865
rect 14735 -1885 14765 -1865
rect 14785 -1885 14815 -1865
rect 14835 -1885 14865 -1865
rect 14885 -1885 14915 -1865
rect 14935 -1885 14965 -1865
rect 14985 -1885 15015 -1865
rect 15035 -1885 15065 -1865
rect 15085 -1885 15115 -1865
rect 15135 -1885 15165 -1865
rect 15185 -1885 15215 -1865
rect 15235 -1885 15265 -1865
rect 15285 -1885 15315 -1865
rect 15335 -1885 15365 -1865
rect 15385 -1885 15415 -1865
rect 15435 -1885 15465 -1865
rect 15485 -1885 15515 -1865
rect 15535 -1885 15565 -1865
rect 15585 -1885 15615 -1865
rect 15635 -1885 15665 -1865
rect 15685 -1885 15715 -1865
rect 15735 -1885 15765 -1865
rect 15785 -1885 15815 -1865
rect 15835 -1885 15865 -1865
rect 15885 -1885 15915 -1865
rect 15935 -1885 15965 -1865
rect 15985 -1885 16015 -1865
rect 16035 -1885 16065 -1865
rect 16085 -1885 16115 -1865
rect 16135 -1885 16165 -1865
rect 16185 -1885 16215 -1865
rect 16235 -1885 16265 -1865
rect 16285 -1885 16315 -1865
rect 16335 -1885 16365 -1865
rect 16385 -1885 16415 -1865
rect 16435 -1885 16465 -1865
rect 16485 -1885 16515 -1865
rect 16535 -1885 16565 -1865
rect 16585 -1885 16615 -1865
rect 16635 -1885 16665 -1865
rect 16685 -1885 16715 -1865
rect 16735 -1885 16765 -1865
rect 16785 -1885 16815 -1865
rect 16835 -1885 16865 -1865
rect 16885 -1885 16915 -1865
rect 16935 -1885 16965 -1865
rect 16985 -1885 17015 -1865
rect 17035 -1885 17065 -1865
rect 17085 -1885 17115 -1865
rect 17135 -1885 17165 -1865
rect 17185 -1885 17215 -1865
rect 17235 -1885 17265 -1865
rect 17285 -1885 17315 -1865
rect 17335 -1885 17365 -1865
rect 17385 -1885 17415 -1865
rect 17435 -1885 17465 -1865
rect 17485 -1885 17515 -1865
rect 17535 -1885 17565 -1865
rect 17585 -1885 17615 -1865
rect 17635 -1885 17665 -1865
rect 17685 -1885 17715 -1865
rect 17735 -1885 17765 -1865
rect 17785 -1885 17815 -1865
rect 17835 -1885 17865 -1865
rect 17885 -1885 17915 -1865
rect 17935 -1885 17965 -1865
rect 17985 -1885 18015 -1865
rect 18035 -1885 18065 -1865
rect 18085 -1885 18115 -1865
rect 18135 -1885 18165 -1865
rect 18185 -1885 18215 -1865
rect 18235 -1885 18265 -1865
rect 18285 -1885 18315 -1865
rect 18335 -1885 18365 -1865
rect 18385 -1885 18415 -1865
rect 18435 -1885 18465 -1865
rect 18485 -1885 18515 -1865
rect 18535 -1885 18565 -1865
rect 18585 -1885 18615 -1865
rect 18635 -1885 18665 -1865
rect 18685 -1885 18715 -1865
rect 18735 -1885 18765 -1865
rect 18785 -1885 18815 -1865
rect 18835 -1885 18865 -1865
rect 18885 -1885 18915 -1865
rect 18935 -1885 18965 -1865
rect 18985 -1885 19015 -1865
rect 19035 -1885 19065 -1865
rect 19085 -1885 19115 -1865
rect 19135 -1885 19165 -1865
rect 19185 -1885 19215 -1865
rect 19235 -1885 19265 -1865
rect 19285 -1885 19315 -1865
rect 19335 -1885 19365 -1865
rect 19385 -1885 19415 -1865
rect 19435 -1885 19465 -1865
rect 19485 -1885 19515 -1865
rect 19535 -1885 19565 -1865
rect 19585 -1885 19615 -1865
rect 19635 -1885 19665 -1865
rect 19685 -1885 19715 -1865
rect 19735 -1885 19765 -1865
rect 19785 -1885 19815 -1865
rect 19835 -1885 19865 -1865
rect 19885 -1885 19915 -1865
rect 19935 -1885 19965 -1865
rect 19985 -1885 20015 -1865
rect 20035 -1885 20065 -1865
rect 20085 -1885 20115 -1865
rect 20135 -1885 20165 -1865
rect 20185 -1885 20215 -1865
rect 20235 -1885 20265 -1865
rect 20285 -1885 20315 -1865
rect 20335 -1885 20365 -1865
rect 20385 -1885 20415 -1865
rect 20435 -1885 20465 -1865
rect 20485 -1885 20515 -1865
rect 20535 -1885 20565 -1865
rect 20585 -1885 20615 -1865
rect 20635 -1885 20665 -1865
rect 20685 -1885 20715 -1865
rect 20735 -1885 20765 -1865
rect 20785 -1885 20815 -1865
rect 20835 -1885 20865 -1865
rect 20885 -1885 20915 -1865
rect 20935 -1885 20965 -1865
rect 20985 -1885 21015 -1865
rect 21035 -1885 21065 -1865
rect 21085 -1885 21115 -1865
rect 21135 -1885 21165 -1865
rect 21185 -1885 21215 -1865
rect 21235 -1885 21265 -1865
rect 21285 -1885 21315 -1865
rect 21335 -1885 21365 -1865
rect 21385 -1885 21415 -1865
rect 21435 -1885 21465 -1865
rect 21485 -1885 21515 -1865
rect 21535 -1885 21565 -1865
rect 21585 -1885 21615 -1865
rect 21635 -1885 21665 -1865
rect 21685 -1885 21715 -1865
rect 21735 -1885 21765 -1865
rect 21785 -1885 21815 -1865
rect 21835 -1885 21865 -1865
rect 21885 -1885 21915 -1865
rect 21935 -1885 21965 -1865
rect 21985 -1885 22015 -1865
rect 22035 -1885 22065 -1865
rect 22085 -1885 22115 -1865
rect 22135 -1885 22165 -1865
rect 22185 -1885 22215 -1865
rect 22235 -1885 22265 -1865
rect 22285 -1885 22315 -1865
rect 22335 -1885 22365 -1865
rect 22385 -1885 22415 -1865
rect 22435 -1885 22465 -1865
rect 22485 -1885 22515 -1865
rect 22535 -1885 22565 -1865
rect 22585 -1885 22615 -1865
rect 22635 -1885 22665 -1865
rect 22685 -1885 22715 -1865
rect 22735 -1885 22765 -1865
rect 22785 -1885 22815 -1865
rect 22835 -1885 22865 -1865
rect 22885 -1885 22915 -1865
rect 22935 -1885 22965 -1865
rect 22985 -1885 23015 -1865
rect 23035 -1885 23065 -1865
rect 23085 -1885 23115 -1865
rect 23135 -1885 23165 -1865
rect 23185 -1885 23215 -1865
rect 23235 -1885 23265 -1865
rect 23285 -1885 23315 -1865
rect 23335 -1885 23365 -1865
rect 23385 -1885 23415 -1865
rect 23435 -1885 23465 -1865
rect 23485 -1885 23515 -1865
rect 23535 -1885 23565 -1865
rect 23585 -1885 23615 -1865
rect 23635 -1885 23665 -1865
rect 23685 -1885 23715 -1865
rect 23735 -1885 23765 -1865
rect 23785 -1885 23815 -1865
rect 23835 -1885 23865 -1865
rect 23885 -1885 23915 -1865
rect 23935 -1885 23965 -1865
rect 23985 -1885 24015 -1865
rect 24035 -1885 24065 -1865
rect 24085 -1885 24115 -1865
rect 24135 -1885 24165 -1865
rect 24185 -1885 24215 -1865
rect 24235 -1885 24265 -1865
rect 24285 -1885 24315 -1865
rect 24335 -1885 24365 -1865
rect 24385 -1885 24415 -1865
rect 24435 -1885 24465 -1865
rect 24485 -1885 24515 -1865
rect 24535 -1885 24565 -1865
rect 24585 -1885 24615 -1865
rect 24635 -1885 24665 -1865
rect 24685 -1885 24715 -1865
rect 24735 -1885 24765 -1865
rect 24785 -1885 24815 -1865
rect 24835 -1885 24865 -1865
rect 24885 -1885 24915 -1865
rect 24935 -1885 24965 -1865
rect 24985 -1885 25015 -1865
rect 25035 -1885 25065 -1865
rect 25085 -1885 25115 -1865
rect 25135 -1885 25165 -1865
rect 25185 -1885 25215 -1865
rect 25235 -1885 25265 -1865
rect 25285 -1885 25315 -1865
rect 25335 -1885 25365 -1865
rect 25385 -1885 25415 -1865
rect 25435 -1885 25465 -1865
rect 25485 -1885 25515 -1865
rect 25535 -1885 25565 -1865
rect 25585 -1885 25615 -1865
rect 25635 -1885 25665 -1865
rect 25685 -1885 25715 -1865
rect 25735 -1885 25765 -1865
rect 25785 -1885 25815 -1865
rect 25835 -1885 25865 -1865
rect 25885 -1885 25915 -1865
rect 25935 -1885 25965 -1865
rect 25985 -1885 26015 -1865
rect 26035 -1885 26065 -1865
rect 26085 -1885 26115 -1865
rect 26135 -1885 26165 -1865
rect 26185 -1885 26215 -1865
rect 26235 -1885 26265 -1865
rect 26285 -1885 26315 -1865
rect 26335 -1885 26365 -1865
rect 26385 -1885 26415 -1865
rect 26435 -1885 26465 -1865
rect 26485 -1885 26515 -1865
rect 26535 -1885 26565 -1865
rect 26585 -1885 26615 -1865
rect 26635 -1885 26665 -1865
rect 26685 -1885 26715 -1865
rect 26735 -1885 26765 -1865
rect 26785 -1885 26815 -1865
rect 26835 -1885 26865 -1865
rect 26885 -1885 26915 -1865
rect 26935 -1885 26965 -1865
rect 26985 -1885 27015 -1865
rect 27035 -1885 27065 -1865
rect 27085 -1885 27115 -1865
rect 27135 -1885 27165 -1865
rect 27185 -1885 27215 -1865
rect 27235 -1885 27265 -1865
rect 27285 -1885 27315 -1865
rect 27335 -1885 27365 -1865
rect 27385 -1885 27415 -1865
rect 27435 -1885 27465 -1865
rect 27485 -1885 27515 -1865
rect 27535 -1885 27565 -1865
rect 27585 -1885 27615 -1865
rect 27635 -1885 27665 -1865
rect 27685 -1885 27715 -1865
rect 27735 -1885 27765 -1865
rect 27785 -1885 27815 -1865
rect 27835 -1885 27865 -1865
rect 27885 -1885 27915 -1865
rect 27935 -1885 27965 -1865
rect 27985 -1885 28015 -1865
rect 28035 -1885 28065 -1865
rect 28085 -1885 28115 -1865
rect 28135 -1885 28165 -1865
rect 28185 -1885 28215 -1865
rect 28235 -1885 28265 -1865
rect 28285 -1885 28315 -1865
rect 28335 -1885 28365 -1865
rect 28385 -1885 28415 -1865
rect 28435 -1885 28465 -1865
rect 28485 -1885 28515 -1865
rect 28535 -1885 28565 -1865
rect 28585 -1885 28615 -1865
rect 28635 -1885 28665 -1865
rect 28685 -1885 28715 -1865
rect 28735 -1885 28765 -1865
rect 28785 -1885 28800 -1865
rect -650 -1900 28800 -1885
<< viali >>
rect -635 5565 -615 5585
rect 8365 5565 8385 5585
rect 8665 5565 8685 5585
rect 8965 5565 8985 5585
rect 9265 5565 9285 5585
rect 9565 5565 9585 5585
rect 9865 5565 9885 5585
rect 10165 5565 10185 5585
rect 10465 5565 10485 5585
rect 10765 5565 10785 5585
rect 11965 5565 11985 5585
rect 13165 5565 13185 5585
rect 14365 5565 14385 5585
rect 15565 5565 15585 5585
rect 20365 5565 20385 5585
rect 22465 5565 22485 5585
rect 24565 5565 24585 5585
rect 26665 5565 26685 5585
rect 28165 5565 28185 5585
rect 28765 5565 28785 5585
rect 32065 5565 32085 5585
rect -635 5465 -615 5485
rect -635 5415 -615 5435
rect -635 5365 -615 5385
rect -635 5315 -615 5335
rect -635 5265 -615 5285
rect -635 5215 -615 5235
rect -635 5165 -615 5185
rect -635 5115 -615 5135
rect -635 5065 -615 5085
rect -635 5015 -615 5035
rect -485 5465 -465 5485
rect -485 5415 -465 5435
rect -485 5365 -465 5385
rect -485 5315 -465 5335
rect -485 5265 -465 5285
rect -485 5215 -465 5235
rect -485 5165 -465 5185
rect -485 5115 -465 5135
rect -485 5065 -465 5085
rect -485 5015 -465 5035
rect -335 5465 -315 5485
rect -335 5415 -315 5435
rect -335 5365 -315 5385
rect -335 5315 -315 5335
rect -335 5265 -315 5285
rect -335 5215 -315 5235
rect -335 5165 -315 5185
rect -335 5115 -315 5135
rect -185 5465 -165 5485
rect -185 5415 -165 5435
rect -185 5365 -165 5385
rect -185 5315 -165 5335
rect -185 5265 -165 5285
rect -185 5215 -165 5235
rect -185 5165 -165 5185
rect -185 5115 -165 5135
rect -185 5065 -165 5085
rect -185 5015 -165 5035
rect -35 5465 -15 5485
rect -35 5415 -15 5435
rect -35 5365 -15 5385
rect -35 5315 -15 5335
rect -35 5265 -15 5285
rect -35 5215 -15 5235
rect -35 5165 -15 5185
rect -35 5115 -15 5135
rect 565 5465 585 5485
rect 565 5415 585 5435
rect 565 5365 585 5385
rect 565 5315 585 5335
rect 565 5265 585 5285
rect 565 5215 585 5235
rect 565 5165 585 5185
rect 565 5115 585 5135
rect 565 5065 585 5085
rect 565 5015 585 5035
rect 715 5365 735 5385
rect 715 5315 735 5335
rect 715 5265 735 5285
rect 715 5215 735 5235
rect 715 5165 735 5185
rect 715 5115 735 5135
rect 715 5065 735 5085
rect 715 5015 735 5035
rect 865 5465 885 5485
rect 865 5415 885 5435
rect 865 5365 885 5385
rect 865 5315 885 5335
rect 865 5265 885 5285
rect 865 5215 885 5235
rect 865 5165 885 5185
rect 865 5115 885 5135
rect 1015 5365 1035 5385
rect 1015 5315 1035 5335
rect 1015 5265 1035 5285
rect 1015 5215 1035 5235
rect 1015 5165 1035 5185
rect 1015 5115 1035 5135
rect 1015 5065 1035 5085
rect 1165 5465 1185 5485
rect 1165 5415 1185 5435
rect 1165 5365 1185 5385
rect 1165 5315 1185 5335
rect 1165 5265 1185 5285
rect 1165 5215 1185 5235
rect 1165 5165 1185 5185
rect 1165 5115 1185 5135
rect 1315 5365 1335 5385
rect 1315 5315 1335 5335
rect 1315 5265 1335 5285
rect 1315 5215 1335 5235
rect 1315 5165 1335 5185
rect 1315 5115 1335 5135
rect 1315 5065 1335 5085
rect 1465 5465 1485 5485
rect 1465 5415 1485 5435
rect 1465 5365 1485 5385
rect 1465 5315 1485 5335
rect 1465 5265 1485 5285
rect 1465 5215 1485 5235
rect 1465 5165 1485 5185
rect 1465 5115 1485 5135
rect 1615 5365 1635 5385
rect 1615 5315 1635 5335
rect 1615 5265 1635 5285
rect 1615 5215 1635 5235
rect 1615 5165 1635 5185
rect 1615 5115 1635 5135
rect 1615 5065 1635 5085
rect 1765 5465 1785 5485
rect 1765 5415 1785 5435
rect 1765 5365 1785 5385
rect 1765 5315 1785 5335
rect 1765 5265 1785 5285
rect 1765 5215 1785 5235
rect 1765 5165 1785 5185
rect 1765 5115 1785 5135
rect 1765 5065 1785 5085
rect 1765 5015 1785 5035
rect 1915 5365 1935 5385
rect 1915 5315 1935 5335
rect 1915 5265 1935 5285
rect 1915 5215 1935 5235
rect 1915 5165 1935 5185
rect 1915 5115 1935 5135
rect 1915 5065 1935 5085
rect 1915 5015 1935 5035
rect 2065 5465 2085 5485
rect 2065 5415 2085 5435
rect 2065 5365 2085 5385
rect 2065 5315 2085 5335
rect 2065 5265 2085 5285
rect 2065 5215 2085 5235
rect 2065 5165 2085 5185
rect 2065 5115 2085 5135
rect 2215 5365 2235 5385
rect 2215 5315 2235 5335
rect 2215 5265 2235 5285
rect 2215 5215 2235 5235
rect 2215 5165 2235 5185
rect 2215 5115 2235 5135
rect 2215 5065 2235 5085
rect 2215 5015 2235 5035
rect 2365 5465 2385 5485
rect 2365 5415 2385 5435
rect 2365 5365 2385 5385
rect 2365 5315 2385 5335
rect 2365 5265 2385 5285
rect 2365 5215 2385 5235
rect 2365 5165 2385 5185
rect 2365 5115 2385 5135
rect 2365 5065 2385 5085
rect 2365 5015 2385 5035
rect 2515 5365 2535 5385
rect 2515 5315 2535 5335
rect 2515 5265 2535 5285
rect 2515 5215 2535 5235
rect 2515 5165 2535 5185
rect 2515 5115 2535 5135
rect 2515 5065 2535 5085
rect 2665 5465 2685 5485
rect 2665 5415 2685 5435
rect 2665 5365 2685 5385
rect 2665 5315 2685 5335
rect 2665 5265 2685 5285
rect 2665 5215 2685 5235
rect 2665 5165 2685 5185
rect 2665 5115 2685 5135
rect 2815 5365 2835 5385
rect 2815 5315 2835 5335
rect 2815 5265 2835 5285
rect 2815 5215 2835 5235
rect 2815 5165 2835 5185
rect 2815 5115 2835 5135
rect 2815 5065 2835 5085
rect 2965 5465 2985 5485
rect 2965 5415 2985 5435
rect 2965 5365 2985 5385
rect 2965 5315 2985 5335
rect 2965 5265 2985 5285
rect 2965 5215 2985 5235
rect 2965 5165 2985 5185
rect 2965 5115 2985 5135
rect 3115 5365 3135 5385
rect 3115 5315 3135 5335
rect 3115 5265 3135 5285
rect 3115 5215 3135 5235
rect 3115 5165 3135 5185
rect 3115 5115 3135 5135
rect 3115 5065 3135 5085
rect 3265 5465 3285 5485
rect 3265 5415 3285 5435
rect 3265 5365 3285 5385
rect 3265 5315 3285 5335
rect 3265 5265 3285 5285
rect 3265 5215 3285 5235
rect 3265 5165 3285 5185
rect 3265 5115 3285 5135
rect 3415 5365 3435 5385
rect 3415 5315 3435 5335
rect 3415 5265 3435 5285
rect 3415 5215 3435 5235
rect 3415 5165 3435 5185
rect 3415 5115 3435 5135
rect 3415 5065 3435 5085
rect 3415 5015 3435 5035
rect 3565 5465 3585 5485
rect 3565 5415 3585 5435
rect 3565 5365 3585 5385
rect 3565 5315 3585 5335
rect 3565 5265 3585 5285
rect 3565 5215 3585 5235
rect 3565 5165 3585 5185
rect 3565 5115 3585 5135
rect 3565 5065 3585 5085
rect 3565 5015 3585 5035
rect 4165 5465 4185 5485
rect 4165 5415 4185 5435
rect 4165 5365 4185 5385
rect 4165 5315 4185 5335
rect 4165 5265 4185 5285
rect 4165 5215 4185 5235
rect 4165 5165 4185 5185
rect 4165 5115 4185 5135
rect 4765 5465 4785 5485
rect 4765 5415 4785 5435
rect 4765 5365 4785 5385
rect 4765 5315 4785 5335
rect 4765 5265 4785 5285
rect 4765 5215 4785 5235
rect 4765 5165 4785 5185
rect 4765 5115 4785 5135
rect 4765 5065 4785 5085
rect 4765 5015 4785 5035
rect 4915 5365 4935 5385
rect 4915 5315 4935 5335
rect 4915 5265 4935 5285
rect 4915 5215 4935 5235
rect 4915 5165 4935 5185
rect 4915 5115 4935 5135
rect 4915 5065 4935 5085
rect 4915 5015 4935 5035
rect 5065 5465 5085 5485
rect 5065 5415 5085 5435
rect 5065 5365 5085 5385
rect 5065 5315 5085 5335
rect 5065 5265 5085 5285
rect 5065 5215 5085 5235
rect 5065 5165 5085 5185
rect 5065 5115 5085 5135
rect 5215 5365 5235 5385
rect 5215 5315 5235 5335
rect 5215 5265 5235 5285
rect 5215 5215 5235 5235
rect 5215 5165 5235 5185
rect 5215 5115 5235 5135
rect 5215 5065 5235 5085
rect 5365 5465 5385 5485
rect 5365 5415 5385 5435
rect 5365 5365 5385 5385
rect 5365 5315 5385 5335
rect 5365 5265 5385 5285
rect 5365 5215 5385 5235
rect 5365 5165 5385 5185
rect 5365 5115 5385 5135
rect 5515 5365 5535 5385
rect 5515 5315 5535 5335
rect 5515 5265 5535 5285
rect 5515 5215 5535 5235
rect 5515 5165 5535 5185
rect 5515 5115 5535 5135
rect 5515 5065 5535 5085
rect 5665 5465 5685 5485
rect 5665 5415 5685 5435
rect 5665 5365 5685 5385
rect 5665 5315 5685 5335
rect 5665 5265 5685 5285
rect 5665 5215 5685 5235
rect 5665 5165 5685 5185
rect 5665 5115 5685 5135
rect 5815 5365 5835 5385
rect 5815 5315 5835 5335
rect 5815 5265 5835 5285
rect 5815 5215 5835 5235
rect 5815 5165 5835 5185
rect 5815 5115 5835 5135
rect 5815 5065 5835 5085
rect 5965 5465 5985 5485
rect 5965 5415 5985 5435
rect 5965 5365 5985 5385
rect 5965 5315 5985 5335
rect 5965 5265 5985 5285
rect 5965 5215 5985 5235
rect 5965 5165 5985 5185
rect 5965 5115 5985 5135
rect 5965 5065 5985 5085
rect 5965 5015 5985 5035
rect 6115 5365 6135 5385
rect 6115 5315 6135 5335
rect 6115 5265 6135 5285
rect 6115 5215 6135 5235
rect 6115 5165 6135 5185
rect 6115 5115 6135 5135
rect 6115 5065 6135 5085
rect 6115 5015 6135 5035
rect 6265 5465 6285 5485
rect 6265 5415 6285 5435
rect 6265 5365 6285 5385
rect 6265 5315 6285 5335
rect 6265 5265 6285 5285
rect 6265 5215 6285 5235
rect 6265 5165 6285 5185
rect 6265 5115 6285 5135
rect 6415 5365 6435 5385
rect 6415 5315 6435 5335
rect 6415 5265 6435 5285
rect 6415 5215 6435 5235
rect 6415 5165 6435 5185
rect 6415 5115 6435 5135
rect 6415 5065 6435 5085
rect 6415 5015 6435 5035
rect 6565 5465 6585 5485
rect 6565 5415 6585 5435
rect 6565 5365 6585 5385
rect 6565 5315 6585 5335
rect 6565 5265 6585 5285
rect 6565 5215 6585 5235
rect 6565 5165 6585 5185
rect 6565 5115 6585 5135
rect 6565 5065 6585 5085
rect 6565 5015 6585 5035
rect 6715 5365 6735 5385
rect 6715 5315 6735 5335
rect 6715 5265 6735 5285
rect 6715 5215 6735 5235
rect 6715 5165 6735 5185
rect 6715 5115 6735 5135
rect 6715 5065 6735 5085
rect 6865 5465 6885 5485
rect 6865 5415 6885 5435
rect 6865 5365 6885 5385
rect 6865 5315 6885 5335
rect 6865 5265 6885 5285
rect 6865 5215 6885 5235
rect 6865 5165 6885 5185
rect 6865 5115 6885 5135
rect 7015 5365 7035 5385
rect 7015 5315 7035 5335
rect 7015 5265 7035 5285
rect 7015 5215 7035 5235
rect 7015 5165 7035 5185
rect 7015 5115 7035 5135
rect 7015 5065 7035 5085
rect 7165 5465 7185 5485
rect 7165 5415 7185 5435
rect 7165 5365 7185 5385
rect 7165 5315 7185 5335
rect 7165 5265 7185 5285
rect 7165 5215 7185 5235
rect 7165 5165 7185 5185
rect 7165 5115 7185 5135
rect 7315 5365 7335 5385
rect 7315 5315 7335 5335
rect 7315 5265 7335 5285
rect 7315 5215 7335 5235
rect 7315 5165 7335 5185
rect 7315 5115 7335 5135
rect 7315 5065 7335 5085
rect 7465 5465 7485 5485
rect 7465 5415 7485 5435
rect 7465 5365 7485 5385
rect 7465 5315 7485 5335
rect 7465 5265 7485 5285
rect 7465 5215 7485 5235
rect 7465 5165 7485 5185
rect 7465 5115 7485 5135
rect 7615 5365 7635 5385
rect 7615 5315 7635 5335
rect 7615 5265 7635 5285
rect 7615 5215 7635 5235
rect 7615 5165 7635 5185
rect 7615 5115 7635 5135
rect 7615 5065 7635 5085
rect 7615 5015 7635 5035
rect 7765 5465 7785 5485
rect 7765 5415 7785 5435
rect 7765 5365 7785 5385
rect 7765 5315 7785 5335
rect 7765 5265 7785 5285
rect 7765 5215 7785 5235
rect 7765 5165 7785 5185
rect 7765 5115 7785 5135
rect 7765 5065 7785 5085
rect 7765 5015 7785 5035
rect 8365 5465 8385 5485
rect 8365 5415 8385 5435
rect 8365 5365 8385 5385
rect 8365 5315 8385 5335
rect 8365 5265 8385 5285
rect 8365 5215 8385 5235
rect 8365 5165 8385 5185
rect 8365 5115 8385 5135
rect 8365 5065 8385 5085
rect 8365 5015 8385 5035
rect 8515 5465 8535 5485
rect 8515 5415 8535 5435
rect 8515 5365 8535 5385
rect 8515 5315 8535 5335
rect 8515 5265 8535 5285
rect 8515 5215 8535 5235
rect 8515 5165 8535 5185
rect 8515 5115 8535 5135
rect 8515 5065 8535 5085
rect 8515 5015 8535 5035
rect 8665 5465 8685 5485
rect 8665 5415 8685 5435
rect 8665 5365 8685 5385
rect 8665 5315 8685 5335
rect 8665 5265 8685 5285
rect 8665 5215 8685 5235
rect 8665 5165 8685 5185
rect 8665 5115 8685 5135
rect 8665 5065 8685 5085
rect 8665 5015 8685 5035
rect 8815 5465 8835 5485
rect 8815 5415 8835 5435
rect 8815 5365 8835 5385
rect 8815 5315 8835 5335
rect 8815 5265 8835 5285
rect 8815 5215 8835 5235
rect 8815 5165 8835 5185
rect 8815 5115 8835 5135
rect 8815 5065 8835 5085
rect 8815 5015 8835 5035
rect 8965 5465 8985 5485
rect 8965 5415 8985 5435
rect 8965 5365 8985 5385
rect 8965 5315 8985 5335
rect 8965 5265 8985 5285
rect 8965 5215 8985 5235
rect 8965 5165 8985 5185
rect 8965 5115 8985 5135
rect 8965 5065 8985 5085
rect 8965 5015 8985 5035
rect 9115 5465 9135 5485
rect 9115 5415 9135 5435
rect 9115 5365 9135 5385
rect 9115 5315 9135 5335
rect 9115 5265 9135 5285
rect 9115 5215 9135 5235
rect 9115 5165 9135 5185
rect 9115 5115 9135 5135
rect 9115 5065 9135 5085
rect 9115 5015 9135 5035
rect 9265 5465 9285 5485
rect 9265 5415 9285 5435
rect 9265 5365 9285 5385
rect 9265 5315 9285 5335
rect 9265 5265 9285 5285
rect 9265 5215 9285 5235
rect 9265 5165 9285 5185
rect 9265 5115 9285 5135
rect 9265 5065 9285 5085
rect 9265 5015 9285 5035
rect 9415 5465 9435 5485
rect 9415 5415 9435 5435
rect 9415 5365 9435 5385
rect 9415 5315 9435 5335
rect 9415 5265 9435 5285
rect 9415 5215 9435 5235
rect 9415 5165 9435 5185
rect 9415 5115 9435 5135
rect 9415 5065 9435 5085
rect 9415 5015 9435 5035
rect 9565 5465 9585 5485
rect 9565 5415 9585 5435
rect 9565 5365 9585 5385
rect 9565 5315 9585 5335
rect 9565 5265 9585 5285
rect 9565 5215 9585 5235
rect 9565 5165 9585 5185
rect 9565 5115 9585 5135
rect 9565 5065 9585 5085
rect 9565 5015 9585 5035
rect 9715 5465 9735 5485
rect 9715 5415 9735 5435
rect 9715 5365 9735 5385
rect 9715 5315 9735 5335
rect 9715 5265 9735 5285
rect 9715 5215 9735 5235
rect 9715 5165 9735 5185
rect 9715 5115 9735 5135
rect 9715 5065 9735 5085
rect 9715 5015 9735 5035
rect 9865 5465 9885 5485
rect 9865 5415 9885 5435
rect 9865 5365 9885 5385
rect 9865 5315 9885 5335
rect 9865 5265 9885 5285
rect 9865 5215 9885 5235
rect 9865 5165 9885 5185
rect 9865 5115 9885 5135
rect 9865 5065 9885 5085
rect 9865 5015 9885 5035
rect 10015 5465 10035 5485
rect 10015 5415 10035 5435
rect 10015 5365 10035 5385
rect 10015 5315 10035 5335
rect 10015 5265 10035 5285
rect 10015 5215 10035 5235
rect 10015 5165 10035 5185
rect 10015 5115 10035 5135
rect 10015 5065 10035 5085
rect 10015 5015 10035 5035
rect 10165 5465 10185 5485
rect 10165 5415 10185 5435
rect 10165 5365 10185 5385
rect 10165 5315 10185 5335
rect 10165 5265 10185 5285
rect 10165 5215 10185 5235
rect 10165 5165 10185 5185
rect 10165 5115 10185 5135
rect 10165 5065 10185 5085
rect 10165 5015 10185 5035
rect 10315 5465 10335 5485
rect 10315 5415 10335 5435
rect 10315 5365 10335 5385
rect 10315 5315 10335 5335
rect 10315 5265 10335 5285
rect 10315 5215 10335 5235
rect 10315 5165 10335 5185
rect 10315 5115 10335 5135
rect 10315 5065 10335 5085
rect 10315 5015 10335 5035
rect 10465 5465 10485 5485
rect 10465 5415 10485 5435
rect 10465 5365 10485 5385
rect 10465 5315 10485 5335
rect 10465 5265 10485 5285
rect 10465 5215 10485 5235
rect 10465 5165 10485 5185
rect 10465 5115 10485 5135
rect 10465 5065 10485 5085
rect 10465 5015 10485 5035
rect 10615 5465 10635 5485
rect 10615 5415 10635 5435
rect 10615 5365 10635 5385
rect 10615 5315 10635 5335
rect 10615 5265 10635 5285
rect 10615 5215 10635 5235
rect 10615 5165 10635 5185
rect 10615 5115 10635 5135
rect 10615 5065 10635 5085
rect 10615 5015 10635 5035
rect 10765 5465 10785 5485
rect 10765 5415 10785 5435
rect 10765 5365 10785 5385
rect 10765 5315 10785 5335
rect 10765 5265 10785 5285
rect 10765 5215 10785 5235
rect 10765 5165 10785 5185
rect 10765 5115 10785 5135
rect 10765 5065 10785 5085
rect 10765 5015 10785 5035
rect 11365 5465 11385 5485
rect 11365 5415 11385 5435
rect 11365 5365 11385 5385
rect 11365 5315 11385 5335
rect 11365 5265 11385 5285
rect 11365 5215 11385 5235
rect 11365 5165 11385 5185
rect 11365 5115 11385 5135
rect 11365 5065 11385 5085
rect 11365 5015 11385 5035
rect 11965 5465 11985 5485
rect 11965 5415 11985 5435
rect 11965 5365 11985 5385
rect 11965 5315 11985 5335
rect 11965 5265 11985 5285
rect 11965 5215 11985 5235
rect 11965 5165 11985 5185
rect 11965 5115 11985 5135
rect 11965 5065 11985 5085
rect 11965 5015 11985 5035
rect 12565 5465 12585 5485
rect 12565 5415 12585 5435
rect 12565 5365 12585 5385
rect 12565 5315 12585 5335
rect 12565 5265 12585 5285
rect 12565 5215 12585 5235
rect 12565 5165 12585 5185
rect 12565 5115 12585 5135
rect 12565 5065 12585 5085
rect 12565 5015 12585 5035
rect 13165 5465 13185 5485
rect 13165 5415 13185 5435
rect 13165 5365 13185 5385
rect 13165 5315 13185 5335
rect 13165 5265 13185 5285
rect 13165 5215 13185 5235
rect 13165 5165 13185 5185
rect 13165 5115 13185 5135
rect 13165 5065 13185 5085
rect 13165 5015 13185 5035
rect 13765 5465 13785 5485
rect 13765 5415 13785 5435
rect 13765 5365 13785 5385
rect 13765 5315 13785 5335
rect 13765 5265 13785 5285
rect 13765 5215 13785 5235
rect 13765 5165 13785 5185
rect 13765 5115 13785 5135
rect 13765 5065 13785 5085
rect 13765 5015 13785 5035
rect 14365 5465 14385 5485
rect 14365 5415 14385 5435
rect 14365 5365 14385 5385
rect 14365 5315 14385 5335
rect 14365 5265 14385 5285
rect 14365 5215 14385 5235
rect 14365 5165 14385 5185
rect 14365 5115 14385 5135
rect 14365 5065 14385 5085
rect 14365 5015 14385 5035
rect 14965 5465 14985 5485
rect 14965 5415 14985 5435
rect 14965 5365 14985 5385
rect 14965 5315 14985 5335
rect 14965 5265 14985 5285
rect 14965 5215 14985 5235
rect 14965 5165 14985 5185
rect 14965 5115 14985 5135
rect 14965 5065 14985 5085
rect 14965 5015 14985 5035
rect 15565 5465 15585 5485
rect 15565 5415 15585 5435
rect 15565 5365 15585 5385
rect 15565 5315 15585 5335
rect 15565 5265 15585 5285
rect 15565 5215 15585 5235
rect 15565 5165 15585 5185
rect 15565 5115 15585 5135
rect 15565 5065 15585 5085
rect 15565 5015 15585 5035
rect 16165 5465 16185 5485
rect 16165 5415 16185 5435
rect 16165 5365 16185 5385
rect 16165 5315 16185 5335
rect 16165 5265 16185 5285
rect 16165 5215 16185 5235
rect 16165 5165 16185 5185
rect 16165 5115 16185 5135
rect 16165 5065 16185 5085
rect 16165 5015 16185 5035
rect 16315 5365 16335 5385
rect 16315 5315 16335 5335
rect 16315 5265 16335 5285
rect 16315 5215 16335 5235
rect 16315 5165 16335 5185
rect 16315 5115 16335 5135
rect 16315 5065 16335 5085
rect 16315 5015 16335 5035
rect 16465 5465 16485 5485
rect 16465 5415 16485 5435
rect 16465 5365 16485 5385
rect 16465 5315 16485 5335
rect 16465 5265 16485 5285
rect 16465 5215 16485 5235
rect 16465 5165 16485 5185
rect 16465 5115 16485 5135
rect 16615 5365 16635 5385
rect 16615 5315 16635 5335
rect 16615 5265 16635 5285
rect 16615 5215 16635 5235
rect 16615 5165 16635 5185
rect 16615 5115 16635 5135
rect 16615 5065 16635 5085
rect 16615 5015 16635 5035
rect 16765 5465 16785 5485
rect 16765 5415 16785 5435
rect 16765 5365 16785 5385
rect 16765 5315 16785 5335
rect 16765 5265 16785 5285
rect 16765 5215 16785 5235
rect 16765 5165 16785 5185
rect 16765 5115 16785 5135
rect 16915 5365 16935 5385
rect 16915 5315 16935 5335
rect 16915 5265 16935 5285
rect 16915 5215 16935 5235
rect 16915 5165 16935 5185
rect 16915 5115 16935 5135
rect 16915 5065 16935 5085
rect 16915 5015 16935 5035
rect 17065 5465 17085 5485
rect 17065 5415 17085 5435
rect 17065 5365 17085 5385
rect 17065 5315 17085 5335
rect 17065 5265 17085 5285
rect 17065 5215 17085 5235
rect 17065 5165 17085 5185
rect 17065 5115 17085 5135
rect 17215 5365 17235 5385
rect 17215 5315 17235 5335
rect 17215 5265 17235 5285
rect 17215 5215 17235 5235
rect 17215 5165 17235 5185
rect 17215 5115 17235 5135
rect 17215 5065 17235 5085
rect 17215 5015 17235 5035
rect 17365 5465 17385 5485
rect 17365 5415 17385 5435
rect 17365 5365 17385 5385
rect 17365 5315 17385 5335
rect 17365 5265 17385 5285
rect 17365 5215 17385 5235
rect 17365 5165 17385 5185
rect 17365 5115 17385 5135
rect 17365 5065 17385 5085
rect 17365 5015 17385 5035
rect 17965 5365 17985 5385
rect 17965 5315 17985 5335
rect 17965 5265 17985 5285
rect 17965 5215 17985 5235
rect 17965 5165 17985 5185
rect 17965 5115 17985 5135
rect 17965 5065 17985 5085
rect 17965 5015 17985 5035
rect 18565 5465 18585 5485
rect 18565 5415 18585 5435
rect 18565 5365 18585 5385
rect 18565 5315 18585 5335
rect 18565 5265 18585 5285
rect 18565 5215 18585 5235
rect 18565 5165 18585 5185
rect 18565 5115 18585 5135
rect 18565 5065 18585 5085
rect 18565 5015 18585 5035
rect 18715 5365 18735 5385
rect 18715 5315 18735 5335
rect 18715 5265 18735 5285
rect 18715 5215 18735 5235
rect 18715 5165 18735 5185
rect 18715 5115 18735 5135
rect 18715 5065 18735 5085
rect 18715 5015 18735 5035
rect 18865 5465 18885 5485
rect 18865 5415 18885 5435
rect 18865 5365 18885 5385
rect 18865 5315 18885 5335
rect 18865 5265 18885 5285
rect 18865 5215 18885 5235
rect 18865 5165 18885 5185
rect 18865 5115 18885 5135
rect 19015 5365 19035 5385
rect 19015 5315 19035 5335
rect 19015 5265 19035 5285
rect 19015 5215 19035 5235
rect 19015 5165 19035 5185
rect 19015 5115 19035 5135
rect 19015 5065 19035 5085
rect 19015 5015 19035 5035
rect 19165 5465 19185 5485
rect 19165 5415 19185 5435
rect 19165 5365 19185 5385
rect 19165 5315 19185 5335
rect 19165 5265 19185 5285
rect 19165 5215 19185 5235
rect 19165 5165 19185 5185
rect 19165 5115 19185 5135
rect 19315 5365 19335 5385
rect 19315 5315 19335 5335
rect 19315 5265 19335 5285
rect 19315 5215 19335 5235
rect 19315 5165 19335 5185
rect 19315 5115 19335 5135
rect 19315 5065 19335 5085
rect 19315 5015 19335 5035
rect 19465 5465 19485 5485
rect 19465 5415 19485 5435
rect 19465 5365 19485 5385
rect 19465 5315 19485 5335
rect 19465 5265 19485 5285
rect 19465 5215 19485 5235
rect 19465 5165 19485 5185
rect 19465 5115 19485 5135
rect 19615 5365 19635 5385
rect 19615 5315 19635 5335
rect 19615 5265 19635 5285
rect 19615 5215 19635 5235
rect 19615 5165 19635 5185
rect 19615 5115 19635 5135
rect 19615 5065 19635 5085
rect 19615 5015 19635 5035
rect 19765 5465 19785 5485
rect 19765 5415 19785 5435
rect 19765 5365 19785 5385
rect 19765 5315 19785 5335
rect 19765 5265 19785 5285
rect 19765 5215 19785 5235
rect 19765 5165 19785 5185
rect 19765 5115 19785 5135
rect 19765 5065 19785 5085
rect 19765 5015 19785 5035
rect 20365 5465 20385 5485
rect 20365 5415 20385 5435
rect 20365 5365 20385 5385
rect 20365 5315 20385 5335
rect 20365 5265 20385 5285
rect 20365 5215 20385 5235
rect 20365 5165 20385 5185
rect 20365 5115 20385 5135
rect 20365 5065 20385 5085
rect 20365 5015 20385 5035
rect 20965 5465 20985 5485
rect 20965 5415 20985 5435
rect 20965 5365 20985 5385
rect 20965 5315 20985 5335
rect 20965 5265 20985 5285
rect 20965 5215 20985 5235
rect 20965 5165 20985 5185
rect 20965 5115 20985 5135
rect 20965 5065 20985 5085
rect 20965 5015 20985 5035
rect 21415 5465 21435 5485
rect 21415 5415 21435 5435
rect 21415 5365 21435 5385
rect 21415 5315 21435 5335
rect 21415 5265 21435 5285
rect 21415 5215 21435 5235
rect 21415 5165 21435 5185
rect 21415 5115 21435 5135
rect 21415 5065 21435 5085
rect 21415 5015 21435 5035
rect 21865 5465 21885 5485
rect 21865 5415 21885 5435
rect 21865 5365 21885 5385
rect 21865 5315 21885 5335
rect 21865 5265 21885 5285
rect 21865 5215 21885 5235
rect 21865 5165 21885 5185
rect 21865 5115 21885 5135
rect 21865 5065 21885 5085
rect 21865 5015 21885 5035
rect 22465 5465 22485 5485
rect 22465 5415 22485 5435
rect 22465 5365 22485 5385
rect 22465 5315 22485 5335
rect 22465 5265 22485 5285
rect 22465 5215 22485 5235
rect 22465 5165 22485 5185
rect 22465 5115 22485 5135
rect 22465 5065 22485 5085
rect 22465 5015 22485 5035
rect 23065 5465 23085 5485
rect 23065 5415 23085 5435
rect 23065 5365 23085 5385
rect 23065 5315 23085 5335
rect 23065 5265 23085 5285
rect 23065 5215 23085 5235
rect 23065 5165 23085 5185
rect 23065 5115 23085 5135
rect 23065 5065 23085 5085
rect 23065 5015 23085 5035
rect 23515 5465 23535 5485
rect 23515 5415 23535 5435
rect 23515 5365 23535 5385
rect 23515 5315 23535 5335
rect 23515 5265 23535 5285
rect 23515 5215 23535 5235
rect 23515 5165 23535 5185
rect 23515 5115 23535 5135
rect 23515 5065 23535 5085
rect 23515 5015 23535 5035
rect 23965 5465 23985 5485
rect 23965 5415 23985 5435
rect 23965 5365 23985 5385
rect 23965 5315 23985 5335
rect 23965 5265 23985 5285
rect 23965 5215 23985 5235
rect 23965 5165 23985 5185
rect 23965 5115 23985 5135
rect 23965 5065 23985 5085
rect 23965 5015 23985 5035
rect 24565 5465 24585 5485
rect 24565 5415 24585 5435
rect 24565 5365 24585 5385
rect 24565 5315 24585 5335
rect 24565 5265 24585 5285
rect 24565 5215 24585 5235
rect 24565 5165 24585 5185
rect 24565 5115 24585 5135
rect 24565 5065 24585 5085
rect 24565 5015 24585 5035
rect 25165 5465 25185 5485
rect 25165 5415 25185 5435
rect 25165 5365 25185 5385
rect 25165 5315 25185 5335
rect 25165 5265 25185 5285
rect 25165 5215 25185 5235
rect 25165 5165 25185 5185
rect 25165 5115 25185 5135
rect 25165 5065 25185 5085
rect 25165 5015 25185 5035
rect 25615 5465 25635 5485
rect 25615 5415 25635 5435
rect 25615 5365 25635 5385
rect 25615 5315 25635 5335
rect 25615 5265 25635 5285
rect 25615 5215 25635 5235
rect 25615 5165 25635 5185
rect 25615 5115 25635 5135
rect 25615 5065 25635 5085
rect 25615 5015 25635 5035
rect 26065 5465 26085 5485
rect 26065 5415 26085 5435
rect 26065 5365 26085 5385
rect 26065 5315 26085 5335
rect 26065 5265 26085 5285
rect 26065 5215 26085 5235
rect 26065 5165 26085 5185
rect 26065 5115 26085 5135
rect 26065 5065 26085 5085
rect 26065 5015 26085 5035
rect 26665 5465 26685 5485
rect 26665 5415 26685 5435
rect 26665 5365 26685 5385
rect 26665 5315 26685 5335
rect 26665 5265 26685 5285
rect 26665 5215 26685 5235
rect 26665 5165 26685 5185
rect 26665 5115 26685 5135
rect 26665 5065 26685 5085
rect 26665 5015 26685 5035
rect 27265 5465 27285 5485
rect 27265 5415 27285 5435
rect 27265 5365 27285 5385
rect 27265 5315 27285 5335
rect 27265 5265 27285 5285
rect 27265 5215 27285 5235
rect 27265 5165 27285 5185
rect 27265 5115 27285 5135
rect 27265 5065 27285 5085
rect 27265 5015 27285 5035
rect 27715 5465 27735 5485
rect 27715 5415 27735 5435
rect 27715 5365 27735 5385
rect 27715 5315 27735 5335
rect 27715 5265 27735 5285
rect 27715 5215 27735 5235
rect 27715 5165 27735 5185
rect 27715 5115 27735 5135
rect 27715 5065 27735 5085
rect 27715 5015 27735 5035
rect 28165 5465 28185 5485
rect 28165 5415 28185 5435
rect 28165 5365 28185 5385
rect 28165 5315 28185 5335
rect 28165 5265 28185 5285
rect 28165 5215 28185 5235
rect 28165 5165 28185 5185
rect 28165 5115 28185 5135
rect 28165 5065 28185 5085
rect 28165 5015 28185 5035
rect 28765 5465 28785 5485
rect 28765 5415 28785 5435
rect 28765 5365 28785 5385
rect 28765 5315 28785 5335
rect 28765 5265 28785 5285
rect 28765 5215 28785 5235
rect 28765 5165 28785 5185
rect 28765 5115 28785 5135
rect 28765 5065 28785 5085
rect 28765 5015 28785 5035
rect 29365 5465 29385 5485
rect 29365 5415 29385 5435
rect 29365 5365 29385 5385
rect 29365 5315 29385 5335
rect 29365 5265 29385 5285
rect 29365 5215 29385 5235
rect 29365 5165 29385 5185
rect 29365 5115 29385 5135
rect 29365 5065 29385 5085
rect 29365 5015 29385 5035
rect 29515 5365 29535 5385
rect 29515 5315 29535 5335
rect 29515 5265 29535 5285
rect 29515 5215 29535 5235
rect 29515 5165 29535 5185
rect 29515 5115 29535 5135
rect 29515 5065 29535 5085
rect 29515 5015 29535 5035
rect 29665 5465 29685 5485
rect 29665 5415 29685 5435
rect 29665 5365 29685 5385
rect 29665 5315 29685 5335
rect 29665 5265 29685 5285
rect 29665 5215 29685 5235
rect 29665 5165 29685 5185
rect 29665 5115 29685 5135
rect 29815 5465 29835 5485
rect 29815 5415 29835 5435
rect 29815 5365 29835 5385
rect 29815 5315 29835 5335
rect 29815 5265 29835 5285
rect 29815 5215 29835 5235
rect 29815 5165 29835 5185
rect 29815 5115 29835 5135
rect 29815 5065 29835 5085
rect 29815 5015 29835 5035
rect 29965 5465 29985 5485
rect 29965 5415 29985 5435
rect 29965 5365 29985 5385
rect 29965 5315 29985 5335
rect 29965 5265 29985 5285
rect 29965 5215 29985 5235
rect 29965 5165 29985 5185
rect 29965 5115 29985 5135
rect 30115 5365 30135 5385
rect 30115 5315 30135 5335
rect 30115 5265 30135 5285
rect 30115 5215 30135 5235
rect 30115 5165 30135 5185
rect 30115 5115 30135 5135
rect 30115 5065 30135 5085
rect 30115 5015 30135 5035
rect 30265 5465 30285 5485
rect 30265 5415 30285 5435
rect 30265 5365 30285 5385
rect 30265 5315 30285 5335
rect 30265 5265 30285 5285
rect 30265 5215 30285 5235
rect 30265 5165 30285 5185
rect 30265 5115 30285 5135
rect 30415 5465 30435 5485
rect 30415 5415 30435 5435
rect 30415 5365 30435 5385
rect 30415 5315 30435 5335
rect 30415 5265 30435 5285
rect 30415 5215 30435 5235
rect 30415 5165 30435 5185
rect 30415 5115 30435 5135
rect 30415 5065 30435 5085
rect 30415 5015 30435 5035
rect 30565 5465 30585 5485
rect 30565 5415 30585 5435
rect 30565 5365 30585 5385
rect 30565 5315 30585 5335
rect 30565 5265 30585 5285
rect 30565 5215 30585 5235
rect 30565 5165 30585 5185
rect 30565 5115 30585 5135
rect 30715 5365 30735 5385
rect 30715 5315 30735 5335
rect 30715 5265 30735 5285
rect 30715 5215 30735 5235
rect 30715 5165 30735 5185
rect 30715 5115 30735 5135
rect 30715 5065 30735 5085
rect 30715 5015 30735 5035
rect 30865 5465 30885 5485
rect 30865 5415 30885 5435
rect 30865 5365 30885 5385
rect 30865 5315 30885 5335
rect 30865 5265 30885 5285
rect 30865 5215 30885 5235
rect 30865 5165 30885 5185
rect 30865 5115 30885 5135
rect 31015 5465 31035 5485
rect 31015 5415 31035 5435
rect 31015 5365 31035 5385
rect 31015 5315 31035 5335
rect 31015 5265 31035 5285
rect 31015 5215 31035 5235
rect 31015 5165 31035 5185
rect 31015 5115 31035 5135
rect 31015 5065 31035 5085
rect 31015 5015 31035 5035
rect 31165 5465 31185 5485
rect 31165 5415 31185 5435
rect 31165 5365 31185 5385
rect 31165 5315 31185 5335
rect 31165 5265 31185 5285
rect 31165 5215 31185 5235
rect 31165 5165 31185 5185
rect 31165 5115 31185 5135
rect 31315 5365 31335 5385
rect 31315 5315 31335 5335
rect 31315 5265 31335 5285
rect 31315 5215 31335 5235
rect 31315 5165 31335 5185
rect 31315 5115 31335 5135
rect 31315 5065 31335 5085
rect 31315 5015 31335 5035
rect 31465 5465 31485 5485
rect 31465 5415 31485 5435
rect 31465 5365 31485 5385
rect 31465 5315 31485 5335
rect 31465 5265 31485 5285
rect 31465 5215 31485 5235
rect 31465 5165 31485 5185
rect 31465 5115 31485 5135
rect 31465 5065 31485 5085
rect 31465 5015 31485 5035
rect 32065 5465 32085 5485
rect 32065 5415 32085 5435
rect 32065 5365 32085 5385
rect 32065 5315 32085 5335
rect 32065 5265 32085 5285
rect 32065 5215 32085 5235
rect 32065 5165 32085 5185
rect 32065 5115 32085 5135
rect 32065 5065 32085 5085
rect 32065 5015 32085 5035
rect -485 4915 -465 4935
rect -185 4915 -165 4935
rect 115 4915 135 4935
rect 415 4915 435 4935
rect 715 4915 735 4935
rect 1015 4915 1035 4935
rect 1315 4915 1335 4935
rect 1615 4915 1635 4935
rect 1915 4915 1935 4935
rect 2215 4915 2235 4935
rect 2515 4915 2535 4935
rect 2815 4915 2835 4935
rect 3115 4915 3135 4935
rect 3415 4915 3435 4935
rect 3715 4915 3735 4935
rect 4015 4915 4035 4935
rect 4315 4915 4335 4935
rect 4615 4915 4635 4935
rect 4915 4915 4935 4935
rect 5215 4915 5235 4935
rect 5515 4915 5535 4935
rect 5815 4915 5835 4935
rect 6115 4915 6135 4935
rect 6415 4915 6435 4935
rect 6715 4915 6735 4935
rect 7015 4915 7035 4935
rect 7315 4915 7335 4935
rect 7615 4915 7635 4935
rect 7915 4915 7935 4935
rect 8215 4915 8235 4935
rect 8515 4915 8535 4935
rect 8815 4915 8835 4935
rect 9115 4915 9135 4935
rect 9415 4915 9435 4935
rect 9715 4915 9735 4935
rect 10015 4915 10035 4935
rect 10315 4915 10335 4935
rect 10615 4915 10635 4935
rect 10915 4915 10935 4935
rect 11215 4915 11235 4935
rect 11515 4915 11535 4935
rect 11815 4915 11835 4935
rect 12115 4915 12135 4935
rect 12415 4915 12435 4935
rect 12715 4915 12735 4935
rect 13015 4915 13035 4935
rect 13315 4915 13335 4935
rect 13615 4915 13635 4935
rect 13915 4915 13935 4935
rect 14215 4915 14235 4935
rect 14515 4915 14535 4935
rect 14815 4915 14835 4935
rect 15115 4915 15135 4935
rect 15415 4915 15435 4935
rect 15715 4915 15735 4935
rect 16015 4915 16035 4935
rect 16315 4915 16335 4935
rect 16615 4915 16635 4935
rect 16915 4915 16935 4935
rect 17215 4915 17235 4935
rect 17515 4915 17535 4935
rect 17815 4915 17835 4935
rect 18115 4915 18135 4935
rect 18415 4915 18435 4935
rect 18715 4915 18735 4935
rect 19015 4915 19035 4935
rect 19315 4915 19335 4935
rect 19615 4915 19635 4935
rect 19915 4915 19935 4935
rect 20215 4915 20235 4935
rect 20515 4915 20535 4935
rect 20815 4915 20835 4935
rect 21115 4915 21135 4935
rect 21715 4915 21735 4935
rect 22015 4915 22035 4935
rect 22315 4915 22335 4935
rect 22615 4915 22635 4935
rect 22915 4915 22935 4935
rect 23215 4915 23235 4935
rect 23365 4915 23385 4935
rect 23665 4915 23685 4935
rect 23815 4915 23835 4935
rect 24115 4915 24135 4935
rect 24415 4915 24435 4935
rect 24715 4915 24735 4935
rect 25015 4915 25035 4935
rect 25465 4915 25485 4935
rect 25765 4915 25785 4935
rect 26215 4915 26235 4935
rect 26515 4915 26535 4935
rect 26815 4915 26835 4935
rect 27115 4915 27135 4935
rect 27565 4915 27585 4935
rect 27865 4915 27885 4935
rect 28315 4915 28335 4935
rect 28615 4915 28635 4935
rect 28915 4915 28935 4935
rect 29215 4915 29235 4935
rect 29665 4915 29685 4935
rect 29965 4915 29985 4935
rect 30265 4915 30285 4935
rect 30565 4915 30585 4935
rect 30865 4915 30885 4935
rect 31165 4915 31185 4935
rect 31615 4915 31635 4935
rect 31915 4915 31935 4935
rect -635 4815 -615 4835
rect -635 4765 -615 4785
rect -635 4715 -615 4735
rect -635 4665 -615 4685
rect -635 4615 -615 4635
rect -635 4565 -615 4585
rect -635 4515 -615 4535
rect -635 4465 -615 4485
rect -635 4415 -615 4435
rect -635 4365 -615 4385
rect -485 4815 -465 4835
rect -485 4765 -465 4785
rect -485 4715 -465 4735
rect -485 4665 -465 4685
rect -485 4615 -465 4635
rect -485 4565 -465 4585
rect -485 4515 -465 4535
rect -485 4465 -465 4485
rect -485 4415 -465 4435
rect -485 4365 -465 4385
rect -335 4715 -315 4735
rect -335 4665 -315 4685
rect -335 4615 -315 4635
rect -335 4565 -315 4585
rect -335 4515 -315 4535
rect -335 4465 -315 4485
rect -335 4415 -315 4435
rect -335 4365 -315 4385
rect -185 4815 -165 4835
rect -185 4765 -165 4785
rect -185 4715 -165 4735
rect -185 4665 -165 4685
rect -185 4615 -165 4635
rect -185 4565 -165 4585
rect -185 4515 -165 4535
rect -185 4465 -165 4485
rect -185 4415 -165 4435
rect -185 4365 -165 4385
rect -35 4715 -15 4735
rect -35 4665 -15 4685
rect -35 4615 -15 4635
rect -35 4565 -15 4585
rect -35 4515 -15 4535
rect -35 4465 -15 4485
rect -35 4415 -15 4435
rect -35 4365 -15 4385
rect 565 4815 585 4835
rect 565 4765 585 4785
rect 565 4715 585 4735
rect 565 4665 585 4685
rect 565 4615 585 4635
rect 565 4565 585 4585
rect 565 4515 585 4535
rect 565 4465 585 4485
rect 565 4415 585 4435
rect 565 4365 585 4385
rect 715 4815 735 4835
rect 715 4765 735 4785
rect 715 4715 735 4735
rect 715 4665 735 4685
rect 715 4615 735 4635
rect 715 4565 735 4585
rect 715 4515 735 4535
rect 715 4465 735 4485
rect 865 4715 885 4735
rect 865 4665 885 4685
rect 865 4615 885 4635
rect 865 4565 885 4585
rect 865 4515 885 4535
rect 865 4465 885 4485
rect 865 4415 885 4435
rect 865 4365 885 4385
rect 1015 4765 1035 4785
rect 1015 4715 1035 4735
rect 1015 4665 1035 4685
rect 1015 4615 1035 4635
rect 1015 4565 1035 4585
rect 1015 4515 1035 4535
rect 1015 4465 1035 4485
rect 1165 4715 1185 4735
rect 1165 4665 1185 4685
rect 1165 4615 1185 4635
rect 1165 4565 1185 4585
rect 1165 4515 1185 4535
rect 1165 4465 1185 4485
rect 1165 4415 1185 4435
rect 1165 4365 1185 4385
rect 1315 4765 1335 4785
rect 1315 4715 1335 4735
rect 1315 4665 1335 4685
rect 1315 4615 1335 4635
rect 1315 4565 1335 4585
rect 1315 4515 1335 4535
rect 1315 4465 1335 4485
rect 1465 4715 1485 4735
rect 1465 4665 1485 4685
rect 1465 4615 1485 4635
rect 1465 4565 1485 4585
rect 1465 4515 1485 4535
rect 1465 4465 1485 4485
rect 1465 4415 1485 4435
rect 1465 4365 1485 4385
rect 1615 4765 1635 4785
rect 1615 4715 1635 4735
rect 1615 4665 1635 4685
rect 1615 4615 1635 4635
rect 1615 4565 1635 4585
rect 1615 4515 1635 4535
rect 1615 4465 1635 4485
rect 1765 4815 1785 4835
rect 1765 4765 1785 4785
rect 1765 4715 1785 4735
rect 1765 4665 1785 4685
rect 1765 4615 1785 4635
rect 1765 4565 1785 4585
rect 1765 4515 1785 4535
rect 1765 4465 1785 4485
rect 1765 4415 1785 4435
rect 1765 4365 1785 4385
rect 1915 4815 1935 4835
rect 1915 4765 1935 4785
rect 1915 4715 1935 4735
rect 1915 4665 1935 4685
rect 1915 4615 1935 4635
rect 1915 4565 1935 4585
rect 1915 4515 1935 4535
rect 1915 4465 1935 4485
rect 2065 4715 2085 4735
rect 2065 4665 2085 4685
rect 2065 4615 2085 4635
rect 2065 4565 2085 4585
rect 2065 4515 2085 4535
rect 2065 4465 2085 4485
rect 2065 4415 2085 4435
rect 2065 4365 2085 4385
rect 2215 4815 2235 4835
rect 2215 4765 2235 4785
rect 2215 4715 2235 4735
rect 2215 4665 2235 4685
rect 2215 4615 2235 4635
rect 2215 4565 2235 4585
rect 2215 4515 2235 4535
rect 2215 4465 2235 4485
rect 2365 4815 2385 4835
rect 2365 4765 2385 4785
rect 2365 4715 2385 4735
rect 2365 4665 2385 4685
rect 2365 4615 2385 4635
rect 2365 4565 2385 4585
rect 2365 4515 2385 4535
rect 2365 4465 2385 4485
rect 2365 4415 2385 4435
rect 2365 4365 2385 4385
rect 2515 4765 2535 4785
rect 2515 4715 2535 4735
rect 2515 4665 2535 4685
rect 2515 4615 2535 4635
rect 2515 4565 2535 4585
rect 2515 4515 2535 4535
rect 2515 4465 2535 4485
rect 2665 4715 2685 4735
rect 2665 4665 2685 4685
rect 2665 4615 2685 4635
rect 2665 4565 2685 4585
rect 2665 4515 2685 4535
rect 2665 4465 2685 4485
rect 2665 4415 2685 4435
rect 2665 4365 2685 4385
rect 2815 4765 2835 4785
rect 2815 4715 2835 4735
rect 2815 4665 2835 4685
rect 2815 4615 2835 4635
rect 2815 4565 2835 4585
rect 2815 4515 2835 4535
rect 2815 4465 2835 4485
rect 2965 4715 2985 4735
rect 2965 4665 2985 4685
rect 2965 4615 2985 4635
rect 2965 4565 2985 4585
rect 2965 4515 2985 4535
rect 2965 4465 2985 4485
rect 2965 4415 2985 4435
rect 2965 4365 2985 4385
rect 3115 4765 3135 4785
rect 3115 4715 3135 4735
rect 3115 4665 3135 4685
rect 3115 4615 3135 4635
rect 3115 4565 3135 4585
rect 3115 4515 3135 4535
rect 3115 4465 3135 4485
rect 3265 4715 3285 4735
rect 3265 4665 3285 4685
rect 3265 4615 3285 4635
rect 3265 4565 3285 4585
rect 3265 4515 3285 4535
rect 3265 4465 3285 4485
rect 3265 4415 3285 4435
rect 3265 4365 3285 4385
rect 3415 4815 3435 4835
rect 3415 4765 3435 4785
rect 3415 4715 3435 4735
rect 3415 4665 3435 4685
rect 3415 4615 3435 4635
rect 3415 4565 3435 4585
rect 3415 4515 3435 4535
rect 3415 4465 3435 4485
rect 3565 4815 3585 4835
rect 3565 4765 3585 4785
rect 3565 4715 3585 4735
rect 3565 4665 3585 4685
rect 3565 4615 3585 4635
rect 3565 4565 3585 4585
rect 3565 4515 3585 4535
rect 3565 4465 3585 4485
rect 3565 4415 3585 4435
rect 3565 4365 3585 4385
rect 4165 4715 4185 4735
rect 4165 4665 4185 4685
rect 4165 4615 4185 4635
rect 4165 4565 4185 4585
rect 4165 4515 4185 4535
rect 4165 4465 4185 4485
rect 4165 4415 4185 4435
rect 4165 4365 4185 4385
rect 4765 4815 4785 4835
rect 4765 4765 4785 4785
rect 4765 4715 4785 4735
rect 4765 4665 4785 4685
rect 4765 4615 4785 4635
rect 4765 4565 4785 4585
rect 4765 4515 4785 4535
rect 4765 4465 4785 4485
rect 4765 4415 4785 4435
rect 4765 4365 4785 4385
rect 4915 4815 4935 4835
rect 4915 4765 4935 4785
rect 4915 4715 4935 4735
rect 4915 4665 4935 4685
rect 4915 4615 4935 4635
rect 4915 4565 4935 4585
rect 4915 4515 4935 4535
rect 4915 4465 4935 4485
rect 5065 4715 5085 4735
rect 5065 4665 5085 4685
rect 5065 4615 5085 4635
rect 5065 4565 5085 4585
rect 5065 4515 5085 4535
rect 5065 4465 5085 4485
rect 5065 4415 5085 4435
rect 5065 4365 5085 4385
rect 5215 4765 5235 4785
rect 5215 4715 5235 4735
rect 5215 4665 5235 4685
rect 5215 4615 5235 4635
rect 5215 4565 5235 4585
rect 5215 4515 5235 4535
rect 5215 4465 5235 4485
rect 5365 4715 5385 4735
rect 5365 4665 5385 4685
rect 5365 4615 5385 4635
rect 5365 4565 5385 4585
rect 5365 4515 5385 4535
rect 5365 4465 5385 4485
rect 5365 4415 5385 4435
rect 5365 4365 5385 4385
rect 5515 4765 5535 4785
rect 5515 4715 5535 4735
rect 5515 4665 5535 4685
rect 5515 4615 5535 4635
rect 5515 4565 5535 4585
rect 5515 4515 5535 4535
rect 5515 4465 5535 4485
rect 5665 4715 5685 4735
rect 5665 4665 5685 4685
rect 5665 4615 5685 4635
rect 5665 4565 5685 4585
rect 5665 4515 5685 4535
rect 5665 4465 5685 4485
rect 5665 4415 5685 4435
rect 5665 4365 5685 4385
rect 5815 4765 5835 4785
rect 5815 4715 5835 4735
rect 5815 4665 5835 4685
rect 5815 4615 5835 4635
rect 5815 4565 5835 4585
rect 5815 4515 5835 4535
rect 5815 4465 5835 4485
rect 5965 4815 5985 4835
rect 5965 4765 5985 4785
rect 5965 4715 5985 4735
rect 5965 4665 5985 4685
rect 5965 4615 5985 4635
rect 5965 4565 5985 4585
rect 5965 4515 5985 4535
rect 5965 4465 5985 4485
rect 5965 4415 5985 4435
rect 5965 4365 5985 4385
rect 6115 4815 6135 4835
rect 6115 4765 6135 4785
rect 6115 4715 6135 4735
rect 6115 4665 6135 4685
rect 6115 4615 6135 4635
rect 6115 4565 6135 4585
rect 6115 4515 6135 4535
rect 6115 4465 6135 4485
rect 6265 4715 6285 4735
rect 6265 4665 6285 4685
rect 6265 4615 6285 4635
rect 6265 4565 6285 4585
rect 6265 4515 6285 4535
rect 6265 4465 6285 4485
rect 6265 4415 6285 4435
rect 6265 4365 6285 4385
rect 6415 4815 6435 4835
rect 6415 4765 6435 4785
rect 6415 4715 6435 4735
rect 6415 4665 6435 4685
rect 6415 4615 6435 4635
rect 6415 4565 6435 4585
rect 6415 4515 6435 4535
rect 6415 4465 6435 4485
rect 6565 4815 6585 4835
rect 6565 4765 6585 4785
rect 6565 4715 6585 4735
rect 6565 4665 6585 4685
rect 6565 4615 6585 4635
rect 6565 4565 6585 4585
rect 6565 4515 6585 4535
rect 6565 4465 6585 4485
rect 6565 4415 6585 4435
rect 6565 4365 6585 4385
rect 6715 4765 6735 4785
rect 6715 4715 6735 4735
rect 6715 4665 6735 4685
rect 6715 4615 6735 4635
rect 6715 4565 6735 4585
rect 6715 4515 6735 4535
rect 6715 4465 6735 4485
rect 6865 4715 6885 4735
rect 6865 4665 6885 4685
rect 6865 4615 6885 4635
rect 6865 4565 6885 4585
rect 6865 4515 6885 4535
rect 6865 4465 6885 4485
rect 6865 4415 6885 4435
rect 6865 4365 6885 4385
rect 7015 4765 7035 4785
rect 7015 4715 7035 4735
rect 7015 4665 7035 4685
rect 7015 4615 7035 4635
rect 7015 4565 7035 4585
rect 7015 4515 7035 4535
rect 7015 4465 7035 4485
rect 7165 4715 7185 4735
rect 7165 4665 7185 4685
rect 7165 4615 7185 4635
rect 7165 4565 7185 4585
rect 7165 4515 7185 4535
rect 7165 4465 7185 4485
rect 7165 4415 7185 4435
rect 7165 4365 7185 4385
rect 7315 4765 7335 4785
rect 7315 4715 7335 4735
rect 7315 4665 7335 4685
rect 7315 4615 7335 4635
rect 7315 4565 7335 4585
rect 7315 4515 7335 4535
rect 7315 4465 7335 4485
rect 7465 4715 7485 4735
rect 7465 4665 7485 4685
rect 7465 4615 7485 4635
rect 7465 4565 7485 4585
rect 7465 4515 7485 4535
rect 7465 4465 7485 4485
rect 7465 4415 7485 4435
rect 7465 4365 7485 4385
rect 7615 4815 7635 4835
rect 7615 4765 7635 4785
rect 7615 4715 7635 4735
rect 7615 4665 7635 4685
rect 7615 4615 7635 4635
rect 7615 4565 7635 4585
rect 7615 4515 7635 4535
rect 7615 4465 7635 4485
rect 7765 4815 7785 4835
rect 7765 4765 7785 4785
rect 7765 4715 7785 4735
rect 7765 4665 7785 4685
rect 7765 4615 7785 4635
rect 7765 4565 7785 4585
rect 7765 4515 7785 4535
rect 7765 4465 7785 4485
rect 7765 4415 7785 4435
rect 7765 4365 7785 4385
rect 8365 4815 8385 4835
rect 8365 4765 8385 4785
rect 8365 4715 8385 4735
rect 8365 4665 8385 4685
rect 8365 4615 8385 4635
rect 8365 4565 8385 4585
rect 8365 4515 8385 4535
rect 8365 4465 8385 4485
rect 8365 4415 8385 4435
rect 8365 4365 8385 4385
rect 8515 4815 8535 4835
rect 8515 4765 8535 4785
rect 8515 4715 8535 4735
rect 8515 4665 8535 4685
rect 8515 4615 8535 4635
rect 8515 4565 8535 4585
rect 8515 4515 8535 4535
rect 8515 4465 8535 4485
rect 8515 4415 8535 4435
rect 8515 4365 8535 4385
rect 8665 4815 8685 4835
rect 8665 4765 8685 4785
rect 8665 4715 8685 4735
rect 8665 4665 8685 4685
rect 8665 4615 8685 4635
rect 8665 4565 8685 4585
rect 8665 4515 8685 4535
rect 8665 4465 8685 4485
rect 8665 4415 8685 4435
rect 8665 4365 8685 4385
rect 8815 4815 8835 4835
rect 8815 4765 8835 4785
rect 8815 4715 8835 4735
rect 8815 4665 8835 4685
rect 8815 4615 8835 4635
rect 8815 4565 8835 4585
rect 8815 4515 8835 4535
rect 8815 4465 8835 4485
rect 8815 4415 8835 4435
rect 8815 4365 8835 4385
rect 8965 4815 8985 4835
rect 8965 4765 8985 4785
rect 8965 4715 8985 4735
rect 8965 4665 8985 4685
rect 8965 4615 8985 4635
rect 8965 4565 8985 4585
rect 8965 4515 8985 4535
rect 8965 4465 8985 4485
rect 8965 4415 8985 4435
rect 8965 4365 8985 4385
rect 9115 4815 9135 4835
rect 9115 4765 9135 4785
rect 9115 4715 9135 4735
rect 9115 4665 9135 4685
rect 9115 4615 9135 4635
rect 9115 4565 9135 4585
rect 9115 4515 9135 4535
rect 9115 4465 9135 4485
rect 9115 4415 9135 4435
rect 9115 4365 9135 4385
rect 9265 4815 9285 4835
rect 9265 4765 9285 4785
rect 9265 4715 9285 4735
rect 9265 4665 9285 4685
rect 9265 4615 9285 4635
rect 9265 4565 9285 4585
rect 9265 4515 9285 4535
rect 9265 4465 9285 4485
rect 9265 4415 9285 4435
rect 9265 4365 9285 4385
rect 9415 4815 9435 4835
rect 9415 4765 9435 4785
rect 9415 4715 9435 4735
rect 9415 4665 9435 4685
rect 9415 4615 9435 4635
rect 9415 4565 9435 4585
rect 9415 4515 9435 4535
rect 9415 4465 9435 4485
rect 9415 4415 9435 4435
rect 9415 4365 9435 4385
rect 9565 4815 9585 4835
rect 9565 4765 9585 4785
rect 9565 4715 9585 4735
rect 9565 4665 9585 4685
rect 9565 4615 9585 4635
rect 9565 4565 9585 4585
rect 9565 4515 9585 4535
rect 9565 4465 9585 4485
rect 9565 4415 9585 4435
rect 9565 4365 9585 4385
rect 9715 4815 9735 4835
rect 9715 4765 9735 4785
rect 9715 4715 9735 4735
rect 9715 4665 9735 4685
rect 9715 4615 9735 4635
rect 9715 4565 9735 4585
rect 9715 4515 9735 4535
rect 9715 4465 9735 4485
rect 9715 4415 9735 4435
rect 9715 4365 9735 4385
rect 9865 4815 9885 4835
rect 9865 4765 9885 4785
rect 9865 4715 9885 4735
rect 9865 4665 9885 4685
rect 9865 4615 9885 4635
rect 9865 4565 9885 4585
rect 9865 4515 9885 4535
rect 9865 4465 9885 4485
rect 9865 4415 9885 4435
rect 9865 4365 9885 4385
rect 10015 4815 10035 4835
rect 10015 4765 10035 4785
rect 10015 4715 10035 4735
rect 10015 4665 10035 4685
rect 10015 4615 10035 4635
rect 10015 4565 10035 4585
rect 10015 4515 10035 4535
rect 10015 4465 10035 4485
rect 10015 4415 10035 4435
rect 10015 4365 10035 4385
rect 10165 4815 10185 4835
rect 10165 4765 10185 4785
rect 10165 4715 10185 4735
rect 10165 4665 10185 4685
rect 10165 4615 10185 4635
rect 10165 4565 10185 4585
rect 10165 4515 10185 4535
rect 10165 4465 10185 4485
rect 10165 4415 10185 4435
rect 10165 4365 10185 4385
rect 10315 4815 10335 4835
rect 10315 4765 10335 4785
rect 10315 4715 10335 4735
rect 10315 4665 10335 4685
rect 10315 4615 10335 4635
rect 10315 4565 10335 4585
rect 10315 4515 10335 4535
rect 10315 4465 10335 4485
rect 10315 4415 10335 4435
rect 10315 4365 10335 4385
rect 10465 4815 10485 4835
rect 10465 4765 10485 4785
rect 10465 4715 10485 4735
rect 10465 4665 10485 4685
rect 10465 4615 10485 4635
rect 10465 4565 10485 4585
rect 10465 4515 10485 4535
rect 10465 4465 10485 4485
rect 10465 4415 10485 4435
rect 10465 4365 10485 4385
rect 10615 4815 10635 4835
rect 10615 4765 10635 4785
rect 10615 4715 10635 4735
rect 10615 4665 10635 4685
rect 10615 4615 10635 4635
rect 10615 4565 10635 4585
rect 10615 4515 10635 4535
rect 10615 4465 10635 4485
rect 10615 4415 10635 4435
rect 10615 4365 10635 4385
rect 10765 4815 10785 4835
rect 10765 4765 10785 4785
rect 10765 4715 10785 4735
rect 10765 4665 10785 4685
rect 10765 4615 10785 4635
rect 10765 4565 10785 4585
rect 10765 4515 10785 4535
rect 10765 4465 10785 4485
rect 10765 4415 10785 4435
rect 10765 4365 10785 4385
rect 11365 4815 11385 4835
rect 11365 4765 11385 4785
rect 11365 4715 11385 4735
rect 11365 4665 11385 4685
rect 11365 4615 11385 4635
rect 11365 4565 11385 4585
rect 11365 4515 11385 4535
rect 11365 4465 11385 4485
rect 11365 4415 11385 4435
rect 11365 4365 11385 4385
rect 11965 4815 11985 4835
rect 11965 4765 11985 4785
rect 11965 4715 11985 4735
rect 11965 4665 11985 4685
rect 11965 4615 11985 4635
rect 11965 4565 11985 4585
rect 11965 4515 11985 4535
rect 11965 4465 11985 4485
rect 11965 4415 11985 4435
rect 11965 4365 11985 4385
rect 12565 4815 12585 4835
rect 12565 4765 12585 4785
rect 12565 4715 12585 4735
rect 12565 4665 12585 4685
rect 12565 4615 12585 4635
rect 12565 4565 12585 4585
rect 12565 4515 12585 4535
rect 12565 4465 12585 4485
rect 12565 4415 12585 4435
rect 12565 4365 12585 4385
rect 13165 4815 13185 4835
rect 13165 4765 13185 4785
rect 13165 4715 13185 4735
rect 13165 4665 13185 4685
rect 13165 4615 13185 4635
rect 13165 4565 13185 4585
rect 13165 4515 13185 4535
rect 13165 4465 13185 4485
rect 13165 4415 13185 4435
rect 13165 4365 13185 4385
rect 13765 4815 13785 4835
rect 13765 4765 13785 4785
rect 13765 4715 13785 4735
rect 13765 4665 13785 4685
rect 13765 4615 13785 4635
rect 13765 4565 13785 4585
rect 13765 4515 13785 4535
rect 13765 4465 13785 4485
rect 13765 4415 13785 4435
rect 13765 4365 13785 4385
rect 14365 4815 14385 4835
rect 14365 4765 14385 4785
rect 14365 4715 14385 4735
rect 14365 4665 14385 4685
rect 14365 4615 14385 4635
rect 14365 4565 14385 4585
rect 14365 4515 14385 4535
rect 14365 4465 14385 4485
rect 14365 4415 14385 4435
rect 14365 4365 14385 4385
rect 14965 4815 14985 4835
rect 14965 4765 14985 4785
rect 14965 4715 14985 4735
rect 14965 4665 14985 4685
rect 14965 4615 14985 4635
rect 14965 4565 14985 4585
rect 14965 4515 14985 4535
rect 14965 4465 14985 4485
rect 14965 4415 14985 4435
rect 14965 4365 14985 4385
rect 15565 4815 15585 4835
rect 15565 4765 15585 4785
rect 15565 4715 15585 4735
rect 15565 4665 15585 4685
rect 15565 4615 15585 4635
rect 15565 4565 15585 4585
rect 15565 4515 15585 4535
rect 15565 4465 15585 4485
rect 15565 4415 15585 4435
rect 15565 4365 15585 4385
rect 16165 4815 16185 4835
rect 16165 4765 16185 4785
rect 16165 4715 16185 4735
rect 16165 4665 16185 4685
rect 16165 4615 16185 4635
rect 16165 4565 16185 4585
rect 16165 4515 16185 4535
rect 16165 4465 16185 4485
rect 16165 4415 16185 4435
rect 16165 4365 16185 4385
rect 16315 4815 16335 4835
rect 16315 4765 16335 4785
rect 16315 4715 16335 4735
rect 16315 4665 16335 4685
rect 16315 4615 16335 4635
rect 16315 4565 16335 4585
rect 16315 4515 16335 4535
rect 16315 4465 16335 4485
rect 16465 4715 16485 4735
rect 16465 4665 16485 4685
rect 16465 4615 16485 4635
rect 16465 4565 16485 4585
rect 16465 4515 16485 4535
rect 16465 4465 16485 4485
rect 16465 4415 16485 4435
rect 16465 4365 16485 4385
rect 16615 4815 16635 4835
rect 16615 4765 16635 4785
rect 16615 4715 16635 4735
rect 16615 4665 16635 4685
rect 16615 4615 16635 4635
rect 16615 4565 16635 4585
rect 16615 4515 16635 4535
rect 16615 4465 16635 4485
rect 16765 4715 16785 4735
rect 16765 4665 16785 4685
rect 16765 4615 16785 4635
rect 16765 4565 16785 4585
rect 16765 4515 16785 4535
rect 16765 4465 16785 4485
rect 16765 4415 16785 4435
rect 16765 4365 16785 4385
rect 16915 4815 16935 4835
rect 16915 4765 16935 4785
rect 16915 4715 16935 4735
rect 16915 4665 16935 4685
rect 16915 4615 16935 4635
rect 16915 4565 16935 4585
rect 16915 4515 16935 4535
rect 16915 4465 16935 4485
rect 17065 4715 17085 4735
rect 17065 4665 17085 4685
rect 17065 4615 17085 4635
rect 17065 4565 17085 4585
rect 17065 4515 17085 4535
rect 17065 4465 17085 4485
rect 17065 4415 17085 4435
rect 17065 4365 17085 4385
rect 17215 4815 17235 4835
rect 17215 4765 17235 4785
rect 17215 4715 17235 4735
rect 17215 4665 17235 4685
rect 17215 4615 17235 4635
rect 17215 4565 17235 4585
rect 17215 4515 17235 4535
rect 17215 4465 17235 4485
rect 17365 4815 17385 4835
rect 17365 4765 17385 4785
rect 17365 4715 17385 4735
rect 17365 4665 17385 4685
rect 17365 4615 17385 4635
rect 17365 4565 17385 4585
rect 17365 4515 17385 4535
rect 17365 4465 17385 4485
rect 17365 4415 17385 4435
rect 17365 4365 17385 4385
rect 17965 4815 17985 4835
rect 17965 4765 17985 4785
rect 17965 4715 17985 4735
rect 17965 4665 17985 4685
rect 17965 4615 17985 4635
rect 17965 4565 17985 4585
rect 17965 4515 17985 4535
rect 17965 4465 17985 4485
rect 18565 4815 18585 4835
rect 18565 4765 18585 4785
rect 18565 4715 18585 4735
rect 18565 4665 18585 4685
rect 18565 4615 18585 4635
rect 18565 4565 18585 4585
rect 18565 4515 18585 4535
rect 18565 4465 18585 4485
rect 18565 4415 18585 4435
rect 18565 4365 18585 4385
rect 18715 4815 18735 4835
rect 18715 4765 18735 4785
rect 18715 4715 18735 4735
rect 18715 4665 18735 4685
rect 18715 4615 18735 4635
rect 18715 4565 18735 4585
rect 18715 4515 18735 4535
rect 18715 4465 18735 4485
rect 18865 4715 18885 4735
rect 18865 4665 18885 4685
rect 18865 4615 18885 4635
rect 18865 4565 18885 4585
rect 18865 4515 18885 4535
rect 18865 4465 18885 4485
rect 18865 4415 18885 4435
rect 18865 4365 18885 4385
rect 19015 4815 19035 4835
rect 19015 4765 19035 4785
rect 19015 4715 19035 4735
rect 19015 4665 19035 4685
rect 19015 4615 19035 4635
rect 19015 4565 19035 4585
rect 19015 4515 19035 4535
rect 19015 4465 19035 4485
rect 19165 4715 19185 4735
rect 19165 4665 19185 4685
rect 19165 4615 19185 4635
rect 19165 4565 19185 4585
rect 19165 4515 19185 4535
rect 19165 4465 19185 4485
rect 19165 4415 19185 4435
rect 19165 4365 19185 4385
rect 19315 4815 19335 4835
rect 19315 4765 19335 4785
rect 19315 4715 19335 4735
rect 19315 4665 19335 4685
rect 19315 4615 19335 4635
rect 19315 4565 19335 4585
rect 19315 4515 19335 4535
rect 19315 4465 19335 4485
rect 19465 4715 19485 4735
rect 19465 4665 19485 4685
rect 19465 4615 19485 4635
rect 19465 4565 19485 4585
rect 19465 4515 19485 4535
rect 19465 4465 19485 4485
rect 19465 4415 19485 4435
rect 19465 4365 19485 4385
rect 19615 4815 19635 4835
rect 19615 4765 19635 4785
rect 19615 4715 19635 4735
rect 19615 4665 19635 4685
rect 19615 4615 19635 4635
rect 19615 4565 19635 4585
rect 19615 4515 19635 4535
rect 19615 4465 19635 4485
rect 19765 4815 19785 4835
rect 19765 4765 19785 4785
rect 19765 4715 19785 4735
rect 19765 4665 19785 4685
rect 19765 4615 19785 4635
rect 19765 4565 19785 4585
rect 19765 4515 19785 4535
rect 19765 4465 19785 4485
rect 19765 4415 19785 4435
rect 19765 4365 19785 4385
rect 20365 4815 20385 4835
rect 20365 4765 20385 4785
rect 20365 4715 20385 4735
rect 20365 4665 20385 4685
rect 20365 4615 20385 4635
rect 20365 4565 20385 4585
rect 20365 4515 20385 4535
rect 20365 4465 20385 4485
rect 20365 4415 20385 4435
rect 20365 4365 20385 4385
rect 20965 4815 20985 4835
rect 20965 4765 20985 4785
rect 20965 4715 20985 4735
rect 20965 4665 20985 4685
rect 20965 4615 20985 4635
rect 20965 4565 20985 4585
rect 20965 4515 20985 4535
rect 20965 4465 20985 4485
rect 20965 4415 20985 4435
rect 20965 4365 20985 4385
rect 21415 4815 21435 4835
rect 21415 4765 21435 4785
rect 21415 4715 21435 4735
rect 21415 4665 21435 4685
rect 21415 4615 21435 4635
rect 21415 4565 21435 4585
rect 21415 4515 21435 4535
rect 21415 4465 21435 4485
rect 21415 4415 21435 4435
rect 21415 4365 21435 4385
rect 21865 4815 21885 4835
rect 21865 4765 21885 4785
rect 21865 4715 21885 4735
rect 21865 4665 21885 4685
rect 21865 4615 21885 4635
rect 21865 4565 21885 4585
rect 21865 4515 21885 4535
rect 21865 4465 21885 4485
rect 21865 4415 21885 4435
rect 21865 4365 21885 4385
rect 22465 4815 22485 4835
rect 22465 4765 22485 4785
rect 22465 4715 22485 4735
rect 22465 4665 22485 4685
rect 22465 4615 22485 4635
rect 22465 4565 22485 4585
rect 22465 4515 22485 4535
rect 22465 4465 22485 4485
rect 22465 4415 22485 4435
rect 22465 4365 22485 4385
rect 23065 4815 23085 4835
rect 23065 4765 23085 4785
rect 23065 4715 23085 4735
rect 23065 4665 23085 4685
rect 23065 4615 23085 4635
rect 23065 4565 23085 4585
rect 23065 4515 23085 4535
rect 23065 4465 23085 4485
rect 23065 4415 23085 4435
rect 23065 4365 23085 4385
rect 23515 4815 23535 4835
rect 23515 4765 23535 4785
rect 23515 4715 23535 4735
rect 23515 4665 23535 4685
rect 23515 4615 23535 4635
rect 23515 4565 23535 4585
rect 23515 4515 23535 4535
rect 23515 4465 23535 4485
rect 23515 4415 23535 4435
rect 23515 4365 23535 4385
rect 23965 4815 23985 4835
rect 23965 4765 23985 4785
rect 23965 4715 23985 4735
rect 23965 4665 23985 4685
rect 23965 4615 23985 4635
rect 23965 4565 23985 4585
rect 23965 4515 23985 4535
rect 23965 4465 23985 4485
rect 23965 4415 23985 4435
rect 23965 4365 23985 4385
rect 24565 4815 24585 4835
rect 24565 4765 24585 4785
rect 24565 4715 24585 4735
rect 24565 4665 24585 4685
rect 24565 4615 24585 4635
rect 24565 4565 24585 4585
rect 24565 4515 24585 4535
rect 24565 4465 24585 4485
rect 24565 4415 24585 4435
rect 24565 4365 24585 4385
rect 25165 4815 25185 4835
rect 25165 4765 25185 4785
rect 25165 4715 25185 4735
rect 25165 4665 25185 4685
rect 25165 4615 25185 4635
rect 25165 4565 25185 4585
rect 25165 4515 25185 4535
rect 25165 4465 25185 4485
rect 25165 4415 25185 4435
rect 25165 4365 25185 4385
rect 25615 4815 25635 4835
rect 25615 4765 25635 4785
rect 25615 4715 25635 4735
rect 25615 4665 25635 4685
rect 25615 4615 25635 4635
rect 25615 4565 25635 4585
rect 25615 4515 25635 4535
rect 25615 4465 25635 4485
rect 25615 4415 25635 4435
rect 25615 4365 25635 4385
rect 26065 4815 26085 4835
rect 26065 4765 26085 4785
rect 26065 4715 26085 4735
rect 26065 4665 26085 4685
rect 26065 4615 26085 4635
rect 26065 4565 26085 4585
rect 26065 4515 26085 4535
rect 26065 4465 26085 4485
rect 26065 4415 26085 4435
rect 26065 4365 26085 4385
rect 26665 4815 26685 4835
rect 26665 4765 26685 4785
rect 26665 4715 26685 4735
rect 26665 4665 26685 4685
rect 26665 4615 26685 4635
rect 26665 4565 26685 4585
rect 26665 4515 26685 4535
rect 26665 4465 26685 4485
rect 26665 4415 26685 4435
rect 26665 4365 26685 4385
rect 27265 4815 27285 4835
rect 27265 4765 27285 4785
rect 27265 4715 27285 4735
rect 27265 4665 27285 4685
rect 27265 4615 27285 4635
rect 27265 4565 27285 4585
rect 27265 4515 27285 4535
rect 27265 4465 27285 4485
rect 27265 4415 27285 4435
rect 27265 4365 27285 4385
rect 27715 4815 27735 4835
rect 27715 4765 27735 4785
rect 27715 4715 27735 4735
rect 27715 4665 27735 4685
rect 27715 4615 27735 4635
rect 27715 4565 27735 4585
rect 27715 4515 27735 4535
rect 27715 4465 27735 4485
rect 27715 4415 27735 4435
rect 27715 4365 27735 4385
rect 28165 4815 28185 4835
rect 28165 4765 28185 4785
rect 28165 4715 28185 4735
rect 28165 4665 28185 4685
rect 28165 4615 28185 4635
rect 28165 4565 28185 4585
rect 28165 4515 28185 4535
rect 28165 4465 28185 4485
rect 28165 4415 28185 4435
rect 28165 4365 28185 4385
rect 28765 4815 28785 4835
rect 28765 4765 28785 4785
rect 28765 4715 28785 4735
rect 28765 4665 28785 4685
rect 28765 4615 28785 4635
rect 28765 4565 28785 4585
rect 28765 4515 28785 4535
rect 28765 4465 28785 4485
rect 28765 4415 28785 4435
rect 28765 4365 28785 4385
rect 29365 4815 29385 4835
rect 29365 4765 29385 4785
rect 29365 4715 29385 4735
rect 29365 4665 29385 4685
rect 29365 4615 29385 4635
rect 29365 4565 29385 4585
rect 29365 4515 29385 4535
rect 29365 4465 29385 4485
rect 29365 4415 29385 4435
rect 29365 4365 29385 4385
rect 29515 4815 29535 4835
rect 29515 4765 29535 4785
rect 29515 4715 29535 4735
rect 29515 4665 29535 4685
rect 29515 4615 29535 4635
rect 29515 4565 29535 4585
rect 29515 4515 29535 4535
rect 29515 4465 29535 4485
rect 29665 4715 29685 4735
rect 29665 4665 29685 4685
rect 29665 4615 29685 4635
rect 29665 4565 29685 4585
rect 29665 4515 29685 4535
rect 29665 4465 29685 4485
rect 29665 4415 29685 4435
rect 29665 4365 29685 4385
rect 29815 4815 29835 4835
rect 29815 4765 29835 4785
rect 29815 4715 29835 4735
rect 29815 4665 29835 4685
rect 29815 4615 29835 4635
rect 29815 4565 29835 4585
rect 29815 4515 29835 4535
rect 29815 4465 29835 4485
rect 29815 4415 29835 4435
rect 29815 4365 29835 4385
rect 29965 4715 29985 4735
rect 29965 4665 29985 4685
rect 29965 4615 29985 4635
rect 29965 4565 29985 4585
rect 29965 4515 29985 4535
rect 29965 4465 29985 4485
rect 29965 4415 29985 4435
rect 29965 4365 29985 4385
rect 30115 4815 30135 4835
rect 30115 4765 30135 4785
rect 30115 4715 30135 4735
rect 30115 4665 30135 4685
rect 30115 4615 30135 4635
rect 30115 4565 30135 4585
rect 30115 4515 30135 4535
rect 30115 4465 30135 4485
rect 30265 4715 30285 4735
rect 30265 4665 30285 4685
rect 30265 4615 30285 4635
rect 30265 4565 30285 4585
rect 30265 4515 30285 4535
rect 30265 4465 30285 4485
rect 30265 4415 30285 4435
rect 30265 4365 30285 4385
rect 30415 4815 30435 4835
rect 30415 4765 30435 4785
rect 30415 4715 30435 4735
rect 30415 4665 30435 4685
rect 30415 4615 30435 4635
rect 30415 4565 30435 4585
rect 30415 4515 30435 4535
rect 30415 4465 30435 4485
rect 30415 4415 30435 4435
rect 30415 4365 30435 4385
rect 30565 4715 30585 4735
rect 30565 4665 30585 4685
rect 30565 4615 30585 4635
rect 30565 4565 30585 4585
rect 30565 4515 30585 4535
rect 30565 4465 30585 4485
rect 30565 4415 30585 4435
rect 30565 4365 30585 4385
rect 30715 4815 30735 4835
rect 30715 4765 30735 4785
rect 30715 4715 30735 4735
rect 30715 4665 30735 4685
rect 30715 4615 30735 4635
rect 30715 4565 30735 4585
rect 30715 4515 30735 4535
rect 30715 4465 30735 4485
rect 30865 4715 30885 4735
rect 30865 4665 30885 4685
rect 30865 4615 30885 4635
rect 30865 4565 30885 4585
rect 30865 4515 30885 4535
rect 30865 4465 30885 4485
rect 30865 4415 30885 4435
rect 30865 4365 30885 4385
rect 31015 4815 31035 4835
rect 31015 4765 31035 4785
rect 31015 4715 31035 4735
rect 31015 4665 31035 4685
rect 31015 4615 31035 4635
rect 31015 4565 31035 4585
rect 31015 4515 31035 4535
rect 31015 4465 31035 4485
rect 31015 4415 31035 4435
rect 31015 4365 31035 4385
rect 31165 4715 31185 4735
rect 31165 4665 31185 4685
rect 31165 4615 31185 4635
rect 31165 4565 31185 4585
rect 31165 4515 31185 4535
rect 31165 4465 31185 4485
rect 31165 4415 31185 4435
rect 31165 4365 31185 4385
rect 31315 4815 31335 4835
rect 31315 4765 31335 4785
rect 31315 4715 31335 4735
rect 31315 4665 31335 4685
rect 31315 4615 31335 4635
rect 31315 4565 31335 4585
rect 31315 4515 31335 4535
rect 31315 4465 31335 4485
rect 31465 4815 31485 4835
rect 31465 4765 31485 4785
rect 31465 4715 31485 4735
rect 31465 4665 31485 4685
rect 31465 4615 31485 4635
rect 31465 4565 31485 4585
rect 31465 4515 31485 4535
rect 31465 4465 31485 4485
rect 31465 4415 31485 4435
rect 31465 4365 31485 4385
rect 32065 4815 32085 4835
rect 32065 4765 32085 4785
rect 32065 4715 32085 4735
rect 32065 4665 32085 4685
rect 32065 4615 32085 4635
rect 32065 4565 32085 4585
rect 32065 4515 32085 4535
rect 32065 4465 32085 4485
rect 32065 4415 32085 4435
rect 32065 4365 32085 4385
rect -635 4265 -615 4285
rect -35 4265 -15 4285
rect 4165 4265 4185 4285
rect 8365 4265 8385 4285
rect 8665 4265 8685 4285
rect 8965 4265 8985 4285
rect 9265 4265 9285 4285
rect 9565 4265 9585 4285
rect 9865 4265 9885 4285
rect 10165 4265 10185 4285
rect 10465 4265 10485 4285
rect 10765 4265 10785 4285
rect 11965 4265 11985 4285
rect 13165 4265 13185 4285
rect 14365 4265 14385 4285
rect 15565 4265 15585 4285
rect 20365 4265 20385 4285
rect 22465 4265 22485 4285
rect 24565 4265 24585 4285
rect 26665 4265 26685 4285
rect 28165 4265 28185 4285
rect 28765 4265 28785 4285
rect 32065 4265 32085 4285
rect -635 4165 -615 4185
rect -635 4115 -615 4135
rect -635 4065 -615 4085
rect -635 4015 -615 4035
rect -635 3965 -615 3985
rect -635 3915 -615 3935
rect -635 3865 -615 3885
rect -635 3815 -615 3835
rect -635 3765 -615 3785
rect -635 3715 -615 3735
rect -485 4165 -465 4185
rect -485 4115 -465 4135
rect -485 4065 -465 4085
rect -485 4015 -465 4035
rect -485 3965 -465 3985
rect -485 3915 -465 3935
rect -485 3865 -465 3885
rect -485 3815 -465 3835
rect -485 3765 -465 3785
rect -485 3715 -465 3735
rect -335 4165 -315 4185
rect -335 4115 -315 4135
rect -335 4065 -315 4085
rect -335 4015 -315 4035
rect -335 3965 -315 3985
rect -335 3915 -315 3935
rect -335 3865 -315 3885
rect -335 3815 -315 3835
rect -185 4165 -165 4185
rect -185 4115 -165 4135
rect -185 4065 -165 4085
rect -185 4015 -165 4035
rect -185 3965 -165 3985
rect -185 3915 -165 3935
rect -185 3865 -165 3885
rect -185 3815 -165 3835
rect -185 3765 -165 3785
rect -185 3715 -165 3735
rect -35 4165 -15 4185
rect -35 4115 -15 4135
rect -35 4065 -15 4085
rect -35 4015 -15 4035
rect -35 3965 -15 3985
rect -35 3915 -15 3935
rect -35 3865 -15 3885
rect -35 3815 -15 3835
rect 565 4165 585 4185
rect 565 4115 585 4135
rect 565 4065 585 4085
rect 565 4015 585 4035
rect 565 3965 585 3985
rect 565 3915 585 3935
rect 565 3865 585 3885
rect 565 3815 585 3835
rect 565 3765 585 3785
rect 565 3715 585 3735
rect 715 4065 735 4085
rect 715 4015 735 4035
rect 715 3965 735 3985
rect 715 3915 735 3935
rect 715 3865 735 3885
rect 715 3815 735 3835
rect 715 3765 735 3785
rect 715 3715 735 3735
rect 865 4165 885 4185
rect 865 4115 885 4135
rect 865 4065 885 4085
rect 865 4015 885 4035
rect 865 3965 885 3985
rect 865 3915 885 3935
rect 865 3865 885 3885
rect 865 3815 885 3835
rect 1015 4065 1035 4085
rect 1015 4015 1035 4035
rect 1015 3965 1035 3985
rect 1015 3915 1035 3935
rect 1015 3865 1035 3885
rect 1015 3815 1035 3835
rect 1015 3765 1035 3785
rect 1165 4165 1185 4185
rect 1165 4115 1185 4135
rect 1165 4065 1185 4085
rect 1165 4015 1185 4035
rect 1165 3965 1185 3985
rect 1165 3915 1185 3935
rect 1165 3865 1185 3885
rect 1165 3815 1185 3835
rect 1315 4065 1335 4085
rect 1315 4015 1335 4035
rect 1315 3965 1335 3985
rect 1315 3915 1335 3935
rect 1315 3865 1335 3885
rect 1315 3815 1335 3835
rect 1315 3765 1335 3785
rect 1465 4165 1485 4185
rect 1465 4115 1485 4135
rect 1465 4065 1485 4085
rect 1465 4015 1485 4035
rect 1465 3965 1485 3985
rect 1465 3915 1485 3935
rect 1465 3865 1485 3885
rect 1465 3815 1485 3835
rect 1615 4065 1635 4085
rect 1615 4015 1635 4035
rect 1615 3965 1635 3985
rect 1615 3915 1635 3935
rect 1615 3865 1635 3885
rect 1615 3815 1635 3835
rect 1615 3765 1635 3785
rect 1765 4165 1785 4185
rect 1765 4115 1785 4135
rect 1765 4065 1785 4085
rect 1765 4015 1785 4035
rect 1765 3965 1785 3985
rect 1765 3915 1785 3935
rect 1765 3865 1785 3885
rect 1765 3815 1785 3835
rect 1765 3765 1785 3785
rect 1765 3715 1785 3735
rect 1915 4065 1935 4085
rect 1915 4015 1935 4035
rect 1915 3965 1935 3985
rect 1915 3915 1935 3935
rect 1915 3865 1935 3885
rect 1915 3815 1935 3835
rect 1915 3765 1935 3785
rect 1915 3715 1935 3735
rect 2065 4165 2085 4185
rect 2065 4115 2085 4135
rect 2065 4065 2085 4085
rect 2065 4015 2085 4035
rect 2065 3965 2085 3985
rect 2065 3915 2085 3935
rect 2065 3865 2085 3885
rect 2065 3815 2085 3835
rect 2215 4065 2235 4085
rect 2215 4015 2235 4035
rect 2215 3965 2235 3985
rect 2215 3915 2235 3935
rect 2215 3865 2235 3885
rect 2215 3815 2235 3835
rect 2215 3765 2235 3785
rect 2215 3715 2235 3735
rect 2365 4165 2385 4185
rect 2365 4115 2385 4135
rect 2365 4065 2385 4085
rect 2365 4015 2385 4035
rect 2365 3965 2385 3985
rect 2365 3915 2385 3935
rect 2365 3865 2385 3885
rect 2365 3815 2385 3835
rect 2365 3765 2385 3785
rect 2365 3715 2385 3735
rect 2515 4065 2535 4085
rect 2515 4015 2535 4035
rect 2515 3965 2535 3985
rect 2515 3915 2535 3935
rect 2515 3865 2535 3885
rect 2515 3815 2535 3835
rect 2515 3765 2535 3785
rect 2665 4165 2685 4185
rect 2665 4115 2685 4135
rect 2665 4065 2685 4085
rect 2665 4015 2685 4035
rect 2665 3965 2685 3985
rect 2665 3915 2685 3935
rect 2665 3865 2685 3885
rect 2665 3815 2685 3835
rect 2815 4065 2835 4085
rect 2815 4015 2835 4035
rect 2815 3965 2835 3985
rect 2815 3915 2835 3935
rect 2815 3865 2835 3885
rect 2815 3815 2835 3835
rect 2815 3765 2835 3785
rect 2965 4165 2985 4185
rect 2965 4115 2985 4135
rect 2965 4065 2985 4085
rect 2965 4015 2985 4035
rect 2965 3965 2985 3985
rect 2965 3915 2985 3935
rect 2965 3865 2985 3885
rect 2965 3815 2985 3835
rect 3115 4065 3135 4085
rect 3115 4015 3135 4035
rect 3115 3965 3135 3985
rect 3115 3915 3135 3935
rect 3115 3865 3135 3885
rect 3115 3815 3135 3835
rect 3115 3765 3135 3785
rect 3265 4165 3285 4185
rect 3265 4115 3285 4135
rect 3265 4065 3285 4085
rect 3265 4015 3285 4035
rect 3265 3965 3285 3985
rect 3265 3915 3285 3935
rect 3265 3865 3285 3885
rect 3265 3815 3285 3835
rect 3415 4065 3435 4085
rect 3415 4015 3435 4035
rect 3415 3965 3435 3985
rect 3415 3915 3435 3935
rect 3415 3865 3435 3885
rect 3415 3815 3435 3835
rect 3415 3765 3435 3785
rect 3415 3715 3435 3735
rect 3565 4165 3585 4185
rect 3565 4115 3585 4135
rect 3565 4065 3585 4085
rect 3565 4015 3585 4035
rect 3565 3965 3585 3985
rect 3565 3915 3585 3935
rect 3565 3865 3585 3885
rect 3565 3815 3585 3835
rect 3565 3765 3585 3785
rect 3565 3715 3585 3735
rect 4165 4165 4185 4185
rect 4165 4115 4185 4135
rect 4165 4065 4185 4085
rect 4165 4015 4185 4035
rect 4165 3965 4185 3985
rect 4165 3915 4185 3935
rect 4165 3865 4185 3885
rect 4165 3815 4185 3835
rect 4765 4165 4785 4185
rect 4765 4115 4785 4135
rect 4765 4065 4785 4085
rect 4765 4015 4785 4035
rect 4765 3965 4785 3985
rect 4765 3915 4785 3935
rect 4765 3865 4785 3885
rect 4765 3815 4785 3835
rect 4765 3765 4785 3785
rect 4765 3715 4785 3735
rect 4915 4065 4935 4085
rect 4915 4015 4935 4035
rect 4915 3965 4935 3985
rect 4915 3915 4935 3935
rect 4915 3865 4935 3885
rect 4915 3815 4935 3835
rect 4915 3765 4935 3785
rect 4915 3715 4935 3735
rect 5065 4165 5085 4185
rect 5065 4115 5085 4135
rect 5065 4065 5085 4085
rect 5065 4015 5085 4035
rect 5065 3965 5085 3985
rect 5065 3915 5085 3935
rect 5065 3865 5085 3885
rect 5065 3815 5085 3835
rect 5215 4065 5235 4085
rect 5215 4015 5235 4035
rect 5215 3965 5235 3985
rect 5215 3915 5235 3935
rect 5215 3865 5235 3885
rect 5215 3815 5235 3835
rect 5215 3765 5235 3785
rect 5365 4165 5385 4185
rect 5365 4115 5385 4135
rect 5365 4065 5385 4085
rect 5365 4015 5385 4035
rect 5365 3965 5385 3985
rect 5365 3915 5385 3935
rect 5365 3865 5385 3885
rect 5365 3815 5385 3835
rect 5515 4065 5535 4085
rect 5515 4015 5535 4035
rect 5515 3965 5535 3985
rect 5515 3915 5535 3935
rect 5515 3865 5535 3885
rect 5515 3815 5535 3835
rect 5515 3765 5535 3785
rect 5665 4165 5685 4185
rect 5665 4115 5685 4135
rect 5665 4065 5685 4085
rect 5665 4015 5685 4035
rect 5665 3965 5685 3985
rect 5665 3915 5685 3935
rect 5665 3865 5685 3885
rect 5665 3815 5685 3835
rect 5815 4065 5835 4085
rect 5815 4015 5835 4035
rect 5815 3965 5835 3985
rect 5815 3915 5835 3935
rect 5815 3865 5835 3885
rect 5815 3815 5835 3835
rect 5815 3765 5835 3785
rect 5965 4165 5985 4185
rect 5965 4115 5985 4135
rect 5965 4065 5985 4085
rect 5965 4015 5985 4035
rect 5965 3965 5985 3985
rect 5965 3915 5985 3935
rect 5965 3865 5985 3885
rect 5965 3815 5985 3835
rect 5965 3765 5985 3785
rect 5965 3715 5985 3735
rect 6115 4065 6135 4085
rect 6115 4015 6135 4035
rect 6115 3965 6135 3985
rect 6115 3915 6135 3935
rect 6115 3865 6135 3885
rect 6115 3815 6135 3835
rect 6115 3765 6135 3785
rect 6115 3715 6135 3735
rect 6265 4165 6285 4185
rect 6265 4115 6285 4135
rect 6265 4065 6285 4085
rect 6265 4015 6285 4035
rect 6265 3965 6285 3985
rect 6265 3915 6285 3935
rect 6265 3865 6285 3885
rect 6265 3815 6285 3835
rect 6415 4065 6435 4085
rect 6415 4015 6435 4035
rect 6415 3965 6435 3985
rect 6415 3915 6435 3935
rect 6415 3865 6435 3885
rect 6415 3815 6435 3835
rect 6415 3765 6435 3785
rect 6415 3715 6435 3735
rect 6565 4165 6585 4185
rect 6565 4115 6585 4135
rect 6565 4065 6585 4085
rect 6565 4015 6585 4035
rect 6565 3965 6585 3985
rect 6565 3915 6585 3935
rect 6565 3865 6585 3885
rect 6565 3815 6585 3835
rect 6565 3765 6585 3785
rect 6565 3715 6585 3735
rect 6715 4065 6735 4085
rect 6715 4015 6735 4035
rect 6715 3965 6735 3985
rect 6715 3915 6735 3935
rect 6715 3865 6735 3885
rect 6715 3815 6735 3835
rect 6715 3765 6735 3785
rect 6865 4165 6885 4185
rect 6865 4115 6885 4135
rect 6865 4065 6885 4085
rect 6865 4015 6885 4035
rect 6865 3965 6885 3985
rect 6865 3915 6885 3935
rect 6865 3865 6885 3885
rect 6865 3815 6885 3835
rect 7015 4065 7035 4085
rect 7015 4015 7035 4035
rect 7015 3965 7035 3985
rect 7015 3915 7035 3935
rect 7015 3865 7035 3885
rect 7015 3815 7035 3835
rect 7015 3765 7035 3785
rect 7165 4165 7185 4185
rect 7165 4115 7185 4135
rect 7165 4065 7185 4085
rect 7165 4015 7185 4035
rect 7165 3965 7185 3985
rect 7165 3915 7185 3935
rect 7165 3865 7185 3885
rect 7165 3815 7185 3835
rect 7315 4065 7335 4085
rect 7315 4015 7335 4035
rect 7315 3965 7335 3985
rect 7315 3915 7335 3935
rect 7315 3865 7335 3885
rect 7315 3815 7335 3835
rect 7315 3765 7335 3785
rect 7465 4165 7485 4185
rect 7465 4115 7485 4135
rect 7465 4065 7485 4085
rect 7465 4015 7485 4035
rect 7465 3965 7485 3985
rect 7465 3915 7485 3935
rect 7465 3865 7485 3885
rect 7465 3815 7485 3835
rect 7615 4065 7635 4085
rect 7615 4015 7635 4035
rect 7615 3965 7635 3985
rect 7615 3915 7635 3935
rect 7615 3865 7635 3885
rect 7615 3815 7635 3835
rect 7615 3765 7635 3785
rect 7615 3715 7635 3735
rect 7765 4165 7785 4185
rect 7765 4115 7785 4135
rect 7765 4065 7785 4085
rect 7765 4015 7785 4035
rect 7765 3965 7785 3985
rect 7765 3915 7785 3935
rect 7765 3865 7785 3885
rect 7765 3815 7785 3835
rect 7765 3765 7785 3785
rect 7765 3715 7785 3735
rect 8365 4165 8385 4185
rect 8365 4115 8385 4135
rect 8365 4065 8385 4085
rect 8365 4015 8385 4035
rect 8365 3965 8385 3985
rect 8365 3915 8385 3935
rect 8365 3865 8385 3885
rect 8365 3815 8385 3835
rect 8365 3765 8385 3785
rect 8365 3715 8385 3735
rect 8515 4165 8535 4185
rect 8515 4115 8535 4135
rect 8515 4065 8535 4085
rect 8515 4015 8535 4035
rect 8515 3965 8535 3985
rect 8515 3915 8535 3935
rect 8515 3865 8535 3885
rect 8515 3815 8535 3835
rect 8515 3765 8535 3785
rect 8515 3715 8535 3735
rect 8665 4165 8685 4185
rect 8665 4115 8685 4135
rect 8665 4065 8685 4085
rect 8665 4015 8685 4035
rect 8665 3965 8685 3985
rect 8665 3915 8685 3935
rect 8665 3865 8685 3885
rect 8665 3815 8685 3835
rect 8665 3765 8685 3785
rect 8665 3715 8685 3735
rect 8815 4165 8835 4185
rect 8815 4115 8835 4135
rect 8815 4065 8835 4085
rect 8815 4015 8835 4035
rect 8815 3965 8835 3985
rect 8815 3915 8835 3935
rect 8815 3865 8835 3885
rect 8815 3815 8835 3835
rect 8815 3765 8835 3785
rect 8815 3715 8835 3735
rect 8965 4165 8985 4185
rect 8965 4115 8985 4135
rect 8965 4065 8985 4085
rect 8965 4015 8985 4035
rect 8965 3965 8985 3985
rect 8965 3915 8985 3935
rect 8965 3865 8985 3885
rect 8965 3815 8985 3835
rect 8965 3765 8985 3785
rect 8965 3715 8985 3735
rect 9115 4165 9135 4185
rect 9115 4115 9135 4135
rect 9115 4065 9135 4085
rect 9115 4015 9135 4035
rect 9115 3965 9135 3985
rect 9115 3915 9135 3935
rect 9115 3865 9135 3885
rect 9115 3815 9135 3835
rect 9115 3765 9135 3785
rect 9115 3715 9135 3735
rect 9265 4165 9285 4185
rect 9265 4115 9285 4135
rect 9265 4065 9285 4085
rect 9265 4015 9285 4035
rect 9265 3965 9285 3985
rect 9265 3915 9285 3935
rect 9265 3865 9285 3885
rect 9265 3815 9285 3835
rect 9265 3765 9285 3785
rect 9265 3715 9285 3735
rect 9415 4165 9435 4185
rect 9415 4115 9435 4135
rect 9415 4065 9435 4085
rect 9415 4015 9435 4035
rect 9415 3965 9435 3985
rect 9415 3915 9435 3935
rect 9415 3865 9435 3885
rect 9415 3815 9435 3835
rect 9415 3765 9435 3785
rect 9415 3715 9435 3735
rect 9565 4165 9585 4185
rect 9565 4115 9585 4135
rect 9565 4065 9585 4085
rect 9565 4015 9585 4035
rect 9565 3965 9585 3985
rect 9565 3915 9585 3935
rect 9565 3865 9585 3885
rect 9565 3815 9585 3835
rect 9565 3765 9585 3785
rect 9565 3715 9585 3735
rect 9715 4165 9735 4185
rect 9715 4115 9735 4135
rect 9715 4065 9735 4085
rect 9715 4015 9735 4035
rect 9715 3965 9735 3985
rect 9715 3915 9735 3935
rect 9715 3865 9735 3885
rect 9715 3815 9735 3835
rect 9715 3765 9735 3785
rect 9715 3715 9735 3735
rect 9865 4165 9885 4185
rect 9865 4115 9885 4135
rect 9865 4065 9885 4085
rect 9865 4015 9885 4035
rect 9865 3965 9885 3985
rect 9865 3915 9885 3935
rect 9865 3865 9885 3885
rect 9865 3815 9885 3835
rect 9865 3765 9885 3785
rect 9865 3715 9885 3735
rect 10015 4165 10035 4185
rect 10015 4115 10035 4135
rect 10015 4065 10035 4085
rect 10015 4015 10035 4035
rect 10015 3965 10035 3985
rect 10015 3915 10035 3935
rect 10015 3865 10035 3885
rect 10015 3815 10035 3835
rect 10015 3765 10035 3785
rect 10015 3715 10035 3735
rect 10165 4165 10185 4185
rect 10165 4115 10185 4135
rect 10165 4065 10185 4085
rect 10165 4015 10185 4035
rect 10165 3965 10185 3985
rect 10165 3915 10185 3935
rect 10165 3865 10185 3885
rect 10165 3815 10185 3835
rect 10165 3765 10185 3785
rect 10165 3715 10185 3735
rect 10315 4165 10335 4185
rect 10315 4115 10335 4135
rect 10315 4065 10335 4085
rect 10315 4015 10335 4035
rect 10315 3965 10335 3985
rect 10315 3915 10335 3935
rect 10315 3865 10335 3885
rect 10315 3815 10335 3835
rect 10315 3765 10335 3785
rect 10315 3715 10335 3735
rect 10465 4165 10485 4185
rect 10465 4115 10485 4135
rect 10465 4065 10485 4085
rect 10465 4015 10485 4035
rect 10465 3965 10485 3985
rect 10465 3915 10485 3935
rect 10465 3865 10485 3885
rect 10465 3815 10485 3835
rect 10465 3765 10485 3785
rect 10465 3715 10485 3735
rect 10615 4165 10635 4185
rect 10615 4115 10635 4135
rect 10615 4065 10635 4085
rect 10615 4015 10635 4035
rect 10615 3965 10635 3985
rect 10615 3915 10635 3935
rect 10615 3865 10635 3885
rect 10615 3815 10635 3835
rect 10615 3765 10635 3785
rect 10615 3715 10635 3735
rect 10765 4165 10785 4185
rect 10765 4115 10785 4135
rect 10765 4065 10785 4085
rect 10765 4015 10785 4035
rect 10765 3965 10785 3985
rect 10765 3915 10785 3935
rect 10765 3865 10785 3885
rect 10765 3815 10785 3835
rect 10765 3765 10785 3785
rect 10765 3715 10785 3735
rect 11365 4165 11385 4185
rect 11365 4115 11385 4135
rect 11365 4065 11385 4085
rect 11365 4015 11385 4035
rect 11365 3965 11385 3985
rect 11365 3915 11385 3935
rect 11365 3865 11385 3885
rect 11365 3815 11385 3835
rect 11365 3765 11385 3785
rect 11365 3715 11385 3735
rect 11965 4165 11985 4185
rect 11965 4115 11985 4135
rect 11965 4065 11985 4085
rect 11965 4015 11985 4035
rect 11965 3965 11985 3985
rect 11965 3915 11985 3935
rect 11965 3865 11985 3885
rect 11965 3815 11985 3835
rect 11965 3765 11985 3785
rect 11965 3715 11985 3735
rect 12565 4165 12585 4185
rect 12565 4115 12585 4135
rect 12565 4065 12585 4085
rect 12565 4015 12585 4035
rect 12565 3965 12585 3985
rect 12565 3915 12585 3935
rect 12565 3865 12585 3885
rect 12565 3815 12585 3835
rect 12565 3765 12585 3785
rect 12565 3715 12585 3735
rect 13165 4165 13185 4185
rect 13165 4115 13185 4135
rect 13165 4065 13185 4085
rect 13165 4015 13185 4035
rect 13165 3965 13185 3985
rect 13165 3915 13185 3935
rect 13165 3865 13185 3885
rect 13165 3815 13185 3835
rect 13165 3765 13185 3785
rect 13165 3715 13185 3735
rect 13765 4165 13785 4185
rect 13765 4115 13785 4135
rect 13765 4065 13785 4085
rect 13765 4015 13785 4035
rect 13765 3965 13785 3985
rect 13765 3915 13785 3935
rect 13765 3865 13785 3885
rect 13765 3815 13785 3835
rect 13765 3765 13785 3785
rect 13765 3715 13785 3735
rect 14365 4165 14385 4185
rect 14365 4115 14385 4135
rect 14365 4065 14385 4085
rect 14365 4015 14385 4035
rect 14365 3965 14385 3985
rect 14365 3915 14385 3935
rect 14365 3865 14385 3885
rect 14365 3815 14385 3835
rect 14365 3765 14385 3785
rect 14365 3715 14385 3735
rect 14965 4165 14985 4185
rect 14965 4115 14985 4135
rect 14965 4065 14985 4085
rect 14965 4015 14985 4035
rect 14965 3965 14985 3985
rect 14965 3915 14985 3935
rect 14965 3865 14985 3885
rect 14965 3815 14985 3835
rect 14965 3765 14985 3785
rect 14965 3715 14985 3735
rect 15565 4165 15585 4185
rect 15565 4115 15585 4135
rect 15565 4065 15585 4085
rect 15565 4015 15585 4035
rect 15565 3965 15585 3985
rect 15565 3915 15585 3935
rect 15565 3865 15585 3885
rect 15565 3815 15585 3835
rect 15565 3765 15585 3785
rect 15565 3715 15585 3735
rect 16165 4165 16185 4185
rect 16165 4115 16185 4135
rect 16165 4065 16185 4085
rect 16165 4015 16185 4035
rect 16165 3965 16185 3985
rect 16165 3915 16185 3935
rect 16165 3865 16185 3885
rect 16165 3815 16185 3835
rect 16165 3765 16185 3785
rect 16165 3715 16185 3735
rect 16315 4065 16335 4085
rect 16315 4015 16335 4035
rect 16315 3965 16335 3985
rect 16315 3915 16335 3935
rect 16315 3865 16335 3885
rect 16315 3815 16335 3835
rect 16315 3765 16335 3785
rect 16315 3715 16335 3735
rect 16465 4165 16485 4185
rect 16465 4115 16485 4135
rect 16465 4065 16485 4085
rect 16465 4015 16485 4035
rect 16465 3965 16485 3985
rect 16465 3915 16485 3935
rect 16465 3865 16485 3885
rect 16465 3815 16485 3835
rect 16615 4065 16635 4085
rect 16615 4015 16635 4035
rect 16615 3965 16635 3985
rect 16615 3915 16635 3935
rect 16615 3865 16635 3885
rect 16615 3815 16635 3835
rect 16615 3765 16635 3785
rect 16615 3715 16635 3735
rect 16765 4165 16785 4185
rect 16765 4115 16785 4135
rect 16765 4065 16785 4085
rect 16765 4015 16785 4035
rect 16765 3965 16785 3985
rect 16765 3915 16785 3935
rect 16765 3865 16785 3885
rect 16765 3815 16785 3835
rect 16915 4065 16935 4085
rect 16915 4015 16935 4035
rect 16915 3965 16935 3985
rect 16915 3915 16935 3935
rect 16915 3865 16935 3885
rect 16915 3815 16935 3835
rect 16915 3765 16935 3785
rect 16915 3715 16935 3735
rect 17065 4165 17085 4185
rect 17065 4115 17085 4135
rect 17065 4065 17085 4085
rect 17065 4015 17085 4035
rect 17065 3965 17085 3985
rect 17065 3915 17085 3935
rect 17065 3865 17085 3885
rect 17065 3815 17085 3835
rect 17215 4065 17235 4085
rect 17215 4015 17235 4035
rect 17215 3965 17235 3985
rect 17215 3915 17235 3935
rect 17215 3865 17235 3885
rect 17215 3815 17235 3835
rect 17215 3765 17235 3785
rect 17215 3715 17235 3735
rect 17365 4165 17385 4185
rect 17365 4115 17385 4135
rect 17365 4065 17385 4085
rect 17365 4015 17385 4035
rect 17365 3965 17385 3985
rect 17365 3915 17385 3935
rect 17365 3865 17385 3885
rect 17365 3815 17385 3835
rect 17365 3765 17385 3785
rect 17365 3715 17385 3735
rect 17965 4065 17985 4085
rect 17965 4015 17985 4035
rect 17965 3965 17985 3985
rect 17965 3915 17985 3935
rect 17965 3865 17985 3885
rect 17965 3815 17985 3835
rect 17965 3765 17985 3785
rect 17965 3715 17985 3735
rect 18565 4165 18585 4185
rect 18565 4115 18585 4135
rect 18565 4065 18585 4085
rect 18565 4015 18585 4035
rect 18565 3965 18585 3985
rect 18565 3915 18585 3935
rect 18565 3865 18585 3885
rect 18565 3815 18585 3835
rect 18565 3765 18585 3785
rect 18565 3715 18585 3735
rect 18715 4065 18735 4085
rect 18715 4015 18735 4035
rect 18715 3965 18735 3985
rect 18715 3915 18735 3935
rect 18715 3865 18735 3885
rect 18715 3815 18735 3835
rect 18715 3765 18735 3785
rect 18715 3715 18735 3735
rect 18865 4165 18885 4185
rect 18865 4115 18885 4135
rect 18865 4065 18885 4085
rect 18865 4015 18885 4035
rect 18865 3965 18885 3985
rect 18865 3915 18885 3935
rect 18865 3865 18885 3885
rect 18865 3815 18885 3835
rect 19015 4065 19035 4085
rect 19015 4015 19035 4035
rect 19015 3965 19035 3985
rect 19015 3915 19035 3935
rect 19015 3865 19035 3885
rect 19015 3815 19035 3835
rect 19015 3765 19035 3785
rect 19015 3715 19035 3735
rect 19165 4165 19185 4185
rect 19165 4115 19185 4135
rect 19165 4065 19185 4085
rect 19165 4015 19185 4035
rect 19165 3965 19185 3985
rect 19165 3915 19185 3935
rect 19165 3865 19185 3885
rect 19165 3815 19185 3835
rect 19315 4065 19335 4085
rect 19315 4015 19335 4035
rect 19315 3965 19335 3985
rect 19315 3915 19335 3935
rect 19315 3865 19335 3885
rect 19315 3815 19335 3835
rect 19315 3765 19335 3785
rect 19315 3715 19335 3735
rect 19465 4165 19485 4185
rect 19465 4115 19485 4135
rect 19465 4065 19485 4085
rect 19465 4015 19485 4035
rect 19465 3965 19485 3985
rect 19465 3915 19485 3935
rect 19465 3865 19485 3885
rect 19465 3815 19485 3835
rect 19615 4065 19635 4085
rect 19615 4015 19635 4035
rect 19615 3965 19635 3985
rect 19615 3915 19635 3935
rect 19615 3865 19635 3885
rect 19615 3815 19635 3835
rect 19615 3765 19635 3785
rect 19615 3715 19635 3735
rect 19765 4165 19785 4185
rect 19765 4115 19785 4135
rect 19765 4065 19785 4085
rect 19765 4015 19785 4035
rect 19765 3965 19785 3985
rect 19765 3915 19785 3935
rect 19765 3865 19785 3885
rect 19765 3815 19785 3835
rect 19765 3765 19785 3785
rect 19765 3715 19785 3735
rect 20365 4165 20385 4185
rect 20365 4115 20385 4135
rect 20365 4065 20385 4085
rect 20365 4015 20385 4035
rect 20365 3965 20385 3985
rect 20365 3915 20385 3935
rect 20365 3865 20385 3885
rect 20365 3815 20385 3835
rect 20365 3765 20385 3785
rect 20365 3715 20385 3735
rect 20965 4165 20985 4185
rect 20965 4115 20985 4135
rect 20965 4065 20985 4085
rect 20965 4015 20985 4035
rect 20965 3965 20985 3985
rect 20965 3915 20985 3935
rect 20965 3865 20985 3885
rect 20965 3815 20985 3835
rect 20965 3765 20985 3785
rect 20965 3715 20985 3735
rect 21415 4165 21435 4185
rect 21415 4115 21435 4135
rect 21415 4065 21435 4085
rect 21415 4015 21435 4035
rect 21415 3965 21435 3985
rect 21415 3915 21435 3935
rect 21415 3865 21435 3885
rect 21415 3815 21435 3835
rect 21415 3765 21435 3785
rect 21415 3715 21435 3735
rect 21865 4165 21885 4185
rect 21865 4115 21885 4135
rect 21865 4065 21885 4085
rect 21865 4015 21885 4035
rect 21865 3965 21885 3985
rect 21865 3915 21885 3935
rect 21865 3865 21885 3885
rect 21865 3815 21885 3835
rect 21865 3765 21885 3785
rect 21865 3715 21885 3735
rect 22465 4165 22485 4185
rect 22465 4115 22485 4135
rect 22465 4065 22485 4085
rect 22465 4015 22485 4035
rect 22465 3965 22485 3985
rect 22465 3915 22485 3935
rect 22465 3865 22485 3885
rect 22465 3815 22485 3835
rect 22465 3765 22485 3785
rect 22465 3715 22485 3735
rect 23065 4165 23085 4185
rect 23065 4115 23085 4135
rect 23065 4065 23085 4085
rect 23065 4015 23085 4035
rect 23065 3965 23085 3985
rect 23065 3915 23085 3935
rect 23065 3865 23085 3885
rect 23065 3815 23085 3835
rect 23065 3765 23085 3785
rect 23065 3715 23085 3735
rect 23515 4165 23535 4185
rect 23515 4115 23535 4135
rect 23515 4065 23535 4085
rect 23515 4015 23535 4035
rect 23515 3965 23535 3985
rect 23515 3915 23535 3935
rect 23515 3865 23535 3885
rect 23515 3815 23535 3835
rect 23515 3765 23535 3785
rect 23515 3715 23535 3735
rect 23965 4165 23985 4185
rect 23965 4115 23985 4135
rect 23965 4065 23985 4085
rect 23965 4015 23985 4035
rect 23965 3965 23985 3985
rect 23965 3915 23985 3935
rect 23965 3865 23985 3885
rect 23965 3815 23985 3835
rect 23965 3765 23985 3785
rect 23965 3715 23985 3735
rect 24565 4165 24585 4185
rect 24565 4115 24585 4135
rect 24565 4065 24585 4085
rect 24565 4015 24585 4035
rect 24565 3965 24585 3985
rect 24565 3915 24585 3935
rect 24565 3865 24585 3885
rect 24565 3815 24585 3835
rect 24565 3765 24585 3785
rect 24565 3715 24585 3735
rect 25165 4165 25185 4185
rect 25165 4115 25185 4135
rect 25165 4065 25185 4085
rect 25165 4015 25185 4035
rect 25165 3965 25185 3985
rect 25165 3915 25185 3935
rect 25165 3865 25185 3885
rect 25165 3815 25185 3835
rect 25165 3765 25185 3785
rect 25165 3715 25185 3735
rect 25615 4165 25635 4185
rect 25615 4115 25635 4135
rect 25615 4065 25635 4085
rect 25615 4015 25635 4035
rect 25615 3965 25635 3985
rect 25615 3915 25635 3935
rect 25615 3865 25635 3885
rect 25615 3815 25635 3835
rect 25615 3765 25635 3785
rect 25615 3715 25635 3735
rect 26065 4165 26085 4185
rect 26065 4115 26085 4135
rect 26065 4065 26085 4085
rect 26065 4015 26085 4035
rect 26065 3965 26085 3985
rect 26065 3915 26085 3935
rect 26065 3865 26085 3885
rect 26065 3815 26085 3835
rect 26065 3765 26085 3785
rect 26065 3715 26085 3735
rect 26665 4165 26685 4185
rect 26665 4115 26685 4135
rect 26665 4065 26685 4085
rect 26665 4015 26685 4035
rect 26665 3965 26685 3985
rect 26665 3915 26685 3935
rect 26665 3865 26685 3885
rect 26665 3815 26685 3835
rect 26665 3765 26685 3785
rect 26665 3715 26685 3735
rect 27265 4165 27285 4185
rect 27265 4115 27285 4135
rect 27265 4065 27285 4085
rect 27265 4015 27285 4035
rect 27265 3965 27285 3985
rect 27265 3915 27285 3935
rect 27265 3865 27285 3885
rect 27265 3815 27285 3835
rect 27265 3765 27285 3785
rect 27265 3715 27285 3735
rect 27715 4165 27735 4185
rect 27715 4115 27735 4135
rect 27715 4065 27735 4085
rect 27715 4015 27735 4035
rect 27715 3965 27735 3985
rect 27715 3915 27735 3935
rect 27715 3865 27735 3885
rect 27715 3815 27735 3835
rect 27715 3765 27735 3785
rect 27715 3715 27735 3735
rect 28165 4165 28185 4185
rect 28165 4115 28185 4135
rect 28165 4065 28185 4085
rect 28165 4015 28185 4035
rect 28165 3965 28185 3985
rect 28165 3915 28185 3935
rect 28165 3865 28185 3885
rect 28165 3815 28185 3835
rect 28165 3765 28185 3785
rect 28165 3715 28185 3735
rect 28765 4165 28785 4185
rect 28765 4115 28785 4135
rect 28765 4065 28785 4085
rect 28765 4015 28785 4035
rect 28765 3965 28785 3985
rect 28765 3915 28785 3935
rect 28765 3865 28785 3885
rect 28765 3815 28785 3835
rect 28765 3765 28785 3785
rect 28765 3715 28785 3735
rect 29365 4165 29385 4185
rect 29365 4115 29385 4135
rect 29365 4065 29385 4085
rect 29365 4015 29385 4035
rect 29365 3965 29385 3985
rect 29365 3915 29385 3935
rect 29365 3865 29385 3885
rect 29365 3815 29385 3835
rect 29365 3765 29385 3785
rect 29365 3715 29385 3735
rect 29515 4065 29535 4085
rect 29515 4015 29535 4035
rect 29515 3965 29535 3985
rect 29515 3915 29535 3935
rect 29515 3865 29535 3885
rect 29515 3815 29535 3835
rect 29515 3765 29535 3785
rect 29515 3715 29535 3735
rect 29665 4165 29685 4185
rect 29665 4115 29685 4135
rect 29665 4065 29685 4085
rect 29665 4015 29685 4035
rect 29665 3965 29685 3985
rect 29665 3915 29685 3935
rect 29665 3865 29685 3885
rect 29665 3815 29685 3835
rect 29815 4165 29835 4185
rect 29815 4115 29835 4135
rect 29815 4065 29835 4085
rect 29815 4015 29835 4035
rect 29815 3965 29835 3985
rect 29815 3915 29835 3935
rect 29815 3865 29835 3885
rect 29815 3815 29835 3835
rect 29815 3765 29835 3785
rect 29815 3715 29835 3735
rect 29965 4165 29985 4185
rect 29965 4115 29985 4135
rect 29965 4065 29985 4085
rect 29965 4015 29985 4035
rect 29965 3965 29985 3985
rect 29965 3915 29985 3935
rect 29965 3865 29985 3885
rect 29965 3815 29985 3835
rect 30115 4065 30135 4085
rect 30115 4015 30135 4035
rect 30115 3965 30135 3985
rect 30115 3915 30135 3935
rect 30115 3865 30135 3885
rect 30115 3815 30135 3835
rect 30115 3765 30135 3785
rect 30115 3715 30135 3735
rect 30265 4165 30285 4185
rect 30265 4115 30285 4135
rect 30265 4065 30285 4085
rect 30265 4015 30285 4035
rect 30265 3965 30285 3985
rect 30265 3915 30285 3935
rect 30265 3865 30285 3885
rect 30265 3815 30285 3835
rect 30415 4165 30435 4185
rect 30415 4115 30435 4135
rect 30415 4065 30435 4085
rect 30415 4015 30435 4035
rect 30415 3965 30435 3985
rect 30415 3915 30435 3935
rect 30415 3865 30435 3885
rect 30415 3815 30435 3835
rect 30415 3765 30435 3785
rect 30415 3715 30435 3735
rect 30565 4165 30585 4185
rect 30565 4115 30585 4135
rect 30565 4065 30585 4085
rect 30565 4015 30585 4035
rect 30565 3965 30585 3985
rect 30565 3915 30585 3935
rect 30565 3865 30585 3885
rect 30565 3815 30585 3835
rect 30715 4065 30735 4085
rect 30715 4015 30735 4035
rect 30715 3965 30735 3985
rect 30715 3915 30735 3935
rect 30715 3865 30735 3885
rect 30715 3815 30735 3835
rect 30715 3765 30735 3785
rect 30715 3715 30735 3735
rect 30865 4165 30885 4185
rect 30865 4115 30885 4135
rect 30865 4065 30885 4085
rect 30865 4015 30885 4035
rect 30865 3965 30885 3985
rect 30865 3915 30885 3935
rect 30865 3865 30885 3885
rect 30865 3815 30885 3835
rect 31015 4165 31035 4185
rect 31015 4115 31035 4135
rect 31015 4065 31035 4085
rect 31015 4015 31035 4035
rect 31015 3965 31035 3985
rect 31015 3915 31035 3935
rect 31015 3865 31035 3885
rect 31015 3815 31035 3835
rect 31015 3765 31035 3785
rect 31015 3715 31035 3735
rect 31165 4165 31185 4185
rect 31165 4115 31185 4135
rect 31165 4065 31185 4085
rect 31165 4015 31185 4035
rect 31165 3965 31185 3985
rect 31165 3915 31185 3935
rect 31165 3865 31185 3885
rect 31165 3815 31185 3835
rect 31315 4065 31335 4085
rect 31315 4015 31335 4035
rect 31315 3965 31335 3985
rect 31315 3915 31335 3935
rect 31315 3865 31335 3885
rect 31315 3815 31335 3835
rect 31315 3765 31335 3785
rect 31315 3715 31335 3735
rect 31465 4165 31485 4185
rect 31465 4115 31485 4135
rect 31465 4065 31485 4085
rect 31465 4015 31485 4035
rect 31465 3965 31485 3985
rect 31465 3915 31485 3935
rect 31465 3865 31485 3885
rect 31465 3815 31485 3835
rect 31465 3765 31485 3785
rect 31465 3715 31485 3735
rect 32065 4165 32085 4185
rect 32065 4115 32085 4135
rect 32065 4065 32085 4085
rect 32065 4015 32085 4035
rect 32065 3965 32085 3985
rect 32065 3915 32085 3935
rect 32065 3865 32085 3885
rect 32065 3815 32085 3835
rect 32065 3765 32085 3785
rect 32065 3715 32085 3735
rect -485 3615 -465 3635
rect -185 3615 -165 3635
rect 115 3615 135 3635
rect 415 3615 435 3635
rect 715 3615 735 3635
rect 1015 3615 1035 3635
rect 1315 3615 1335 3635
rect 1615 3615 1635 3635
rect 1915 3615 1935 3635
rect 2215 3615 2235 3635
rect 2515 3615 2535 3635
rect 2815 3615 2835 3635
rect 3115 3615 3135 3635
rect 3415 3615 3435 3635
rect 3715 3615 3735 3635
rect 4015 3615 4035 3635
rect 4315 3615 4335 3635
rect 4615 3615 4635 3635
rect 4915 3615 4935 3635
rect 5215 3615 5235 3635
rect 5515 3615 5535 3635
rect 5815 3615 5835 3635
rect 6115 3615 6135 3635
rect 6415 3615 6435 3635
rect 6715 3615 6735 3635
rect 7015 3615 7035 3635
rect 7315 3615 7335 3635
rect 7615 3615 7635 3635
rect 7915 3615 7935 3635
rect 8215 3615 8235 3635
rect 8515 3615 8535 3635
rect 8815 3615 8835 3635
rect 9115 3615 9135 3635
rect 9415 3615 9435 3635
rect 9715 3615 9735 3635
rect 10015 3615 10035 3635
rect 10315 3615 10335 3635
rect 10615 3615 10635 3635
rect 10915 3615 10935 3635
rect 11215 3615 11235 3635
rect 11515 3615 11535 3635
rect 11815 3615 11835 3635
rect 12115 3615 12135 3635
rect 12415 3615 12435 3635
rect 12715 3615 12735 3635
rect 13015 3615 13035 3635
rect 13315 3615 13335 3635
rect 13615 3615 13635 3635
rect 13915 3615 13935 3635
rect 14215 3615 14235 3635
rect 14515 3615 14535 3635
rect 14815 3615 14835 3635
rect 15115 3615 15135 3635
rect 15415 3615 15435 3635
rect 15715 3615 15735 3635
rect 16015 3615 16035 3635
rect 16315 3615 16335 3635
rect 16615 3615 16635 3635
rect 16915 3615 16935 3635
rect 17215 3615 17235 3635
rect 17515 3615 17535 3635
rect 17815 3615 17835 3635
rect 18115 3615 18135 3635
rect 18415 3615 18435 3635
rect 18715 3615 18735 3635
rect 19015 3615 19035 3635
rect 19315 3615 19335 3635
rect 19615 3615 19635 3635
rect 19915 3615 19935 3635
rect 20215 3615 20235 3635
rect 20515 3615 20535 3635
rect 20815 3615 20835 3635
rect 21115 3615 21135 3635
rect 21715 3615 21735 3635
rect 22015 3615 22035 3635
rect 22315 3615 22335 3635
rect 22615 3615 22635 3635
rect 22915 3615 22935 3635
rect 23215 3615 23235 3635
rect 23365 3615 23385 3635
rect 23665 3615 23685 3635
rect 23815 3615 23835 3635
rect 24115 3615 24135 3635
rect 24415 3615 24435 3635
rect 24715 3615 24735 3635
rect 25015 3615 25035 3635
rect 25465 3615 25485 3635
rect 25765 3615 25785 3635
rect 26215 3615 26235 3635
rect 26515 3615 26535 3635
rect 26815 3615 26835 3635
rect 27115 3615 27135 3635
rect 27565 3615 27585 3635
rect 27865 3615 27885 3635
rect 28315 3615 28335 3635
rect 28615 3615 28635 3635
rect 28915 3615 28935 3635
rect 29215 3615 29235 3635
rect 29665 3615 29685 3635
rect 29965 3615 29985 3635
rect 30265 3615 30285 3635
rect 30565 3615 30585 3635
rect 30865 3615 30885 3635
rect 31165 3615 31185 3635
rect 31615 3615 31635 3635
rect 31915 3615 31935 3635
rect -635 3515 -615 3535
rect -635 3465 -615 3485
rect -635 3415 -615 3435
rect -635 3365 -615 3385
rect -635 3315 -615 3335
rect -635 3265 -615 3285
rect -635 3215 -615 3235
rect -635 3165 -615 3185
rect -635 3115 -615 3135
rect -635 3065 -615 3085
rect -485 3515 -465 3535
rect -485 3465 -465 3485
rect -485 3415 -465 3435
rect -485 3365 -465 3385
rect -485 3315 -465 3335
rect -485 3265 -465 3285
rect -485 3215 -465 3235
rect -485 3165 -465 3185
rect -485 3115 -465 3135
rect -485 3065 -465 3085
rect -335 3415 -315 3435
rect -335 3365 -315 3385
rect -335 3315 -315 3335
rect -335 3265 -315 3285
rect -335 3215 -315 3235
rect -335 3165 -315 3185
rect -335 3115 -315 3135
rect -335 3065 -315 3085
rect -185 3515 -165 3535
rect -185 3465 -165 3485
rect -185 3415 -165 3435
rect -185 3365 -165 3385
rect -185 3315 -165 3335
rect -185 3265 -165 3285
rect -185 3215 -165 3235
rect -185 3165 -165 3185
rect -185 3115 -165 3135
rect -185 3065 -165 3085
rect -35 3415 -15 3435
rect -35 3365 -15 3385
rect -35 3315 -15 3335
rect -35 3265 -15 3285
rect -35 3215 -15 3235
rect -35 3165 -15 3185
rect -35 3115 -15 3135
rect -35 3065 -15 3085
rect 565 3515 585 3535
rect 565 3465 585 3485
rect 565 3415 585 3435
rect 565 3365 585 3385
rect 565 3315 585 3335
rect 565 3265 585 3285
rect 565 3215 585 3235
rect 565 3165 585 3185
rect 565 3115 585 3135
rect 565 3065 585 3085
rect 715 3515 735 3535
rect 715 3465 735 3485
rect 715 3415 735 3435
rect 715 3365 735 3385
rect 715 3315 735 3335
rect 715 3265 735 3285
rect 715 3215 735 3235
rect 715 3165 735 3185
rect 865 3415 885 3435
rect 865 3365 885 3385
rect 865 3315 885 3335
rect 865 3265 885 3285
rect 865 3215 885 3235
rect 865 3165 885 3185
rect 865 3115 885 3135
rect 865 3065 885 3085
rect 1015 3515 1035 3535
rect 1015 3465 1035 3485
rect 1015 3415 1035 3435
rect 1015 3365 1035 3385
rect 1015 3315 1035 3335
rect 1015 3265 1035 3285
rect 1015 3215 1035 3235
rect 1015 3165 1035 3185
rect 1165 3415 1185 3435
rect 1165 3365 1185 3385
rect 1165 3315 1185 3335
rect 1165 3265 1185 3285
rect 1165 3215 1185 3235
rect 1165 3165 1185 3185
rect 1165 3115 1185 3135
rect 1165 3065 1185 3085
rect 1315 3515 1335 3535
rect 1315 3465 1335 3485
rect 1315 3415 1335 3435
rect 1315 3365 1335 3385
rect 1315 3315 1335 3335
rect 1315 3265 1335 3285
rect 1315 3215 1335 3235
rect 1315 3165 1335 3185
rect 1465 3415 1485 3435
rect 1465 3365 1485 3385
rect 1465 3315 1485 3335
rect 1465 3265 1485 3285
rect 1465 3215 1485 3235
rect 1465 3165 1485 3185
rect 1465 3115 1485 3135
rect 1465 3065 1485 3085
rect 1615 3515 1635 3535
rect 1615 3465 1635 3485
rect 1615 3415 1635 3435
rect 1615 3365 1635 3385
rect 1615 3315 1635 3335
rect 1615 3265 1635 3285
rect 1615 3215 1635 3235
rect 1615 3165 1635 3185
rect 1765 3515 1785 3535
rect 1765 3465 1785 3485
rect 1765 3415 1785 3435
rect 1765 3365 1785 3385
rect 1765 3315 1785 3335
rect 1765 3265 1785 3285
rect 1765 3215 1785 3235
rect 1765 3165 1785 3185
rect 1765 3115 1785 3135
rect 1765 3065 1785 3085
rect 1915 3515 1935 3535
rect 1915 3465 1935 3485
rect 1915 3415 1935 3435
rect 1915 3365 1935 3385
rect 1915 3315 1935 3335
rect 1915 3265 1935 3285
rect 1915 3215 1935 3235
rect 1915 3165 1935 3185
rect 2065 3415 2085 3435
rect 2065 3365 2085 3385
rect 2065 3315 2085 3335
rect 2065 3265 2085 3285
rect 2065 3215 2085 3235
rect 2065 3165 2085 3185
rect 2065 3115 2085 3135
rect 2065 3065 2085 3085
rect 2215 3515 2235 3535
rect 2215 3465 2235 3485
rect 2215 3415 2235 3435
rect 2215 3365 2235 3385
rect 2215 3315 2235 3335
rect 2215 3265 2235 3285
rect 2215 3215 2235 3235
rect 2215 3165 2235 3185
rect 2365 3515 2385 3535
rect 2365 3465 2385 3485
rect 2365 3415 2385 3435
rect 2365 3365 2385 3385
rect 2365 3315 2385 3335
rect 2365 3265 2385 3285
rect 2365 3215 2385 3235
rect 2365 3165 2385 3185
rect 2365 3115 2385 3135
rect 2365 3065 2385 3085
rect 2515 3515 2535 3535
rect 2515 3465 2535 3485
rect 2515 3415 2535 3435
rect 2515 3365 2535 3385
rect 2515 3315 2535 3335
rect 2515 3265 2535 3285
rect 2515 3215 2535 3235
rect 2515 3165 2535 3185
rect 2665 3415 2685 3435
rect 2665 3365 2685 3385
rect 2665 3315 2685 3335
rect 2665 3265 2685 3285
rect 2665 3215 2685 3235
rect 2665 3165 2685 3185
rect 2665 3115 2685 3135
rect 2665 3065 2685 3085
rect 2815 3515 2835 3535
rect 2815 3465 2835 3485
rect 2815 3415 2835 3435
rect 2815 3365 2835 3385
rect 2815 3315 2835 3335
rect 2815 3265 2835 3285
rect 2815 3215 2835 3235
rect 2815 3165 2835 3185
rect 2965 3415 2985 3435
rect 2965 3365 2985 3385
rect 2965 3315 2985 3335
rect 2965 3265 2985 3285
rect 2965 3215 2985 3235
rect 2965 3165 2985 3185
rect 2965 3115 2985 3135
rect 2965 3065 2985 3085
rect 3115 3515 3135 3535
rect 3115 3465 3135 3485
rect 3115 3415 3135 3435
rect 3115 3365 3135 3385
rect 3115 3315 3135 3335
rect 3115 3265 3135 3285
rect 3115 3215 3135 3235
rect 3115 3165 3135 3185
rect 3265 3415 3285 3435
rect 3265 3365 3285 3385
rect 3265 3315 3285 3335
rect 3265 3265 3285 3285
rect 3265 3215 3285 3235
rect 3265 3165 3285 3185
rect 3265 3115 3285 3135
rect 3265 3065 3285 3085
rect 3415 3515 3435 3535
rect 3415 3465 3435 3485
rect 3415 3415 3435 3435
rect 3415 3365 3435 3385
rect 3415 3315 3435 3335
rect 3415 3265 3435 3285
rect 3415 3215 3435 3235
rect 3415 3165 3435 3185
rect 3565 3515 3585 3535
rect 3565 3465 3585 3485
rect 3565 3415 3585 3435
rect 3565 3365 3585 3385
rect 3565 3315 3585 3335
rect 3565 3265 3585 3285
rect 3565 3215 3585 3235
rect 3565 3165 3585 3185
rect 3565 3115 3585 3135
rect 3565 3065 3585 3085
rect 4165 3415 4185 3435
rect 4165 3365 4185 3385
rect 4165 3315 4185 3335
rect 4165 3265 4185 3285
rect 4165 3215 4185 3235
rect 4165 3165 4185 3185
rect 4165 3115 4185 3135
rect 4165 3065 4185 3085
rect 4765 3515 4785 3535
rect 4765 3465 4785 3485
rect 4765 3415 4785 3435
rect 4765 3365 4785 3385
rect 4765 3315 4785 3335
rect 4765 3265 4785 3285
rect 4765 3215 4785 3235
rect 4765 3165 4785 3185
rect 4765 3115 4785 3135
rect 4765 3065 4785 3085
rect 4915 3515 4935 3535
rect 4915 3465 4935 3485
rect 4915 3415 4935 3435
rect 4915 3365 4935 3385
rect 4915 3315 4935 3335
rect 4915 3265 4935 3285
rect 4915 3215 4935 3235
rect 4915 3165 4935 3185
rect 5065 3415 5085 3435
rect 5065 3365 5085 3385
rect 5065 3315 5085 3335
rect 5065 3265 5085 3285
rect 5065 3215 5085 3235
rect 5065 3165 5085 3185
rect 5065 3115 5085 3135
rect 5065 3065 5085 3085
rect 5215 3515 5235 3535
rect 5215 3465 5235 3485
rect 5215 3415 5235 3435
rect 5215 3365 5235 3385
rect 5215 3315 5235 3335
rect 5215 3265 5235 3285
rect 5215 3215 5235 3235
rect 5215 3165 5235 3185
rect 5365 3415 5385 3435
rect 5365 3365 5385 3385
rect 5365 3315 5385 3335
rect 5365 3265 5385 3285
rect 5365 3215 5385 3235
rect 5365 3165 5385 3185
rect 5365 3115 5385 3135
rect 5365 3065 5385 3085
rect 5515 3515 5535 3535
rect 5515 3465 5535 3485
rect 5515 3415 5535 3435
rect 5515 3365 5535 3385
rect 5515 3315 5535 3335
rect 5515 3265 5535 3285
rect 5515 3215 5535 3235
rect 5515 3165 5535 3185
rect 5665 3415 5685 3435
rect 5665 3365 5685 3385
rect 5665 3315 5685 3335
rect 5665 3265 5685 3285
rect 5665 3215 5685 3235
rect 5665 3165 5685 3185
rect 5665 3115 5685 3135
rect 5665 3065 5685 3085
rect 5815 3515 5835 3535
rect 5815 3465 5835 3485
rect 5815 3415 5835 3435
rect 5815 3365 5835 3385
rect 5815 3315 5835 3335
rect 5815 3265 5835 3285
rect 5815 3215 5835 3235
rect 5815 3165 5835 3185
rect 5965 3515 5985 3535
rect 5965 3465 5985 3485
rect 5965 3415 5985 3435
rect 5965 3365 5985 3385
rect 5965 3315 5985 3335
rect 5965 3265 5985 3285
rect 5965 3215 5985 3235
rect 5965 3165 5985 3185
rect 5965 3115 5985 3135
rect 5965 3065 5985 3085
rect 6115 3515 6135 3535
rect 6115 3465 6135 3485
rect 6115 3415 6135 3435
rect 6115 3365 6135 3385
rect 6115 3315 6135 3335
rect 6115 3265 6135 3285
rect 6115 3215 6135 3235
rect 6115 3165 6135 3185
rect 6265 3415 6285 3435
rect 6265 3365 6285 3385
rect 6265 3315 6285 3335
rect 6265 3265 6285 3285
rect 6265 3215 6285 3235
rect 6265 3165 6285 3185
rect 6265 3115 6285 3135
rect 6265 3065 6285 3085
rect 6415 3515 6435 3535
rect 6415 3465 6435 3485
rect 6415 3415 6435 3435
rect 6415 3365 6435 3385
rect 6415 3315 6435 3335
rect 6415 3265 6435 3285
rect 6415 3215 6435 3235
rect 6415 3165 6435 3185
rect 6565 3515 6585 3535
rect 6565 3465 6585 3485
rect 6565 3415 6585 3435
rect 6565 3365 6585 3385
rect 6565 3315 6585 3335
rect 6565 3265 6585 3285
rect 6565 3215 6585 3235
rect 6565 3165 6585 3185
rect 6565 3115 6585 3135
rect 6565 3065 6585 3085
rect 6715 3515 6735 3535
rect 6715 3465 6735 3485
rect 6715 3415 6735 3435
rect 6715 3365 6735 3385
rect 6715 3315 6735 3335
rect 6715 3265 6735 3285
rect 6715 3215 6735 3235
rect 6715 3165 6735 3185
rect 6865 3415 6885 3435
rect 6865 3365 6885 3385
rect 6865 3315 6885 3335
rect 6865 3265 6885 3285
rect 6865 3215 6885 3235
rect 6865 3165 6885 3185
rect 6865 3115 6885 3135
rect 6865 3065 6885 3085
rect 7015 3515 7035 3535
rect 7015 3465 7035 3485
rect 7015 3415 7035 3435
rect 7015 3365 7035 3385
rect 7015 3315 7035 3335
rect 7015 3265 7035 3285
rect 7015 3215 7035 3235
rect 7015 3165 7035 3185
rect 7165 3415 7185 3435
rect 7165 3365 7185 3385
rect 7165 3315 7185 3335
rect 7165 3265 7185 3285
rect 7165 3215 7185 3235
rect 7165 3165 7185 3185
rect 7165 3115 7185 3135
rect 7165 3065 7185 3085
rect 7315 3515 7335 3535
rect 7315 3465 7335 3485
rect 7315 3415 7335 3435
rect 7315 3365 7335 3385
rect 7315 3315 7335 3335
rect 7315 3265 7335 3285
rect 7315 3215 7335 3235
rect 7315 3165 7335 3185
rect 7465 3415 7485 3435
rect 7465 3365 7485 3385
rect 7465 3315 7485 3335
rect 7465 3265 7485 3285
rect 7465 3215 7485 3235
rect 7465 3165 7485 3185
rect 7465 3115 7485 3135
rect 7465 3065 7485 3085
rect 7615 3515 7635 3535
rect 7615 3465 7635 3485
rect 7615 3415 7635 3435
rect 7615 3365 7635 3385
rect 7615 3315 7635 3335
rect 7615 3265 7635 3285
rect 7615 3215 7635 3235
rect 7615 3165 7635 3185
rect 7765 3515 7785 3535
rect 7765 3465 7785 3485
rect 7765 3415 7785 3435
rect 7765 3365 7785 3385
rect 7765 3315 7785 3335
rect 7765 3265 7785 3285
rect 7765 3215 7785 3235
rect 7765 3165 7785 3185
rect 7765 3115 7785 3135
rect 7765 3065 7785 3085
rect 8365 3515 8385 3535
rect 8365 3465 8385 3485
rect 8365 3415 8385 3435
rect 8365 3365 8385 3385
rect 8365 3315 8385 3335
rect 8365 3265 8385 3285
rect 8365 3215 8385 3235
rect 8365 3165 8385 3185
rect 8365 3115 8385 3135
rect 8365 3065 8385 3085
rect 8515 3515 8535 3535
rect 8515 3465 8535 3485
rect 8515 3415 8535 3435
rect 8515 3365 8535 3385
rect 8515 3315 8535 3335
rect 8515 3265 8535 3285
rect 8515 3215 8535 3235
rect 8515 3165 8535 3185
rect 8515 3115 8535 3135
rect 8515 3065 8535 3085
rect 8665 3515 8685 3535
rect 8665 3465 8685 3485
rect 8665 3415 8685 3435
rect 8665 3365 8685 3385
rect 8665 3315 8685 3335
rect 8665 3265 8685 3285
rect 8665 3215 8685 3235
rect 8665 3165 8685 3185
rect 8665 3115 8685 3135
rect 8665 3065 8685 3085
rect 8815 3515 8835 3535
rect 8815 3465 8835 3485
rect 8815 3415 8835 3435
rect 8815 3365 8835 3385
rect 8815 3315 8835 3335
rect 8815 3265 8835 3285
rect 8815 3215 8835 3235
rect 8815 3165 8835 3185
rect 8815 3115 8835 3135
rect 8815 3065 8835 3085
rect 8965 3515 8985 3535
rect 8965 3465 8985 3485
rect 8965 3415 8985 3435
rect 8965 3365 8985 3385
rect 8965 3315 8985 3335
rect 8965 3265 8985 3285
rect 8965 3215 8985 3235
rect 8965 3165 8985 3185
rect 8965 3115 8985 3135
rect 8965 3065 8985 3085
rect 9115 3515 9135 3535
rect 9115 3465 9135 3485
rect 9115 3415 9135 3435
rect 9115 3365 9135 3385
rect 9115 3315 9135 3335
rect 9115 3265 9135 3285
rect 9115 3215 9135 3235
rect 9115 3165 9135 3185
rect 9115 3115 9135 3135
rect 9115 3065 9135 3085
rect 9265 3515 9285 3535
rect 9265 3465 9285 3485
rect 9265 3415 9285 3435
rect 9265 3365 9285 3385
rect 9265 3315 9285 3335
rect 9265 3265 9285 3285
rect 9265 3215 9285 3235
rect 9265 3165 9285 3185
rect 9265 3115 9285 3135
rect 9265 3065 9285 3085
rect 9415 3515 9435 3535
rect 9415 3465 9435 3485
rect 9415 3415 9435 3435
rect 9415 3365 9435 3385
rect 9415 3315 9435 3335
rect 9415 3265 9435 3285
rect 9415 3215 9435 3235
rect 9415 3165 9435 3185
rect 9415 3115 9435 3135
rect 9415 3065 9435 3085
rect 9565 3515 9585 3535
rect 9565 3465 9585 3485
rect 9565 3415 9585 3435
rect 9565 3365 9585 3385
rect 9565 3315 9585 3335
rect 9565 3265 9585 3285
rect 9565 3215 9585 3235
rect 9565 3165 9585 3185
rect 9565 3115 9585 3135
rect 9565 3065 9585 3085
rect 9715 3515 9735 3535
rect 9715 3465 9735 3485
rect 9715 3415 9735 3435
rect 9715 3365 9735 3385
rect 9715 3315 9735 3335
rect 9715 3265 9735 3285
rect 9715 3215 9735 3235
rect 9715 3165 9735 3185
rect 9715 3115 9735 3135
rect 9715 3065 9735 3085
rect 9865 3515 9885 3535
rect 9865 3465 9885 3485
rect 9865 3415 9885 3435
rect 9865 3365 9885 3385
rect 9865 3315 9885 3335
rect 9865 3265 9885 3285
rect 9865 3215 9885 3235
rect 9865 3165 9885 3185
rect 9865 3115 9885 3135
rect 9865 3065 9885 3085
rect 10015 3515 10035 3535
rect 10015 3465 10035 3485
rect 10015 3415 10035 3435
rect 10015 3365 10035 3385
rect 10015 3315 10035 3335
rect 10015 3265 10035 3285
rect 10015 3215 10035 3235
rect 10015 3165 10035 3185
rect 10015 3115 10035 3135
rect 10015 3065 10035 3085
rect 10165 3515 10185 3535
rect 10165 3465 10185 3485
rect 10165 3415 10185 3435
rect 10165 3365 10185 3385
rect 10165 3315 10185 3335
rect 10165 3265 10185 3285
rect 10165 3215 10185 3235
rect 10165 3165 10185 3185
rect 10165 3115 10185 3135
rect 10165 3065 10185 3085
rect 10315 3515 10335 3535
rect 10315 3465 10335 3485
rect 10315 3415 10335 3435
rect 10315 3365 10335 3385
rect 10315 3315 10335 3335
rect 10315 3265 10335 3285
rect 10315 3215 10335 3235
rect 10315 3165 10335 3185
rect 10315 3115 10335 3135
rect 10315 3065 10335 3085
rect 10465 3515 10485 3535
rect 10465 3465 10485 3485
rect 10465 3415 10485 3435
rect 10465 3365 10485 3385
rect 10465 3315 10485 3335
rect 10465 3265 10485 3285
rect 10465 3215 10485 3235
rect 10465 3165 10485 3185
rect 10465 3115 10485 3135
rect 10465 3065 10485 3085
rect 10615 3515 10635 3535
rect 10615 3465 10635 3485
rect 10615 3415 10635 3435
rect 10615 3365 10635 3385
rect 10615 3315 10635 3335
rect 10615 3265 10635 3285
rect 10615 3215 10635 3235
rect 10615 3165 10635 3185
rect 10615 3115 10635 3135
rect 10615 3065 10635 3085
rect 10765 3515 10785 3535
rect 10765 3465 10785 3485
rect 10765 3415 10785 3435
rect 10765 3365 10785 3385
rect 10765 3315 10785 3335
rect 10765 3265 10785 3285
rect 10765 3215 10785 3235
rect 10765 3165 10785 3185
rect 10765 3115 10785 3135
rect 10765 3065 10785 3085
rect 11365 3515 11385 3535
rect 11365 3465 11385 3485
rect 11365 3415 11385 3435
rect 11365 3365 11385 3385
rect 11365 3315 11385 3335
rect 11365 3265 11385 3285
rect 11365 3215 11385 3235
rect 11365 3165 11385 3185
rect 11365 3115 11385 3135
rect 11365 3065 11385 3085
rect 11965 3515 11985 3535
rect 11965 3465 11985 3485
rect 11965 3415 11985 3435
rect 11965 3365 11985 3385
rect 11965 3315 11985 3335
rect 11965 3265 11985 3285
rect 11965 3215 11985 3235
rect 11965 3165 11985 3185
rect 11965 3115 11985 3135
rect 11965 3065 11985 3085
rect 12565 3515 12585 3535
rect 12565 3465 12585 3485
rect 12565 3415 12585 3435
rect 12565 3365 12585 3385
rect 12565 3315 12585 3335
rect 12565 3265 12585 3285
rect 12565 3215 12585 3235
rect 12565 3165 12585 3185
rect 12565 3115 12585 3135
rect 12565 3065 12585 3085
rect 13165 3515 13185 3535
rect 13165 3465 13185 3485
rect 13165 3415 13185 3435
rect 13165 3365 13185 3385
rect 13165 3315 13185 3335
rect 13165 3265 13185 3285
rect 13165 3215 13185 3235
rect 13165 3165 13185 3185
rect 13165 3115 13185 3135
rect 13165 3065 13185 3085
rect 13765 3515 13785 3535
rect 13765 3465 13785 3485
rect 13765 3415 13785 3435
rect 13765 3365 13785 3385
rect 13765 3315 13785 3335
rect 13765 3265 13785 3285
rect 13765 3215 13785 3235
rect 13765 3165 13785 3185
rect 13765 3115 13785 3135
rect 13765 3065 13785 3085
rect 14365 3515 14385 3535
rect 14365 3465 14385 3485
rect 14365 3415 14385 3435
rect 14365 3365 14385 3385
rect 14365 3315 14385 3335
rect 14365 3265 14385 3285
rect 14365 3215 14385 3235
rect 14365 3165 14385 3185
rect 14365 3115 14385 3135
rect 14365 3065 14385 3085
rect 14965 3515 14985 3535
rect 14965 3465 14985 3485
rect 14965 3415 14985 3435
rect 14965 3365 14985 3385
rect 14965 3315 14985 3335
rect 14965 3265 14985 3285
rect 14965 3215 14985 3235
rect 14965 3165 14985 3185
rect 14965 3115 14985 3135
rect 14965 3065 14985 3085
rect 15565 3515 15585 3535
rect 15565 3465 15585 3485
rect 15565 3415 15585 3435
rect 15565 3365 15585 3385
rect 15565 3315 15585 3335
rect 15565 3265 15585 3285
rect 15565 3215 15585 3235
rect 15565 3165 15585 3185
rect 15565 3115 15585 3135
rect 15565 3065 15585 3085
rect 16165 3515 16185 3535
rect 16165 3465 16185 3485
rect 16165 3415 16185 3435
rect 16165 3365 16185 3385
rect 16165 3315 16185 3335
rect 16165 3265 16185 3285
rect 16165 3215 16185 3235
rect 16165 3165 16185 3185
rect 16165 3115 16185 3135
rect 16165 3065 16185 3085
rect 16315 3515 16335 3535
rect 16315 3465 16335 3485
rect 16315 3415 16335 3435
rect 16315 3365 16335 3385
rect 16315 3315 16335 3335
rect 16315 3265 16335 3285
rect 16315 3215 16335 3235
rect 16315 3165 16335 3185
rect 16465 3415 16485 3435
rect 16465 3365 16485 3385
rect 16465 3315 16485 3335
rect 16465 3265 16485 3285
rect 16465 3215 16485 3235
rect 16465 3165 16485 3185
rect 16465 3115 16485 3135
rect 16465 3065 16485 3085
rect 16615 3515 16635 3535
rect 16615 3465 16635 3485
rect 16615 3415 16635 3435
rect 16615 3365 16635 3385
rect 16615 3315 16635 3335
rect 16615 3265 16635 3285
rect 16615 3215 16635 3235
rect 16615 3165 16635 3185
rect 16765 3415 16785 3435
rect 16765 3365 16785 3385
rect 16765 3315 16785 3335
rect 16765 3265 16785 3285
rect 16765 3215 16785 3235
rect 16765 3165 16785 3185
rect 16765 3115 16785 3135
rect 16765 3065 16785 3085
rect 16915 3515 16935 3535
rect 16915 3465 16935 3485
rect 16915 3415 16935 3435
rect 16915 3365 16935 3385
rect 16915 3315 16935 3335
rect 16915 3265 16935 3285
rect 16915 3215 16935 3235
rect 16915 3165 16935 3185
rect 17065 3415 17085 3435
rect 17065 3365 17085 3385
rect 17065 3315 17085 3335
rect 17065 3265 17085 3285
rect 17065 3215 17085 3235
rect 17065 3165 17085 3185
rect 17065 3115 17085 3135
rect 17065 3065 17085 3085
rect 17215 3515 17235 3535
rect 17215 3465 17235 3485
rect 17215 3415 17235 3435
rect 17215 3365 17235 3385
rect 17215 3315 17235 3335
rect 17215 3265 17235 3285
rect 17215 3215 17235 3235
rect 17215 3165 17235 3185
rect 17365 3515 17385 3535
rect 17365 3465 17385 3485
rect 17365 3415 17385 3435
rect 17365 3365 17385 3385
rect 17365 3315 17385 3335
rect 17365 3265 17385 3285
rect 17365 3215 17385 3235
rect 17365 3165 17385 3185
rect 17365 3115 17385 3135
rect 17365 3065 17385 3085
rect 17965 3515 17985 3535
rect 17965 3465 17985 3485
rect 17965 3415 17985 3435
rect 17965 3365 17985 3385
rect 17965 3315 17985 3335
rect 17965 3265 17985 3285
rect 17965 3215 17985 3235
rect 17965 3165 17985 3185
rect 18565 3515 18585 3535
rect 18565 3465 18585 3485
rect 18565 3415 18585 3435
rect 18565 3365 18585 3385
rect 18565 3315 18585 3335
rect 18565 3265 18585 3285
rect 18565 3215 18585 3235
rect 18565 3165 18585 3185
rect 18565 3115 18585 3135
rect 18565 3065 18585 3085
rect 18715 3515 18735 3535
rect 18715 3465 18735 3485
rect 18715 3415 18735 3435
rect 18715 3365 18735 3385
rect 18715 3315 18735 3335
rect 18715 3265 18735 3285
rect 18715 3215 18735 3235
rect 18715 3165 18735 3185
rect 18865 3415 18885 3435
rect 18865 3365 18885 3385
rect 18865 3315 18885 3335
rect 18865 3265 18885 3285
rect 18865 3215 18885 3235
rect 18865 3165 18885 3185
rect 18865 3115 18885 3135
rect 18865 3065 18885 3085
rect 19015 3515 19035 3535
rect 19015 3465 19035 3485
rect 19015 3415 19035 3435
rect 19015 3365 19035 3385
rect 19015 3315 19035 3335
rect 19015 3265 19035 3285
rect 19015 3215 19035 3235
rect 19015 3165 19035 3185
rect 19165 3415 19185 3435
rect 19165 3365 19185 3385
rect 19165 3315 19185 3335
rect 19165 3265 19185 3285
rect 19165 3215 19185 3235
rect 19165 3165 19185 3185
rect 19165 3115 19185 3135
rect 19165 3065 19185 3085
rect 19315 3515 19335 3535
rect 19315 3465 19335 3485
rect 19315 3415 19335 3435
rect 19315 3365 19335 3385
rect 19315 3315 19335 3335
rect 19315 3265 19335 3285
rect 19315 3215 19335 3235
rect 19315 3165 19335 3185
rect 19465 3415 19485 3435
rect 19465 3365 19485 3385
rect 19465 3315 19485 3335
rect 19465 3265 19485 3285
rect 19465 3215 19485 3235
rect 19465 3165 19485 3185
rect 19465 3115 19485 3135
rect 19465 3065 19485 3085
rect 19615 3515 19635 3535
rect 19615 3465 19635 3485
rect 19615 3415 19635 3435
rect 19615 3365 19635 3385
rect 19615 3315 19635 3335
rect 19615 3265 19635 3285
rect 19615 3215 19635 3235
rect 19615 3165 19635 3185
rect 19765 3515 19785 3535
rect 19765 3465 19785 3485
rect 19765 3415 19785 3435
rect 19765 3365 19785 3385
rect 19765 3315 19785 3335
rect 19765 3265 19785 3285
rect 19765 3215 19785 3235
rect 19765 3165 19785 3185
rect 19765 3115 19785 3135
rect 19765 3065 19785 3085
rect 20365 3515 20385 3535
rect 20365 3465 20385 3485
rect 20365 3415 20385 3435
rect 20365 3365 20385 3385
rect 20365 3315 20385 3335
rect 20365 3265 20385 3285
rect 20365 3215 20385 3235
rect 20365 3165 20385 3185
rect 20365 3115 20385 3135
rect 20365 3065 20385 3085
rect 20965 3515 20985 3535
rect 20965 3465 20985 3485
rect 20965 3415 20985 3435
rect 20965 3365 20985 3385
rect 20965 3315 20985 3335
rect 20965 3265 20985 3285
rect 20965 3215 20985 3235
rect 20965 3165 20985 3185
rect 20965 3115 20985 3135
rect 20965 3065 20985 3085
rect 21415 3515 21435 3535
rect 21415 3465 21435 3485
rect 21415 3415 21435 3435
rect 21415 3365 21435 3385
rect 21415 3315 21435 3335
rect 21415 3265 21435 3285
rect 21415 3215 21435 3235
rect 21415 3165 21435 3185
rect 21415 3115 21435 3135
rect 21415 3065 21435 3085
rect 21865 3515 21885 3535
rect 21865 3465 21885 3485
rect 21865 3415 21885 3435
rect 21865 3365 21885 3385
rect 21865 3315 21885 3335
rect 21865 3265 21885 3285
rect 21865 3215 21885 3235
rect 21865 3165 21885 3185
rect 21865 3115 21885 3135
rect 21865 3065 21885 3085
rect 22465 3515 22485 3535
rect 22465 3465 22485 3485
rect 22465 3415 22485 3435
rect 22465 3365 22485 3385
rect 22465 3315 22485 3335
rect 22465 3265 22485 3285
rect 22465 3215 22485 3235
rect 22465 3165 22485 3185
rect 22465 3115 22485 3135
rect 22465 3065 22485 3085
rect 23065 3515 23085 3535
rect 23065 3465 23085 3485
rect 23065 3415 23085 3435
rect 23065 3365 23085 3385
rect 23065 3315 23085 3335
rect 23065 3265 23085 3285
rect 23065 3215 23085 3235
rect 23065 3165 23085 3185
rect 23065 3115 23085 3135
rect 23065 3065 23085 3085
rect 23515 3515 23535 3535
rect 23515 3465 23535 3485
rect 23515 3415 23535 3435
rect 23515 3365 23535 3385
rect 23515 3315 23535 3335
rect 23515 3265 23535 3285
rect 23515 3215 23535 3235
rect 23515 3165 23535 3185
rect 23515 3115 23535 3135
rect 23515 3065 23535 3085
rect 23965 3515 23985 3535
rect 23965 3465 23985 3485
rect 23965 3415 23985 3435
rect 23965 3365 23985 3385
rect 23965 3315 23985 3335
rect 23965 3265 23985 3285
rect 23965 3215 23985 3235
rect 23965 3165 23985 3185
rect 23965 3115 23985 3135
rect 23965 3065 23985 3085
rect 24565 3515 24585 3535
rect 24565 3465 24585 3485
rect 24565 3415 24585 3435
rect 24565 3365 24585 3385
rect 24565 3315 24585 3335
rect 24565 3265 24585 3285
rect 24565 3215 24585 3235
rect 24565 3165 24585 3185
rect 24565 3115 24585 3135
rect 24565 3065 24585 3085
rect 25165 3515 25185 3535
rect 25165 3465 25185 3485
rect 25165 3415 25185 3435
rect 25165 3365 25185 3385
rect 25165 3315 25185 3335
rect 25165 3265 25185 3285
rect 25165 3215 25185 3235
rect 25165 3165 25185 3185
rect 25165 3115 25185 3135
rect 25165 3065 25185 3085
rect 25615 3515 25635 3535
rect 25615 3465 25635 3485
rect 25615 3415 25635 3435
rect 25615 3365 25635 3385
rect 25615 3315 25635 3335
rect 25615 3265 25635 3285
rect 25615 3215 25635 3235
rect 25615 3165 25635 3185
rect 25615 3115 25635 3135
rect 25615 3065 25635 3085
rect 26065 3515 26085 3535
rect 26065 3465 26085 3485
rect 26065 3415 26085 3435
rect 26065 3365 26085 3385
rect 26065 3315 26085 3335
rect 26065 3265 26085 3285
rect 26065 3215 26085 3235
rect 26065 3165 26085 3185
rect 26065 3115 26085 3135
rect 26065 3065 26085 3085
rect 26665 3515 26685 3535
rect 26665 3465 26685 3485
rect 26665 3415 26685 3435
rect 26665 3365 26685 3385
rect 26665 3315 26685 3335
rect 26665 3265 26685 3285
rect 26665 3215 26685 3235
rect 26665 3165 26685 3185
rect 26665 3115 26685 3135
rect 26665 3065 26685 3085
rect 27265 3515 27285 3535
rect 27265 3465 27285 3485
rect 27265 3415 27285 3435
rect 27265 3365 27285 3385
rect 27265 3315 27285 3335
rect 27265 3265 27285 3285
rect 27265 3215 27285 3235
rect 27265 3165 27285 3185
rect 27265 3115 27285 3135
rect 27265 3065 27285 3085
rect 27715 3515 27735 3535
rect 27715 3465 27735 3485
rect 27715 3415 27735 3435
rect 27715 3365 27735 3385
rect 27715 3315 27735 3335
rect 27715 3265 27735 3285
rect 27715 3215 27735 3235
rect 27715 3165 27735 3185
rect 27715 3115 27735 3135
rect 27715 3065 27735 3085
rect 28165 3515 28185 3535
rect 28165 3465 28185 3485
rect 28165 3415 28185 3435
rect 28165 3365 28185 3385
rect 28165 3315 28185 3335
rect 28165 3265 28185 3285
rect 28165 3215 28185 3235
rect 28165 3165 28185 3185
rect 28165 3115 28185 3135
rect 28165 3065 28185 3085
rect 28765 3515 28785 3535
rect 28765 3465 28785 3485
rect 28765 3415 28785 3435
rect 28765 3365 28785 3385
rect 28765 3315 28785 3335
rect 28765 3265 28785 3285
rect 28765 3215 28785 3235
rect 28765 3165 28785 3185
rect 28765 3115 28785 3135
rect 28765 3065 28785 3085
rect 29365 3515 29385 3535
rect 29365 3465 29385 3485
rect 29365 3415 29385 3435
rect 29365 3365 29385 3385
rect 29365 3315 29385 3335
rect 29365 3265 29385 3285
rect 29365 3215 29385 3235
rect 29365 3165 29385 3185
rect 29365 3115 29385 3135
rect 29365 3065 29385 3085
rect 29515 3515 29535 3535
rect 29515 3465 29535 3485
rect 29515 3415 29535 3435
rect 29515 3365 29535 3385
rect 29515 3315 29535 3335
rect 29515 3265 29535 3285
rect 29515 3215 29535 3235
rect 29515 3165 29535 3185
rect 29665 3415 29685 3435
rect 29665 3365 29685 3385
rect 29665 3315 29685 3335
rect 29665 3265 29685 3285
rect 29665 3215 29685 3235
rect 29665 3165 29685 3185
rect 29665 3115 29685 3135
rect 29665 3065 29685 3085
rect 29815 3515 29835 3535
rect 29815 3465 29835 3485
rect 29815 3415 29835 3435
rect 29815 3365 29835 3385
rect 29815 3315 29835 3335
rect 29815 3265 29835 3285
rect 29815 3215 29835 3235
rect 29815 3165 29835 3185
rect 29815 3115 29835 3135
rect 29815 3065 29835 3085
rect 29965 3415 29985 3435
rect 29965 3365 29985 3385
rect 29965 3315 29985 3335
rect 29965 3265 29985 3285
rect 29965 3215 29985 3235
rect 29965 3165 29985 3185
rect 29965 3115 29985 3135
rect 29965 3065 29985 3085
rect 30115 3515 30135 3535
rect 30115 3465 30135 3485
rect 30115 3415 30135 3435
rect 30115 3365 30135 3385
rect 30115 3315 30135 3335
rect 30115 3265 30135 3285
rect 30115 3215 30135 3235
rect 30115 3165 30135 3185
rect 30265 3415 30285 3435
rect 30265 3365 30285 3385
rect 30265 3315 30285 3335
rect 30265 3265 30285 3285
rect 30265 3215 30285 3235
rect 30265 3165 30285 3185
rect 30265 3115 30285 3135
rect 30265 3065 30285 3085
rect 30415 3515 30435 3535
rect 30415 3465 30435 3485
rect 30415 3415 30435 3435
rect 30415 3365 30435 3385
rect 30415 3315 30435 3335
rect 30415 3265 30435 3285
rect 30415 3215 30435 3235
rect 30415 3165 30435 3185
rect 30565 3415 30585 3435
rect 30565 3365 30585 3385
rect 30565 3315 30585 3335
rect 30565 3265 30585 3285
rect 30565 3215 30585 3235
rect 30565 3165 30585 3185
rect 30565 3115 30585 3135
rect 30565 3065 30585 3085
rect 30715 3515 30735 3535
rect 30715 3465 30735 3485
rect 30715 3415 30735 3435
rect 30715 3365 30735 3385
rect 30715 3315 30735 3335
rect 30715 3265 30735 3285
rect 30715 3215 30735 3235
rect 30715 3165 30735 3185
rect 30865 3415 30885 3435
rect 30865 3365 30885 3385
rect 30865 3315 30885 3335
rect 30865 3265 30885 3285
rect 30865 3215 30885 3235
rect 30865 3165 30885 3185
rect 30865 3115 30885 3135
rect 30865 3065 30885 3085
rect 31015 3515 31035 3535
rect 31015 3465 31035 3485
rect 31015 3415 31035 3435
rect 31015 3365 31035 3385
rect 31015 3315 31035 3335
rect 31015 3265 31035 3285
rect 31015 3215 31035 3235
rect 31015 3165 31035 3185
rect 31015 3115 31035 3135
rect 31015 3065 31035 3085
rect 31165 3415 31185 3435
rect 31165 3365 31185 3385
rect 31165 3315 31185 3335
rect 31165 3265 31185 3285
rect 31165 3215 31185 3235
rect 31165 3165 31185 3185
rect 31165 3115 31185 3135
rect 31165 3065 31185 3085
rect 31315 3515 31335 3535
rect 31315 3465 31335 3485
rect 31315 3415 31335 3435
rect 31315 3365 31335 3385
rect 31315 3315 31335 3335
rect 31315 3265 31335 3285
rect 31315 3215 31335 3235
rect 31315 3165 31335 3185
rect 31465 3515 31485 3535
rect 31465 3465 31485 3485
rect 31465 3415 31485 3435
rect 31465 3365 31485 3385
rect 31465 3315 31485 3335
rect 31465 3265 31485 3285
rect 31465 3215 31485 3235
rect 31465 3165 31485 3185
rect 31465 3115 31485 3135
rect 31465 3065 31485 3085
rect 32065 3515 32085 3535
rect 32065 3465 32085 3485
rect 32065 3415 32085 3435
rect 32065 3365 32085 3385
rect 32065 3315 32085 3335
rect 32065 3265 32085 3285
rect 32065 3215 32085 3235
rect 32065 3165 32085 3185
rect 32065 3115 32085 3135
rect 32065 3065 32085 3085
rect -635 2965 -615 2985
rect -35 2965 -15 2985
rect 4165 2965 4185 2985
rect 8365 2965 8385 2985
rect 8665 2965 8685 2985
rect 8965 2965 8985 2985
rect 9265 2965 9285 2985
rect 9565 2965 9585 2985
rect 9865 2965 9885 2985
rect 10165 2965 10185 2985
rect 10465 2965 10485 2985
rect 10765 2965 10785 2985
rect 11965 2965 11985 2985
rect 13165 2965 13185 2985
rect 14365 2965 14385 2985
rect 15565 2965 15585 2985
rect 20365 2965 20385 2985
rect 24565 2965 24585 2985
rect 28165 2965 28185 2985
rect 28765 2965 28785 2985
rect 32065 2965 32085 2985
rect -635 1665 -615 1685
rect -35 1665 -15 1685
rect 8365 1665 8385 1685
rect 10765 1665 10785 1685
rect 15565 1665 15585 1685
rect 17965 1665 17985 1685
rect 20365 1665 20385 1685
rect 24565 1665 24585 1685
rect 28765 1665 28785 1685
rect -635 1565 -615 1585
rect -635 1515 -615 1535
rect -635 1465 -615 1485
rect -635 1415 -615 1435
rect -635 1365 -615 1385
rect -635 1315 -615 1335
rect -635 1265 -615 1285
rect -635 1215 -615 1235
rect -635 1165 -615 1185
rect -635 1115 -615 1135
rect -635 1065 -615 1085
rect -635 1015 -615 1035
rect -635 965 -615 985
rect -635 915 -615 935
rect -485 1565 -465 1585
rect -485 1515 -465 1535
rect -485 1465 -465 1485
rect -485 1415 -465 1435
rect -485 1365 -465 1385
rect -485 1315 -465 1335
rect -485 1265 -465 1285
rect -485 1215 -465 1235
rect -485 1165 -465 1185
rect -485 1115 -465 1135
rect -485 1065 -465 1085
rect -485 1015 -465 1035
rect -485 965 -465 985
rect -485 915 -465 935
rect -335 1565 -315 1585
rect -335 1515 -315 1535
rect -335 1465 -315 1485
rect -335 1415 -315 1435
rect -335 1365 -315 1385
rect -335 1315 -315 1335
rect -335 1265 -315 1285
rect -335 1215 -315 1235
rect -335 1165 -315 1185
rect -335 1115 -315 1135
rect -335 1065 -315 1085
rect -335 1015 -315 1035
rect -335 965 -315 985
rect -335 915 -315 935
rect -185 1565 -165 1585
rect -185 1515 -165 1535
rect -185 1465 -165 1485
rect -185 1415 -165 1435
rect -185 1365 -165 1385
rect -185 1315 -165 1335
rect -185 1265 -165 1285
rect -185 1215 -165 1235
rect -185 1165 -165 1185
rect -185 1115 -165 1135
rect -185 1065 -165 1085
rect -185 1015 -165 1035
rect -185 965 -165 985
rect -185 915 -165 935
rect -35 1565 -15 1585
rect -35 1515 -15 1535
rect -35 1465 -15 1485
rect -35 1415 -15 1435
rect -35 1365 -15 1385
rect -35 1315 -15 1335
rect -35 1265 -15 1285
rect -35 1215 -15 1235
rect -35 1165 -15 1185
rect -35 1115 -15 1135
rect -35 1065 -15 1085
rect -35 1015 -15 1035
rect -35 965 -15 985
rect -35 915 -15 935
rect 1165 1565 1185 1585
rect 1165 1515 1185 1535
rect 1165 1465 1185 1485
rect 1165 1415 1185 1435
rect 1165 1365 1185 1385
rect 1165 1315 1185 1335
rect 1165 1265 1185 1285
rect 1165 1215 1185 1235
rect 1165 1165 1185 1185
rect 1165 1115 1185 1135
rect 1165 1065 1185 1085
rect 1165 1015 1185 1035
rect 1165 965 1185 985
rect 1165 915 1185 935
rect 1465 1465 1485 1485
rect 1465 1415 1485 1435
rect 1465 1365 1485 1385
rect 1465 1315 1485 1335
rect 1465 1265 1485 1285
rect 1465 1215 1485 1235
rect 1465 1165 1485 1185
rect 1465 1115 1485 1135
rect 1465 1065 1485 1085
rect 1465 1015 1485 1035
rect 1465 965 1485 985
rect 1465 915 1485 935
rect 1765 1565 1785 1585
rect 1765 1515 1785 1535
rect 1765 1465 1785 1485
rect 1765 1415 1785 1435
rect 1765 1365 1785 1385
rect 1765 1315 1785 1335
rect 1765 1265 1785 1285
rect 1765 1215 1785 1235
rect 1765 1165 1785 1185
rect 1765 1115 1785 1135
rect 1765 1065 1785 1085
rect 1765 1015 1785 1035
rect 2065 1465 2085 1485
rect 2065 1415 2085 1435
rect 2065 1365 2085 1385
rect 2065 1315 2085 1335
rect 2065 1265 2085 1285
rect 2065 1215 2085 1235
rect 2065 1165 2085 1185
rect 2065 1115 2085 1135
rect 2065 1065 2085 1085
rect 2065 1015 2085 1035
rect 2065 965 2085 985
rect 2065 915 2085 935
rect 2365 1565 2385 1585
rect 2365 1515 2385 1535
rect 2365 1465 2385 1485
rect 2365 1415 2385 1435
rect 2365 1365 2385 1385
rect 2365 1315 2385 1335
rect 2365 1265 2385 1285
rect 2365 1215 2385 1235
rect 2365 1165 2385 1185
rect 2365 1115 2385 1135
rect 2365 1065 2385 1085
rect 2365 1015 2385 1035
rect 2665 1465 2685 1485
rect 2665 1415 2685 1435
rect 2665 1365 2685 1385
rect 2665 1315 2685 1335
rect 2665 1265 2685 1285
rect 2665 1215 2685 1235
rect 2665 1165 2685 1185
rect 2665 1115 2685 1135
rect 2665 1065 2685 1085
rect 2665 1015 2685 1035
rect 2665 965 2685 985
rect 2665 915 2685 935
rect 2965 1565 2985 1585
rect 2965 1515 2985 1535
rect 2965 1465 2985 1485
rect 2965 1415 2985 1435
rect 2965 1365 2985 1385
rect 2965 1315 2985 1335
rect 2965 1265 2985 1285
rect 2965 1215 2985 1235
rect 2965 1165 2985 1185
rect 2965 1115 2985 1135
rect 2965 1065 2985 1085
rect 2965 1015 2985 1035
rect 3265 1465 3285 1485
rect 3265 1415 3285 1435
rect 3265 1365 3285 1385
rect 3265 1315 3285 1335
rect 3265 1265 3285 1285
rect 3265 1215 3285 1235
rect 3265 1165 3285 1185
rect 3265 1115 3285 1135
rect 3265 1065 3285 1085
rect 3265 1015 3285 1035
rect 3265 965 3285 985
rect 3265 915 3285 935
rect 3565 1565 3585 1585
rect 3565 1515 3585 1535
rect 3565 1465 3585 1485
rect 3565 1415 3585 1435
rect 3565 1365 3585 1385
rect 3565 1315 3585 1335
rect 3565 1265 3585 1285
rect 3565 1215 3585 1235
rect 3565 1165 3585 1185
rect 3565 1115 3585 1135
rect 3565 1065 3585 1085
rect 3565 1015 3585 1035
rect 3565 965 3585 985
rect 3565 915 3585 935
rect 3715 1465 3735 1485
rect 3715 1415 3735 1435
rect 3715 1365 3735 1385
rect 3715 1315 3735 1335
rect 3715 1265 3735 1285
rect 3715 1215 3735 1235
rect 3715 1165 3735 1185
rect 3715 1115 3735 1135
rect 3715 1065 3735 1085
rect 3715 1015 3735 1035
rect 3715 965 3735 985
rect 3715 915 3735 935
rect 3865 1565 3885 1585
rect 3865 1515 3885 1535
rect 3865 1465 3885 1485
rect 3865 1415 3885 1435
rect 3865 1365 3885 1385
rect 3865 1315 3885 1335
rect 3865 1265 3885 1285
rect 3865 1215 3885 1235
rect 3865 1165 3885 1185
rect 3865 1115 3885 1135
rect 3865 1065 3885 1085
rect 3865 1015 3885 1035
rect 4015 1465 4035 1485
rect 4015 1415 4035 1435
rect 4015 1365 4035 1385
rect 4015 1315 4035 1335
rect 4015 1265 4035 1285
rect 4015 1215 4035 1235
rect 4015 1165 4035 1185
rect 4015 1115 4035 1135
rect 4015 1065 4035 1085
rect 4015 1015 4035 1035
rect 4015 965 4035 985
rect 4015 915 4035 935
rect 4165 1565 4185 1585
rect 4165 1515 4185 1535
rect 4165 1465 4185 1485
rect 4165 1415 4185 1435
rect 4165 1365 4185 1385
rect 4165 1315 4185 1335
rect 4165 1265 4185 1285
rect 4165 1215 4185 1235
rect 4165 1165 4185 1185
rect 4165 1115 4185 1135
rect 4165 1065 4185 1085
rect 4165 1015 4185 1035
rect 4165 965 4185 985
rect 4165 915 4185 935
rect 4315 1465 4335 1485
rect 4315 1415 4335 1435
rect 4315 1365 4335 1385
rect 4315 1315 4335 1335
rect 4315 1265 4335 1285
rect 4315 1215 4335 1235
rect 4315 1165 4335 1185
rect 4315 1115 4335 1135
rect 4315 1065 4335 1085
rect 4315 1015 4335 1035
rect 4315 965 4335 985
rect 4315 915 4335 935
rect 4465 1565 4485 1585
rect 4465 1515 4485 1535
rect 4465 1465 4485 1485
rect 4465 1415 4485 1435
rect 4465 1365 4485 1385
rect 4465 1315 4485 1335
rect 4465 1265 4485 1285
rect 4465 1215 4485 1235
rect 4465 1165 4485 1185
rect 4465 1115 4485 1135
rect 4465 1065 4485 1085
rect 4465 1015 4485 1035
rect 4615 1465 4635 1485
rect 4615 1415 4635 1435
rect 4615 1365 4635 1385
rect 4615 1315 4635 1335
rect 4615 1265 4635 1285
rect 4615 1215 4635 1235
rect 4615 1165 4635 1185
rect 4615 1115 4635 1135
rect 4615 1065 4635 1085
rect 4615 1015 4635 1035
rect 4615 965 4635 985
rect 4615 915 4635 935
rect 4765 1565 4785 1585
rect 4765 1515 4785 1535
rect 4765 1465 4785 1485
rect 4765 1415 4785 1435
rect 4765 1365 4785 1385
rect 4765 1315 4785 1335
rect 4765 1265 4785 1285
rect 4765 1215 4785 1235
rect 4765 1165 4785 1185
rect 4765 1115 4785 1135
rect 4765 1065 4785 1085
rect 4765 1015 4785 1035
rect 4765 965 4785 985
rect 4765 915 4785 935
rect 5065 1465 5085 1485
rect 5065 1415 5085 1435
rect 5065 1365 5085 1385
rect 5065 1315 5085 1335
rect 5065 1265 5085 1285
rect 5065 1215 5085 1235
rect 5065 1165 5085 1185
rect 5065 1115 5085 1135
rect 5065 1065 5085 1085
rect 5065 1015 5085 1035
rect 5065 965 5085 985
rect 5065 915 5085 935
rect 5365 1565 5385 1585
rect 5365 1515 5385 1535
rect 5365 1465 5385 1485
rect 5365 1415 5385 1435
rect 5365 1365 5385 1385
rect 5365 1315 5385 1335
rect 5365 1265 5385 1285
rect 5365 1215 5385 1235
rect 5365 1165 5385 1185
rect 5365 1115 5385 1135
rect 5365 1065 5385 1085
rect 5365 1015 5385 1035
rect 5665 1465 5685 1485
rect 5665 1415 5685 1435
rect 5665 1365 5685 1385
rect 5665 1315 5685 1335
rect 5665 1265 5685 1285
rect 5665 1215 5685 1235
rect 5665 1165 5685 1185
rect 5665 1115 5685 1135
rect 5665 1065 5685 1085
rect 5665 1015 5685 1035
rect 5665 965 5685 985
rect 5665 915 5685 935
rect 5965 1565 5985 1585
rect 5965 1515 5985 1535
rect 5965 1465 5985 1485
rect 5965 1415 5985 1435
rect 5965 1365 5985 1385
rect 5965 1315 5985 1335
rect 5965 1265 5985 1285
rect 5965 1215 5985 1235
rect 5965 1165 5985 1185
rect 5965 1115 5985 1135
rect 5965 1065 5985 1085
rect 5965 1015 5985 1035
rect 6265 1465 6285 1485
rect 6265 1415 6285 1435
rect 6265 1365 6285 1385
rect 6265 1315 6285 1335
rect 6265 1265 6285 1285
rect 6265 1215 6285 1235
rect 6265 1165 6285 1185
rect 6265 1115 6285 1135
rect 6265 1065 6285 1085
rect 6265 1015 6285 1035
rect 6265 965 6285 985
rect 6265 915 6285 935
rect 6565 1565 6585 1585
rect 6565 1515 6585 1535
rect 6565 1465 6585 1485
rect 6565 1415 6585 1435
rect 6565 1365 6585 1385
rect 6565 1315 6585 1335
rect 6565 1265 6585 1285
rect 6565 1215 6585 1235
rect 6565 1165 6585 1185
rect 6565 1115 6585 1135
rect 6565 1065 6585 1085
rect 6565 1015 6585 1035
rect 6865 1465 6885 1485
rect 6865 1415 6885 1435
rect 6865 1365 6885 1385
rect 6865 1315 6885 1335
rect 6865 1265 6885 1285
rect 6865 1215 6885 1235
rect 6865 1165 6885 1185
rect 6865 1115 6885 1135
rect 6865 1065 6885 1085
rect 6865 1015 6885 1035
rect 6865 965 6885 985
rect 6865 915 6885 935
rect 7165 1565 7185 1585
rect 7165 1515 7185 1535
rect 7165 1465 7185 1485
rect 7165 1415 7185 1435
rect 7165 1365 7185 1385
rect 7165 1315 7185 1335
rect 7165 1265 7185 1285
rect 7165 1215 7185 1235
rect 7165 1165 7185 1185
rect 7165 1115 7185 1135
rect 7165 1065 7185 1085
rect 7165 1015 7185 1035
rect 7165 965 7185 985
rect 7165 915 7185 935
rect 8365 1565 8385 1585
rect 8365 1515 8385 1535
rect 8365 1465 8385 1485
rect 8365 1415 8385 1435
rect 8365 1365 8385 1385
rect 8365 1315 8385 1335
rect 8365 1265 8385 1285
rect 8365 1215 8385 1235
rect 8365 1165 8385 1185
rect 8365 1115 8385 1135
rect 8365 1065 8385 1085
rect 8365 1015 8385 1035
rect 8365 965 8385 985
rect 8365 915 8385 935
rect 9565 1565 9585 1585
rect 9565 1515 9585 1535
rect 9565 1465 9585 1485
rect 9565 1415 9585 1435
rect 9565 1365 9585 1385
rect 9565 1315 9585 1335
rect 9565 1265 9585 1285
rect 9565 1215 9585 1235
rect 9565 1165 9585 1185
rect 9565 1115 9585 1135
rect 9565 1065 9585 1085
rect 9565 1015 9585 1035
rect 9565 965 9585 985
rect 9565 915 9585 935
rect 10765 1565 10785 1585
rect 10765 1515 10785 1535
rect 10765 1465 10785 1485
rect 10765 1415 10785 1435
rect 10765 1365 10785 1385
rect 10765 1315 10785 1335
rect 10765 1265 10785 1285
rect 10765 1215 10785 1235
rect 10765 1165 10785 1185
rect 10765 1115 10785 1135
rect 10765 1065 10785 1085
rect 10765 1015 10785 1035
rect 10765 965 10785 985
rect 10765 915 10785 935
rect 11965 1565 11985 1585
rect 11965 1515 11985 1535
rect 11965 1465 11985 1485
rect 11965 1415 11985 1435
rect 11965 1365 11985 1385
rect 11965 1315 11985 1335
rect 11965 1265 11985 1285
rect 11965 1215 11985 1235
rect 11965 1165 11985 1185
rect 11965 1115 11985 1135
rect 11965 1065 11985 1085
rect 11965 1015 11985 1035
rect 11965 965 11985 985
rect 11965 915 11985 935
rect 12265 1465 12285 1485
rect 12265 1415 12285 1435
rect 12265 1365 12285 1385
rect 12265 1315 12285 1335
rect 12265 1265 12285 1285
rect 12265 1215 12285 1235
rect 12265 1165 12285 1185
rect 12265 1115 12285 1135
rect 12265 1065 12285 1085
rect 12265 1015 12285 1035
rect 12265 965 12285 985
rect 12265 915 12285 935
rect 12565 1565 12585 1585
rect 12565 1515 12585 1535
rect 12565 1465 12585 1485
rect 12565 1415 12585 1435
rect 12565 1365 12585 1385
rect 12565 1315 12585 1335
rect 12565 1265 12585 1285
rect 12565 1215 12585 1235
rect 12565 1165 12585 1185
rect 12565 1115 12585 1135
rect 12565 1065 12585 1085
rect 12565 1015 12585 1035
rect 12865 1465 12885 1485
rect 12865 1415 12885 1435
rect 12865 1365 12885 1385
rect 12865 1315 12885 1335
rect 12865 1265 12885 1285
rect 12865 1215 12885 1235
rect 12865 1165 12885 1185
rect 12865 1115 12885 1135
rect 12865 1065 12885 1085
rect 12865 1015 12885 1035
rect 12865 965 12885 985
rect 12865 915 12885 935
rect 13165 1565 13185 1585
rect 13165 1515 13185 1535
rect 13165 1465 13185 1485
rect 13165 1415 13185 1435
rect 13165 1365 13185 1385
rect 13165 1315 13185 1335
rect 13165 1265 13185 1285
rect 13165 1215 13185 1235
rect 13165 1165 13185 1185
rect 13165 1115 13185 1135
rect 13165 1065 13185 1085
rect 13165 1015 13185 1035
rect 13465 1465 13485 1485
rect 13465 1415 13485 1435
rect 13465 1365 13485 1385
rect 13465 1315 13485 1335
rect 13465 1265 13485 1285
rect 13465 1215 13485 1235
rect 13465 1165 13485 1185
rect 13465 1115 13485 1135
rect 13465 1065 13485 1085
rect 13465 1015 13485 1035
rect 13465 965 13485 985
rect 13465 915 13485 935
rect 13765 1565 13785 1585
rect 13765 1515 13785 1535
rect 13765 1465 13785 1485
rect 13765 1415 13785 1435
rect 13765 1365 13785 1385
rect 13765 1315 13785 1335
rect 13765 1265 13785 1285
rect 13765 1215 13785 1235
rect 13765 1165 13785 1185
rect 13765 1115 13785 1135
rect 13765 1065 13785 1085
rect 13765 1015 13785 1035
rect 14065 1465 14085 1485
rect 14065 1415 14085 1435
rect 14065 1365 14085 1385
rect 14065 1315 14085 1335
rect 14065 1265 14085 1285
rect 14065 1215 14085 1235
rect 14065 1165 14085 1185
rect 14065 1115 14085 1135
rect 14065 1065 14085 1085
rect 14065 1015 14085 1035
rect 14065 965 14085 985
rect 14065 915 14085 935
rect 14365 1565 14385 1585
rect 14365 1515 14385 1535
rect 14365 1465 14385 1485
rect 14365 1415 14385 1435
rect 14365 1365 14385 1385
rect 14365 1315 14385 1335
rect 14365 1265 14385 1285
rect 14365 1215 14385 1235
rect 14365 1165 14385 1185
rect 14365 1115 14385 1135
rect 14365 1065 14385 1085
rect 14365 1015 14385 1035
rect 14365 965 14385 985
rect 14365 915 14385 935
rect 15565 1565 15585 1585
rect 15565 1515 15585 1535
rect 15565 1465 15585 1485
rect 15565 1415 15585 1435
rect 15565 1365 15585 1385
rect 15565 1315 15585 1335
rect 15565 1265 15585 1285
rect 15565 1215 15585 1235
rect 15565 1165 15585 1185
rect 15565 1115 15585 1135
rect 15565 1065 15585 1085
rect 15565 1015 15585 1035
rect 15565 965 15585 985
rect 15565 915 15585 935
rect 16765 1565 16785 1585
rect 16765 1515 16785 1535
rect 16765 1465 16785 1485
rect 16765 1415 16785 1435
rect 16765 1365 16785 1385
rect 16765 1315 16785 1335
rect 16765 1265 16785 1285
rect 16765 1215 16785 1235
rect 16765 1165 16785 1185
rect 16765 1115 16785 1135
rect 16765 1065 16785 1085
rect 16765 1015 16785 1035
rect 16765 965 16785 985
rect 16765 915 16785 935
rect 17965 1565 17985 1585
rect 17965 1515 17985 1535
rect 17965 1465 17985 1485
rect 17965 1415 17985 1435
rect 17965 1365 17985 1385
rect 17965 1315 17985 1335
rect 17965 1265 17985 1285
rect 17965 1215 17985 1235
rect 17965 1165 17985 1185
rect 17965 1115 17985 1135
rect 17965 1065 17985 1085
rect 17965 1015 17985 1035
rect 17965 965 17985 985
rect 17965 915 17985 935
rect 19165 1565 19185 1585
rect 19165 1515 19185 1535
rect 19165 1465 19185 1485
rect 19165 1415 19185 1435
rect 19165 1365 19185 1385
rect 19165 1315 19185 1335
rect 19165 1265 19185 1285
rect 19165 1215 19185 1235
rect 19165 1165 19185 1185
rect 19165 1115 19185 1135
rect 19165 1065 19185 1085
rect 19165 1015 19185 1035
rect 19165 965 19185 985
rect 19165 915 19185 935
rect 20365 1565 20385 1585
rect 20365 1515 20385 1535
rect 20365 1465 20385 1485
rect 20365 1415 20385 1435
rect 20365 1365 20385 1385
rect 20365 1315 20385 1335
rect 20365 1265 20385 1285
rect 20365 1215 20385 1235
rect 20365 1165 20385 1185
rect 20365 1115 20385 1135
rect 20365 1065 20385 1085
rect 20365 1015 20385 1035
rect 20365 965 20385 985
rect 20365 915 20385 935
rect 21565 1565 21585 1585
rect 21565 1515 21585 1535
rect 21565 1465 21585 1485
rect 21565 1415 21585 1435
rect 21565 1365 21585 1385
rect 21565 1315 21585 1335
rect 21565 1265 21585 1285
rect 21565 1215 21585 1235
rect 21565 1165 21585 1185
rect 21565 1115 21585 1135
rect 21565 1065 21585 1085
rect 21565 1015 21585 1035
rect 21565 965 21585 985
rect 21565 915 21585 935
rect 22465 1565 22485 1585
rect 22465 1515 22485 1535
rect 22465 1465 22485 1485
rect 22465 1415 22485 1435
rect 22465 1365 22485 1385
rect 22465 1315 22485 1335
rect 22465 1265 22485 1285
rect 22465 1215 22485 1235
rect 22465 1165 22485 1185
rect 22465 1115 22485 1135
rect 22465 1065 22485 1085
rect 22465 1015 22485 1035
rect 22465 965 22485 985
rect 22465 915 22485 935
rect 23365 1565 23385 1585
rect 23365 1515 23385 1535
rect 23365 1465 23385 1485
rect 23365 1415 23385 1435
rect 23365 1365 23385 1385
rect 23365 1315 23385 1335
rect 23365 1265 23385 1285
rect 23365 1215 23385 1235
rect 23365 1165 23385 1185
rect 23365 1115 23385 1135
rect 23365 1065 23385 1085
rect 23365 1015 23385 1035
rect 23365 965 23385 985
rect 23365 915 23385 935
rect 24565 1565 24585 1585
rect 24565 1515 24585 1535
rect 24565 1465 24585 1485
rect 24565 1415 24585 1435
rect 24565 1365 24585 1385
rect 24565 1315 24585 1335
rect 24565 1265 24585 1285
rect 24565 1215 24585 1235
rect 24565 1165 24585 1185
rect 24565 1115 24585 1135
rect 24565 1065 24585 1085
rect 24565 1015 24585 1035
rect 24565 965 24585 985
rect 24565 915 24585 935
rect 25765 1565 25785 1585
rect 25765 1515 25785 1535
rect 25765 1465 25785 1485
rect 25765 1415 25785 1435
rect 25765 1365 25785 1385
rect 25765 1315 25785 1335
rect 25765 1265 25785 1285
rect 25765 1215 25785 1235
rect 25765 1165 25785 1185
rect 25765 1115 25785 1135
rect 25765 1065 25785 1085
rect 25765 1015 25785 1035
rect 25765 965 25785 985
rect 25765 915 25785 935
rect 26665 1565 26685 1585
rect 26665 1515 26685 1535
rect 26665 1465 26685 1485
rect 26665 1415 26685 1435
rect 26665 1365 26685 1385
rect 26665 1315 26685 1335
rect 26665 1265 26685 1285
rect 26665 1215 26685 1235
rect 26665 1165 26685 1185
rect 26665 1115 26685 1135
rect 26665 1065 26685 1085
rect 26665 1015 26685 1035
rect 26665 965 26685 985
rect 26665 915 26685 935
rect 27565 1565 27585 1585
rect 27565 1515 27585 1535
rect 27565 1465 27585 1485
rect 27565 1415 27585 1435
rect 27565 1365 27585 1385
rect 27565 1315 27585 1335
rect 27565 1265 27585 1285
rect 27565 1215 27585 1235
rect 27565 1165 27585 1185
rect 27565 1115 27585 1135
rect 27565 1065 27585 1085
rect 27565 1015 27585 1035
rect 27565 965 27585 985
rect 27565 915 27585 935
rect 28765 1565 28785 1585
rect 28765 1515 28785 1535
rect 28765 1465 28785 1485
rect 28765 1415 28785 1435
rect 28765 1365 28785 1385
rect 28765 1315 28785 1335
rect 28765 1265 28785 1285
rect 28765 1215 28785 1235
rect 28765 1165 28785 1185
rect 28765 1115 28785 1135
rect 28765 1065 28785 1085
rect 28765 1015 28785 1035
rect 28765 965 28785 985
rect 28765 915 28785 935
rect -485 815 -465 835
rect -185 815 -165 835
rect 115 815 135 835
rect 415 815 435 835
rect 715 815 735 835
rect 1015 815 1035 835
rect 1315 815 1335 835
rect 1615 815 1635 835
rect 1915 815 1935 835
rect 2215 815 2235 835
rect 2515 815 2535 835
rect 2815 815 2835 835
rect 3115 815 3135 835
rect 3415 815 3435 835
rect 3715 815 3735 835
rect 4015 815 4035 835
rect 4315 815 4335 835
rect 4615 815 4635 835
rect 4915 815 4935 835
rect 5215 815 5235 835
rect 5515 815 5535 835
rect 5815 815 5835 835
rect 6115 815 6135 835
rect 6415 815 6435 835
rect 6715 815 6735 835
rect 7015 815 7035 835
rect 7315 815 7335 835
rect 7615 815 7635 835
rect 7915 815 7935 835
rect 8215 815 8235 835
rect 8515 815 8535 835
rect 8815 815 8835 835
rect 9115 815 9135 835
rect 9415 815 9435 835
rect 9715 815 9735 835
rect 10015 815 10035 835
rect 10315 815 10335 835
rect 10615 815 10635 835
rect 10915 815 10935 835
rect 11215 815 11235 835
rect 11515 815 11535 835
rect 11815 815 11835 835
rect 12115 815 12135 835
rect 12415 815 12435 835
rect 12715 815 12735 835
rect 13015 815 13035 835
rect 13315 815 13335 835
rect 13615 815 13635 835
rect 13915 815 13935 835
rect 14215 815 14235 835
rect 14515 815 14535 835
rect 14815 815 14835 835
rect 15115 815 15135 835
rect 15415 815 15435 835
rect 15715 815 15735 835
rect 16015 815 16035 835
rect 16315 815 16335 835
rect 16615 815 16635 835
rect 16915 815 16935 835
rect 17215 815 17235 835
rect 17515 815 17535 835
rect 17815 815 17835 835
rect 18115 815 18135 835
rect 18415 815 18435 835
rect 18715 815 18735 835
rect 19015 815 19035 835
rect 19315 815 19335 835
rect 19615 815 19635 835
rect 19915 815 19935 835
rect 20215 815 20235 835
rect 20515 815 20535 835
rect 20815 815 20835 835
rect 21115 815 21135 835
rect 21415 815 21435 835
rect 21715 815 21735 835
rect 22015 815 22035 835
rect 22315 815 22335 835
rect 22615 815 22635 835
rect 22915 815 22935 835
rect 23215 815 23235 835
rect 23515 815 23535 835
rect 23815 815 23835 835
rect 24115 815 24135 835
rect 24415 815 24435 835
rect 24715 815 24735 835
rect 25015 815 25035 835
rect 25315 815 25335 835
rect 25615 815 25635 835
rect 25915 815 25935 835
rect 26215 815 26235 835
rect 26515 815 26535 835
rect 26815 815 26835 835
rect 27115 815 27135 835
rect 27415 815 27435 835
rect 27715 815 27735 835
rect 28015 815 28035 835
rect 28315 815 28335 835
rect 28615 815 28635 835
rect -635 715 -615 735
rect -635 665 -615 685
rect -635 615 -615 635
rect -635 565 -615 585
rect -635 515 -615 535
rect -635 465 -615 485
rect -635 415 -615 435
rect -635 365 -615 385
rect -635 315 -615 335
rect -635 265 -615 285
rect -635 215 -615 235
rect -635 165 -615 185
rect -635 115 -615 135
rect -635 65 -615 85
rect -485 715 -465 735
rect -485 665 -465 685
rect -485 615 -465 635
rect -485 565 -465 585
rect -485 515 -465 535
rect -485 465 -465 485
rect -485 415 -465 435
rect -485 365 -465 385
rect -485 315 -465 335
rect -485 265 -465 285
rect -485 215 -465 235
rect -485 165 -465 185
rect -485 115 -465 135
rect -485 65 -465 85
rect -335 715 -315 735
rect -335 665 -315 685
rect -335 615 -315 635
rect -335 565 -315 585
rect -335 515 -315 535
rect -335 465 -315 485
rect -335 415 -315 435
rect -335 365 -315 385
rect -335 315 -315 335
rect -335 265 -315 285
rect -335 215 -315 235
rect -335 165 -315 185
rect -335 115 -315 135
rect -335 65 -315 85
rect -185 715 -165 735
rect -185 665 -165 685
rect -185 615 -165 635
rect -185 565 -165 585
rect -185 515 -165 535
rect -185 465 -165 485
rect -185 415 -165 435
rect -185 365 -165 385
rect -185 315 -165 335
rect -185 265 -165 285
rect -185 215 -165 235
rect -185 165 -165 185
rect -185 115 -165 135
rect -185 65 -165 85
rect -35 715 -15 735
rect -35 665 -15 685
rect -35 615 -15 635
rect -35 565 -15 585
rect -35 515 -15 535
rect -35 465 -15 485
rect -35 415 -15 435
rect -35 365 -15 385
rect -35 315 -15 335
rect -35 265 -15 285
rect -35 215 -15 235
rect -35 165 -15 185
rect -35 115 -15 135
rect -35 65 -15 85
rect 1165 715 1185 735
rect 1165 665 1185 685
rect 1165 615 1185 635
rect 1165 565 1185 585
rect 1165 515 1185 535
rect 1165 465 1185 485
rect 1165 415 1185 435
rect 1165 365 1185 385
rect 1165 315 1185 335
rect 1165 265 1185 285
rect 1165 215 1185 235
rect 1165 165 1185 185
rect 1165 115 1185 135
rect 1165 65 1185 85
rect 1465 715 1485 735
rect 1465 665 1485 685
rect 1465 615 1485 635
rect 1465 565 1485 585
rect 1465 515 1485 535
rect 1465 465 1485 485
rect 1465 415 1485 435
rect 1465 365 1485 385
rect 1465 315 1485 335
rect 1465 265 1485 285
rect 1465 215 1485 235
rect 1465 165 1485 185
rect 1765 615 1785 635
rect 1765 565 1785 585
rect 1765 515 1785 535
rect 1765 465 1785 485
rect 1765 415 1785 435
rect 1765 365 1785 385
rect 1765 315 1785 335
rect 1765 265 1785 285
rect 1765 215 1785 235
rect 1765 165 1785 185
rect 1765 115 1785 135
rect 1765 65 1785 85
rect 2065 715 2085 735
rect 2065 665 2085 685
rect 2065 615 2085 635
rect 2065 565 2085 585
rect 2065 515 2085 535
rect 2065 465 2085 485
rect 2065 415 2085 435
rect 2065 365 2085 385
rect 2065 315 2085 335
rect 2065 265 2085 285
rect 2065 215 2085 235
rect 2065 165 2085 185
rect 2365 615 2385 635
rect 2365 565 2385 585
rect 2365 515 2385 535
rect 2365 465 2385 485
rect 2365 415 2385 435
rect 2365 365 2385 385
rect 2365 315 2385 335
rect 2365 265 2385 285
rect 2365 215 2385 235
rect 2365 165 2385 185
rect 2365 115 2385 135
rect 2365 65 2385 85
rect 2665 715 2685 735
rect 2665 665 2685 685
rect 2665 615 2685 635
rect 2665 565 2685 585
rect 2665 515 2685 535
rect 2665 465 2685 485
rect 2665 415 2685 435
rect 2665 365 2685 385
rect 2665 315 2685 335
rect 2665 265 2685 285
rect 2665 215 2685 235
rect 2665 165 2685 185
rect 2965 615 2985 635
rect 2965 565 2985 585
rect 2965 515 2985 535
rect 2965 465 2985 485
rect 2965 415 2985 435
rect 2965 365 2985 385
rect 2965 315 2985 335
rect 2965 265 2985 285
rect 2965 215 2985 235
rect 2965 165 2985 185
rect 2965 115 2985 135
rect 2965 65 2985 85
rect 3265 715 3285 735
rect 3265 665 3285 685
rect 3265 615 3285 635
rect 3265 565 3285 585
rect 3265 515 3285 535
rect 3265 465 3285 485
rect 3265 415 3285 435
rect 3265 365 3285 385
rect 3265 315 3285 335
rect 3265 265 3285 285
rect 3265 215 3285 235
rect 3265 165 3285 185
rect 3565 715 3585 735
rect 3565 665 3585 685
rect 3565 615 3585 635
rect 3565 565 3585 585
rect 3565 515 3585 535
rect 3565 465 3585 485
rect 3565 415 3585 435
rect 3565 365 3585 385
rect 3565 315 3585 335
rect 3565 265 3585 285
rect 3565 215 3585 235
rect 3565 165 3585 185
rect 3565 115 3585 135
rect 3565 65 3585 85
rect 3715 715 3735 735
rect 3715 665 3735 685
rect 3715 615 3735 635
rect 3715 565 3735 585
rect 3715 515 3735 535
rect 3715 465 3735 485
rect 3715 415 3735 435
rect 3715 365 3735 385
rect 3715 315 3735 335
rect 3715 265 3735 285
rect 3715 215 3735 235
rect 3715 165 3735 185
rect 3865 615 3885 635
rect 3865 565 3885 585
rect 3865 515 3885 535
rect 3865 465 3885 485
rect 3865 415 3885 435
rect 3865 365 3885 385
rect 3865 315 3885 335
rect 3865 265 3885 285
rect 3865 215 3885 235
rect 3865 165 3885 185
rect 3865 115 3885 135
rect 3865 65 3885 85
rect 4015 715 4035 735
rect 4015 665 4035 685
rect 4015 615 4035 635
rect 4015 565 4035 585
rect 4015 515 4035 535
rect 4015 465 4035 485
rect 4015 415 4035 435
rect 4015 365 4035 385
rect 4015 315 4035 335
rect 4015 265 4035 285
rect 4015 215 4035 235
rect 4015 165 4035 185
rect 4165 715 4185 735
rect 4165 665 4185 685
rect 4165 615 4185 635
rect 4165 565 4185 585
rect 4165 515 4185 535
rect 4165 465 4185 485
rect 4165 415 4185 435
rect 4165 365 4185 385
rect 4165 315 4185 335
rect 4165 265 4185 285
rect 4165 215 4185 235
rect 4165 165 4185 185
rect 4165 115 4185 135
rect 4165 65 4185 85
rect 4315 715 4335 735
rect 4315 665 4335 685
rect 4315 615 4335 635
rect 4315 565 4335 585
rect 4315 515 4335 535
rect 4315 465 4335 485
rect 4315 415 4335 435
rect 4315 365 4335 385
rect 4315 315 4335 335
rect 4315 265 4335 285
rect 4315 215 4335 235
rect 4315 165 4335 185
rect 4465 615 4485 635
rect 4465 565 4485 585
rect 4465 515 4485 535
rect 4465 465 4485 485
rect 4465 415 4485 435
rect 4465 365 4485 385
rect 4465 315 4485 335
rect 4465 265 4485 285
rect 4465 215 4485 235
rect 4465 165 4485 185
rect 4465 115 4485 135
rect 4465 65 4485 85
rect 4615 715 4635 735
rect 4615 665 4635 685
rect 4615 615 4635 635
rect 4615 565 4635 585
rect 4615 515 4635 535
rect 4615 465 4635 485
rect 4615 415 4635 435
rect 4615 365 4635 385
rect 4615 315 4635 335
rect 4615 265 4635 285
rect 4615 215 4635 235
rect 4615 165 4635 185
rect 4765 715 4785 735
rect 4765 665 4785 685
rect 4765 615 4785 635
rect 4765 565 4785 585
rect 4765 515 4785 535
rect 4765 465 4785 485
rect 4765 415 4785 435
rect 4765 365 4785 385
rect 4765 315 4785 335
rect 4765 265 4785 285
rect 4765 215 4785 235
rect 4765 165 4785 185
rect 4765 115 4785 135
rect 4765 65 4785 85
rect 5065 715 5085 735
rect 5065 665 5085 685
rect 5065 615 5085 635
rect 5065 565 5085 585
rect 5065 515 5085 535
rect 5065 465 5085 485
rect 5065 415 5085 435
rect 5065 365 5085 385
rect 5065 315 5085 335
rect 5065 265 5085 285
rect 5065 215 5085 235
rect 5065 165 5085 185
rect 5365 615 5385 635
rect 5365 565 5385 585
rect 5365 515 5385 535
rect 5365 465 5385 485
rect 5365 415 5385 435
rect 5365 365 5385 385
rect 5365 315 5385 335
rect 5365 265 5385 285
rect 5365 215 5385 235
rect 5365 165 5385 185
rect 5365 115 5385 135
rect 5365 65 5385 85
rect 5665 715 5685 735
rect 5665 665 5685 685
rect 5665 615 5685 635
rect 5665 565 5685 585
rect 5665 515 5685 535
rect 5665 465 5685 485
rect 5665 415 5685 435
rect 5665 365 5685 385
rect 5665 315 5685 335
rect 5665 265 5685 285
rect 5665 215 5685 235
rect 5665 165 5685 185
rect 5965 615 5985 635
rect 5965 565 5985 585
rect 5965 515 5985 535
rect 5965 465 5985 485
rect 5965 415 5985 435
rect 5965 365 5985 385
rect 5965 315 5985 335
rect 5965 265 5985 285
rect 5965 215 5985 235
rect 5965 165 5985 185
rect 5965 115 5985 135
rect 5965 65 5985 85
rect 6265 715 6285 735
rect 6265 665 6285 685
rect 6265 615 6285 635
rect 6265 565 6285 585
rect 6265 515 6285 535
rect 6265 465 6285 485
rect 6265 415 6285 435
rect 6265 365 6285 385
rect 6265 315 6285 335
rect 6265 265 6285 285
rect 6265 215 6285 235
rect 6265 165 6285 185
rect 6565 615 6585 635
rect 6565 565 6585 585
rect 6565 515 6585 535
rect 6565 465 6585 485
rect 6565 415 6585 435
rect 6565 365 6585 385
rect 6565 315 6585 335
rect 6565 265 6585 285
rect 6565 215 6585 235
rect 6565 165 6585 185
rect 6565 115 6585 135
rect 6565 65 6585 85
rect 6865 715 6885 735
rect 6865 665 6885 685
rect 6865 615 6885 635
rect 6865 565 6885 585
rect 6865 515 6885 535
rect 6865 465 6885 485
rect 6865 415 6885 435
rect 6865 365 6885 385
rect 6865 315 6885 335
rect 6865 265 6885 285
rect 6865 215 6885 235
rect 6865 165 6885 185
rect 7165 715 7185 735
rect 7165 665 7185 685
rect 7165 615 7185 635
rect 7165 565 7185 585
rect 7165 515 7185 535
rect 7165 465 7185 485
rect 7165 415 7185 435
rect 7165 365 7185 385
rect 7165 315 7185 335
rect 7165 265 7185 285
rect 7165 215 7185 235
rect 7165 165 7185 185
rect 7165 115 7185 135
rect 7165 65 7185 85
rect 8365 715 8385 735
rect 8365 665 8385 685
rect 8365 615 8385 635
rect 8365 565 8385 585
rect 8365 515 8385 535
rect 8365 465 8385 485
rect 8365 415 8385 435
rect 8365 365 8385 385
rect 8365 315 8385 335
rect 8365 265 8385 285
rect 8365 215 8385 235
rect 8365 165 8385 185
rect 8365 115 8385 135
rect 8365 65 8385 85
rect 9565 715 9585 735
rect 9565 665 9585 685
rect 9565 615 9585 635
rect 9565 565 9585 585
rect 9565 515 9585 535
rect 9565 465 9585 485
rect 9565 415 9585 435
rect 9565 365 9585 385
rect 9565 315 9585 335
rect 9565 265 9585 285
rect 9565 215 9585 235
rect 9565 165 9585 185
rect 9565 115 9585 135
rect 9565 65 9585 85
rect 10765 715 10785 735
rect 10765 665 10785 685
rect 10765 615 10785 635
rect 10765 565 10785 585
rect 10765 515 10785 535
rect 10765 465 10785 485
rect 10765 415 10785 435
rect 10765 365 10785 385
rect 10765 315 10785 335
rect 10765 265 10785 285
rect 10765 215 10785 235
rect 10765 165 10785 185
rect 10765 115 10785 135
rect 10765 65 10785 85
rect 11965 715 11985 735
rect 11965 665 11985 685
rect 11965 615 11985 635
rect 11965 565 11985 585
rect 11965 515 11985 535
rect 11965 465 11985 485
rect 11965 415 11985 435
rect 11965 365 11985 385
rect 11965 315 11985 335
rect 11965 265 11985 285
rect 11965 215 11985 235
rect 11965 165 11985 185
rect 11965 115 11985 135
rect 11965 65 11985 85
rect 12265 715 12285 735
rect 12265 665 12285 685
rect 12265 615 12285 635
rect 12265 565 12285 585
rect 12265 515 12285 535
rect 12265 465 12285 485
rect 12265 415 12285 435
rect 12265 365 12285 385
rect 12265 315 12285 335
rect 12265 265 12285 285
rect 12265 215 12285 235
rect 12265 165 12285 185
rect 12565 615 12585 635
rect 12565 565 12585 585
rect 12565 515 12585 535
rect 12565 465 12585 485
rect 12565 415 12585 435
rect 12565 365 12585 385
rect 12565 315 12585 335
rect 12565 265 12585 285
rect 12565 215 12585 235
rect 12565 165 12585 185
rect 12565 115 12585 135
rect 12565 65 12585 85
rect 12865 715 12885 735
rect 12865 665 12885 685
rect 12865 615 12885 635
rect 12865 565 12885 585
rect 12865 515 12885 535
rect 12865 465 12885 485
rect 12865 415 12885 435
rect 12865 365 12885 385
rect 12865 315 12885 335
rect 12865 265 12885 285
rect 12865 215 12885 235
rect 12865 165 12885 185
rect 13165 615 13185 635
rect 13165 565 13185 585
rect 13165 515 13185 535
rect 13165 465 13185 485
rect 13165 415 13185 435
rect 13165 365 13185 385
rect 13165 315 13185 335
rect 13165 265 13185 285
rect 13165 215 13185 235
rect 13165 165 13185 185
rect 13165 115 13185 135
rect 13165 65 13185 85
rect 13465 715 13485 735
rect 13465 665 13485 685
rect 13465 615 13485 635
rect 13465 565 13485 585
rect 13465 515 13485 535
rect 13465 465 13485 485
rect 13465 415 13485 435
rect 13465 365 13485 385
rect 13465 315 13485 335
rect 13465 265 13485 285
rect 13465 215 13485 235
rect 13465 165 13485 185
rect 13765 615 13785 635
rect 13765 565 13785 585
rect 13765 515 13785 535
rect 13765 465 13785 485
rect 13765 415 13785 435
rect 13765 365 13785 385
rect 13765 315 13785 335
rect 13765 265 13785 285
rect 13765 215 13785 235
rect 13765 165 13785 185
rect 13765 115 13785 135
rect 13765 65 13785 85
rect 14065 715 14085 735
rect 14065 665 14085 685
rect 14065 615 14085 635
rect 14065 565 14085 585
rect 14065 515 14085 535
rect 14065 465 14085 485
rect 14065 415 14085 435
rect 14065 365 14085 385
rect 14065 315 14085 335
rect 14065 265 14085 285
rect 14065 215 14085 235
rect 14065 165 14085 185
rect 14365 715 14385 735
rect 14365 665 14385 685
rect 14365 615 14385 635
rect 14365 565 14385 585
rect 14365 515 14385 535
rect 14365 465 14385 485
rect 14365 415 14385 435
rect 14365 365 14385 385
rect 14365 315 14385 335
rect 14365 265 14385 285
rect 14365 215 14385 235
rect 14365 165 14385 185
rect 14365 115 14385 135
rect 14365 65 14385 85
rect 15565 715 15585 735
rect 15565 665 15585 685
rect 15565 615 15585 635
rect 15565 565 15585 585
rect 15565 515 15585 535
rect 15565 465 15585 485
rect 15565 415 15585 435
rect 15565 365 15585 385
rect 15565 315 15585 335
rect 15565 265 15585 285
rect 15565 215 15585 235
rect 15565 165 15585 185
rect 15565 115 15585 135
rect 15565 65 15585 85
rect 16765 715 16785 735
rect 16765 665 16785 685
rect 16765 615 16785 635
rect 16765 565 16785 585
rect 16765 515 16785 535
rect 16765 465 16785 485
rect 16765 415 16785 435
rect 16765 365 16785 385
rect 16765 315 16785 335
rect 16765 265 16785 285
rect 16765 215 16785 235
rect 16765 165 16785 185
rect 16765 115 16785 135
rect 16765 65 16785 85
rect 17965 715 17985 735
rect 17965 665 17985 685
rect 17965 615 17985 635
rect 17965 565 17985 585
rect 17965 515 17985 535
rect 17965 465 17985 485
rect 17965 415 17985 435
rect 17965 365 17985 385
rect 17965 315 17985 335
rect 17965 265 17985 285
rect 17965 215 17985 235
rect 17965 165 17985 185
rect 17965 115 17985 135
rect 17965 65 17985 85
rect 19165 715 19185 735
rect 19165 665 19185 685
rect 19165 615 19185 635
rect 19165 565 19185 585
rect 19165 515 19185 535
rect 19165 465 19185 485
rect 19165 415 19185 435
rect 19165 365 19185 385
rect 19165 315 19185 335
rect 19165 265 19185 285
rect 19165 215 19185 235
rect 19165 165 19185 185
rect 19165 115 19185 135
rect 19165 65 19185 85
rect 20365 715 20385 735
rect 20365 665 20385 685
rect 20365 615 20385 635
rect 20365 565 20385 585
rect 20365 515 20385 535
rect 20365 465 20385 485
rect 20365 415 20385 435
rect 20365 365 20385 385
rect 20365 315 20385 335
rect 20365 265 20385 285
rect 20365 215 20385 235
rect 20365 165 20385 185
rect 20365 115 20385 135
rect 20365 65 20385 85
rect 21565 715 21585 735
rect 21565 665 21585 685
rect 21565 615 21585 635
rect 21565 565 21585 585
rect 21565 515 21585 535
rect 21565 465 21585 485
rect 21565 415 21585 435
rect 21565 365 21585 385
rect 21565 315 21585 335
rect 21565 265 21585 285
rect 21565 215 21585 235
rect 21565 165 21585 185
rect 21565 115 21585 135
rect 21565 65 21585 85
rect 22465 715 22485 735
rect 22465 665 22485 685
rect 22465 615 22485 635
rect 22465 565 22485 585
rect 22465 515 22485 535
rect 22465 465 22485 485
rect 22465 415 22485 435
rect 22465 365 22485 385
rect 22465 315 22485 335
rect 22465 265 22485 285
rect 22465 215 22485 235
rect 22465 165 22485 185
rect 22465 115 22485 135
rect 22465 65 22485 85
rect 23365 715 23385 735
rect 23365 665 23385 685
rect 23365 615 23385 635
rect 23365 565 23385 585
rect 23365 515 23385 535
rect 23365 465 23385 485
rect 23365 415 23385 435
rect 23365 365 23385 385
rect 23365 315 23385 335
rect 23365 265 23385 285
rect 23365 215 23385 235
rect 23365 165 23385 185
rect 23365 115 23385 135
rect 23365 65 23385 85
rect 24565 715 24585 735
rect 24565 665 24585 685
rect 24565 615 24585 635
rect 24565 565 24585 585
rect 24565 515 24585 535
rect 24565 465 24585 485
rect 24565 415 24585 435
rect 24565 365 24585 385
rect 24565 315 24585 335
rect 24565 265 24585 285
rect 24565 215 24585 235
rect 24565 165 24585 185
rect 24565 115 24585 135
rect 24565 65 24585 85
rect 25765 715 25785 735
rect 25765 665 25785 685
rect 25765 615 25785 635
rect 25765 565 25785 585
rect 25765 515 25785 535
rect 25765 465 25785 485
rect 25765 415 25785 435
rect 25765 365 25785 385
rect 25765 315 25785 335
rect 25765 265 25785 285
rect 25765 215 25785 235
rect 25765 165 25785 185
rect 25765 115 25785 135
rect 25765 65 25785 85
rect 26665 715 26685 735
rect 26665 665 26685 685
rect 26665 615 26685 635
rect 26665 565 26685 585
rect 26665 515 26685 535
rect 26665 465 26685 485
rect 26665 415 26685 435
rect 26665 365 26685 385
rect 26665 315 26685 335
rect 26665 265 26685 285
rect 26665 215 26685 235
rect 26665 165 26685 185
rect 26665 115 26685 135
rect 26665 65 26685 85
rect 27565 715 27585 735
rect 27565 665 27585 685
rect 27565 615 27585 635
rect 27565 565 27585 585
rect 27565 515 27585 535
rect 27565 465 27585 485
rect 27565 415 27585 435
rect 27565 365 27585 385
rect 27565 315 27585 335
rect 27565 265 27585 285
rect 27565 215 27585 235
rect 27565 165 27585 185
rect 27565 115 27585 135
rect 27565 65 27585 85
rect 28765 715 28785 735
rect 28765 665 28785 685
rect 28765 615 28785 635
rect 28765 565 28785 585
rect 28765 515 28785 535
rect 28765 465 28785 485
rect 28765 415 28785 435
rect 28765 365 28785 385
rect 28765 315 28785 335
rect 28765 265 28785 285
rect 28765 215 28785 235
rect 28765 165 28785 185
rect 28765 115 28785 135
rect 28765 65 28785 85
rect -635 -35 -615 -15
rect -35 -35 -15 -15
rect 8365 -35 8385 -15
rect 10765 -35 10785 -15
rect 15565 -35 15585 -15
rect 17965 -35 17985 -15
rect 20365 -35 20385 -15
rect 24565 -35 24585 -15
rect 28765 -35 28785 -15
rect -635 -135 -615 -115
rect -635 -185 -615 -165
rect -635 -235 -615 -215
rect -635 -285 -615 -265
rect -635 -335 -615 -315
rect -635 -385 -615 -365
rect -635 -435 -615 -415
rect -635 -485 -615 -465
rect -635 -535 -615 -515
rect -635 -585 -615 -565
rect -635 -635 -615 -615
rect -635 -685 -615 -665
rect -635 -735 -615 -715
rect -635 -785 -615 -765
rect -485 -135 -465 -115
rect -485 -185 -465 -165
rect -485 -235 -465 -215
rect -485 -285 -465 -265
rect -485 -335 -465 -315
rect -485 -385 -465 -365
rect -485 -435 -465 -415
rect -485 -485 -465 -465
rect -485 -535 -465 -515
rect -485 -585 -465 -565
rect -485 -635 -465 -615
rect -485 -685 -465 -665
rect -485 -735 -465 -715
rect -485 -785 -465 -765
rect -335 -135 -315 -115
rect -335 -185 -315 -165
rect -335 -235 -315 -215
rect -335 -285 -315 -265
rect -335 -335 -315 -315
rect -335 -385 -315 -365
rect -335 -435 -315 -415
rect -335 -485 -315 -465
rect -335 -535 -315 -515
rect -335 -585 -315 -565
rect -335 -635 -315 -615
rect -335 -685 -315 -665
rect -335 -735 -315 -715
rect -335 -785 -315 -765
rect -185 -135 -165 -115
rect -185 -185 -165 -165
rect -185 -235 -165 -215
rect -185 -285 -165 -265
rect -185 -335 -165 -315
rect -185 -385 -165 -365
rect -185 -435 -165 -415
rect -185 -485 -165 -465
rect -185 -535 -165 -515
rect -185 -585 -165 -565
rect -185 -635 -165 -615
rect -185 -685 -165 -665
rect -185 -735 -165 -715
rect -185 -785 -165 -765
rect -35 -135 -15 -115
rect -35 -185 -15 -165
rect -35 -235 -15 -215
rect -35 -285 -15 -265
rect -35 -335 -15 -315
rect -35 -385 -15 -365
rect -35 -435 -15 -415
rect -35 -485 -15 -465
rect -35 -535 -15 -515
rect -35 -585 -15 -565
rect -35 -635 -15 -615
rect -35 -685 -15 -665
rect -35 -735 -15 -715
rect -35 -785 -15 -765
rect 1165 -135 1185 -115
rect 1165 -185 1185 -165
rect 1165 -235 1185 -215
rect 1165 -285 1185 -265
rect 1165 -335 1185 -315
rect 1165 -385 1185 -365
rect 1165 -435 1185 -415
rect 1165 -485 1185 -465
rect 1165 -535 1185 -515
rect 1165 -585 1185 -565
rect 1165 -635 1185 -615
rect 1165 -685 1185 -665
rect 1165 -735 1185 -715
rect 1165 -785 1185 -765
rect 1465 -235 1485 -215
rect 1465 -285 1485 -265
rect 1465 -335 1485 -315
rect 1465 -385 1485 -365
rect 1465 -435 1485 -415
rect 1465 -485 1485 -465
rect 1465 -535 1485 -515
rect 1465 -585 1485 -565
rect 1465 -635 1485 -615
rect 1465 -685 1485 -665
rect 1465 -735 1485 -715
rect 1465 -785 1485 -765
rect 1765 -135 1785 -115
rect 1765 -185 1785 -165
rect 1765 -235 1785 -215
rect 1765 -285 1785 -265
rect 1765 -335 1785 -315
rect 1765 -385 1785 -365
rect 1765 -435 1785 -415
rect 1765 -485 1785 -465
rect 1765 -535 1785 -515
rect 1765 -585 1785 -565
rect 1765 -635 1785 -615
rect 1765 -685 1785 -665
rect 2065 -235 2085 -215
rect 2065 -285 2085 -265
rect 2065 -335 2085 -315
rect 2065 -385 2085 -365
rect 2065 -435 2085 -415
rect 2065 -485 2085 -465
rect 2065 -535 2085 -515
rect 2065 -585 2085 -565
rect 2065 -635 2085 -615
rect 2065 -685 2085 -665
rect 2065 -735 2085 -715
rect 2065 -785 2085 -765
rect 2365 -135 2385 -115
rect 2365 -185 2385 -165
rect 2365 -235 2385 -215
rect 2365 -285 2385 -265
rect 2365 -335 2385 -315
rect 2365 -385 2385 -365
rect 2365 -435 2385 -415
rect 2365 -485 2385 -465
rect 2365 -535 2385 -515
rect 2365 -585 2385 -565
rect 2365 -635 2385 -615
rect 2365 -685 2385 -665
rect 2665 -235 2685 -215
rect 2665 -285 2685 -265
rect 2665 -335 2685 -315
rect 2665 -385 2685 -365
rect 2665 -435 2685 -415
rect 2665 -485 2685 -465
rect 2665 -535 2685 -515
rect 2665 -585 2685 -565
rect 2665 -635 2685 -615
rect 2665 -685 2685 -665
rect 2665 -735 2685 -715
rect 2665 -785 2685 -765
rect 2965 -135 2985 -115
rect 2965 -185 2985 -165
rect 2965 -235 2985 -215
rect 2965 -285 2985 -265
rect 2965 -335 2985 -315
rect 2965 -385 2985 -365
rect 2965 -435 2985 -415
rect 2965 -485 2985 -465
rect 2965 -535 2985 -515
rect 2965 -585 2985 -565
rect 2965 -635 2985 -615
rect 2965 -685 2985 -665
rect 3265 -235 3285 -215
rect 3265 -285 3285 -265
rect 3265 -335 3285 -315
rect 3265 -385 3285 -365
rect 3265 -435 3285 -415
rect 3265 -485 3285 -465
rect 3265 -535 3285 -515
rect 3265 -585 3285 -565
rect 3265 -635 3285 -615
rect 3265 -685 3285 -665
rect 3265 -735 3285 -715
rect 3265 -785 3285 -765
rect 3565 -135 3585 -115
rect 3565 -185 3585 -165
rect 3565 -235 3585 -215
rect 3565 -285 3585 -265
rect 3565 -335 3585 -315
rect 3565 -385 3585 -365
rect 3565 -435 3585 -415
rect 3565 -485 3585 -465
rect 3565 -535 3585 -515
rect 3565 -585 3585 -565
rect 3565 -635 3585 -615
rect 3565 -685 3585 -665
rect 3565 -735 3585 -715
rect 3565 -785 3585 -765
rect 3715 -235 3735 -215
rect 3715 -285 3735 -265
rect 3715 -335 3735 -315
rect 3715 -385 3735 -365
rect 3715 -435 3735 -415
rect 3715 -485 3735 -465
rect 3715 -535 3735 -515
rect 3715 -585 3735 -565
rect 3715 -635 3735 -615
rect 3715 -685 3735 -665
rect 3715 -735 3735 -715
rect 3715 -785 3735 -765
rect 3865 -135 3885 -115
rect 3865 -185 3885 -165
rect 3865 -235 3885 -215
rect 3865 -285 3885 -265
rect 3865 -335 3885 -315
rect 3865 -385 3885 -365
rect 3865 -435 3885 -415
rect 3865 -485 3885 -465
rect 3865 -535 3885 -515
rect 3865 -585 3885 -565
rect 3865 -635 3885 -615
rect 3865 -685 3885 -665
rect 4015 -235 4035 -215
rect 4015 -285 4035 -265
rect 4015 -335 4035 -315
rect 4015 -385 4035 -365
rect 4015 -435 4035 -415
rect 4015 -485 4035 -465
rect 4015 -535 4035 -515
rect 4015 -585 4035 -565
rect 4015 -635 4035 -615
rect 4015 -685 4035 -665
rect 4015 -735 4035 -715
rect 4015 -785 4035 -765
rect 4165 -135 4185 -115
rect 4165 -185 4185 -165
rect 4165 -235 4185 -215
rect 4165 -285 4185 -265
rect 4165 -335 4185 -315
rect 4165 -385 4185 -365
rect 4165 -435 4185 -415
rect 4165 -485 4185 -465
rect 4165 -535 4185 -515
rect 4165 -585 4185 -565
rect 4165 -635 4185 -615
rect 4165 -685 4185 -665
rect 4165 -735 4185 -715
rect 4165 -785 4185 -765
rect 4315 -235 4335 -215
rect 4315 -285 4335 -265
rect 4315 -335 4335 -315
rect 4315 -385 4335 -365
rect 4315 -435 4335 -415
rect 4315 -485 4335 -465
rect 4315 -535 4335 -515
rect 4315 -585 4335 -565
rect 4315 -635 4335 -615
rect 4315 -685 4335 -665
rect 4315 -735 4335 -715
rect 4315 -785 4335 -765
rect 4465 -135 4485 -115
rect 4465 -185 4485 -165
rect 4465 -235 4485 -215
rect 4465 -285 4485 -265
rect 4465 -335 4485 -315
rect 4465 -385 4485 -365
rect 4465 -435 4485 -415
rect 4465 -485 4485 -465
rect 4465 -535 4485 -515
rect 4465 -585 4485 -565
rect 4465 -635 4485 -615
rect 4465 -685 4485 -665
rect 4615 -235 4635 -215
rect 4615 -285 4635 -265
rect 4615 -335 4635 -315
rect 4615 -385 4635 -365
rect 4615 -435 4635 -415
rect 4615 -485 4635 -465
rect 4615 -535 4635 -515
rect 4615 -585 4635 -565
rect 4615 -635 4635 -615
rect 4615 -685 4635 -665
rect 4615 -735 4635 -715
rect 4615 -785 4635 -765
rect 4765 -135 4785 -115
rect 4765 -185 4785 -165
rect 4765 -235 4785 -215
rect 4765 -285 4785 -265
rect 4765 -335 4785 -315
rect 4765 -385 4785 -365
rect 4765 -435 4785 -415
rect 4765 -485 4785 -465
rect 4765 -535 4785 -515
rect 4765 -585 4785 -565
rect 4765 -635 4785 -615
rect 4765 -685 4785 -665
rect 4765 -735 4785 -715
rect 4765 -785 4785 -765
rect 5065 -235 5085 -215
rect 5065 -285 5085 -265
rect 5065 -335 5085 -315
rect 5065 -385 5085 -365
rect 5065 -435 5085 -415
rect 5065 -485 5085 -465
rect 5065 -535 5085 -515
rect 5065 -585 5085 -565
rect 5065 -635 5085 -615
rect 5065 -685 5085 -665
rect 5065 -735 5085 -715
rect 5065 -785 5085 -765
rect 5365 -135 5385 -115
rect 5365 -185 5385 -165
rect 5365 -235 5385 -215
rect 5365 -285 5385 -265
rect 5365 -335 5385 -315
rect 5365 -385 5385 -365
rect 5365 -435 5385 -415
rect 5365 -485 5385 -465
rect 5365 -535 5385 -515
rect 5365 -585 5385 -565
rect 5365 -635 5385 -615
rect 5365 -685 5385 -665
rect 5665 -235 5685 -215
rect 5665 -285 5685 -265
rect 5665 -335 5685 -315
rect 5665 -385 5685 -365
rect 5665 -435 5685 -415
rect 5665 -485 5685 -465
rect 5665 -535 5685 -515
rect 5665 -585 5685 -565
rect 5665 -635 5685 -615
rect 5665 -685 5685 -665
rect 5665 -735 5685 -715
rect 5665 -785 5685 -765
rect 5965 -135 5985 -115
rect 5965 -185 5985 -165
rect 5965 -235 5985 -215
rect 5965 -285 5985 -265
rect 5965 -335 5985 -315
rect 5965 -385 5985 -365
rect 5965 -435 5985 -415
rect 5965 -485 5985 -465
rect 5965 -535 5985 -515
rect 5965 -585 5985 -565
rect 5965 -635 5985 -615
rect 5965 -685 5985 -665
rect 6265 -235 6285 -215
rect 6265 -285 6285 -265
rect 6265 -335 6285 -315
rect 6265 -385 6285 -365
rect 6265 -435 6285 -415
rect 6265 -485 6285 -465
rect 6265 -535 6285 -515
rect 6265 -585 6285 -565
rect 6265 -635 6285 -615
rect 6265 -685 6285 -665
rect 6265 -735 6285 -715
rect 6265 -785 6285 -765
rect 6565 -135 6585 -115
rect 6565 -185 6585 -165
rect 6565 -235 6585 -215
rect 6565 -285 6585 -265
rect 6565 -335 6585 -315
rect 6565 -385 6585 -365
rect 6565 -435 6585 -415
rect 6565 -485 6585 -465
rect 6565 -535 6585 -515
rect 6565 -585 6585 -565
rect 6565 -635 6585 -615
rect 6565 -685 6585 -665
rect 6865 -235 6885 -215
rect 6865 -285 6885 -265
rect 6865 -335 6885 -315
rect 6865 -385 6885 -365
rect 6865 -435 6885 -415
rect 6865 -485 6885 -465
rect 6865 -535 6885 -515
rect 6865 -585 6885 -565
rect 6865 -635 6885 -615
rect 6865 -685 6885 -665
rect 6865 -735 6885 -715
rect 6865 -785 6885 -765
rect 7165 -135 7185 -115
rect 7165 -185 7185 -165
rect 7165 -235 7185 -215
rect 7165 -285 7185 -265
rect 7165 -335 7185 -315
rect 7165 -385 7185 -365
rect 7165 -435 7185 -415
rect 7165 -485 7185 -465
rect 7165 -535 7185 -515
rect 7165 -585 7185 -565
rect 7165 -635 7185 -615
rect 7165 -685 7185 -665
rect 7165 -735 7185 -715
rect 7165 -785 7185 -765
rect 8365 -135 8385 -115
rect 8365 -185 8385 -165
rect 8365 -235 8385 -215
rect 8365 -285 8385 -265
rect 8365 -335 8385 -315
rect 8365 -385 8385 -365
rect 8365 -435 8385 -415
rect 8365 -485 8385 -465
rect 8365 -535 8385 -515
rect 8365 -585 8385 -565
rect 8365 -635 8385 -615
rect 8365 -685 8385 -665
rect 8365 -735 8385 -715
rect 8365 -785 8385 -765
rect 9565 -135 9585 -115
rect 9565 -185 9585 -165
rect 9565 -235 9585 -215
rect 9565 -285 9585 -265
rect 9565 -335 9585 -315
rect 9565 -385 9585 -365
rect 9565 -435 9585 -415
rect 9565 -485 9585 -465
rect 9565 -535 9585 -515
rect 9565 -585 9585 -565
rect 9565 -635 9585 -615
rect 9565 -685 9585 -665
rect 9565 -735 9585 -715
rect 9565 -785 9585 -765
rect 10765 -135 10785 -115
rect 10765 -185 10785 -165
rect 10765 -235 10785 -215
rect 10765 -285 10785 -265
rect 10765 -335 10785 -315
rect 10765 -385 10785 -365
rect 10765 -435 10785 -415
rect 10765 -485 10785 -465
rect 10765 -535 10785 -515
rect 10765 -585 10785 -565
rect 10765 -635 10785 -615
rect 10765 -685 10785 -665
rect 10765 -735 10785 -715
rect 10765 -785 10785 -765
rect 11965 -135 11985 -115
rect 11965 -185 11985 -165
rect 11965 -235 11985 -215
rect 11965 -285 11985 -265
rect 11965 -335 11985 -315
rect 11965 -385 11985 -365
rect 11965 -435 11985 -415
rect 11965 -485 11985 -465
rect 11965 -535 11985 -515
rect 11965 -585 11985 -565
rect 11965 -635 11985 -615
rect 11965 -685 11985 -665
rect 11965 -735 11985 -715
rect 11965 -785 11985 -765
rect 12265 -235 12285 -215
rect 12265 -285 12285 -265
rect 12265 -335 12285 -315
rect 12265 -385 12285 -365
rect 12265 -435 12285 -415
rect 12265 -485 12285 -465
rect 12265 -535 12285 -515
rect 12265 -585 12285 -565
rect 12265 -635 12285 -615
rect 12265 -685 12285 -665
rect 12265 -735 12285 -715
rect 12265 -785 12285 -765
rect 12565 -135 12585 -115
rect 12565 -185 12585 -165
rect 12565 -235 12585 -215
rect 12565 -285 12585 -265
rect 12565 -335 12585 -315
rect 12565 -385 12585 -365
rect 12565 -435 12585 -415
rect 12565 -485 12585 -465
rect 12565 -535 12585 -515
rect 12565 -585 12585 -565
rect 12565 -635 12585 -615
rect 12565 -685 12585 -665
rect 12865 -235 12885 -215
rect 12865 -285 12885 -265
rect 12865 -335 12885 -315
rect 12865 -385 12885 -365
rect 12865 -435 12885 -415
rect 12865 -485 12885 -465
rect 12865 -535 12885 -515
rect 12865 -585 12885 -565
rect 12865 -635 12885 -615
rect 12865 -685 12885 -665
rect 12865 -735 12885 -715
rect 12865 -785 12885 -765
rect 13165 -135 13185 -115
rect 13165 -185 13185 -165
rect 13165 -235 13185 -215
rect 13165 -285 13185 -265
rect 13165 -335 13185 -315
rect 13165 -385 13185 -365
rect 13165 -435 13185 -415
rect 13165 -485 13185 -465
rect 13165 -535 13185 -515
rect 13165 -585 13185 -565
rect 13165 -635 13185 -615
rect 13165 -685 13185 -665
rect 13465 -235 13485 -215
rect 13465 -285 13485 -265
rect 13465 -335 13485 -315
rect 13465 -385 13485 -365
rect 13465 -435 13485 -415
rect 13465 -485 13485 -465
rect 13465 -535 13485 -515
rect 13465 -585 13485 -565
rect 13465 -635 13485 -615
rect 13465 -685 13485 -665
rect 13465 -735 13485 -715
rect 13465 -785 13485 -765
rect 13765 -135 13785 -115
rect 13765 -185 13785 -165
rect 13765 -235 13785 -215
rect 13765 -285 13785 -265
rect 13765 -335 13785 -315
rect 13765 -385 13785 -365
rect 13765 -435 13785 -415
rect 13765 -485 13785 -465
rect 13765 -535 13785 -515
rect 13765 -585 13785 -565
rect 13765 -635 13785 -615
rect 13765 -685 13785 -665
rect 14065 -235 14085 -215
rect 14065 -285 14085 -265
rect 14065 -335 14085 -315
rect 14065 -385 14085 -365
rect 14065 -435 14085 -415
rect 14065 -485 14085 -465
rect 14065 -535 14085 -515
rect 14065 -585 14085 -565
rect 14065 -635 14085 -615
rect 14065 -685 14085 -665
rect 14065 -735 14085 -715
rect 14065 -785 14085 -765
rect 14365 -135 14385 -115
rect 14365 -185 14385 -165
rect 14365 -235 14385 -215
rect 14365 -285 14385 -265
rect 14365 -335 14385 -315
rect 14365 -385 14385 -365
rect 14365 -435 14385 -415
rect 14365 -485 14385 -465
rect 14365 -535 14385 -515
rect 14365 -585 14385 -565
rect 14365 -635 14385 -615
rect 14365 -685 14385 -665
rect 14365 -735 14385 -715
rect 14365 -785 14385 -765
rect 15565 -135 15585 -115
rect 15565 -185 15585 -165
rect 15565 -235 15585 -215
rect 15565 -285 15585 -265
rect 15565 -335 15585 -315
rect 15565 -385 15585 -365
rect 15565 -435 15585 -415
rect 15565 -485 15585 -465
rect 15565 -535 15585 -515
rect 15565 -585 15585 -565
rect 15565 -635 15585 -615
rect 15565 -685 15585 -665
rect 15565 -735 15585 -715
rect 15565 -785 15585 -765
rect 16765 -135 16785 -115
rect 16765 -185 16785 -165
rect 16765 -235 16785 -215
rect 16765 -285 16785 -265
rect 16765 -335 16785 -315
rect 16765 -385 16785 -365
rect 16765 -435 16785 -415
rect 16765 -485 16785 -465
rect 16765 -535 16785 -515
rect 16765 -585 16785 -565
rect 16765 -635 16785 -615
rect 16765 -685 16785 -665
rect 16765 -735 16785 -715
rect 16765 -785 16785 -765
rect 17965 -135 17985 -115
rect 17965 -185 17985 -165
rect 17965 -235 17985 -215
rect 17965 -285 17985 -265
rect 17965 -335 17985 -315
rect 17965 -385 17985 -365
rect 17965 -435 17985 -415
rect 17965 -485 17985 -465
rect 17965 -535 17985 -515
rect 17965 -585 17985 -565
rect 17965 -635 17985 -615
rect 17965 -685 17985 -665
rect 17965 -735 17985 -715
rect 17965 -785 17985 -765
rect 19165 -135 19185 -115
rect 19165 -185 19185 -165
rect 19165 -235 19185 -215
rect 19165 -285 19185 -265
rect 19165 -335 19185 -315
rect 19165 -385 19185 -365
rect 19165 -435 19185 -415
rect 19165 -485 19185 -465
rect 19165 -535 19185 -515
rect 19165 -585 19185 -565
rect 19165 -635 19185 -615
rect 19165 -685 19185 -665
rect 19165 -735 19185 -715
rect 19165 -785 19185 -765
rect 20365 -135 20385 -115
rect 20365 -185 20385 -165
rect 20365 -235 20385 -215
rect 20365 -285 20385 -265
rect 20365 -335 20385 -315
rect 20365 -385 20385 -365
rect 20365 -435 20385 -415
rect 20365 -485 20385 -465
rect 20365 -535 20385 -515
rect 20365 -585 20385 -565
rect 20365 -635 20385 -615
rect 20365 -685 20385 -665
rect 20365 -735 20385 -715
rect 20365 -785 20385 -765
rect 21565 -135 21585 -115
rect 21565 -185 21585 -165
rect 21565 -235 21585 -215
rect 21565 -285 21585 -265
rect 21565 -335 21585 -315
rect 21565 -385 21585 -365
rect 21565 -435 21585 -415
rect 21565 -485 21585 -465
rect 21565 -535 21585 -515
rect 21565 -585 21585 -565
rect 21565 -635 21585 -615
rect 21565 -685 21585 -665
rect 21565 -735 21585 -715
rect 21565 -785 21585 -765
rect 22465 -135 22485 -115
rect 22465 -185 22485 -165
rect 22465 -235 22485 -215
rect 22465 -285 22485 -265
rect 22465 -335 22485 -315
rect 22465 -385 22485 -365
rect 22465 -435 22485 -415
rect 22465 -485 22485 -465
rect 22465 -535 22485 -515
rect 22465 -585 22485 -565
rect 22465 -635 22485 -615
rect 22465 -685 22485 -665
rect 22465 -735 22485 -715
rect 22465 -785 22485 -765
rect 23365 -135 23385 -115
rect 23365 -185 23385 -165
rect 23365 -235 23385 -215
rect 23365 -285 23385 -265
rect 23365 -335 23385 -315
rect 23365 -385 23385 -365
rect 23365 -435 23385 -415
rect 23365 -485 23385 -465
rect 23365 -535 23385 -515
rect 23365 -585 23385 -565
rect 23365 -635 23385 -615
rect 23365 -685 23385 -665
rect 23365 -735 23385 -715
rect 23365 -785 23385 -765
rect 24565 -135 24585 -115
rect 24565 -185 24585 -165
rect 24565 -235 24585 -215
rect 24565 -285 24585 -265
rect 24565 -335 24585 -315
rect 24565 -385 24585 -365
rect 24565 -435 24585 -415
rect 24565 -485 24585 -465
rect 24565 -535 24585 -515
rect 24565 -585 24585 -565
rect 24565 -635 24585 -615
rect 24565 -685 24585 -665
rect 24565 -735 24585 -715
rect 24565 -785 24585 -765
rect 25765 -135 25785 -115
rect 25765 -185 25785 -165
rect 25765 -235 25785 -215
rect 25765 -285 25785 -265
rect 25765 -335 25785 -315
rect 25765 -385 25785 -365
rect 25765 -435 25785 -415
rect 25765 -485 25785 -465
rect 25765 -535 25785 -515
rect 25765 -585 25785 -565
rect 25765 -635 25785 -615
rect 25765 -685 25785 -665
rect 25765 -735 25785 -715
rect 25765 -785 25785 -765
rect 26665 -135 26685 -115
rect 26665 -185 26685 -165
rect 26665 -235 26685 -215
rect 26665 -285 26685 -265
rect 26665 -335 26685 -315
rect 26665 -385 26685 -365
rect 26665 -435 26685 -415
rect 26665 -485 26685 -465
rect 26665 -535 26685 -515
rect 26665 -585 26685 -565
rect 26665 -635 26685 -615
rect 26665 -685 26685 -665
rect 26665 -735 26685 -715
rect 26665 -785 26685 -765
rect 27565 -135 27585 -115
rect 27565 -185 27585 -165
rect 27565 -235 27585 -215
rect 27565 -285 27585 -265
rect 27565 -335 27585 -315
rect 27565 -385 27585 -365
rect 27565 -435 27585 -415
rect 27565 -485 27585 -465
rect 27565 -535 27585 -515
rect 27565 -585 27585 -565
rect 27565 -635 27585 -615
rect 27565 -685 27585 -665
rect 27565 -735 27585 -715
rect 27565 -785 27585 -765
rect 28765 -135 28785 -115
rect 28765 -185 28785 -165
rect 28765 -235 28785 -215
rect 28765 -285 28785 -265
rect 28765 -335 28785 -315
rect 28765 -385 28785 -365
rect 28765 -435 28785 -415
rect 28765 -485 28785 -465
rect 28765 -535 28785 -515
rect 28765 -585 28785 -565
rect 28765 -635 28785 -615
rect 28765 -685 28785 -665
rect 28765 -735 28785 -715
rect 28765 -785 28785 -765
rect -485 -885 -465 -865
rect -185 -885 -165 -865
rect 115 -885 135 -865
rect 415 -885 435 -865
rect 715 -885 735 -865
rect 1015 -885 1035 -865
rect 1315 -885 1335 -865
rect 1615 -885 1635 -865
rect 1915 -885 1935 -865
rect 2215 -885 2235 -865
rect 2515 -885 2535 -865
rect 2815 -885 2835 -865
rect 3115 -885 3135 -865
rect 3415 -885 3435 -865
rect 3715 -885 3735 -865
rect 4015 -885 4035 -865
rect 4315 -885 4335 -865
rect 4615 -885 4635 -865
rect 4915 -885 4935 -865
rect 5215 -885 5235 -865
rect 5515 -885 5535 -865
rect 5815 -885 5835 -865
rect 6115 -885 6135 -865
rect 6415 -885 6435 -865
rect 6715 -885 6735 -865
rect 7015 -885 7035 -865
rect 7315 -885 7335 -865
rect 7615 -885 7635 -865
rect 7915 -885 7935 -865
rect 8215 -885 8235 -865
rect 8515 -885 8535 -865
rect 8815 -885 8835 -865
rect 9115 -885 9135 -865
rect 9415 -885 9435 -865
rect 9715 -885 9735 -865
rect 10015 -885 10035 -865
rect 10315 -885 10335 -865
rect 10615 -885 10635 -865
rect 10915 -885 10935 -865
rect 11215 -885 11235 -865
rect 11515 -885 11535 -865
rect 11815 -885 11835 -865
rect 12115 -885 12135 -865
rect 12415 -885 12435 -865
rect 12715 -885 12735 -865
rect 13015 -885 13035 -865
rect 13315 -885 13335 -865
rect 13615 -885 13635 -865
rect 13915 -885 13935 -865
rect 14215 -885 14235 -865
rect 14515 -885 14535 -865
rect 14815 -885 14835 -865
rect 15115 -885 15135 -865
rect 15415 -885 15435 -865
rect 15715 -885 15735 -865
rect 16015 -885 16035 -865
rect 16315 -885 16335 -865
rect 16615 -885 16635 -865
rect 16915 -885 16935 -865
rect 17215 -885 17235 -865
rect 17515 -885 17535 -865
rect 17815 -885 17835 -865
rect 18115 -885 18135 -865
rect 18415 -885 18435 -865
rect 18715 -885 18735 -865
rect 19015 -885 19035 -865
rect 19315 -885 19335 -865
rect 19615 -885 19635 -865
rect 19915 -885 19935 -865
rect 20215 -885 20235 -865
rect 20515 -885 20535 -865
rect 20815 -885 20835 -865
rect 21115 -885 21135 -865
rect 21415 -885 21435 -865
rect 21715 -885 21735 -865
rect 22015 -885 22035 -865
rect 22315 -885 22335 -865
rect 22615 -885 22635 -865
rect 22915 -885 22935 -865
rect 23215 -885 23235 -865
rect 23515 -885 23535 -865
rect 23815 -885 23835 -865
rect 24115 -885 24135 -865
rect 24415 -885 24435 -865
rect 24715 -885 24735 -865
rect 25015 -885 25035 -865
rect 25315 -885 25335 -865
rect 25615 -885 25635 -865
rect 25915 -885 25935 -865
rect 26215 -885 26235 -865
rect 26515 -885 26535 -865
rect 26815 -885 26835 -865
rect 27115 -885 27135 -865
rect 27415 -885 27435 -865
rect 27715 -885 27735 -865
rect 28015 -885 28035 -865
rect 28315 -885 28335 -865
rect 28615 -885 28635 -865
rect -635 -985 -615 -965
rect -635 -1035 -615 -1015
rect -635 -1085 -615 -1065
rect -635 -1135 -615 -1115
rect -635 -1185 -615 -1165
rect -635 -1235 -615 -1215
rect -635 -1285 -615 -1265
rect -635 -1335 -615 -1315
rect -635 -1385 -615 -1365
rect -635 -1435 -615 -1415
rect -635 -1485 -615 -1465
rect -635 -1535 -615 -1515
rect -635 -1585 -615 -1565
rect -635 -1635 -615 -1615
rect -485 -985 -465 -965
rect -485 -1035 -465 -1015
rect -485 -1085 -465 -1065
rect -485 -1135 -465 -1115
rect -485 -1185 -465 -1165
rect -485 -1235 -465 -1215
rect -485 -1285 -465 -1265
rect -485 -1335 -465 -1315
rect -485 -1385 -465 -1365
rect -485 -1435 -465 -1415
rect -485 -1485 -465 -1465
rect -485 -1535 -465 -1515
rect -485 -1585 -465 -1565
rect -485 -1635 -465 -1615
rect -335 -985 -315 -965
rect -335 -1035 -315 -1015
rect -335 -1085 -315 -1065
rect -335 -1135 -315 -1115
rect -335 -1185 -315 -1165
rect -335 -1235 -315 -1215
rect -335 -1285 -315 -1265
rect -335 -1335 -315 -1315
rect -335 -1385 -315 -1365
rect -335 -1435 -315 -1415
rect -335 -1485 -315 -1465
rect -335 -1535 -315 -1515
rect -335 -1585 -315 -1565
rect -335 -1635 -315 -1615
rect -185 -985 -165 -965
rect -185 -1035 -165 -1015
rect -185 -1085 -165 -1065
rect -185 -1135 -165 -1115
rect -185 -1185 -165 -1165
rect -185 -1235 -165 -1215
rect -185 -1285 -165 -1265
rect -185 -1335 -165 -1315
rect -185 -1385 -165 -1365
rect -185 -1435 -165 -1415
rect -185 -1485 -165 -1465
rect -185 -1535 -165 -1515
rect -185 -1585 -165 -1565
rect -185 -1635 -165 -1615
rect -35 -985 -15 -965
rect -35 -1035 -15 -1015
rect -35 -1085 -15 -1065
rect -35 -1135 -15 -1115
rect -35 -1185 -15 -1165
rect -35 -1235 -15 -1215
rect -35 -1285 -15 -1265
rect -35 -1335 -15 -1315
rect -35 -1385 -15 -1365
rect -35 -1435 -15 -1415
rect -35 -1485 -15 -1465
rect -35 -1535 -15 -1515
rect -35 -1585 -15 -1565
rect -35 -1635 -15 -1615
rect 1165 -985 1185 -965
rect 1165 -1035 1185 -1015
rect 1165 -1085 1185 -1065
rect 1165 -1135 1185 -1115
rect 1165 -1185 1185 -1165
rect 1165 -1235 1185 -1215
rect 1165 -1285 1185 -1265
rect 1165 -1335 1185 -1315
rect 1165 -1385 1185 -1365
rect 1165 -1435 1185 -1415
rect 1165 -1485 1185 -1465
rect 1165 -1535 1185 -1515
rect 1165 -1585 1185 -1565
rect 1165 -1635 1185 -1615
rect 1465 -985 1485 -965
rect 1465 -1035 1485 -1015
rect 1465 -1085 1485 -1065
rect 1465 -1135 1485 -1115
rect 1465 -1185 1485 -1165
rect 1465 -1235 1485 -1215
rect 1465 -1285 1485 -1265
rect 1465 -1335 1485 -1315
rect 1465 -1385 1485 -1365
rect 1465 -1435 1485 -1415
rect 1465 -1485 1485 -1465
rect 1465 -1535 1485 -1515
rect 1765 -1085 1785 -1065
rect 1765 -1135 1785 -1115
rect 1765 -1185 1785 -1165
rect 1765 -1235 1785 -1215
rect 1765 -1285 1785 -1265
rect 1765 -1335 1785 -1315
rect 1765 -1385 1785 -1365
rect 1765 -1435 1785 -1415
rect 1765 -1485 1785 -1465
rect 1765 -1535 1785 -1515
rect 1765 -1585 1785 -1565
rect 1765 -1635 1785 -1615
rect 2065 -985 2085 -965
rect 2065 -1035 2085 -1015
rect 2065 -1085 2085 -1065
rect 2065 -1135 2085 -1115
rect 2065 -1185 2085 -1165
rect 2065 -1235 2085 -1215
rect 2065 -1285 2085 -1265
rect 2065 -1335 2085 -1315
rect 2065 -1385 2085 -1365
rect 2065 -1435 2085 -1415
rect 2065 -1485 2085 -1465
rect 2065 -1535 2085 -1515
rect 2365 -1085 2385 -1065
rect 2365 -1135 2385 -1115
rect 2365 -1185 2385 -1165
rect 2365 -1235 2385 -1215
rect 2365 -1285 2385 -1265
rect 2365 -1335 2385 -1315
rect 2365 -1385 2385 -1365
rect 2365 -1435 2385 -1415
rect 2365 -1485 2385 -1465
rect 2365 -1535 2385 -1515
rect 2365 -1585 2385 -1565
rect 2365 -1635 2385 -1615
rect 2665 -985 2685 -965
rect 2665 -1035 2685 -1015
rect 2665 -1085 2685 -1065
rect 2665 -1135 2685 -1115
rect 2665 -1185 2685 -1165
rect 2665 -1235 2685 -1215
rect 2665 -1285 2685 -1265
rect 2665 -1335 2685 -1315
rect 2665 -1385 2685 -1365
rect 2665 -1435 2685 -1415
rect 2665 -1485 2685 -1465
rect 2665 -1535 2685 -1515
rect 2965 -1085 2985 -1065
rect 2965 -1135 2985 -1115
rect 2965 -1185 2985 -1165
rect 2965 -1235 2985 -1215
rect 2965 -1285 2985 -1265
rect 2965 -1335 2985 -1315
rect 2965 -1385 2985 -1365
rect 2965 -1435 2985 -1415
rect 2965 -1485 2985 -1465
rect 2965 -1535 2985 -1515
rect 2965 -1585 2985 -1565
rect 2965 -1635 2985 -1615
rect 3265 -985 3285 -965
rect 3265 -1035 3285 -1015
rect 3265 -1085 3285 -1065
rect 3265 -1135 3285 -1115
rect 3265 -1185 3285 -1165
rect 3265 -1235 3285 -1215
rect 3265 -1285 3285 -1265
rect 3265 -1335 3285 -1315
rect 3265 -1385 3285 -1365
rect 3265 -1435 3285 -1415
rect 3265 -1485 3285 -1465
rect 3265 -1535 3285 -1515
rect 3565 -985 3585 -965
rect 3565 -1035 3585 -1015
rect 3565 -1085 3585 -1065
rect 3565 -1135 3585 -1115
rect 3565 -1185 3585 -1165
rect 3565 -1235 3585 -1215
rect 3565 -1285 3585 -1265
rect 3565 -1335 3585 -1315
rect 3565 -1385 3585 -1365
rect 3565 -1435 3585 -1415
rect 3565 -1485 3585 -1465
rect 3565 -1535 3585 -1515
rect 3565 -1585 3585 -1565
rect 3565 -1635 3585 -1615
rect 3715 -985 3735 -965
rect 3715 -1035 3735 -1015
rect 3715 -1085 3735 -1065
rect 3715 -1135 3735 -1115
rect 3715 -1185 3735 -1165
rect 3715 -1235 3735 -1215
rect 3715 -1285 3735 -1265
rect 3715 -1335 3735 -1315
rect 3715 -1385 3735 -1365
rect 3715 -1435 3735 -1415
rect 3715 -1485 3735 -1465
rect 3715 -1535 3735 -1515
rect 3865 -1085 3885 -1065
rect 3865 -1135 3885 -1115
rect 3865 -1185 3885 -1165
rect 3865 -1235 3885 -1215
rect 3865 -1285 3885 -1265
rect 3865 -1335 3885 -1315
rect 3865 -1385 3885 -1365
rect 3865 -1435 3885 -1415
rect 3865 -1485 3885 -1465
rect 3865 -1535 3885 -1515
rect 3865 -1585 3885 -1565
rect 3865 -1635 3885 -1615
rect 4015 -985 4035 -965
rect 4015 -1035 4035 -1015
rect 4015 -1085 4035 -1065
rect 4015 -1135 4035 -1115
rect 4015 -1185 4035 -1165
rect 4015 -1235 4035 -1215
rect 4015 -1285 4035 -1265
rect 4015 -1335 4035 -1315
rect 4015 -1385 4035 -1365
rect 4015 -1435 4035 -1415
rect 4015 -1485 4035 -1465
rect 4015 -1535 4035 -1515
rect 4165 -985 4185 -965
rect 4165 -1035 4185 -1015
rect 4165 -1085 4185 -1065
rect 4165 -1135 4185 -1115
rect 4165 -1185 4185 -1165
rect 4165 -1235 4185 -1215
rect 4165 -1285 4185 -1265
rect 4165 -1335 4185 -1315
rect 4165 -1385 4185 -1365
rect 4165 -1435 4185 -1415
rect 4165 -1485 4185 -1465
rect 4165 -1535 4185 -1515
rect 4165 -1585 4185 -1565
rect 4165 -1635 4185 -1615
rect 4315 -985 4335 -965
rect 4315 -1035 4335 -1015
rect 4315 -1085 4335 -1065
rect 4315 -1135 4335 -1115
rect 4315 -1185 4335 -1165
rect 4315 -1235 4335 -1215
rect 4315 -1285 4335 -1265
rect 4315 -1335 4335 -1315
rect 4315 -1385 4335 -1365
rect 4315 -1435 4335 -1415
rect 4315 -1485 4335 -1465
rect 4315 -1535 4335 -1515
rect 4465 -1085 4485 -1065
rect 4465 -1135 4485 -1115
rect 4465 -1185 4485 -1165
rect 4465 -1235 4485 -1215
rect 4465 -1285 4485 -1265
rect 4465 -1335 4485 -1315
rect 4465 -1385 4485 -1365
rect 4465 -1435 4485 -1415
rect 4465 -1485 4485 -1465
rect 4465 -1535 4485 -1515
rect 4465 -1585 4485 -1565
rect 4465 -1635 4485 -1615
rect 4615 -985 4635 -965
rect 4615 -1035 4635 -1015
rect 4615 -1085 4635 -1065
rect 4615 -1135 4635 -1115
rect 4615 -1185 4635 -1165
rect 4615 -1235 4635 -1215
rect 4615 -1285 4635 -1265
rect 4615 -1335 4635 -1315
rect 4615 -1385 4635 -1365
rect 4615 -1435 4635 -1415
rect 4615 -1485 4635 -1465
rect 4615 -1535 4635 -1515
rect 4765 -985 4785 -965
rect 4765 -1035 4785 -1015
rect 4765 -1085 4785 -1065
rect 4765 -1135 4785 -1115
rect 4765 -1185 4785 -1165
rect 4765 -1235 4785 -1215
rect 4765 -1285 4785 -1265
rect 4765 -1335 4785 -1315
rect 4765 -1385 4785 -1365
rect 4765 -1435 4785 -1415
rect 4765 -1485 4785 -1465
rect 4765 -1535 4785 -1515
rect 4765 -1585 4785 -1565
rect 4765 -1635 4785 -1615
rect 5065 -985 5085 -965
rect 5065 -1035 5085 -1015
rect 5065 -1085 5085 -1065
rect 5065 -1135 5085 -1115
rect 5065 -1185 5085 -1165
rect 5065 -1235 5085 -1215
rect 5065 -1285 5085 -1265
rect 5065 -1335 5085 -1315
rect 5065 -1385 5085 -1365
rect 5065 -1435 5085 -1415
rect 5065 -1485 5085 -1465
rect 5065 -1535 5085 -1515
rect 5365 -1085 5385 -1065
rect 5365 -1135 5385 -1115
rect 5365 -1185 5385 -1165
rect 5365 -1235 5385 -1215
rect 5365 -1285 5385 -1265
rect 5365 -1335 5385 -1315
rect 5365 -1385 5385 -1365
rect 5365 -1435 5385 -1415
rect 5365 -1485 5385 -1465
rect 5365 -1535 5385 -1515
rect 5365 -1585 5385 -1565
rect 5365 -1635 5385 -1615
rect 5665 -985 5685 -965
rect 5665 -1035 5685 -1015
rect 5665 -1085 5685 -1065
rect 5665 -1135 5685 -1115
rect 5665 -1185 5685 -1165
rect 5665 -1235 5685 -1215
rect 5665 -1285 5685 -1265
rect 5665 -1335 5685 -1315
rect 5665 -1385 5685 -1365
rect 5665 -1435 5685 -1415
rect 5665 -1485 5685 -1465
rect 5665 -1535 5685 -1515
rect 5965 -1085 5985 -1065
rect 5965 -1135 5985 -1115
rect 5965 -1185 5985 -1165
rect 5965 -1235 5985 -1215
rect 5965 -1285 5985 -1265
rect 5965 -1335 5985 -1315
rect 5965 -1385 5985 -1365
rect 5965 -1435 5985 -1415
rect 5965 -1485 5985 -1465
rect 5965 -1535 5985 -1515
rect 5965 -1585 5985 -1565
rect 5965 -1635 5985 -1615
rect 6265 -985 6285 -965
rect 6265 -1035 6285 -1015
rect 6265 -1085 6285 -1065
rect 6265 -1135 6285 -1115
rect 6265 -1185 6285 -1165
rect 6265 -1235 6285 -1215
rect 6265 -1285 6285 -1265
rect 6265 -1335 6285 -1315
rect 6265 -1385 6285 -1365
rect 6265 -1435 6285 -1415
rect 6265 -1485 6285 -1465
rect 6265 -1535 6285 -1515
rect 6565 -1085 6585 -1065
rect 6565 -1135 6585 -1115
rect 6565 -1185 6585 -1165
rect 6565 -1235 6585 -1215
rect 6565 -1285 6585 -1265
rect 6565 -1335 6585 -1315
rect 6565 -1385 6585 -1365
rect 6565 -1435 6585 -1415
rect 6565 -1485 6585 -1465
rect 6565 -1535 6585 -1515
rect 6565 -1585 6585 -1565
rect 6565 -1635 6585 -1615
rect 6865 -985 6885 -965
rect 6865 -1035 6885 -1015
rect 6865 -1085 6885 -1065
rect 6865 -1135 6885 -1115
rect 6865 -1185 6885 -1165
rect 6865 -1235 6885 -1215
rect 6865 -1285 6885 -1265
rect 6865 -1335 6885 -1315
rect 6865 -1385 6885 -1365
rect 6865 -1435 6885 -1415
rect 6865 -1485 6885 -1465
rect 6865 -1535 6885 -1515
rect 7165 -985 7185 -965
rect 7165 -1035 7185 -1015
rect 7165 -1085 7185 -1065
rect 7165 -1135 7185 -1115
rect 7165 -1185 7185 -1165
rect 7165 -1235 7185 -1215
rect 7165 -1285 7185 -1265
rect 7165 -1335 7185 -1315
rect 7165 -1385 7185 -1365
rect 7165 -1435 7185 -1415
rect 7165 -1485 7185 -1465
rect 7165 -1535 7185 -1515
rect 7165 -1585 7185 -1565
rect 7165 -1635 7185 -1615
rect 8365 -985 8385 -965
rect 8365 -1035 8385 -1015
rect 8365 -1085 8385 -1065
rect 8365 -1135 8385 -1115
rect 8365 -1185 8385 -1165
rect 8365 -1235 8385 -1215
rect 8365 -1285 8385 -1265
rect 8365 -1335 8385 -1315
rect 8365 -1385 8385 -1365
rect 8365 -1435 8385 -1415
rect 8365 -1485 8385 -1465
rect 8365 -1535 8385 -1515
rect 8365 -1585 8385 -1565
rect 8365 -1635 8385 -1615
rect 9565 -985 9585 -965
rect 9565 -1035 9585 -1015
rect 9565 -1085 9585 -1065
rect 9565 -1135 9585 -1115
rect 9565 -1185 9585 -1165
rect 9565 -1235 9585 -1215
rect 9565 -1285 9585 -1265
rect 9565 -1335 9585 -1315
rect 9565 -1385 9585 -1365
rect 9565 -1435 9585 -1415
rect 9565 -1485 9585 -1465
rect 9565 -1535 9585 -1515
rect 9565 -1585 9585 -1565
rect 9565 -1635 9585 -1615
rect 10765 -985 10785 -965
rect 10765 -1035 10785 -1015
rect 10765 -1085 10785 -1065
rect 10765 -1135 10785 -1115
rect 10765 -1185 10785 -1165
rect 10765 -1235 10785 -1215
rect 10765 -1285 10785 -1265
rect 10765 -1335 10785 -1315
rect 10765 -1385 10785 -1365
rect 10765 -1435 10785 -1415
rect 10765 -1485 10785 -1465
rect 10765 -1535 10785 -1515
rect 10765 -1585 10785 -1565
rect 10765 -1635 10785 -1615
rect 11965 -985 11985 -965
rect 11965 -1035 11985 -1015
rect 11965 -1085 11985 -1065
rect 11965 -1135 11985 -1115
rect 11965 -1185 11985 -1165
rect 11965 -1235 11985 -1215
rect 11965 -1285 11985 -1265
rect 11965 -1335 11985 -1315
rect 11965 -1385 11985 -1365
rect 11965 -1435 11985 -1415
rect 11965 -1485 11985 -1465
rect 11965 -1535 11985 -1515
rect 11965 -1585 11985 -1565
rect 11965 -1635 11985 -1615
rect 12265 -985 12285 -965
rect 12265 -1035 12285 -1015
rect 12265 -1085 12285 -1065
rect 12265 -1135 12285 -1115
rect 12265 -1185 12285 -1165
rect 12265 -1235 12285 -1215
rect 12265 -1285 12285 -1265
rect 12265 -1335 12285 -1315
rect 12265 -1385 12285 -1365
rect 12265 -1435 12285 -1415
rect 12265 -1485 12285 -1465
rect 12265 -1535 12285 -1515
rect 12565 -1085 12585 -1065
rect 12565 -1135 12585 -1115
rect 12565 -1185 12585 -1165
rect 12565 -1235 12585 -1215
rect 12565 -1285 12585 -1265
rect 12565 -1335 12585 -1315
rect 12565 -1385 12585 -1365
rect 12565 -1435 12585 -1415
rect 12565 -1485 12585 -1465
rect 12565 -1535 12585 -1515
rect 12565 -1585 12585 -1565
rect 12565 -1635 12585 -1615
rect 12865 -985 12885 -965
rect 12865 -1035 12885 -1015
rect 12865 -1085 12885 -1065
rect 12865 -1135 12885 -1115
rect 12865 -1185 12885 -1165
rect 12865 -1235 12885 -1215
rect 12865 -1285 12885 -1265
rect 12865 -1335 12885 -1315
rect 12865 -1385 12885 -1365
rect 12865 -1435 12885 -1415
rect 12865 -1485 12885 -1465
rect 12865 -1535 12885 -1515
rect 13165 -1085 13185 -1065
rect 13165 -1135 13185 -1115
rect 13165 -1185 13185 -1165
rect 13165 -1235 13185 -1215
rect 13165 -1285 13185 -1265
rect 13165 -1335 13185 -1315
rect 13165 -1385 13185 -1365
rect 13165 -1435 13185 -1415
rect 13165 -1485 13185 -1465
rect 13165 -1535 13185 -1515
rect 13165 -1585 13185 -1565
rect 13165 -1635 13185 -1615
rect 13465 -985 13485 -965
rect 13465 -1035 13485 -1015
rect 13465 -1085 13485 -1065
rect 13465 -1135 13485 -1115
rect 13465 -1185 13485 -1165
rect 13465 -1235 13485 -1215
rect 13465 -1285 13485 -1265
rect 13465 -1335 13485 -1315
rect 13465 -1385 13485 -1365
rect 13465 -1435 13485 -1415
rect 13465 -1485 13485 -1465
rect 13465 -1535 13485 -1515
rect 13765 -1085 13785 -1065
rect 13765 -1135 13785 -1115
rect 13765 -1185 13785 -1165
rect 13765 -1235 13785 -1215
rect 13765 -1285 13785 -1265
rect 13765 -1335 13785 -1315
rect 13765 -1385 13785 -1365
rect 13765 -1435 13785 -1415
rect 13765 -1485 13785 -1465
rect 13765 -1535 13785 -1515
rect 13765 -1585 13785 -1565
rect 13765 -1635 13785 -1615
rect 14065 -985 14085 -965
rect 14065 -1035 14085 -1015
rect 14065 -1085 14085 -1065
rect 14065 -1135 14085 -1115
rect 14065 -1185 14085 -1165
rect 14065 -1235 14085 -1215
rect 14065 -1285 14085 -1265
rect 14065 -1335 14085 -1315
rect 14065 -1385 14085 -1365
rect 14065 -1435 14085 -1415
rect 14065 -1485 14085 -1465
rect 14065 -1535 14085 -1515
rect 14365 -985 14385 -965
rect 14365 -1035 14385 -1015
rect 14365 -1085 14385 -1065
rect 14365 -1135 14385 -1115
rect 14365 -1185 14385 -1165
rect 14365 -1235 14385 -1215
rect 14365 -1285 14385 -1265
rect 14365 -1335 14385 -1315
rect 14365 -1385 14385 -1365
rect 14365 -1435 14385 -1415
rect 14365 -1485 14385 -1465
rect 14365 -1535 14385 -1515
rect 14365 -1585 14385 -1565
rect 14365 -1635 14385 -1615
rect 15565 -985 15585 -965
rect 15565 -1035 15585 -1015
rect 15565 -1085 15585 -1065
rect 15565 -1135 15585 -1115
rect 15565 -1185 15585 -1165
rect 15565 -1235 15585 -1215
rect 15565 -1285 15585 -1265
rect 15565 -1335 15585 -1315
rect 15565 -1385 15585 -1365
rect 15565 -1435 15585 -1415
rect 15565 -1485 15585 -1465
rect 15565 -1535 15585 -1515
rect 15565 -1585 15585 -1565
rect 15565 -1635 15585 -1615
rect 16765 -985 16785 -965
rect 16765 -1035 16785 -1015
rect 16765 -1085 16785 -1065
rect 16765 -1135 16785 -1115
rect 16765 -1185 16785 -1165
rect 16765 -1235 16785 -1215
rect 16765 -1285 16785 -1265
rect 16765 -1335 16785 -1315
rect 16765 -1385 16785 -1365
rect 16765 -1435 16785 -1415
rect 16765 -1485 16785 -1465
rect 16765 -1535 16785 -1515
rect 16765 -1585 16785 -1565
rect 16765 -1635 16785 -1615
rect 17965 -985 17985 -965
rect 17965 -1035 17985 -1015
rect 17965 -1085 17985 -1065
rect 17965 -1135 17985 -1115
rect 17965 -1185 17985 -1165
rect 17965 -1235 17985 -1215
rect 17965 -1285 17985 -1265
rect 17965 -1335 17985 -1315
rect 17965 -1385 17985 -1365
rect 17965 -1435 17985 -1415
rect 17965 -1485 17985 -1465
rect 17965 -1535 17985 -1515
rect 17965 -1585 17985 -1565
rect 17965 -1635 17985 -1615
rect 19165 -985 19185 -965
rect 19165 -1035 19185 -1015
rect 19165 -1085 19185 -1065
rect 19165 -1135 19185 -1115
rect 19165 -1185 19185 -1165
rect 19165 -1235 19185 -1215
rect 19165 -1285 19185 -1265
rect 19165 -1335 19185 -1315
rect 19165 -1385 19185 -1365
rect 19165 -1435 19185 -1415
rect 19165 -1485 19185 -1465
rect 19165 -1535 19185 -1515
rect 19165 -1585 19185 -1565
rect 19165 -1635 19185 -1615
rect 20365 -985 20385 -965
rect 20365 -1035 20385 -1015
rect 20365 -1085 20385 -1065
rect 20365 -1135 20385 -1115
rect 20365 -1185 20385 -1165
rect 20365 -1235 20385 -1215
rect 20365 -1285 20385 -1265
rect 20365 -1335 20385 -1315
rect 20365 -1385 20385 -1365
rect 20365 -1435 20385 -1415
rect 20365 -1485 20385 -1465
rect 20365 -1535 20385 -1515
rect 20365 -1585 20385 -1565
rect 20365 -1635 20385 -1615
rect 21565 -985 21585 -965
rect 21565 -1035 21585 -1015
rect 21565 -1085 21585 -1065
rect 21565 -1135 21585 -1115
rect 21565 -1185 21585 -1165
rect 21565 -1235 21585 -1215
rect 21565 -1285 21585 -1265
rect 21565 -1335 21585 -1315
rect 21565 -1385 21585 -1365
rect 21565 -1435 21585 -1415
rect 21565 -1485 21585 -1465
rect 21565 -1535 21585 -1515
rect 21565 -1585 21585 -1565
rect 21565 -1635 21585 -1615
rect 22465 -985 22485 -965
rect 22465 -1035 22485 -1015
rect 22465 -1085 22485 -1065
rect 22465 -1135 22485 -1115
rect 22465 -1185 22485 -1165
rect 22465 -1235 22485 -1215
rect 22465 -1285 22485 -1265
rect 22465 -1335 22485 -1315
rect 22465 -1385 22485 -1365
rect 22465 -1435 22485 -1415
rect 22465 -1485 22485 -1465
rect 22465 -1535 22485 -1515
rect 22465 -1585 22485 -1565
rect 22465 -1635 22485 -1615
rect 23365 -985 23385 -965
rect 23365 -1035 23385 -1015
rect 23365 -1085 23385 -1065
rect 23365 -1135 23385 -1115
rect 23365 -1185 23385 -1165
rect 23365 -1235 23385 -1215
rect 23365 -1285 23385 -1265
rect 23365 -1335 23385 -1315
rect 23365 -1385 23385 -1365
rect 23365 -1435 23385 -1415
rect 23365 -1485 23385 -1465
rect 23365 -1535 23385 -1515
rect 23365 -1585 23385 -1565
rect 23365 -1635 23385 -1615
rect 24565 -985 24585 -965
rect 24565 -1035 24585 -1015
rect 24565 -1085 24585 -1065
rect 24565 -1135 24585 -1115
rect 24565 -1185 24585 -1165
rect 24565 -1235 24585 -1215
rect 24565 -1285 24585 -1265
rect 24565 -1335 24585 -1315
rect 24565 -1385 24585 -1365
rect 24565 -1435 24585 -1415
rect 24565 -1485 24585 -1465
rect 24565 -1535 24585 -1515
rect 24565 -1585 24585 -1565
rect 24565 -1635 24585 -1615
rect 25765 -985 25785 -965
rect 25765 -1035 25785 -1015
rect 25765 -1085 25785 -1065
rect 25765 -1135 25785 -1115
rect 25765 -1185 25785 -1165
rect 25765 -1235 25785 -1215
rect 25765 -1285 25785 -1265
rect 25765 -1335 25785 -1315
rect 25765 -1385 25785 -1365
rect 25765 -1435 25785 -1415
rect 25765 -1485 25785 -1465
rect 25765 -1535 25785 -1515
rect 25765 -1585 25785 -1565
rect 25765 -1635 25785 -1615
rect 26665 -985 26685 -965
rect 26665 -1035 26685 -1015
rect 26665 -1085 26685 -1065
rect 26665 -1135 26685 -1115
rect 26665 -1185 26685 -1165
rect 26665 -1235 26685 -1215
rect 26665 -1285 26685 -1265
rect 26665 -1335 26685 -1315
rect 26665 -1385 26685 -1365
rect 26665 -1435 26685 -1415
rect 26665 -1485 26685 -1465
rect 26665 -1535 26685 -1515
rect 26665 -1585 26685 -1565
rect 26665 -1635 26685 -1615
rect 27565 -985 27585 -965
rect 27565 -1035 27585 -1015
rect 27565 -1085 27585 -1065
rect 27565 -1135 27585 -1115
rect 27565 -1185 27585 -1165
rect 27565 -1235 27585 -1215
rect 27565 -1285 27585 -1265
rect 27565 -1335 27585 -1315
rect 27565 -1385 27585 -1365
rect 27565 -1435 27585 -1415
rect 27565 -1485 27585 -1465
rect 27565 -1535 27585 -1515
rect 27565 -1585 27585 -1565
rect 27565 -1635 27585 -1615
rect 28765 -985 28785 -965
rect 28765 -1035 28785 -1015
rect 28765 -1085 28785 -1065
rect 28765 -1135 28785 -1115
rect 28765 -1185 28785 -1165
rect 28765 -1235 28785 -1215
rect 28765 -1285 28785 -1265
rect 28765 -1335 28785 -1315
rect 28765 -1385 28785 -1365
rect 28765 -1435 28785 -1415
rect 28765 -1485 28785 -1465
rect 28765 -1535 28785 -1515
rect 28765 -1585 28785 -1565
rect 28765 -1635 28785 -1615
rect -635 -1735 -615 -1715
rect -35 -1735 -15 -1715
rect 8365 -1735 8385 -1715
rect 10765 -1735 10785 -1715
rect 15565 -1735 15585 -1715
rect 17965 -1735 17985 -1715
rect 20365 -1735 20385 -1715
rect 24565 -1735 24585 -1715
rect 28765 -1735 28785 -1715
<< metal1 >>
rect -650 5590 -600 5600
rect -650 5560 -640 5590
rect -610 5560 -600 5590
rect -650 5485 -600 5560
rect -50 5590 0 5600
rect -50 5560 -40 5590
rect -10 5560 0 5590
rect -650 5465 -635 5485
rect -615 5465 -600 5485
rect -650 5440 -600 5465
rect -650 5410 -640 5440
rect -610 5410 -600 5440
rect -650 5385 -600 5410
rect -650 5365 -635 5385
rect -615 5365 -600 5385
rect -650 5340 -600 5365
rect -650 5310 -640 5340
rect -610 5310 -600 5340
rect -650 5285 -600 5310
rect -650 5265 -635 5285
rect -615 5265 -600 5285
rect -650 5240 -600 5265
rect -650 5210 -640 5240
rect -610 5210 -600 5240
rect -650 5185 -600 5210
rect -650 5165 -635 5185
rect -615 5165 -600 5185
rect -650 5140 -600 5165
rect -650 5110 -640 5140
rect -610 5110 -600 5140
rect -650 5085 -600 5110
rect -650 5065 -635 5085
rect -615 5065 -600 5085
rect -650 5040 -600 5065
rect -650 5010 -640 5040
rect -610 5010 -600 5040
rect -650 4840 -600 5010
rect -500 5485 -450 5500
rect -500 5465 -485 5485
rect -465 5465 -450 5485
rect -500 5435 -450 5465
rect -500 5415 -485 5435
rect -465 5415 -450 5435
rect -500 5385 -450 5415
rect -500 5365 -485 5385
rect -465 5365 -450 5385
rect -500 5335 -450 5365
rect -500 5315 -485 5335
rect -465 5315 -450 5335
rect -500 5285 -450 5315
rect -500 5265 -485 5285
rect -465 5265 -450 5285
rect -500 5235 -450 5265
rect -500 5215 -485 5235
rect -465 5215 -450 5235
rect -500 5185 -450 5215
rect -500 5165 -485 5185
rect -465 5165 -450 5185
rect -500 5135 -450 5165
rect -500 5115 -485 5135
rect -465 5115 -450 5135
rect -500 5085 -450 5115
rect -350 5485 -300 5500
rect -350 5465 -335 5485
rect -315 5465 -300 5485
rect -350 5435 -300 5465
rect -350 5415 -335 5435
rect -315 5415 -300 5435
rect -350 5385 -300 5415
rect -350 5365 -335 5385
rect -315 5365 -300 5385
rect -350 5335 -300 5365
rect -350 5315 -335 5335
rect -315 5315 -300 5335
rect -350 5285 -300 5315
rect -350 5265 -335 5285
rect -315 5265 -300 5285
rect -350 5235 -300 5265
rect -350 5215 -335 5235
rect -315 5215 -300 5235
rect -350 5185 -300 5215
rect -350 5165 -335 5185
rect -315 5165 -300 5185
rect -350 5135 -300 5165
rect -350 5115 -335 5135
rect -315 5115 -300 5135
rect -350 5100 -300 5115
rect -200 5485 -150 5500
rect -200 5465 -185 5485
rect -165 5465 -150 5485
rect -200 5435 -150 5465
rect -200 5415 -185 5435
rect -165 5415 -150 5435
rect -200 5385 -150 5415
rect -200 5365 -185 5385
rect -165 5365 -150 5385
rect -200 5335 -150 5365
rect -200 5315 -185 5335
rect -165 5315 -150 5335
rect -200 5285 -150 5315
rect -200 5265 -185 5285
rect -165 5265 -150 5285
rect -200 5235 -150 5265
rect -200 5215 -185 5235
rect -165 5215 -150 5235
rect -200 5185 -150 5215
rect -200 5165 -185 5185
rect -165 5165 -150 5185
rect -200 5135 -150 5165
rect -200 5115 -185 5135
rect -165 5115 -150 5135
rect -500 5065 -485 5085
rect -465 5065 -450 5085
rect -500 5050 -450 5065
rect -200 5085 -150 5115
rect -200 5065 -185 5085
rect -165 5065 -150 5085
rect -200 5050 -150 5065
rect -500 5035 -150 5050
rect -500 5015 -485 5035
rect -465 5015 -185 5035
rect -165 5015 -150 5035
rect -500 5000 -150 5015
rect -50 5485 0 5560
rect 4150 5590 4200 5600
rect 4150 5560 4160 5590
rect 4190 5560 4200 5590
rect -50 5465 -35 5485
rect -15 5465 0 5485
rect -50 5435 0 5465
rect -50 5415 -35 5435
rect -15 5415 0 5435
rect -50 5385 0 5415
rect -50 5365 -35 5385
rect -15 5365 0 5385
rect -50 5335 0 5365
rect -50 5315 -35 5335
rect -15 5315 0 5335
rect -50 5285 0 5315
rect -50 5265 -35 5285
rect -15 5265 0 5285
rect -50 5235 0 5265
rect -50 5215 -35 5235
rect -15 5215 0 5235
rect -50 5185 0 5215
rect -50 5165 -35 5185
rect -15 5165 0 5185
rect -50 5135 0 5165
rect -50 5115 -35 5135
rect -15 5115 0 5135
rect -500 4940 -450 4950
rect -500 4910 -490 4940
rect -460 4910 -450 4940
rect -500 4900 -450 4910
rect -350 4940 -300 5000
rect -350 4910 -340 4940
rect -310 4910 -300 4940
rect -350 4850 -300 4910
rect -200 4940 -150 4950
rect -200 4910 -190 4940
rect -160 4910 -150 4940
rect -200 4900 -150 4910
rect -650 4810 -640 4840
rect -610 4810 -600 4840
rect -650 4785 -600 4810
rect -650 4765 -635 4785
rect -615 4765 -600 4785
rect -650 4740 -600 4765
rect -650 4710 -640 4740
rect -610 4710 -600 4740
rect -650 4685 -600 4710
rect -650 4665 -635 4685
rect -615 4665 -600 4685
rect -650 4640 -600 4665
rect -650 4610 -640 4640
rect -610 4610 -600 4640
rect -650 4585 -600 4610
rect -650 4565 -635 4585
rect -615 4565 -600 4585
rect -650 4540 -600 4565
rect -650 4510 -640 4540
rect -610 4510 -600 4540
rect -650 4485 -600 4510
rect -650 4465 -635 4485
rect -615 4465 -600 4485
rect -650 4440 -600 4465
rect -650 4410 -640 4440
rect -610 4410 -600 4440
rect -650 4385 -600 4410
rect -650 4365 -635 4385
rect -615 4365 -600 4385
rect -650 4290 -600 4365
rect -500 4835 -150 4850
rect -500 4815 -485 4835
rect -465 4815 -185 4835
rect -165 4815 -150 4835
rect -500 4800 -150 4815
rect -500 4785 -450 4800
rect -500 4765 -485 4785
rect -465 4765 -450 4785
rect -500 4735 -450 4765
rect -200 4785 -150 4800
rect -200 4765 -185 4785
rect -165 4765 -150 4785
rect -500 4715 -485 4735
rect -465 4715 -450 4735
rect -500 4685 -450 4715
rect -500 4665 -485 4685
rect -465 4665 -450 4685
rect -500 4635 -450 4665
rect -500 4615 -485 4635
rect -465 4615 -450 4635
rect -500 4585 -450 4615
rect -500 4565 -485 4585
rect -465 4565 -450 4585
rect -500 4535 -450 4565
rect -500 4515 -485 4535
rect -465 4515 -450 4535
rect -500 4485 -450 4515
rect -500 4465 -485 4485
rect -465 4465 -450 4485
rect -500 4435 -450 4465
rect -500 4415 -485 4435
rect -465 4415 -450 4435
rect -500 4385 -450 4415
rect -500 4365 -485 4385
rect -465 4365 -450 4385
rect -500 4350 -450 4365
rect -350 4735 -300 4750
rect -350 4715 -335 4735
rect -315 4715 -300 4735
rect -350 4685 -300 4715
rect -350 4665 -335 4685
rect -315 4665 -300 4685
rect -350 4635 -300 4665
rect -350 4615 -335 4635
rect -315 4615 -300 4635
rect -350 4585 -300 4615
rect -350 4565 -335 4585
rect -315 4565 -300 4585
rect -350 4535 -300 4565
rect -350 4515 -335 4535
rect -315 4515 -300 4535
rect -350 4485 -300 4515
rect -350 4465 -335 4485
rect -315 4465 -300 4485
rect -350 4435 -300 4465
rect -350 4415 -335 4435
rect -315 4415 -300 4435
rect -350 4385 -300 4415
rect -350 4365 -335 4385
rect -315 4365 -300 4385
rect -350 4350 -300 4365
rect -200 4735 -150 4765
rect -200 4715 -185 4735
rect -165 4715 -150 4735
rect -200 4685 -150 4715
rect -200 4665 -185 4685
rect -165 4665 -150 4685
rect -200 4635 -150 4665
rect -200 4615 -185 4635
rect -165 4615 -150 4635
rect -200 4585 -150 4615
rect -200 4565 -185 4585
rect -165 4565 -150 4585
rect -200 4535 -150 4565
rect -200 4515 -185 4535
rect -165 4515 -150 4535
rect -200 4485 -150 4515
rect -200 4465 -185 4485
rect -165 4465 -150 4485
rect -200 4435 -150 4465
rect -200 4415 -185 4435
rect -165 4415 -150 4435
rect -200 4385 -150 4415
rect -200 4365 -185 4385
rect -165 4365 -150 4385
rect -200 4350 -150 4365
rect -50 4840 0 5115
rect 550 5485 3600 5500
rect 550 5465 565 5485
rect 585 5465 865 5485
rect 885 5465 1165 5485
rect 1185 5465 1465 5485
rect 1485 5465 1765 5485
rect 1785 5465 2065 5485
rect 2085 5465 2365 5485
rect 2385 5465 2665 5485
rect 2685 5465 2965 5485
rect 2985 5465 3265 5485
rect 3285 5465 3565 5485
rect 3585 5465 3600 5485
rect 550 5450 3600 5465
rect 550 5435 600 5450
rect 550 5415 565 5435
rect 585 5415 600 5435
rect 550 5385 600 5415
rect 850 5435 900 5450
rect 850 5415 865 5435
rect 885 5415 900 5435
rect 550 5365 565 5385
rect 585 5365 600 5385
rect 550 5335 600 5365
rect 550 5315 565 5335
rect 585 5315 600 5335
rect 550 5285 600 5315
rect 550 5265 565 5285
rect 585 5265 600 5285
rect 550 5235 600 5265
rect 550 5215 565 5235
rect 585 5215 600 5235
rect 550 5185 600 5215
rect 550 5165 565 5185
rect 585 5165 600 5185
rect 550 5135 600 5165
rect 550 5115 565 5135
rect 585 5115 600 5135
rect 550 5085 600 5115
rect 550 5065 565 5085
rect 585 5065 600 5085
rect 550 5035 600 5065
rect 550 5015 565 5035
rect 585 5015 600 5035
rect 550 5000 600 5015
rect 700 5385 750 5400
rect 700 5365 715 5385
rect 735 5365 750 5385
rect 700 5335 750 5365
rect 700 5315 715 5335
rect 735 5315 750 5335
rect 700 5285 750 5315
rect 700 5265 715 5285
rect 735 5265 750 5285
rect 700 5235 750 5265
rect 700 5215 715 5235
rect 735 5215 750 5235
rect 700 5185 750 5215
rect 700 5165 715 5185
rect 735 5165 750 5185
rect 700 5135 750 5165
rect 700 5115 715 5135
rect 735 5115 750 5135
rect 700 5085 750 5115
rect 850 5385 900 5415
rect 1150 5435 1200 5450
rect 1150 5415 1165 5435
rect 1185 5415 1200 5435
rect 850 5365 865 5385
rect 885 5365 900 5385
rect 850 5335 900 5365
rect 850 5315 865 5335
rect 885 5315 900 5335
rect 850 5285 900 5315
rect 850 5265 865 5285
rect 885 5265 900 5285
rect 850 5235 900 5265
rect 850 5215 865 5235
rect 885 5215 900 5235
rect 850 5185 900 5215
rect 850 5165 865 5185
rect 885 5165 900 5185
rect 850 5135 900 5165
rect 850 5115 865 5135
rect 885 5115 900 5135
rect 850 5100 900 5115
rect 1000 5385 1050 5400
rect 1000 5365 1015 5385
rect 1035 5365 1050 5385
rect 1000 5335 1050 5365
rect 1000 5315 1015 5335
rect 1035 5315 1050 5335
rect 1000 5285 1050 5315
rect 1000 5265 1015 5285
rect 1035 5265 1050 5285
rect 1000 5235 1050 5265
rect 1000 5215 1015 5235
rect 1035 5215 1050 5235
rect 1000 5185 1050 5215
rect 1000 5165 1015 5185
rect 1035 5165 1050 5185
rect 1000 5135 1050 5165
rect 1000 5115 1015 5135
rect 1035 5115 1050 5135
rect 700 5065 715 5085
rect 735 5065 750 5085
rect 700 5050 750 5065
rect 1000 5085 1050 5115
rect 1150 5385 1200 5415
rect 1450 5435 1500 5450
rect 1450 5415 1465 5435
rect 1485 5415 1500 5435
rect 1150 5365 1165 5385
rect 1185 5365 1200 5385
rect 1150 5335 1200 5365
rect 1150 5315 1165 5335
rect 1185 5315 1200 5335
rect 1150 5285 1200 5315
rect 1150 5265 1165 5285
rect 1185 5265 1200 5285
rect 1150 5235 1200 5265
rect 1150 5215 1165 5235
rect 1185 5215 1200 5235
rect 1150 5185 1200 5215
rect 1150 5165 1165 5185
rect 1185 5165 1200 5185
rect 1150 5135 1200 5165
rect 1150 5115 1165 5135
rect 1185 5115 1200 5135
rect 1150 5100 1200 5115
rect 1300 5385 1350 5400
rect 1300 5365 1315 5385
rect 1335 5365 1350 5385
rect 1300 5335 1350 5365
rect 1300 5315 1315 5335
rect 1335 5315 1350 5335
rect 1300 5285 1350 5315
rect 1300 5265 1315 5285
rect 1335 5265 1350 5285
rect 1300 5235 1350 5265
rect 1300 5215 1315 5235
rect 1335 5215 1350 5235
rect 1300 5185 1350 5215
rect 1300 5165 1315 5185
rect 1335 5165 1350 5185
rect 1300 5135 1350 5165
rect 1300 5115 1315 5135
rect 1335 5115 1350 5135
rect 1000 5065 1015 5085
rect 1035 5065 1050 5085
rect 1000 5050 1050 5065
rect 1300 5085 1350 5115
rect 1450 5385 1500 5415
rect 1750 5435 1800 5450
rect 1750 5415 1765 5435
rect 1785 5415 1800 5435
rect 1450 5365 1465 5385
rect 1485 5365 1500 5385
rect 1450 5335 1500 5365
rect 1450 5315 1465 5335
rect 1485 5315 1500 5335
rect 1450 5285 1500 5315
rect 1450 5265 1465 5285
rect 1485 5265 1500 5285
rect 1450 5235 1500 5265
rect 1450 5215 1465 5235
rect 1485 5215 1500 5235
rect 1450 5185 1500 5215
rect 1450 5165 1465 5185
rect 1485 5165 1500 5185
rect 1450 5135 1500 5165
rect 1450 5115 1465 5135
rect 1485 5115 1500 5135
rect 1450 5100 1500 5115
rect 1600 5385 1650 5400
rect 1600 5365 1615 5385
rect 1635 5365 1650 5385
rect 1600 5335 1650 5365
rect 1600 5315 1615 5335
rect 1635 5315 1650 5335
rect 1600 5285 1650 5315
rect 1600 5265 1615 5285
rect 1635 5265 1650 5285
rect 1600 5235 1650 5265
rect 1600 5215 1615 5235
rect 1635 5215 1650 5235
rect 1600 5185 1650 5215
rect 1600 5165 1615 5185
rect 1635 5165 1650 5185
rect 1600 5135 1650 5165
rect 1600 5115 1615 5135
rect 1635 5115 1650 5135
rect 1300 5065 1315 5085
rect 1335 5065 1350 5085
rect 1300 5050 1350 5065
rect 1600 5085 1650 5115
rect 1600 5065 1615 5085
rect 1635 5065 1650 5085
rect 1600 5050 1650 5065
rect 700 5035 1650 5050
rect 700 5015 715 5035
rect 735 5015 1650 5035
rect 700 5000 1650 5015
rect 1750 5385 1800 5415
rect 2050 5435 2100 5450
rect 2050 5415 2065 5435
rect 2085 5415 2100 5435
rect 1750 5365 1765 5385
rect 1785 5365 1800 5385
rect 1750 5335 1800 5365
rect 1750 5315 1765 5335
rect 1785 5315 1800 5335
rect 1750 5285 1800 5315
rect 1750 5265 1765 5285
rect 1785 5265 1800 5285
rect 1750 5235 1800 5265
rect 1750 5215 1765 5235
rect 1785 5215 1800 5235
rect 1750 5185 1800 5215
rect 1750 5165 1765 5185
rect 1785 5165 1800 5185
rect 1750 5135 1800 5165
rect 1750 5115 1765 5135
rect 1785 5115 1800 5135
rect 1750 5085 1800 5115
rect 1750 5065 1765 5085
rect 1785 5065 1800 5085
rect 1750 5035 1800 5065
rect 1750 5015 1765 5035
rect 1785 5015 1800 5035
rect 100 4940 150 4950
rect 100 4910 110 4940
rect 140 4910 150 4940
rect 100 4900 150 4910
rect 400 4940 450 4950
rect 400 4910 410 4940
rect 440 4910 450 4940
rect 400 4900 450 4910
rect 700 4940 750 4950
rect 700 4910 710 4940
rect 740 4910 750 4940
rect 700 4900 750 4910
rect 1000 4940 1050 4950
rect 1000 4910 1010 4940
rect 1040 4910 1050 4940
rect 1000 4900 1050 4910
rect 1150 4940 1200 4950
rect 1150 4910 1160 4940
rect 1190 4910 1200 4940
rect 1150 4900 1200 4910
rect 1300 4940 1350 4950
rect 1300 4910 1310 4940
rect 1340 4910 1350 4940
rect 1300 4900 1350 4910
rect 1600 4940 1650 4950
rect 1600 4910 1610 4940
rect 1640 4910 1650 4940
rect 1600 4900 1650 4910
rect -50 4810 -40 4840
rect -10 4810 0 4840
rect -50 4740 0 4810
rect -50 4710 -40 4740
rect -10 4710 0 4740
rect -50 4685 0 4710
rect -50 4665 -35 4685
rect -15 4665 0 4685
rect -50 4640 0 4665
rect -50 4610 -40 4640
rect -10 4610 0 4640
rect -50 4585 0 4610
rect -50 4565 -35 4585
rect -15 4565 0 4585
rect -50 4540 0 4565
rect -50 4510 -40 4540
rect -10 4510 0 4540
rect -50 4485 0 4510
rect -50 4465 -35 4485
rect -15 4465 0 4485
rect -50 4440 0 4465
rect -50 4410 -40 4440
rect -10 4410 0 4440
rect -50 4385 0 4410
rect -50 4365 -35 4385
rect -15 4365 0 4385
rect -650 4260 -640 4290
rect -610 4260 -600 4290
rect -650 4185 -600 4260
rect -50 4290 0 4365
rect 550 4835 600 4850
rect 550 4815 565 4835
rect 585 4815 600 4835
rect 550 4785 600 4815
rect 550 4765 565 4785
rect 585 4765 600 4785
rect 550 4735 600 4765
rect 550 4715 565 4735
rect 585 4715 600 4735
rect 550 4685 600 4715
rect 550 4665 565 4685
rect 585 4665 600 4685
rect 550 4635 600 4665
rect 550 4615 565 4635
rect 585 4615 600 4635
rect 550 4585 600 4615
rect 550 4565 565 4585
rect 585 4565 600 4585
rect 550 4535 600 4565
rect 550 4515 565 4535
rect 585 4515 600 4535
rect 550 4485 600 4515
rect 550 4465 565 4485
rect 585 4465 600 4485
rect 550 4435 600 4465
rect 700 4835 1650 4850
rect 700 4815 715 4835
rect 735 4815 1650 4835
rect 700 4800 1650 4815
rect 700 4785 750 4800
rect 700 4765 715 4785
rect 735 4765 750 4785
rect 700 4735 750 4765
rect 1000 4785 1050 4800
rect 1000 4765 1015 4785
rect 1035 4765 1050 4785
rect 700 4715 715 4735
rect 735 4715 750 4735
rect 700 4685 750 4715
rect 700 4665 715 4685
rect 735 4665 750 4685
rect 700 4635 750 4665
rect 700 4615 715 4635
rect 735 4615 750 4635
rect 700 4585 750 4615
rect 700 4565 715 4585
rect 735 4565 750 4585
rect 700 4535 750 4565
rect 700 4515 715 4535
rect 735 4515 750 4535
rect 700 4485 750 4515
rect 700 4465 715 4485
rect 735 4465 750 4485
rect 700 4450 750 4465
rect 850 4735 900 4750
rect 850 4715 865 4735
rect 885 4715 900 4735
rect 850 4685 900 4715
rect 850 4665 865 4685
rect 885 4665 900 4685
rect 850 4635 900 4665
rect 850 4615 865 4635
rect 885 4615 900 4635
rect 850 4585 900 4615
rect 850 4565 865 4585
rect 885 4565 900 4585
rect 850 4535 900 4565
rect 850 4515 865 4535
rect 885 4515 900 4535
rect 850 4485 900 4515
rect 850 4465 865 4485
rect 885 4465 900 4485
rect 550 4415 565 4435
rect 585 4415 600 4435
rect 550 4400 600 4415
rect 850 4435 900 4465
rect 1000 4735 1050 4765
rect 1300 4785 1350 4800
rect 1300 4765 1315 4785
rect 1335 4765 1350 4785
rect 1000 4715 1015 4735
rect 1035 4715 1050 4735
rect 1000 4685 1050 4715
rect 1000 4665 1015 4685
rect 1035 4665 1050 4685
rect 1000 4635 1050 4665
rect 1000 4615 1015 4635
rect 1035 4615 1050 4635
rect 1000 4585 1050 4615
rect 1000 4565 1015 4585
rect 1035 4565 1050 4585
rect 1000 4535 1050 4565
rect 1000 4515 1015 4535
rect 1035 4515 1050 4535
rect 1000 4485 1050 4515
rect 1000 4465 1015 4485
rect 1035 4465 1050 4485
rect 1000 4450 1050 4465
rect 1150 4735 1200 4750
rect 1150 4715 1165 4735
rect 1185 4715 1200 4735
rect 1150 4685 1200 4715
rect 1150 4665 1165 4685
rect 1185 4665 1200 4685
rect 1150 4635 1200 4665
rect 1150 4615 1165 4635
rect 1185 4615 1200 4635
rect 1150 4585 1200 4615
rect 1150 4565 1165 4585
rect 1185 4565 1200 4585
rect 1150 4535 1200 4565
rect 1150 4515 1165 4535
rect 1185 4515 1200 4535
rect 1150 4485 1200 4515
rect 1150 4465 1165 4485
rect 1185 4465 1200 4485
rect 850 4415 865 4435
rect 885 4415 900 4435
rect 850 4400 900 4415
rect 1150 4435 1200 4465
rect 1300 4735 1350 4765
rect 1600 4785 1650 4800
rect 1600 4765 1615 4785
rect 1635 4765 1650 4785
rect 1300 4715 1315 4735
rect 1335 4715 1350 4735
rect 1300 4685 1350 4715
rect 1300 4665 1315 4685
rect 1335 4665 1350 4685
rect 1300 4635 1350 4665
rect 1300 4615 1315 4635
rect 1335 4615 1350 4635
rect 1300 4585 1350 4615
rect 1300 4565 1315 4585
rect 1335 4565 1350 4585
rect 1300 4535 1350 4565
rect 1300 4515 1315 4535
rect 1335 4515 1350 4535
rect 1300 4485 1350 4515
rect 1300 4465 1315 4485
rect 1335 4465 1350 4485
rect 1300 4450 1350 4465
rect 1450 4735 1500 4750
rect 1450 4715 1465 4735
rect 1485 4715 1500 4735
rect 1450 4685 1500 4715
rect 1450 4665 1465 4685
rect 1485 4665 1500 4685
rect 1450 4635 1500 4665
rect 1450 4615 1465 4635
rect 1485 4615 1500 4635
rect 1450 4585 1500 4615
rect 1450 4565 1465 4585
rect 1485 4565 1500 4585
rect 1450 4535 1500 4565
rect 1450 4515 1465 4535
rect 1485 4515 1500 4535
rect 1450 4485 1500 4515
rect 1450 4465 1465 4485
rect 1485 4465 1500 4485
rect 1150 4415 1165 4435
rect 1185 4415 1200 4435
rect 1150 4400 1200 4415
rect 1450 4435 1500 4465
rect 1600 4735 1650 4765
rect 1600 4715 1615 4735
rect 1635 4715 1650 4735
rect 1600 4685 1650 4715
rect 1600 4665 1615 4685
rect 1635 4665 1650 4685
rect 1600 4635 1650 4665
rect 1600 4615 1615 4635
rect 1635 4615 1650 4635
rect 1600 4585 1650 4615
rect 1600 4565 1615 4585
rect 1635 4565 1650 4585
rect 1600 4535 1650 4565
rect 1600 4515 1615 4535
rect 1635 4515 1650 4535
rect 1600 4485 1650 4515
rect 1600 4465 1615 4485
rect 1635 4465 1650 4485
rect 1600 4450 1650 4465
rect 1750 4835 1800 5015
rect 1900 5385 1950 5400
rect 1900 5365 1915 5385
rect 1935 5365 1950 5385
rect 1900 5335 1950 5365
rect 1900 5315 1915 5335
rect 1935 5315 1950 5335
rect 1900 5285 1950 5315
rect 1900 5265 1915 5285
rect 1935 5265 1950 5285
rect 1900 5235 1950 5265
rect 1900 5215 1915 5235
rect 1935 5215 1950 5235
rect 1900 5185 1950 5215
rect 1900 5165 1915 5185
rect 1935 5165 1950 5185
rect 1900 5135 1950 5165
rect 1900 5115 1915 5135
rect 1935 5115 1950 5135
rect 1900 5085 1950 5115
rect 2050 5385 2100 5415
rect 2350 5435 2400 5450
rect 2350 5415 2365 5435
rect 2385 5415 2400 5435
rect 2050 5365 2065 5385
rect 2085 5365 2100 5385
rect 2050 5335 2100 5365
rect 2050 5315 2065 5335
rect 2085 5315 2100 5335
rect 2050 5285 2100 5315
rect 2050 5265 2065 5285
rect 2085 5265 2100 5285
rect 2050 5235 2100 5265
rect 2050 5215 2065 5235
rect 2085 5215 2100 5235
rect 2050 5185 2100 5215
rect 2050 5165 2065 5185
rect 2085 5165 2100 5185
rect 2050 5135 2100 5165
rect 2050 5115 2065 5135
rect 2085 5115 2100 5135
rect 2050 5100 2100 5115
rect 2200 5385 2250 5400
rect 2200 5365 2215 5385
rect 2235 5365 2250 5385
rect 2200 5335 2250 5365
rect 2200 5315 2215 5335
rect 2235 5315 2250 5335
rect 2200 5285 2250 5315
rect 2200 5265 2215 5285
rect 2235 5265 2250 5285
rect 2200 5235 2250 5265
rect 2200 5215 2215 5235
rect 2235 5215 2250 5235
rect 2200 5185 2250 5215
rect 2200 5165 2215 5185
rect 2235 5165 2250 5185
rect 2200 5135 2250 5165
rect 2200 5115 2215 5135
rect 2235 5115 2250 5135
rect 1900 5065 1915 5085
rect 1935 5065 1950 5085
rect 1900 5050 1950 5065
rect 2200 5085 2250 5115
rect 2200 5065 2215 5085
rect 2235 5065 2250 5085
rect 2200 5050 2250 5065
rect 1900 5035 2250 5050
rect 1900 5015 1915 5035
rect 1935 5015 2215 5035
rect 2235 5015 2250 5035
rect 1900 5000 2250 5015
rect 2350 5385 2400 5415
rect 2650 5435 2700 5450
rect 2650 5415 2665 5435
rect 2685 5415 2700 5435
rect 2350 5365 2365 5385
rect 2385 5365 2400 5385
rect 2350 5335 2400 5365
rect 2350 5315 2365 5335
rect 2385 5315 2400 5335
rect 2350 5285 2400 5315
rect 2350 5265 2365 5285
rect 2385 5265 2400 5285
rect 2350 5235 2400 5265
rect 2350 5215 2365 5235
rect 2385 5215 2400 5235
rect 2350 5185 2400 5215
rect 2350 5165 2365 5185
rect 2385 5165 2400 5185
rect 2350 5135 2400 5165
rect 2350 5115 2365 5135
rect 2385 5115 2400 5135
rect 2350 5085 2400 5115
rect 2350 5065 2365 5085
rect 2385 5065 2400 5085
rect 2350 5035 2400 5065
rect 2350 5015 2365 5035
rect 2385 5015 2400 5035
rect 1900 4940 1950 4950
rect 1900 4910 1910 4940
rect 1940 4910 1950 4940
rect 1900 4900 1950 4910
rect 2050 4940 2100 5000
rect 2050 4910 2060 4940
rect 2090 4910 2100 4940
rect 2050 4850 2100 4910
rect 2200 4940 2250 4950
rect 2200 4910 2210 4940
rect 2240 4910 2250 4940
rect 2200 4900 2250 4910
rect 1750 4815 1765 4835
rect 1785 4815 1800 4835
rect 1750 4785 1800 4815
rect 1750 4765 1765 4785
rect 1785 4765 1800 4785
rect 1750 4735 1800 4765
rect 1750 4715 1765 4735
rect 1785 4715 1800 4735
rect 1750 4685 1800 4715
rect 1750 4665 1765 4685
rect 1785 4665 1800 4685
rect 1750 4635 1800 4665
rect 1750 4615 1765 4635
rect 1785 4615 1800 4635
rect 1750 4585 1800 4615
rect 1750 4565 1765 4585
rect 1785 4565 1800 4585
rect 1750 4535 1800 4565
rect 1750 4515 1765 4535
rect 1785 4515 1800 4535
rect 1750 4485 1800 4515
rect 1750 4465 1765 4485
rect 1785 4465 1800 4485
rect 1450 4415 1465 4435
rect 1485 4415 1500 4435
rect 1450 4400 1500 4415
rect 1750 4435 1800 4465
rect 1900 4835 2250 4850
rect 1900 4815 1915 4835
rect 1935 4815 2215 4835
rect 2235 4815 2250 4835
rect 1900 4800 2250 4815
rect 1900 4785 1950 4800
rect 1900 4765 1915 4785
rect 1935 4765 1950 4785
rect 1900 4735 1950 4765
rect 2200 4785 2250 4800
rect 2200 4765 2215 4785
rect 2235 4765 2250 4785
rect 1900 4715 1915 4735
rect 1935 4715 1950 4735
rect 1900 4685 1950 4715
rect 1900 4665 1915 4685
rect 1935 4665 1950 4685
rect 1900 4635 1950 4665
rect 1900 4615 1915 4635
rect 1935 4615 1950 4635
rect 1900 4585 1950 4615
rect 1900 4565 1915 4585
rect 1935 4565 1950 4585
rect 1900 4535 1950 4565
rect 1900 4515 1915 4535
rect 1935 4515 1950 4535
rect 1900 4485 1950 4515
rect 1900 4465 1915 4485
rect 1935 4465 1950 4485
rect 1900 4450 1950 4465
rect 2050 4735 2100 4750
rect 2050 4715 2065 4735
rect 2085 4715 2100 4735
rect 2050 4685 2100 4715
rect 2050 4665 2065 4685
rect 2085 4665 2100 4685
rect 2050 4635 2100 4665
rect 2050 4615 2065 4635
rect 2085 4615 2100 4635
rect 2050 4585 2100 4615
rect 2050 4565 2065 4585
rect 2085 4565 2100 4585
rect 2050 4535 2100 4565
rect 2050 4515 2065 4535
rect 2085 4515 2100 4535
rect 2050 4485 2100 4515
rect 2050 4465 2065 4485
rect 2085 4465 2100 4485
rect 1750 4415 1765 4435
rect 1785 4415 1800 4435
rect 1750 4400 1800 4415
rect 2050 4435 2100 4465
rect 2200 4735 2250 4765
rect 2200 4715 2215 4735
rect 2235 4715 2250 4735
rect 2200 4685 2250 4715
rect 2200 4665 2215 4685
rect 2235 4665 2250 4685
rect 2200 4635 2250 4665
rect 2200 4615 2215 4635
rect 2235 4615 2250 4635
rect 2200 4585 2250 4615
rect 2200 4565 2215 4585
rect 2235 4565 2250 4585
rect 2200 4535 2250 4565
rect 2200 4515 2215 4535
rect 2235 4515 2250 4535
rect 2200 4485 2250 4515
rect 2200 4465 2215 4485
rect 2235 4465 2250 4485
rect 2200 4450 2250 4465
rect 2350 4835 2400 5015
rect 2500 5385 2550 5400
rect 2500 5365 2515 5385
rect 2535 5365 2550 5385
rect 2500 5335 2550 5365
rect 2500 5315 2515 5335
rect 2535 5315 2550 5335
rect 2500 5285 2550 5315
rect 2500 5265 2515 5285
rect 2535 5265 2550 5285
rect 2500 5235 2550 5265
rect 2500 5215 2515 5235
rect 2535 5215 2550 5235
rect 2500 5185 2550 5215
rect 2500 5165 2515 5185
rect 2535 5165 2550 5185
rect 2500 5135 2550 5165
rect 2500 5115 2515 5135
rect 2535 5115 2550 5135
rect 2500 5085 2550 5115
rect 2650 5385 2700 5415
rect 2950 5435 3000 5450
rect 2950 5415 2965 5435
rect 2985 5415 3000 5435
rect 2650 5365 2665 5385
rect 2685 5365 2700 5385
rect 2650 5335 2700 5365
rect 2650 5315 2665 5335
rect 2685 5315 2700 5335
rect 2650 5285 2700 5315
rect 2650 5265 2665 5285
rect 2685 5265 2700 5285
rect 2650 5235 2700 5265
rect 2650 5215 2665 5235
rect 2685 5215 2700 5235
rect 2650 5185 2700 5215
rect 2650 5165 2665 5185
rect 2685 5165 2700 5185
rect 2650 5135 2700 5165
rect 2650 5115 2665 5135
rect 2685 5115 2700 5135
rect 2650 5100 2700 5115
rect 2800 5385 2850 5400
rect 2800 5365 2815 5385
rect 2835 5365 2850 5385
rect 2800 5335 2850 5365
rect 2800 5315 2815 5335
rect 2835 5315 2850 5335
rect 2800 5285 2850 5315
rect 2800 5265 2815 5285
rect 2835 5265 2850 5285
rect 2800 5235 2850 5265
rect 2800 5215 2815 5235
rect 2835 5215 2850 5235
rect 2800 5185 2850 5215
rect 2800 5165 2815 5185
rect 2835 5165 2850 5185
rect 2800 5135 2850 5165
rect 2800 5115 2815 5135
rect 2835 5115 2850 5135
rect 2500 5065 2515 5085
rect 2535 5065 2550 5085
rect 2500 5050 2550 5065
rect 2800 5085 2850 5115
rect 2950 5385 3000 5415
rect 3250 5435 3300 5450
rect 3250 5415 3265 5435
rect 3285 5415 3300 5435
rect 2950 5365 2965 5385
rect 2985 5365 3000 5385
rect 2950 5335 3000 5365
rect 2950 5315 2965 5335
rect 2985 5315 3000 5335
rect 2950 5285 3000 5315
rect 2950 5265 2965 5285
rect 2985 5265 3000 5285
rect 2950 5235 3000 5265
rect 2950 5215 2965 5235
rect 2985 5215 3000 5235
rect 2950 5185 3000 5215
rect 2950 5165 2965 5185
rect 2985 5165 3000 5185
rect 2950 5135 3000 5165
rect 2950 5115 2965 5135
rect 2985 5115 3000 5135
rect 2950 5100 3000 5115
rect 3100 5385 3150 5400
rect 3100 5365 3115 5385
rect 3135 5365 3150 5385
rect 3100 5335 3150 5365
rect 3100 5315 3115 5335
rect 3135 5315 3150 5335
rect 3100 5285 3150 5315
rect 3100 5265 3115 5285
rect 3135 5265 3150 5285
rect 3100 5235 3150 5265
rect 3100 5215 3115 5235
rect 3135 5215 3150 5235
rect 3100 5185 3150 5215
rect 3100 5165 3115 5185
rect 3135 5165 3150 5185
rect 3100 5135 3150 5165
rect 3100 5115 3115 5135
rect 3135 5115 3150 5135
rect 2800 5065 2815 5085
rect 2835 5065 2850 5085
rect 2800 5050 2850 5065
rect 3100 5085 3150 5115
rect 3250 5385 3300 5415
rect 3550 5435 3600 5450
rect 3550 5415 3565 5435
rect 3585 5415 3600 5435
rect 3250 5365 3265 5385
rect 3285 5365 3300 5385
rect 3250 5335 3300 5365
rect 3250 5315 3265 5335
rect 3285 5315 3300 5335
rect 3250 5285 3300 5315
rect 3250 5265 3265 5285
rect 3285 5265 3300 5285
rect 3250 5235 3300 5265
rect 3250 5215 3265 5235
rect 3285 5215 3300 5235
rect 3250 5185 3300 5215
rect 3250 5165 3265 5185
rect 3285 5165 3300 5185
rect 3250 5135 3300 5165
rect 3250 5115 3265 5135
rect 3285 5115 3300 5135
rect 3250 5100 3300 5115
rect 3400 5385 3450 5400
rect 3400 5365 3415 5385
rect 3435 5365 3450 5385
rect 3400 5335 3450 5365
rect 3400 5315 3415 5335
rect 3435 5315 3450 5335
rect 3400 5285 3450 5315
rect 3400 5265 3415 5285
rect 3435 5265 3450 5285
rect 3400 5235 3450 5265
rect 3400 5215 3415 5235
rect 3435 5215 3450 5235
rect 3400 5185 3450 5215
rect 3400 5165 3415 5185
rect 3435 5165 3450 5185
rect 3400 5135 3450 5165
rect 3400 5115 3415 5135
rect 3435 5115 3450 5135
rect 3100 5065 3115 5085
rect 3135 5065 3150 5085
rect 3100 5050 3150 5065
rect 3400 5085 3450 5115
rect 3400 5065 3415 5085
rect 3435 5065 3450 5085
rect 3400 5050 3450 5065
rect 2500 5035 3450 5050
rect 2500 5015 3415 5035
rect 3435 5015 3450 5035
rect 2500 5000 3450 5015
rect 3550 5385 3600 5415
rect 3550 5365 3565 5385
rect 3585 5365 3600 5385
rect 3550 5335 3600 5365
rect 3550 5315 3565 5335
rect 3585 5315 3600 5335
rect 3550 5285 3600 5315
rect 3550 5265 3565 5285
rect 3585 5265 3600 5285
rect 3550 5235 3600 5265
rect 3550 5215 3565 5235
rect 3585 5215 3600 5235
rect 3550 5185 3600 5215
rect 3550 5165 3565 5185
rect 3585 5165 3600 5185
rect 3550 5135 3600 5165
rect 3550 5115 3565 5135
rect 3585 5115 3600 5135
rect 3550 5085 3600 5115
rect 3550 5065 3565 5085
rect 3585 5065 3600 5085
rect 3550 5035 3600 5065
rect 3550 5015 3565 5035
rect 3585 5015 3600 5035
rect 3550 5000 3600 5015
rect 4150 5485 4200 5560
rect 8350 5590 8400 5600
rect 8350 5560 8360 5590
rect 8390 5560 8400 5590
rect 4150 5465 4165 5485
rect 4185 5465 4200 5485
rect 4150 5435 4200 5465
rect 4150 5415 4165 5435
rect 4185 5415 4200 5435
rect 4150 5385 4200 5415
rect 4150 5365 4165 5385
rect 4185 5365 4200 5385
rect 4150 5335 4200 5365
rect 4150 5315 4165 5335
rect 4185 5315 4200 5335
rect 4150 5285 4200 5315
rect 4150 5265 4165 5285
rect 4185 5265 4200 5285
rect 4150 5235 4200 5265
rect 4150 5215 4165 5235
rect 4185 5215 4200 5235
rect 4150 5185 4200 5215
rect 4150 5165 4165 5185
rect 4185 5165 4200 5185
rect 4150 5135 4200 5165
rect 4150 5115 4165 5135
rect 4185 5115 4200 5135
rect 2500 4940 2550 4950
rect 2500 4910 2510 4940
rect 2540 4910 2550 4940
rect 2500 4900 2550 4910
rect 2800 4940 2850 4950
rect 2800 4910 2810 4940
rect 2840 4910 2850 4940
rect 2800 4900 2850 4910
rect 2950 4940 3000 4950
rect 2950 4910 2960 4940
rect 2990 4910 3000 4940
rect 2950 4900 3000 4910
rect 3100 4940 3150 4950
rect 3100 4910 3110 4940
rect 3140 4910 3150 4940
rect 3100 4900 3150 4910
rect 3400 4940 3450 4950
rect 3400 4910 3410 4940
rect 3440 4910 3450 4940
rect 3400 4900 3450 4910
rect 3700 4940 3750 4950
rect 3700 4910 3710 4940
rect 3740 4910 3750 4940
rect 3700 4900 3750 4910
rect 4000 4940 4050 4950
rect 4000 4910 4010 4940
rect 4040 4910 4050 4940
rect 4000 4900 4050 4910
rect 2350 4815 2365 4835
rect 2385 4815 2400 4835
rect 2350 4785 2400 4815
rect 2350 4765 2365 4785
rect 2385 4765 2400 4785
rect 2350 4735 2400 4765
rect 2350 4715 2365 4735
rect 2385 4715 2400 4735
rect 2350 4685 2400 4715
rect 2350 4665 2365 4685
rect 2385 4665 2400 4685
rect 2350 4635 2400 4665
rect 2350 4615 2365 4635
rect 2385 4615 2400 4635
rect 2350 4585 2400 4615
rect 2350 4565 2365 4585
rect 2385 4565 2400 4585
rect 2350 4535 2400 4565
rect 2350 4515 2365 4535
rect 2385 4515 2400 4535
rect 2350 4485 2400 4515
rect 2350 4465 2365 4485
rect 2385 4465 2400 4485
rect 2050 4415 2065 4435
rect 2085 4415 2100 4435
rect 2050 4400 2100 4415
rect 2350 4435 2400 4465
rect 2500 4835 3450 4850
rect 2500 4815 3415 4835
rect 3435 4815 3450 4835
rect 2500 4800 3450 4815
rect 2500 4785 2550 4800
rect 2500 4765 2515 4785
rect 2535 4765 2550 4785
rect 2500 4735 2550 4765
rect 2800 4785 2850 4800
rect 2800 4765 2815 4785
rect 2835 4765 2850 4785
rect 2500 4715 2515 4735
rect 2535 4715 2550 4735
rect 2500 4685 2550 4715
rect 2500 4665 2515 4685
rect 2535 4665 2550 4685
rect 2500 4635 2550 4665
rect 2500 4615 2515 4635
rect 2535 4615 2550 4635
rect 2500 4585 2550 4615
rect 2500 4565 2515 4585
rect 2535 4565 2550 4585
rect 2500 4535 2550 4565
rect 2500 4515 2515 4535
rect 2535 4515 2550 4535
rect 2500 4485 2550 4515
rect 2500 4465 2515 4485
rect 2535 4465 2550 4485
rect 2500 4450 2550 4465
rect 2650 4735 2700 4750
rect 2650 4715 2665 4735
rect 2685 4715 2700 4735
rect 2650 4685 2700 4715
rect 2650 4665 2665 4685
rect 2685 4665 2700 4685
rect 2650 4635 2700 4665
rect 2650 4615 2665 4635
rect 2685 4615 2700 4635
rect 2650 4585 2700 4615
rect 2650 4565 2665 4585
rect 2685 4565 2700 4585
rect 2650 4535 2700 4565
rect 2650 4515 2665 4535
rect 2685 4515 2700 4535
rect 2650 4485 2700 4515
rect 2650 4465 2665 4485
rect 2685 4465 2700 4485
rect 2350 4415 2365 4435
rect 2385 4415 2400 4435
rect 2350 4400 2400 4415
rect 2650 4435 2700 4465
rect 2800 4735 2850 4765
rect 3100 4785 3150 4800
rect 3100 4765 3115 4785
rect 3135 4765 3150 4785
rect 2800 4715 2815 4735
rect 2835 4715 2850 4735
rect 2800 4685 2850 4715
rect 2800 4665 2815 4685
rect 2835 4665 2850 4685
rect 2800 4635 2850 4665
rect 2800 4615 2815 4635
rect 2835 4615 2850 4635
rect 2800 4585 2850 4615
rect 2800 4565 2815 4585
rect 2835 4565 2850 4585
rect 2800 4535 2850 4565
rect 2800 4515 2815 4535
rect 2835 4515 2850 4535
rect 2800 4485 2850 4515
rect 2800 4465 2815 4485
rect 2835 4465 2850 4485
rect 2800 4450 2850 4465
rect 2950 4735 3000 4750
rect 2950 4715 2965 4735
rect 2985 4715 3000 4735
rect 2950 4685 3000 4715
rect 2950 4665 2965 4685
rect 2985 4665 3000 4685
rect 2950 4635 3000 4665
rect 2950 4615 2965 4635
rect 2985 4615 3000 4635
rect 2950 4585 3000 4615
rect 2950 4565 2965 4585
rect 2985 4565 3000 4585
rect 2950 4535 3000 4565
rect 2950 4515 2965 4535
rect 2985 4515 3000 4535
rect 2950 4485 3000 4515
rect 2950 4465 2965 4485
rect 2985 4465 3000 4485
rect 2650 4415 2665 4435
rect 2685 4415 2700 4435
rect 2650 4400 2700 4415
rect 2950 4435 3000 4465
rect 3100 4735 3150 4765
rect 3400 4785 3450 4800
rect 3400 4765 3415 4785
rect 3435 4765 3450 4785
rect 3100 4715 3115 4735
rect 3135 4715 3150 4735
rect 3100 4685 3150 4715
rect 3100 4665 3115 4685
rect 3135 4665 3150 4685
rect 3100 4635 3150 4665
rect 3100 4615 3115 4635
rect 3135 4615 3150 4635
rect 3100 4585 3150 4615
rect 3100 4565 3115 4585
rect 3135 4565 3150 4585
rect 3100 4535 3150 4565
rect 3100 4515 3115 4535
rect 3135 4515 3150 4535
rect 3100 4485 3150 4515
rect 3100 4465 3115 4485
rect 3135 4465 3150 4485
rect 3100 4450 3150 4465
rect 3250 4735 3300 4750
rect 3250 4715 3265 4735
rect 3285 4715 3300 4735
rect 3250 4685 3300 4715
rect 3250 4665 3265 4685
rect 3285 4665 3300 4685
rect 3250 4635 3300 4665
rect 3250 4615 3265 4635
rect 3285 4615 3300 4635
rect 3250 4585 3300 4615
rect 3250 4565 3265 4585
rect 3285 4565 3300 4585
rect 3250 4535 3300 4565
rect 3250 4515 3265 4535
rect 3285 4515 3300 4535
rect 3250 4485 3300 4515
rect 3250 4465 3265 4485
rect 3285 4465 3300 4485
rect 2950 4415 2965 4435
rect 2985 4415 3000 4435
rect 2950 4400 3000 4415
rect 3250 4435 3300 4465
rect 3400 4735 3450 4765
rect 3400 4715 3415 4735
rect 3435 4715 3450 4735
rect 3400 4685 3450 4715
rect 3400 4665 3415 4685
rect 3435 4665 3450 4685
rect 3400 4635 3450 4665
rect 3400 4615 3415 4635
rect 3435 4615 3450 4635
rect 3400 4585 3450 4615
rect 3400 4565 3415 4585
rect 3435 4565 3450 4585
rect 3400 4535 3450 4565
rect 3400 4515 3415 4535
rect 3435 4515 3450 4535
rect 3400 4485 3450 4515
rect 3400 4465 3415 4485
rect 3435 4465 3450 4485
rect 3400 4450 3450 4465
rect 3550 4835 3600 4850
rect 3550 4815 3565 4835
rect 3585 4815 3600 4835
rect 3550 4785 3600 4815
rect 3550 4765 3565 4785
rect 3585 4765 3600 4785
rect 3550 4735 3600 4765
rect 3550 4715 3565 4735
rect 3585 4715 3600 4735
rect 3550 4685 3600 4715
rect 3550 4665 3565 4685
rect 3585 4665 3600 4685
rect 3550 4635 3600 4665
rect 3550 4615 3565 4635
rect 3585 4615 3600 4635
rect 3550 4585 3600 4615
rect 3550 4565 3565 4585
rect 3585 4565 3600 4585
rect 3550 4535 3600 4565
rect 3550 4515 3565 4535
rect 3585 4515 3600 4535
rect 3550 4485 3600 4515
rect 3550 4465 3565 4485
rect 3585 4465 3600 4485
rect 3250 4415 3265 4435
rect 3285 4415 3300 4435
rect 3250 4400 3300 4415
rect 3550 4435 3600 4465
rect 3550 4415 3565 4435
rect 3585 4415 3600 4435
rect 3550 4400 3600 4415
rect 550 4385 3600 4400
rect 550 4365 565 4385
rect 585 4365 865 4385
rect 885 4365 1165 4385
rect 1185 4365 1465 4385
rect 1485 4365 1765 4385
rect 1785 4365 2065 4385
rect 2085 4365 2365 4385
rect 2385 4365 2665 4385
rect 2685 4365 2965 4385
rect 2985 4365 3265 4385
rect 3285 4365 3565 4385
rect 3585 4365 3600 4385
rect 550 4350 3600 4365
rect 4150 4840 4200 5115
rect 4750 5485 7800 5500
rect 4750 5465 4765 5485
rect 4785 5465 5065 5485
rect 5085 5465 5365 5485
rect 5385 5465 5665 5485
rect 5685 5465 5965 5485
rect 5985 5465 6265 5485
rect 6285 5465 6565 5485
rect 6585 5465 6865 5485
rect 6885 5465 7165 5485
rect 7185 5465 7465 5485
rect 7485 5465 7765 5485
rect 7785 5465 7800 5485
rect 4750 5450 7800 5465
rect 4750 5435 4800 5450
rect 4750 5415 4765 5435
rect 4785 5415 4800 5435
rect 4750 5385 4800 5415
rect 5050 5435 5100 5450
rect 5050 5415 5065 5435
rect 5085 5415 5100 5435
rect 4750 5365 4765 5385
rect 4785 5365 4800 5385
rect 4750 5335 4800 5365
rect 4750 5315 4765 5335
rect 4785 5315 4800 5335
rect 4750 5285 4800 5315
rect 4750 5265 4765 5285
rect 4785 5265 4800 5285
rect 4750 5235 4800 5265
rect 4750 5215 4765 5235
rect 4785 5215 4800 5235
rect 4750 5185 4800 5215
rect 4750 5165 4765 5185
rect 4785 5165 4800 5185
rect 4750 5135 4800 5165
rect 4750 5115 4765 5135
rect 4785 5115 4800 5135
rect 4750 5085 4800 5115
rect 4750 5065 4765 5085
rect 4785 5065 4800 5085
rect 4750 5035 4800 5065
rect 4750 5015 4765 5035
rect 4785 5015 4800 5035
rect 4750 5000 4800 5015
rect 4900 5385 4950 5400
rect 4900 5365 4915 5385
rect 4935 5365 4950 5385
rect 4900 5335 4950 5365
rect 4900 5315 4915 5335
rect 4935 5315 4950 5335
rect 4900 5285 4950 5315
rect 4900 5265 4915 5285
rect 4935 5265 4950 5285
rect 4900 5235 4950 5265
rect 4900 5215 4915 5235
rect 4935 5215 4950 5235
rect 4900 5185 4950 5215
rect 4900 5165 4915 5185
rect 4935 5165 4950 5185
rect 4900 5135 4950 5165
rect 4900 5115 4915 5135
rect 4935 5115 4950 5135
rect 4900 5085 4950 5115
rect 5050 5385 5100 5415
rect 5350 5435 5400 5450
rect 5350 5415 5365 5435
rect 5385 5415 5400 5435
rect 5050 5365 5065 5385
rect 5085 5365 5100 5385
rect 5050 5335 5100 5365
rect 5050 5315 5065 5335
rect 5085 5315 5100 5335
rect 5050 5285 5100 5315
rect 5050 5265 5065 5285
rect 5085 5265 5100 5285
rect 5050 5235 5100 5265
rect 5050 5215 5065 5235
rect 5085 5215 5100 5235
rect 5050 5185 5100 5215
rect 5050 5165 5065 5185
rect 5085 5165 5100 5185
rect 5050 5135 5100 5165
rect 5050 5115 5065 5135
rect 5085 5115 5100 5135
rect 5050 5100 5100 5115
rect 5200 5385 5250 5400
rect 5200 5365 5215 5385
rect 5235 5365 5250 5385
rect 5200 5335 5250 5365
rect 5200 5315 5215 5335
rect 5235 5315 5250 5335
rect 5200 5285 5250 5315
rect 5200 5265 5215 5285
rect 5235 5265 5250 5285
rect 5200 5235 5250 5265
rect 5200 5215 5215 5235
rect 5235 5215 5250 5235
rect 5200 5185 5250 5215
rect 5200 5165 5215 5185
rect 5235 5165 5250 5185
rect 5200 5135 5250 5165
rect 5200 5115 5215 5135
rect 5235 5115 5250 5135
rect 4900 5065 4915 5085
rect 4935 5065 4950 5085
rect 4900 5050 4950 5065
rect 5200 5085 5250 5115
rect 5350 5385 5400 5415
rect 5650 5435 5700 5450
rect 5650 5415 5665 5435
rect 5685 5415 5700 5435
rect 5350 5365 5365 5385
rect 5385 5365 5400 5385
rect 5350 5335 5400 5365
rect 5350 5315 5365 5335
rect 5385 5315 5400 5335
rect 5350 5285 5400 5315
rect 5350 5265 5365 5285
rect 5385 5265 5400 5285
rect 5350 5235 5400 5265
rect 5350 5215 5365 5235
rect 5385 5215 5400 5235
rect 5350 5185 5400 5215
rect 5350 5165 5365 5185
rect 5385 5165 5400 5185
rect 5350 5135 5400 5165
rect 5350 5115 5365 5135
rect 5385 5115 5400 5135
rect 5350 5100 5400 5115
rect 5500 5385 5550 5400
rect 5500 5365 5515 5385
rect 5535 5365 5550 5385
rect 5500 5335 5550 5365
rect 5500 5315 5515 5335
rect 5535 5315 5550 5335
rect 5500 5285 5550 5315
rect 5500 5265 5515 5285
rect 5535 5265 5550 5285
rect 5500 5235 5550 5265
rect 5500 5215 5515 5235
rect 5535 5215 5550 5235
rect 5500 5185 5550 5215
rect 5500 5165 5515 5185
rect 5535 5165 5550 5185
rect 5500 5135 5550 5165
rect 5500 5115 5515 5135
rect 5535 5115 5550 5135
rect 5200 5065 5215 5085
rect 5235 5065 5250 5085
rect 5200 5050 5250 5065
rect 5500 5085 5550 5115
rect 5650 5385 5700 5415
rect 5950 5435 6000 5450
rect 5950 5415 5965 5435
rect 5985 5415 6000 5435
rect 5650 5365 5665 5385
rect 5685 5365 5700 5385
rect 5650 5335 5700 5365
rect 5650 5315 5665 5335
rect 5685 5315 5700 5335
rect 5650 5285 5700 5315
rect 5650 5265 5665 5285
rect 5685 5265 5700 5285
rect 5650 5235 5700 5265
rect 5650 5215 5665 5235
rect 5685 5215 5700 5235
rect 5650 5185 5700 5215
rect 5650 5165 5665 5185
rect 5685 5165 5700 5185
rect 5650 5135 5700 5165
rect 5650 5115 5665 5135
rect 5685 5115 5700 5135
rect 5650 5100 5700 5115
rect 5800 5385 5850 5400
rect 5800 5365 5815 5385
rect 5835 5365 5850 5385
rect 5800 5335 5850 5365
rect 5800 5315 5815 5335
rect 5835 5315 5850 5335
rect 5800 5285 5850 5315
rect 5800 5265 5815 5285
rect 5835 5265 5850 5285
rect 5800 5235 5850 5265
rect 5800 5215 5815 5235
rect 5835 5215 5850 5235
rect 5800 5185 5850 5215
rect 5800 5165 5815 5185
rect 5835 5165 5850 5185
rect 5800 5135 5850 5165
rect 5800 5115 5815 5135
rect 5835 5115 5850 5135
rect 5500 5065 5515 5085
rect 5535 5065 5550 5085
rect 5500 5050 5550 5065
rect 5800 5085 5850 5115
rect 5800 5065 5815 5085
rect 5835 5065 5850 5085
rect 5800 5050 5850 5065
rect 4900 5035 5850 5050
rect 4900 5015 4915 5035
rect 4935 5015 5850 5035
rect 4900 5000 5850 5015
rect 5950 5385 6000 5415
rect 6250 5435 6300 5450
rect 6250 5415 6265 5435
rect 6285 5415 6300 5435
rect 5950 5365 5965 5385
rect 5985 5365 6000 5385
rect 5950 5335 6000 5365
rect 5950 5315 5965 5335
rect 5985 5315 6000 5335
rect 5950 5285 6000 5315
rect 5950 5265 5965 5285
rect 5985 5265 6000 5285
rect 5950 5235 6000 5265
rect 5950 5215 5965 5235
rect 5985 5215 6000 5235
rect 5950 5185 6000 5215
rect 5950 5165 5965 5185
rect 5985 5165 6000 5185
rect 5950 5135 6000 5165
rect 5950 5115 5965 5135
rect 5985 5115 6000 5135
rect 5950 5085 6000 5115
rect 5950 5065 5965 5085
rect 5985 5065 6000 5085
rect 5950 5035 6000 5065
rect 5950 5015 5965 5035
rect 5985 5015 6000 5035
rect 4300 4940 4350 4950
rect 4300 4910 4310 4940
rect 4340 4910 4350 4940
rect 4300 4900 4350 4910
rect 4600 4940 4650 4950
rect 4600 4910 4610 4940
rect 4640 4910 4650 4940
rect 4600 4900 4650 4910
rect 4900 4940 4950 4950
rect 4900 4910 4910 4940
rect 4940 4910 4950 4940
rect 4900 4900 4950 4910
rect 5200 4940 5250 4950
rect 5200 4910 5210 4940
rect 5240 4910 5250 4940
rect 5200 4900 5250 4910
rect 5350 4940 5400 4950
rect 5350 4910 5360 4940
rect 5390 4910 5400 4940
rect 5350 4900 5400 4910
rect 5500 4940 5550 4950
rect 5500 4910 5510 4940
rect 5540 4910 5550 4940
rect 5500 4900 5550 4910
rect 5800 4940 5850 4950
rect 5800 4910 5810 4940
rect 5840 4910 5850 4940
rect 5800 4900 5850 4910
rect 4150 4810 4160 4840
rect 4190 4810 4200 4840
rect 4150 4740 4200 4810
rect 4150 4710 4160 4740
rect 4190 4710 4200 4740
rect 4150 4685 4200 4710
rect 4150 4665 4165 4685
rect 4185 4665 4200 4685
rect 4150 4640 4200 4665
rect 4150 4610 4160 4640
rect 4190 4610 4200 4640
rect 4150 4585 4200 4610
rect 4150 4565 4165 4585
rect 4185 4565 4200 4585
rect 4150 4540 4200 4565
rect 4150 4510 4160 4540
rect 4190 4510 4200 4540
rect 4150 4485 4200 4510
rect 4150 4465 4165 4485
rect 4185 4465 4200 4485
rect 4150 4440 4200 4465
rect 4150 4410 4160 4440
rect 4190 4410 4200 4440
rect 4150 4385 4200 4410
rect 4150 4365 4165 4385
rect 4185 4365 4200 4385
rect -50 4260 -40 4290
rect -10 4260 0 4290
rect -650 4165 -635 4185
rect -615 4165 -600 4185
rect -650 4140 -600 4165
rect -650 4110 -640 4140
rect -610 4110 -600 4140
rect -650 4085 -600 4110
rect -650 4065 -635 4085
rect -615 4065 -600 4085
rect -650 4040 -600 4065
rect -650 4010 -640 4040
rect -610 4010 -600 4040
rect -650 3985 -600 4010
rect -650 3965 -635 3985
rect -615 3965 -600 3985
rect -650 3940 -600 3965
rect -650 3910 -640 3940
rect -610 3910 -600 3940
rect -650 3885 -600 3910
rect -650 3865 -635 3885
rect -615 3865 -600 3885
rect -650 3840 -600 3865
rect -650 3810 -640 3840
rect -610 3810 -600 3840
rect -650 3785 -600 3810
rect -650 3765 -635 3785
rect -615 3765 -600 3785
rect -650 3740 -600 3765
rect -650 3710 -640 3740
rect -610 3710 -600 3740
rect -650 3540 -600 3710
rect -500 4185 -450 4200
rect -500 4165 -485 4185
rect -465 4165 -450 4185
rect -500 4135 -450 4165
rect -500 4115 -485 4135
rect -465 4115 -450 4135
rect -500 4085 -450 4115
rect -500 4065 -485 4085
rect -465 4065 -450 4085
rect -500 4035 -450 4065
rect -500 4015 -485 4035
rect -465 4015 -450 4035
rect -500 3985 -450 4015
rect -500 3965 -485 3985
rect -465 3965 -450 3985
rect -500 3935 -450 3965
rect -500 3915 -485 3935
rect -465 3915 -450 3935
rect -500 3885 -450 3915
rect -500 3865 -485 3885
rect -465 3865 -450 3885
rect -500 3835 -450 3865
rect -500 3815 -485 3835
rect -465 3815 -450 3835
rect -500 3785 -450 3815
rect -350 4185 -300 4200
rect -350 4165 -335 4185
rect -315 4165 -300 4185
rect -350 4135 -300 4165
rect -350 4115 -335 4135
rect -315 4115 -300 4135
rect -350 4085 -300 4115
rect -350 4065 -335 4085
rect -315 4065 -300 4085
rect -350 4035 -300 4065
rect -350 4015 -335 4035
rect -315 4015 -300 4035
rect -350 3985 -300 4015
rect -350 3965 -335 3985
rect -315 3965 -300 3985
rect -350 3935 -300 3965
rect -350 3915 -335 3935
rect -315 3915 -300 3935
rect -350 3885 -300 3915
rect -350 3865 -335 3885
rect -315 3865 -300 3885
rect -350 3835 -300 3865
rect -350 3815 -335 3835
rect -315 3815 -300 3835
rect -350 3800 -300 3815
rect -200 4185 -150 4200
rect -200 4165 -185 4185
rect -165 4165 -150 4185
rect -200 4135 -150 4165
rect -200 4115 -185 4135
rect -165 4115 -150 4135
rect -200 4085 -150 4115
rect -200 4065 -185 4085
rect -165 4065 -150 4085
rect -200 4035 -150 4065
rect -200 4015 -185 4035
rect -165 4015 -150 4035
rect -200 3985 -150 4015
rect -200 3965 -185 3985
rect -165 3965 -150 3985
rect -200 3935 -150 3965
rect -200 3915 -185 3935
rect -165 3915 -150 3935
rect -200 3885 -150 3915
rect -200 3865 -185 3885
rect -165 3865 -150 3885
rect -200 3835 -150 3865
rect -200 3815 -185 3835
rect -165 3815 -150 3835
rect -500 3765 -485 3785
rect -465 3765 -450 3785
rect -500 3750 -450 3765
rect -200 3785 -150 3815
rect -200 3765 -185 3785
rect -165 3765 -150 3785
rect -200 3750 -150 3765
rect -500 3735 -150 3750
rect -500 3715 -485 3735
rect -465 3715 -185 3735
rect -165 3715 -150 3735
rect -500 3700 -150 3715
rect -50 4185 0 4260
rect 4150 4290 4200 4365
rect 4750 4835 4800 4850
rect 4750 4815 4765 4835
rect 4785 4815 4800 4835
rect 4750 4785 4800 4815
rect 4750 4765 4765 4785
rect 4785 4765 4800 4785
rect 4750 4735 4800 4765
rect 4750 4715 4765 4735
rect 4785 4715 4800 4735
rect 4750 4685 4800 4715
rect 4750 4665 4765 4685
rect 4785 4665 4800 4685
rect 4750 4635 4800 4665
rect 4750 4615 4765 4635
rect 4785 4615 4800 4635
rect 4750 4585 4800 4615
rect 4750 4565 4765 4585
rect 4785 4565 4800 4585
rect 4750 4535 4800 4565
rect 4750 4515 4765 4535
rect 4785 4515 4800 4535
rect 4750 4485 4800 4515
rect 4750 4465 4765 4485
rect 4785 4465 4800 4485
rect 4750 4435 4800 4465
rect 4900 4835 5850 4850
rect 4900 4815 4915 4835
rect 4935 4815 5850 4835
rect 4900 4800 5850 4815
rect 4900 4785 4950 4800
rect 4900 4765 4915 4785
rect 4935 4765 4950 4785
rect 4900 4735 4950 4765
rect 5200 4785 5250 4800
rect 5200 4765 5215 4785
rect 5235 4765 5250 4785
rect 4900 4715 4915 4735
rect 4935 4715 4950 4735
rect 4900 4685 4950 4715
rect 4900 4665 4915 4685
rect 4935 4665 4950 4685
rect 4900 4635 4950 4665
rect 4900 4615 4915 4635
rect 4935 4615 4950 4635
rect 4900 4585 4950 4615
rect 4900 4565 4915 4585
rect 4935 4565 4950 4585
rect 4900 4535 4950 4565
rect 4900 4515 4915 4535
rect 4935 4515 4950 4535
rect 4900 4485 4950 4515
rect 4900 4465 4915 4485
rect 4935 4465 4950 4485
rect 4900 4450 4950 4465
rect 5050 4735 5100 4750
rect 5050 4715 5065 4735
rect 5085 4715 5100 4735
rect 5050 4685 5100 4715
rect 5050 4665 5065 4685
rect 5085 4665 5100 4685
rect 5050 4635 5100 4665
rect 5050 4615 5065 4635
rect 5085 4615 5100 4635
rect 5050 4585 5100 4615
rect 5050 4565 5065 4585
rect 5085 4565 5100 4585
rect 5050 4535 5100 4565
rect 5050 4515 5065 4535
rect 5085 4515 5100 4535
rect 5050 4485 5100 4515
rect 5050 4465 5065 4485
rect 5085 4465 5100 4485
rect 4750 4415 4765 4435
rect 4785 4415 4800 4435
rect 4750 4400 4800 4415
rect 5050 4435 5100 4465
rect 5200 4735 5250 4765
rect 5500 4785 5550 4800
rect 5500 4765 5515 4785
rect 5535 4765 5550 4785
rect 5200 4715 5215 4735
rect 5235 4715 5250 4735
rect 5200 4685 5250 4715
rect 5200 4665 5215 4685
rect 5235 4665 5250 4685
rect 5200 4635 5250 4665
rect 5200 4615 5215 4635
rect 5235 4615 5250 4635
rect 5200 4585 5250 4615
rect 5200 4565 5215 4585
rect 5235 4565 5250 4585
rect 5200 4535 5250 4565
rect 5200 4515 5215 4535
rect 5235 4515 5250 4535
rect 5200 4485 5250 4515
rect 5200 4465 5215 4485
rect 5235 4465 5250 4485
rect 5200 4450 5250 4465
rect 5350 4735 5400 4750
rect 5350 4715 5365 4735
rect 5385 4715 5400 4735
rect 5350 4685 5400 4715
rect 5350 4665 5365 4685
rect 5385 4665 5400 4685
rect 5350 4635 5400 4665
rect 5350 4615 5365 4635
rect 5385 4615 5400 4635
rect 5350 4585 5400 4615
rect 5350 4565 5365 4585
rect 5385 4565 5400 4585
rect 5350 4535 5400 4565
rect 5350 4515 5365 4535
rect 5385 4515 5400 4535
rect 5350 4485 5400 4515
rect 5350 4465 5365 4485
rect 5385 4465 5400 4485
rect 5050 4415 5065 4435
rect 5085 4415 5100 4435
rect 5050 4400 5100 4415
rect 5350 4435 5400 4465
rect 5500 4735 5550 4765
rect 5800 4785 5850 4800
rect 5800 4765 5815 4785
rect 5835 4765 5850 4785
rect 5500 4715 5515 4735
rect 5535 4715 5550 4735
rect 5500 4685 5550 4715
rect 5500 4665 5515 4685
rect 5535 4665 5550 4685
rect 5500 4635 5550 4665
rect 5500 4615 5515 4635
rect 5535 4615 5550 4635
rect 5500 4585 5550 4615
rect 5500 4565 5515 4585
rect 5535 4565 5550 4585
rect 5500 4535 5550 4565
rect 5500 4515 5515 4535
rect 5535 4515 5550 4535
rect 5500 4485 5550 4515
rect 5500 4465 5515 4485
rect 5535 4465 5550 4485
rect 5500 4450 5550 4465
rect 5650 4735 5700 4750
rect 5650 4715 5665 4735
rect 5685 4715 5700 4735
rect 5650 4685 5700 4715
rect 5650 4665 5665 4685
rect 5685 4665 5700 4685
rect 5650 4635 5700 4665
rect 5650 4615 5665 4635
rect 5685 4615 5700 4635
rect 5650 4585 5700 4615
rect 5650 4565 5665 4585
rect 5685 4565 5700 4585
rect 5650 4535 5700 4565
rect 5650 4515 5665 4535
rect 5685 4515 5700 4535
rect 5650 4485 5700 4515
rect 5650 4465 5665 4485
rect 5685 4465 5700 4485
rect 5350 4415 5365 4435
rect 5385 4415 5400 4435
rect 5350 4400 5400 4415
rect 5650 4435 5700 4465
rect 5800 4735 5850 4765
rect 5800 4715 5815 4735
rect 5835 4715 5850 4735
rect 5800 4685 5850 4715
rect 5800 4665 5815 4685
rect 5835 4665 5850 4685
rect 5800 4635 5850 4665
rect 5800 4615 5815 4635
rect 5835 4615 5850 4635
rect 5800 4585 5850 4615
rect 5800 4565 5815 4585
rect 5835 4565 5850 4585
rect 5800 4535 5850 4565
rect 5800 4515 5815 4535
rect 5835 4515 5850 4535
rect 5800 4485 5850 4515
rect 5800 4465 5815 4485
rect 5835 4465 5850 4485
rect 5800 4450 5850 4465
rect 5950 4835 6000 5015
rect 6100 5385 6150 5400
rect 6100 5365 6115 5385
rect 6135 5365 6150 5385
rect 6100 5335 6150 5365
rect 6100 5315 6115 5335
rect 6135 5315 6150 5335
rect 6100 5285 6150 5315
rect 6100 5265 6115 5285
rect 6135 5265 6150 5285
rect 6100 5235 6150 5265
rect 6100 5215 6115 5235
rect 6135 5215 6150 5235
rect 6100 5185 6150 5215
rect 6100 5165 6115 5185
rect 6135 5165 6150 5185
rect 6100 5135 6150 5165
rect 6100 5115 6115 5135
rect 6135 5115 6150 5135
rect 6100 5085 6150 5115
rect 6250 5385 6300 5415
rect 6550 5435 6600 5450
rect 6550 5415 6565 5435
rect 6585 5415 6600 5435
rect 6250 5365 6265 5385
rect 6285 5365 6300 5385
rect 6250 5335 6300 5365
rect 6250 5315 6265 5335
rect 6285 5315 6300 5335
rect 6250 5285 6300 5315
rect 6250 5265 6265 5285
rect 6285 5265 6300 5285
rect 6250 5235 6300 5265
rect 6250 5215 6265 5235
rect 6285 5215 6300 5235
rect 6250 5185 6300 5215
rect 6250 5165 6265 5185
rect 6285 5165 6300 5185
rect 6250 5135 6300 5165
rect 6250 5115 6265 5135
rect 6285 5115 6300 5135
rect 6250 5100 6300 5115
rect 6400 5385 6450 5400
rect 6400 5365 6415 5385
rect 6435 5365 6450 5385
rect 6400 5335 6450 5365
rect 6400 5315 6415 5335
rect 6435 5315 6450 5335
rect 6400 5285 6450 5315
rect 6400 5265 6415 5285
rect 6435 5265 6450 5285
rect 6400 5235 6450 5265
rect 6400 5215 6415 5235
rect 6435 5215 6450 5235
rect 6400 5185 6450 5215
rect 6400 5165 6415 5185
rect 6435 5165 6450 5185
rect 6400 5135 6450 5165
rect 6400 5115 6415 5135
rect 6435 5115 6450 5135
rect 6100 5065 6115 5085
rect 6135 5065 6150 5085
rect 6100 5050 6150 5065
rect 6400 5085 6450 5115
rect 6400 5065 6415 5085
rect 6435 5065 6450 5085
rect 6400 5050 6450 5065
rect 6100 5035 6450 5050
rect 6100 5015 6115 5035
rect 6135 5015 6415 5035
rect 6435 5015 6450 5035
rect 6100 5000 6450 5015
rect 6550 5385 6600 5415
rect 6850 5435 6900 5450
rect 6850 5415 6865 5435
rect 6885 5415 6900 5435
rect 6550 5365 6565 5385
rect 6585 5365 6600 5385
rect 6550 5335 6600 5365
rect 6550 5315 6565 5335
rect 6585 5315 6600 5335
rect 6550 5285 6600 5315
rect 6550 5265 6565 5285
rect 6585 5265 6600 5285
rect 6550 5235 6600 5265
rect 6550 5215 6565 5235
rect 6585 5215 6600 5235
rect 6550 5185 6600 5215
rect 6550 5165 6565 5185
rect 6585 5165 6600 5185
rect 6550 5135 6600 5165
rect 6550 5115 6565 5135
rect 6585 5115 6600 5135
rect 6550 5085 6600 5115
rect 6550 5065 6565 5085
rect 6585 5065 6600 5085
rect 6550 5035 6600 5065
rect 6550 5015 6565 5035
rect 6585 5015 6600 5035
rect 6100 4940 6150 4950
rect 6100 4910 6110 4940
rect 6140 4910 6150 4940
rect 6100 4900 6150 4910
rect 6250 4940 6300 5000
rect 6250 4910 6260 4940
rect 6290 4910 6300 4940
rect 6250 4850 6300 4910
rect 6400 4940 6450 4950
rect 6400 4910 6410 4940
rect 6440 4910 6450 4940
rect 6400 4900 6450 4910
rect 5950 4815 5965 4835
rect 5985 4815 6000 4835
rect 5950 4785 6000 4815
rect 5950 4765 5965 4785
rect 5985 4765 6000 4785
rect 5950 4735 6000 4765
rect 5950 4715 5965 4735
rect 5985 4715 6000 4735
rect 5950 4685 6000 4715
rect 5950 4665 5965 4685
rect 5985 4665 6000 4685
rect 5950 4635 6000 4665
rect 5950 4615 5965 4635
rect 5985 4615 6000 4635
rect 5950 4585 6000 4615
rect 5950 4565 5965 4585
rect 5985 4565 6000 4585
rect 5950 4535 6000 4565
rect 5950 4515 5965 4535
rect 5985 4515 6000 4535
rect 5950 4485 6000 4515
rect 5950 4465 5965 4485
rect 5985 4465 6000 4485
rect 5650 4415 5665 4435
rect 5685 4415 5700 4435
rect 5650 4400 5700 4415
rect 5950 4435 6000 4465
rect 6100 4835 6450 4850
rect 6100 4815 6115 4835
rect 6135 4815 6415 4835
rect 6435 4815 6450 4835
rect 6100 4800 6450 4815
rect 6100 4785 6150 4800
rect 6100 4765 6115 4785
rect 6135 4765 6150 4785
rect 6100 4735 6150 4765
rect 6400 4785 6450 4800
rect 6400 4765 6415 4785
rect 6435 4765 6450 4785
rect 6100 4715 6115 4735
rect 6135 4715 6150 4735
rect 6100 4685 6150 4715
rect 6100 4665 6115 4685
rect 6135 4665 6150 4685
rect 6100 4635 6150 4665
rect 6100 4615 6115 4635
rect 6135 4615 6150 4635
rect 6100 4585 6150 4615
rect 6100 4565 6115 4585
rect 6135 4565 6150 4585
rect 6100 4535 6150 4565
rect 6100 4515 6115 4535
rect 6135 4515 6150 4535
rect 6100 4485 6150 4515
rect 6100 4465 6115 4485
rect 6135 4465 6150 4485
rect 6100 4450 6150 4465
rect 6250 4735 6300 4750
rect 6250 4715 6265 4735
rect 6285 4715 6300 4735
rect 6250 4685 6300 4715
rect 6250 4665 6265 4685
rect 6285 4665 6300 4685
rect 6250 4635 6300 4665
rect 6250 4615 6265 4635
rect 6285 4615 6300 4635
rect 6250 4585 6300 4615
rect 6250 4565 6265 4585
rect 6285 4565 6300 4585
rect 6250 4535 6300 4565
rect 6250 4515 6265 4535
rect 6285 4515 6300 4535
rect 6250 4485 6300 4515
rect 6250 4465 6265 4485
rect 6285 4465 6300 4485
rect 5950 4415 5965 4435
rect 5985 4415 6000 4435
rect 5950 4400 6000 4415
rect 6250 4435 6300 4465
rect 6400 4735 6450 4765
rect 6400 4715 6415 4735
rect 6435 4715 6450 4735
rect 6400 4685 6450 4715
rect 6400 4665 6415 4685
rect 6435 4665 6450 4685
rect 6400 4635 6450 4665
rect 6400 4615 6415 4635
rect 6435 4615 6450 4635
rect 6400 4585 6450 4615
rect 6400 4565 6415 4585
rect 6435 4565 6450 4585
rect 6400 4535 6450 4565
rect 6400 4515 6415 4535
rect 6435 4515 6450 4535
rect 6400 4485 6450 4515
rect 6400 4465 6415 4485
rect 6435 4465 6450 4485
rect 6400 4450 6450 4465
rect 6550 4835 6600 5015
rect 6700 5385 6750 5400
rect 6700 5365 6715 5385
rect 6735 5365 6750 5385
rect 6700 5335 6750 5365
rect 6700 5315 6715 5335
rect 6735 5315 6750 5335
rect 6700 5285 6750 5315
rect 6700 5265 6715 5285
rect 6735 5265 6750 5285
rect 6700 5235 6750 5265
rect 6700 5215 6715 5235
rect 6735 5215 6750 5235
rect 6700 5185 6750 5215
rect 6700 5165 6715 5185
rect 6735 5165 6750 5185
rect 6700 5135 6750 5165
rect 6700 5115 6715 5135
rect 6735 5115 6750 5135
rect 6700 5085 6750 5115
rect 6850 5385 6900 5415
rect 7150 5435 7200 5450
rect 7150 5415 7165 5435
rect 7185 5415 7200 5435
rect 6850 5365 6865 5385
rect 6885 5365 6900 5385
rect 6850 5335 6900 5365
rect 6850 5315 6865 5335
rect 6885 5315 6900 5335
rect 6850 5285 6900 5315
rect 6850 5265 6865 5285
rect 6885 5265 6900 5285
rect 6850 5235 6900 5265
rect 6850 5215 6865 5235
rect 6885 5215 6900 5235
rect 6850 5185 6900 5215
rect 6850 5165 6865 5185
rect 6885 5165 6900 5185
rect 6850 5135 6900 5165
rect 6850 5115 6865 5135
rect 6885 5115 6900 5135
rect 6850 5100 6900 5115
rect 7000 5385 7050 5400
rect 7000 5365 7015 5385
rect 7035 5365 7050 5385
rect 7000 5335 7050 5365
rect 7000 5315 7015 5335
rect 7035 5315 7050 5335
rect 7000 5285 7050 5315
rect 7000 5265 7015 5285
rect 7035 5265 7050 5285
rect 7000 5235 7050 5265
rect 7000 5215 7015 5235
rect 7035 5215 7050 5235
rect 7000 5185 7050 5215
rect 7000 5165 7015 5185
rect 7035 5165 7050 5185
rect 7000 5135 7050 5165
rect 7000 5115 7015 5135
rect 7035 5115 7050 5135
rect 6700 5065 6715 5085
rect 6735 5065 6750 5085
rect 6700 5050 6750 5065
rect 7000 5085 7050 5115
rect 7150 5385 7200 5415
rect 7450 5435 7500 5450
rect 7450 5415 7465 5435
rect 7485 5415 7500 5435
rect 7150 5365 7165 5385
rect 7185 5365 7200 5385
rect 7150 5335 7200 5365
rect 7150 5315 7165 5335
rect 7185 5315 7200 5335
rect 7150 5285 7200 5315
rect 7150 5265 7165 5285
rect 7185 5265 7200 5285
rect 7150 5235 7200 5265
rect 7150 5215 7165 5235
rect 7185 5215 7200 5235
rect 7150 5185 7200 5215
rect 7150 5165 7165 5185
rect 7185 5165 7200 5185
rect 7150 5135 7200 5165
rect 7150 5115 7165 5135
rect 7185 5115 7200 5135
rect 7150 5100 7200 5115
rect 7300 5385 7350 5400
rect 7300 5365 7315 5385
rect 7335 5365 7350 5385
rect 7300 5335 7350 5365
rect 7300 5315 7315 5335
rect 7335 5315 7350 5335
rect 7300 5285 7350 5315
rect 7300 5265 7315 5285
rect 7335 5265 7350 5285
rect 7300 5235 7350 5265
rect 7300 5215 7315 5235
rect 7335 5215 7350 5235
rect 7300 5185 7350 5215
rect 7300 5165 7315 5185
rect 7335 5165 7350 5185
rect 7300 5135 7350 5165
rect 7300 5115 7315 5135
rect 7335 5115 7350 5135
rect 7000 5065 7015 5085
rect 7035 5065 7050 5085
rect 7000 5050 7050 5065
rect 7300 5085 7350 5115
rect 7450 5385 7500 5415
rect 7750 5435 7800 5450
rect 7750 5415 7765 5435
rect 7785 5415 7800 5435
rect 7450 5365 7465 5385
rect 7485 5365 7500 5385
rect 7450 5335 7500 5365
rect 7450 5315 7465 5335
rect 7485 5315 7500 5335
rect 7450 5285 7500 5315
rect 7450 5265 7465 5285
rect 7485 5265 7500 5285
rect 7450 5235 7500 5265
rect 7450 5215 7465 5235
rect 7485 5215 7500 5235
rect 7450 5185 7500 5215
rect 7450 5165 7465 5185
rect 7485 5165 7500 5185
rect 7450 5135 7500 5165
rect 7450 5115 7465 5135
rect 7485 5115 7500 5135
rect 7450 5100 7500 5115
rect 7600 5385 7650 5400
rect 7600 5365 7615 5385
rect 7635 5365 7650 5385
rect 7600 5335 7650 5365
rect 7600 5315 7615 5335
rect 7635 5315 7650 5335
rect 7600 5285 7650 5315
rect 7600 5265 7615 5285
rect 7635 5265 7650 5285
rect 7600 5235 7650 5265
rect 7600 5215 7615 5235
rect 7635 5215 7650 5235
rect 7600 5185 7650 5215
rect 7600 5165 7615 5185
rect 7635 5165 7650 5185
rect 7600 5135 7650 5165
rect 7600 5115 7615 5135
rect 7635 5115 7650 5135
rect 7300 5065 7315 5085
rect 7335 5065 7350 5085
rect 7300 5050 7350 5065
rect 7600 5085 7650 5115
rect 7600 5065 7615 5085
rect 7635 5065 7650 5085
rect 7600 5050 7650 5065
rect 6700 5035 7650 5050
rect 6700 5015 7615 5035
rect 7635 5015 7650 5035
rect 6700 5000 7650 5015
rect 7750 5385 7800 5415
rect 7750 5365 7765 5385
rect 7785 5365 7800 5385
rect 7750 5335 7800 5365
rect 7750 5315 7765 5335
rect 7785 5315 7800 5335
rect 7750 5285 7800 5315
rect 7750 5265 7765 5285
rect 7785 5265 7800 5285
rect 7750 5235 7800 5265
rect 7750 5215 7765 5235
rect 7785 5215 7800 5235
rect 7750 5185 7800 5215
rect 7750 5165 7765 5185
rect 7785 5165 7800 5185
rect 7750 5135 7800 5165
rect 7750 5115 7765 5135
rect 7785 5115 7800 5135
rect 7750 5085 7800 5115
rect 7750 5065 7765 5085
rect 7785 5065 7800 5085
rect 7750 5035 7800 5065
rect 7750 5015 7765 5035
rect 7785 5015 7800 5035
rect 7750 5000 7800 5015
rect 8350 5485 8400 5560
rect 8650 5590 8700 5600
rect 8650 5560 8660 5590
rect 8690 5560 8700 5590
rect 8350 5465 8365 5485
rect 8385 5465 8400 5485
rect 8350 5440 8400 5465
rect 8350 5410 8360 5440
rect 8390 5410 8400 5440
rect 8350 5385 8400 5410
rect 8350 5365 8365 5385
rect 8385 5365 8400 5385
rect 8350 5340 8400 5365
rect 8350 5310 8360 5340
rect 8390 5310 8400 5340
rect 8350 5285 8400 5310
rect 8350 5265 8365 5285
rect 8385 5265 8400 5285
rect 8350 5240 8400 5265
rect 8350 5210 8360 5240
rect 8390 5210 8400 5240
rect 8350 5185 8400 5210
rect 8350 5165 8365 5185
rect 8385 5165 8400 5185
rect 8350 5140 8400 5165
rect 8350 5110 8360 5140
rect 8390 5110 8400 5140
rect 8350 5085 8400 5110
rect 8350 5065 8365 5085
rect 8385 5065 8400 5085
rect 8350 5040 8400 5065
rect 8350 5010 8360 5040
rect 8390 5010 8400 5040
rect 6700 4940 6750 4950
rect 6700 4910 6710 4940
rect 6740 4910 6750 4940
rect 6700 4900 6750 4910
rect 7000 4940 7050 4950
rect 7000 4910 7010 4940
rect 7040 4910 7050 4940
rect 7000 4900 7050 4910
rect 7150 4940 7200 4950
rect 7150 4910 7160 4940
rect 7190 4910 7200 4940
rect 7150 4900 7200 4910
rect 7300 4940 7350 4950
rect 7300 4910 7310 4940
rect 7340 4910 7350 4940
rect 7300 4900 7350 4910
rect 7600 4940 7650 4950
rect 7600 4910 7610 4940
rect 7640 4910 7650 4940
rect 7600 4900 7650 4910
rect 7900 4940 7950 4950
rect 7900 4910 7910 4940
rect 7940 4910 7950 4940
rect 7900 4900 7950 4910
rect 8200 4940 8250 4950
rect 8200 4910 8210 4940
rect 8240 4910 8250 4940
rect 8200 4900 8250 4910
rect 6550 4815 6565 4835
rect 6585 4815 6600 4835
rect 6550 4785 6600 4815
rect 6550 4765 6565 4785
rect 6585 4765 6600 4785
rect 6550 4735 6600 4765
rect 6550 4715 6565 4735
rect 6585 4715 6600 4735
rect 6550 4685 6600 4715
rect 6550 4665 6565 4685
rect 6585 4665 6600 4685
rect 6550 4635 6600 4665
rect 6550 4615 6565 4635
rect 6585 4615 6600 4635
rect 6550 4585 6600 4615
rect 6550 4565 6565 4585
rect 6585 4565 6600 4585
rect 6550 4535 6600 4565
rect 6550 4515 6565 4535
rect 6585 4515 6600 4535
rect 6550 4485 6600 4515
rect 6550 4465 6565 4485
rect 6585 4465 6600 4485
rect 6250 4415 6265 4435
rect 6285 4415 6300 4435
rect 6250 4400 6300 4415
rect 6550 4435 6600 4465
rect 6700 4835 7650 4850
rect 6700 4815 7615 4835
rect 7635 4815 7650 4835
rect 6700 4800 7650 4815
rect 6700 4785 6750 4800
rect 6700 4765 6715 4785
rect 6735 4765 6750 4785
rect 6700 4735 6750 4765
rect 7000 4785 7050 4800
rect 7000 4765 7015 4785
rect 7035 4765 7050 4785
rect 6700 4715 6715 4735
rect 6735 4715 6750 4735
rect 6700 4685 6750 4715
rect 6700 4665 6715 4685
rect 6735 4665 6750 4685
rect 6700 4635 6750 4665
rect 6700 4615 6715 4635
rect 6735 4615 6750 4635
rect 6700 4585 6750 4615
rect 6700 4565 6715 4585
rect 6735 4565 6750 4585
rect 6700 4535 6750 4565
rect 6700 4515 6715 4535
rect 6735 4515 6750 4535
rect 6700 4485 6750 4515
rect 6700 4465 6715 4485
rect 6735 4465 6750 4485
rect 6700 4450 6750 4465
rect 6850 4735 6900 4750
rect 6850 4715 6865 4735
rect 6885 4715 6900 4735
rect 6850 4685 6900 4715
rect 6850 4665 6865 4685
rect 6885 4665 6900 4685
rect 6850 4635 6900 4665
rect 6850 4615 6865 4635
rect 6885 4615 6900 4635
rect 6850 4585 6900 4615
rect 6850 4565 6865 4585
rect 6885 4565 6900 4585
rect 6850 4535 6900 4565
rect 6850 4515 6865 4535
rect 6885 4515 6900 4535
rect 6850 4485 6900 4515
rect 6850 4465 6865 4485
rect 6885 4465 6900 4485
rect 6550 4415 6565 4435
rect 6585 4415 6600 4435
rect 6550 4400 6600 4415
rect 6850 4435 6900 4465
rect 7000 4735 7050 4765
rect 7300 4785 7350 4800
rect 7300 4765 7315 4785
rect 7335 4765 7350 4785
rect 7000 4715 7015 4735
rect 7035 4715 7050 4735
rect 7000 4685 7050 4715
rect 7000 4665 7015 4685
rect 7035 4665 7050 4685
rect 7000 4635 7050 4665
rect 7000 4615 7015 4635
rect 7035 4615 7050 4635
rect 7000 4585 7050 4615
rect 7000 4565 7015 4585
rect 7035 4565 7050 4585
rect 7000 4535 7050 4565
rect 7000 4515 7015 4535
rect 7035 4515 7050 4535
rect 7000 4485 7050 4515
rect 7000 4465 7015 4485
rect 7035 4465 7050 4485
rect 7000 4450 7050 4465
rect 7150 4735 7200 4750
rect 7150 4715 7165 4735
rect 7185 4715 7200 4735
rect 7150 4685 7200 4715
rect 7150 4665 7165 4685
rect 7185 4665 7200 4685
rect 7150 4635 7200 4665
rect 7150 4615 7165 4635
rect 7185 4615 7200 4635
rect 7150 4585 7200 4615
rect 7150 4565 7165 4585
rect 7185 4565 7200 4585
rect 7150 4535 7200 4565
rect 7150 4515 7165 4535
rect 7185 4515 7200 4535
rect 7150 4485 7200 4515
rect 7150 4465 7165 4485
rect 7185 4465 7200 4485
rect 6850 4415 6865 4435
rect 6885 4415 6900 4435
rect 6850 4400 6900 4415
rect 7150 4435 7200 4465
rect 7300 4735 7350 4765
rect 7600 4785 7650 4800
rect 7600 4765 7615 4785
rect 7635 4765 7650 4785
rect 7300 4715 7315 4735
rect 7335 4715 7350 4735
rect 7300 4685 7350 4715
rect 7300 4665 7315 4685
rect 7335 4665 7350 4685
rect 7300 4635 7350 4665
rect 7300 4615 7315 4635
rect 7335 4615 7350 4635
rect 7300 4585 7350 4615
rect 7300 4565 7315 4585
rect 7335 4565 7350 4585
rect 7300 4535 7350 4565
rect 7300 4515 7315 4535
rect 7335 4515 7350 4535
rect 7300 4485 7350 4515
rect 7300 4465 7315 4485
rect 7335 4465 7350 4485
rect 7300 4450 7350 4465
rect 7450 4735 7500 4750
rect 7450 4715 7465 4735
rect 7485 4715 7500 4735
rect 7450 4685 7500 4715
rect 7450 4665 7465 4685
rect 7485 4665 7500 4685
rect 7450 4635 7500 4665
rect 7450 4615 7465 4635
rect 7485 4615 7500 4635
rect 7450 4585 7500 4615
rect 7450 4565 7465 4585
rect 7485 4565 7500 4585
rect 7450 4535 7500 4565
rect 7450 4515 7465 4535
rect 7485 4515 7500 4535
rect 7450 4485 7500 4515
rect 7450 4465 7465 4485
rect 7485 4465 7500 4485
rect 7150 4415 7165 4435
rect 7185 4415 7200 4435
rect 7150 4400 7200 4415
rect 7450 4435 7500 4465
rect 7600 4735 7650 4765
rect 7600 4715 7615 4735
rect 7635 4715 7650 4735
rect 7600 4685 7650 4715
rect 7600 4665 7615 4685
rect 7635 4665 7650 4685
rect 7600 4635 7650 4665
rect 7600 4615 7615 4635
rect 7635 4615 7650 4635
rect 7600 4585 7650 4615
rect 7600 4565 7615 4585
rect 7635 4565 7650 4585
rect 7600 4535 7650 4565
rect 7600 4515 7615 4535
rect 7635 4515 7650 4535
rect 7600 4485 7650 4515
rect 7600 4465 7615 4485
rect 7635 4465 7650 4485
rect 7600 4450 7650 4465
rect 7750 4835 7800 4850
rect 7750 4815 7765 4835
rect 7785 4815 7800 4835
rect 7750 4785 7800 4815
rect 7750 4765 7765 4785
rect 7785 4765 7800 4785
rect 7750 4735 7800 4765
rect 7750 4715 7765 4735
rect 7785 4715 7800 4735
rect 7750 4685 7800 4715
rect 7750 4665 7765 4685
rect 7785 4665 7800 4685
rect 7750 4635 7800 4665
rect 7750 4615 7765 4635
rect 7785 4615 7800 4635
rect 7750 4585 7800 4615
rect 7750 4565 7765 4585
rect 7785 4565 7800 4585
rect 7750 4535 7800 4565
rect 7750 4515 7765 4535
rect 7785 4515 7800 4535
rect 7750 4485 7800 4515
rect 7750 4465 7765 4485
rect 7785 4465 7800 4485
rect 7450 4415 7465 4435
rect 7485 4415 7500 4435
rect 7450 4400 7500 4415
rect 7750 4435 7800 4465
rect 7750 4415 7765 4435
rect 7785 4415 7800 4435
rect 7750 4400 7800 4415
rect 4750 4385 7800 4400
rect 4750 4365 4765 4385
rect 4785 4365 5065 4385
rect 5085 4365 5365 4385
rect 5385 4365 5665 4385
rect 5685 4365 5965 4385
rect 5985 4365 6265 4385
rect 6285 4365 6565 4385
rect 6585 4365 6865 4385
rect 6885 4365 7165 4385
rect 7185 4365 7465 4385
rect 7485 4365 7765 4385
rect 7785 4365 7800 4385
rect 4750 4350 7800 4365
rect 8350 4840 8400 5010
rect 8500 5485 8550 5500
rect 8500 5465 8515 5485
rect 8535 5465 8550 5485
rect 8500 5435 8550 5465
rect 8500 5415 8515 5435
rect 8535 5415 8550 5435
rect 8500 5385 8550 5415
rect 8500 5365 8515 5385
rect 8535 5365 8550 5385
rect 8500 5335 8550 5365
rect 8500 5315 8515 5335
rect 8535 5315 8550 5335
rect 8500 5285 8550 5315
rect 8500 5265 8515 5285
rect 8535 5265 8550 5285
rect 8500 5235 8550 5265
rect 8500 5215 8515 5235
rect 8535 5215 8550 5235
rect 8500 5185 8550 5215
rect 8500 5165 8515 5185
rect 8535 5165 8550 5185
rect 8500 5135 8550 5165
rect 8500 5115 8515 5135
rect 8535 5115 8550 5135
rect 8500 5085 8550 5115
rect 8500 5065 8515 5085
rect 8535 5065 8550 5085
rect 8500 5035 8550 5065
rect 8500 5015 8515 5035
rect 8535 5015 8550 5035
rect 8500 5000 8550 5015
rect 8650 5485 8700 5560
rect 8950 5590 9000 5600
rect 8950 5560 8960 5590
rect 8990 5560 9000 5590
rect 8650 5465 8665 5485
rect 8685 5465 8700 5485
rect 8650 5440 8700 5465
rect 8650 5410 8660 5440
rect 8690 5410 8700 5440
rect 8650 5385 8700 5410
rect 8650 5365 8665 5385
rect 8685 5365 8700 5385
rect 8650 5340 8700 5365
rect 8650 5310 8660 5340
rect 8690 5310 8700 5340
rect 8650 5285 8700 5310
rect 8650 5265 8665 5285
rect 8685 5265 8700 5285
rect 8650 5240 8700 5265
rect 8650 5210 8660 5240
rect 8690 5210 8700 5240
rect 8650 5185 8700 5210
rect 8650 5165 8665 5185
rect 8685 5165 8700 5185
rect 8650 5140 8700 5165
rect 8650 5110 8660 5140
rect 8690 5110 8700 5140
rect 8650 5085 8700 5110
rect 8650 5065 8665 5085
rect 8685 5065 8700 5085
rect 8650 5040 8700 5065
rect 8650 5010 8660 5040
rect 8690 5010 8700 5040
rect 8500 4940 8550 4950
rect 8500 4910 8510 4940
rect 8540 4910 8550 4940
rect 8500 4900 8550 4910
rect 8350 4810 8360 4840
rect 8390 4810 8400 4840
rect 8350 4785 8400 4810
rect 8350 4765 8365 4785
rect 8385 4765 8400 4785
rect 8350 4740 8400 4765
rect 8350 4710 8360 4740
rect 8390 4710 8400 4740
rect 8350 4685 8400 4710
rect 8350 4665 8365 4685
rect 8385 4665 8400 4685
rect 8350 4640 8400 4665
rect 8350 4610 8360 4640
rect 8390 4610 8400 4640
rect 8350 4585 8400 4610
rect 8350 4565 8365 4585
rect 8385 4565 8400 4585
rect 8350 4540 8400 4565
rect 8350 4510 8360 4540
rect 8390 4510 8400 4540
rect 8350 4485 8400 4510
rect 8350 4465 8365 4485
rect 8385 4465 8400 4485
rect 8350 4440 8400 4465
rect 8350 4410 8360 4440
rect 8390 4410 8400 4440
rect 8350 4385 8400 4410
rect 8350 4365 8365 4385
rect 8385 4365 8400 4385
rect 4150 4260 4160 4290
rect 4190 4260 4200 4290
rect -50 4165 -35 4185
rect -15 4165 0 4185
rect -50 4135 0 4165
rect -50 4115 -35 4135
rect -15 4115 0 4135
rect -50 4085 0 4115
rect -50 4065 -35 4085
rect -15 4065 0 4085
rect -50 4035 0 4065
rect -50 4015 -35 4035
rect -15 4015 0 4035
rect -50 3985 0 4015
rect -50 3965 -35 3985
rect -15 3965 0 3985
rect -50 3935 0 3965
rect -50 3915 -35 3935
rect -15 3915 0 3935
rect -50 3885 0 3915
rect -50 3865 -35 3885
rect -15 3865 0 3885
rect -50 3835 0 3865
rect -50 3815 -35 3835
rect -15 3815 0 3835
rect -500 3640 -450 3650
rect -500 3610 -490 3640
rect -460 3610 -450 3640
rect -500 3600 -450 3610
rect -350 3640 -300 3700
rect -350 3610 -340 3640
rect -310 3610 -300 3640
rect -350 3550 -300 3610
rect -200 3640 -150 3650
rect -200 3610 -190 3640
rect -160 3610 -150 3640
rect -200 3600 -150 3610
rect -650 3510 -640 3540
rect -610 3510 -600 3540
rect -650 3485 -600 3510
rect -650 3465 -635 3485
rect -615 3465 -600 3485
rect -650 3440 -600 3465
rect -650 3410 -640 3440
rect -610 3410 -600 3440
rect -650 3385 -600 3410
rect -650 3365 -635 3385
rect -615 3365 -600 3385
rect -650 3340 -600 3365
rect -650 3310 -640 3340
rect -610 3310 -600 3340
rect -650 3285 -600 3310
rect -650 3265 -635 3285
rect -615 3265 -600 3285
rect -650 3240 -600 3265
rect -650 3210 -640 3240
rect -610 3210 -600 3240
rect -650 3185 -600 3210
rect -650 3165 -635 3185
rect -615 3165 -600 3185
rect -650 3140 -600 3165
rect -650 3110 -640 3140
rect -610 3110 -600 3140
rect -650 3085 -600 3110
rect -650 3065 -635 3085
rect -615 3065 -600 3085
rect -650 2990 -600 3065
rect -500 3535 -150 3550
rect -500 3515 -485 3535
rect -465 3515 -185 3535
rect -165 3515 -150 3535
rect -500 3500 -150 3515
rect -500 3485 -450 3500
rect -500 3465 -485 3485
rect -465 3465 -450 3485
rect -500 3435 -450 3465
rect -200 3485 -150 3500
rect -200 3465 -185 3485
rect -165 3465 -150 3485
rect -500 3415 -485 3435
rect -465 3415 -450 3435
rect -500 3385 -450 3415
rect -500 3365 -485 3385
rect -465 3365 -450 3385
rect -500 3335 -450 3365
rect -500 3315 -485 3335
rect -465 3315 -450 3335
rect -500 3285 -450 3315
rect -500 3265 -485 3285
rect -465 3265 -450 3285
rect -500 3235 -450 3265
rect -500 3215 -485 3235
rect -465 3215 -450 3235
rect -500 3185 -450 3215
rect -500 3165 -485 3185
rect -465 3165 -450 3185
rect -500 3135 -450 3165
rect -500 3115 -485 3135
rect -465 3115 -450 3135
rect -500 3085 -450 3115
rect -500 3065 -485 3085
rect -465 3065 -450 3085
rect -500 3050 -450 3065
rect -350 3435 -300 3450
rect -350 3415 -335 3435
rect -315 3415 -300 3435
rect -350 3385 -300 3415
rect -350 3365 -335 3385
rect -315 3365 -300 3385
rect -350 3335 -300 3365
rect -350 3315 -335 3335
rect -315 3315 -300 3335
rect -350 3285 -300 3315
rect -350 3265 -335 3285
rect -315 3265 -300 3285
rect -350 3235 -300 3265
rect -350 3215 -335 3235
rect -315 3215 -300 3235
rect -350 3185 -300 3215
rect -350 3165 -335 3185
rect -315 3165 -300 3185
rect -350 3135 -300 3165
rect -350 3115 -335 3135
rect -315 3115 -300 3135
rect -350 3085 -300 3115
rect -350 3065 -335 3085
rect -315 3065 -300 3085
rect -350 3050 -300 3065
rect -200 3435 -150 3465
rect -200 3415 -185 3435
rect -165 3415 -150 3435
rect -200 3385 -150 3415
rect -200 3365 -185 3385
rect -165 3365 -150 3385
rect -200 3335 -150 3365
rect -200 3315 -185 3335
rect -165 3315 -150 3335
rect -200 3285 -150 3315
rect -200 3265 -185 3285
rect -165 3265 -150 3285
rect -200 3235 -150 3265
rect -200 3215 -185 3235
rect -165 3215 -150 3235
rect -200 3185 -150 3215
rect -200 3165 -185 3185
rect -165 3165 -150 3185
rect -200 3135 -150 3165
rect -200 3115 -185 3135
rect -165 3115 -150 3135
rect -200 3085 -150 3115
rect -200 3065 -185 3085
rect -165 3065 -150 3085
rect -200 3050 -150 3065
rect -50 3540 0 3815
rect 550 4185 3600 4200
rect 550 4165 565 4185
rect 585 4165 865 4185
rect 885 4165 1165 4185
rect 1185 4165 1465 4185
rect 1485 4165 1765 4185
rect 1785 4165 2065 4185
rect 2085 4165 2365 4185
rect 2385 4165 2665 4185
rect 2685 4165 2965 4185
rect 2985 4165 3265 4185
rect 3285 4165 3565 4185
rect 3585 4165 3600 4185
rect 550 4150 3600 4165
rect 550 4135 600 4150
rect 550 4115 565 4135
rect 585 4115 600 4135
rect 550 4085 600 4115
rect 850 4135 900 4150
rect 850 4115 865 4135
rect 885 4115 900 4135
rect 550 4065 565 4085
rect 585 4065 600 4085
rect 550 4035 600 4065
rect 550 4015 565 4035
rect 585 4015 600 4035
rect 550 3985 600 4015
rect 550 3965 565 3985
rect 585 3965 600 3985
rect 550 3935 600 3965
rect 550 3915 565 3935
rect 585 3915 600 3935
rect 550 3885 600 3915
rect 550 3865 565 3885
rect 585 3865 600 3885
rect 550 3835 600 3865
rect 550 3815 565 3835
rect 585 3815 600 3835
rect 550 3785 600 3815
rect 550 3765 565 3785
rect 585 3765 600 3785
rect 550 3735 600 3765
rect 550 3715 565 3735
rect 585 3715 600 3735
rect 100 3640 150 3650
rect 100 3610 110 3640
rect 140 3610 150 3640
rect 100 3600 150 3610
rect 400 3640 450 3650
rect 400 3610 410 3640
rect 440 3610 450 3640
rect 400 3600 450 3610
rect -50 3510 -40 3540
rect -10 3510 0 3540
rect -50 3440 0 3510
rect -50 3410 -40 3440
rect -10 3410 0 3440
rect -50 3385 0 3410
rect -50 3365 -35 3385
rect -15 3365 0 3385
rect -50 3340 0 3365
rect -50 3310 -40 3340
rect -10 3310 0 3340
rect -50 3285 0 3310
rect -50 3265 -35 3285
rect -15 3265 0 3285
rect -50 3240 0 3265
rect -50 3210 -40 3240
rect -10 3210 0 3240
rect -50 3185 0 3210
rect -50 3165 -35 3185
rect -15 3165 0 3185
rect -50 3140 0 3165
rect -50 3110 -40 3140
rect -10 3110 0 3140
rect -50 3085 0 3110
rect -50 3065 -35 3085
rect -15 3065 0 3085
rect -650 2960 -640 2990
rect -610 2960 -600 2990
rect -650 2950 -600 2960
rect -50 2990 0 3065
rect 550 3535 600 3715
rect 700 4085 750 4100
rect 700 4065 715 4085
rect 735 4065 750 4085
rect 700 4035 750 4065
rect 700 4015 715 4035
rect 735 4015 750 4035
rect 700 3985 750 4015
rect 700 3965 715 3985
rect 735 3965 750 3985
rect 700 3935 750 3965
rect 700 3915 715 3935
rect 735 3915 750 3935
rect 700 3885 750 3915
rect 700 3865 715 3885
rect 735 3865 750 3885
rect 700 3835 750 3865
rect 700 3815 715 3835
rect 735 3815 750 3835
rect 700 3785 750 3815
rect 850 4085 900 4115
rect 1150 4135 1200 4150
rect 1150 4115 1165 4135
rect 1185 4115 1200 4135
rect 850 4065 865 4085
rect 885 4065 900 4085
rect 850 4035 900 4065
rect 850 4015 865 4035
rect 885 4015 900 4035
rect 850 3985 900 4015
rect 850 3965 865 3985
rect 885 3965 900 3985
rect 850 3935 900 3965
rect 850 3915 865 3935
rect 885 3915 900 3935
rect 850 3885 900 3915
rect 850 3865 865 3885
rect 885 3865 900 3885
rect 850 3835 900 3865
rect 850 3815 865 3835
rect 885 3815 900 3835
rect 850 3800 900 3815
rect 1000 4085 1050 4100
rect 1000 4065 1015 4085
rect 1035 4065 1050 4085
rect 1000 4035 1050 4065
rect 1000 4015 1015 4035
rect 1035 4015 1050 4035
rect 1000 3985 1050 4015
rect 1000 3965 1015 3985
rect 1035 3965 1050 3985
rect 1000 3935 1050 3965
rect 1000 3915 1015 3935
rect 1035 3915 1050 3935
rect 1000 3885 1050 3915
rect 1000 3865 1015 3885
rect 1035 3865 1050 3885
rect 1000 3835 1050 3865
rect 1000 3815 1015 3835
rect 1035 3815 1050 3835
rect 700 3765 715 3785
rect 735 3765 750 3785
rect 700 3750 750 3765
rect 1000 3785 1050 3815
rect 1150 4085 1200 4115
rect 1450 4135 1500 4150
rect 1450 4115 1465 4135
rect 1485 4115 1500 4135
rect 1150 4065 1165 4085
rect 1185 4065 1200 4085
rect 1150 4035 1200 4065
rect 1150 4015 1165 4035
rect 1185 4015 1200 4035
rect 1150 3985 1200 4015
rect 1150 3965 1165 3985
rect 1185 3965 1200 3985
rect 1150 3935 1200 3965
rect 1150 3915 1165 3935
rect 1185 3915 1200 3935
rect 1150 3885 1200 3915
rect 1150 3865 1165 3885
rect 1185 3865 1200 3885
rect 1150 3835 1200 3865
rect 1150 3815 1165 3835
rect 1185 3815 1200 3835
rect 1150 3800 1200 3815
rect 1300 4085 1350 4100
rect 1300 4065 1315 4085
rect 1335 4065 1350 4085
rect 1300 4035 1350 4065
rect 1300 4015 1315 4035
rect 1335 4015 1350 4035
rect 1300 3985 1350 4015
rect 1300 3965 1315 3985
rect 1335 3965 1350 3985
rect 1300 3935 1350 3965
rect 1300 3915 1315 3935
rect 1335 3915 1350 3935
rect 1300 3885 1350 3915
rect 1300 3865 1315 3885
rect 1335 3865 1350 3885
rect 1300 3835 1350 3865
rect 1300 3815 1315 3835
rect 1335 3815 1350 3835
rect 1000 3765 1015 3785
rect 1035 3765 1050 3785
rect 1000 3750 1050 3765
rect 1300 3785 1350 3815
rect 1450 4085 1500 4115
rect 1750 4135 1800 4150
rect 1750 4115 1765 4135
rect 1785 4115 1800 4135
rect 1450 4065 1465 4085
rect 1485 4065 1500 4085
rect 1450 4035 1500 4065
rect 1450 4015 1465 4035
rect 1485 4015 1500 4035
rect 1450 3985 1500 4015
rect 1450 3965 1465 3985
rect 1485 3965 1500 3985
rect 1450 3935 1500 3965
rect 1450 3915 1465 3935
rect 1485 3915 1500 3935
rect 1450 3885 1500 3915
rect 1450 3865 1465 3885
rect 1485 3865 1500 3885
rect 1450 3835 1500 3865
rect 1450 3815 1465 3835
rect 1485 3815 1500 3835
rect 1450 3800 1500 3815
rect 1600 4085 1650 4100
rect 1600 4065 1615 4085
rect 1635 4065 1650 4085
rect 1600 4035 1650 4065
rect 1600 4015 1615 4035
rect 1635 4015 1650 4035
rect 1600 3985 1650 4015
rect 1600 3965 1615 3985
rect 1635 3965 1650 3985
rect 1600 3935 1650 3965
rect 1600 3915 1615 3935
rect 1635 3915 1650 3935
rect 1600 3885 1650 3915
rect 1600 3865 1615 3885
rect 1635 3865 1650 3885
rect 1600 3835 1650 3865
rect 1600 3815 1615 3835
rect 1635 3815 1650 3835
rect 1300 3765 1315 3785
rect 1335 3765 1350 3785
rect 1300 3750 1350 3765
rect 1600 3785 1650 3815
rect 1600 3765 1615 3785
rect 1635 3765 1650 3785
rect 1600 3750 1650 3765
rect 700 3735 1650 3750
rect 700 3715 715 3735
rect 735 3715 1650 3735
rect 700 3700 1650 3715
rect 1750 4085 1800 4115
rect 2050 4135 2100 4150
rect 2050 4115 2065 4135
rect 2085 4115 2100 4135
rect 1750 4065 1765 4085
rect 1785 4065 1800 4085
rect 1750 4035 1800 4065
rect 1750 4015 1765 4035
rect 1785 4015 1800 4035
rect 1750 3985 1800 4015
rect 1750 3965 1765 3985
rect 1785 3965 1800 3985
rect 1750 3935 1800 3965
rect 1750 3915 1765 3935
rect 1785 3915 1800 3935
rect 1750 3885 1800 3915
rect 1750 3865 1765 3885
rect 1785 3865 1800 3885
rect 1750 3835 1800 3865
rect 1750 3815 1765 3835
rect 1785 3815 1800 3835
rect 1750 3785 1800 3815
rect 1750 3765 1765 3785
rect 1785 3765 1800 3785
rect 1750 3735 1800 3765
rect 1750 3715 1765 3735
rect 1785 3715 1800 3735
rect 700 3640 750 3650
rect 700 3610 710 3640
rect 740 3610 750 3640
rect 700 3600 750 3610
rect 1000 3640 1050 3650
rect 1000 3610 1010 3640
rect 1040 3610 1050 3640
rect 1000 3600 1050 3610
rect 1150 3640 1200 3700
rect 1150 3610 1160 3640
rect 1190 3610 1200 3640
rect 1150 3550 1200 3610
rect 1300 3640 1350 3650
rect 1300 3610 1310 3640
rect 1340 3610 1350 3640
rect 1300 3600 1350 3610
rect 1600 3640 1650 3650
rect 1600 3610 1610 3640
rect 1640 3610 1650 3640
rect 1600 3600 1650 3610
rect 550 3515 565 3535
rect 585 3515 600 3535
rect 550 3485 600 3515
rect 550 3465 565 3485
rect 585 3465 600 3485
rect 550 3435 600 3465
rect 550 3415 565 3435
rect 585 3415 600 3435
rect 550 3385 600 3415
rect 550 3365 565 3385
rect 585 3365 600 3385
rect 550 3335 600 3365
rect 550 3315 565 3335
rect 585 3315 600 3335
rect 550 3285 600 3315
rect 550 3265 565 3285
rect 585 3265 600 3285
rect 550 3235 600 3265
rect 550 3215 565 3235
rect 585 3215 600 3235
rect 550 3185 600 3215
rect 550 3165 565 3185
rect 585 3165 600 3185
rect 550 3135 600 3165
rect 700 3535 1650 3550
rect 700 3515 715 3535
rect 735 3515 1015 3535
rect 1035 3515 1315 3535
rect 1335 3515 1615 3535
rect 1635 3515 1650 3535
rect 700 3500 1650 3515
rect 700 3485 750 3500
rect 700 3465 715 3485
rect 735 3465 750 3485
rect 700 3435 750 3465
rect 1000 3485 1050 3500
rect 1000 3465 1015 3485
rect 1035 3465 1050 3485
rect 700 3415 715 3435
rect 735 3415 750 3435
rect 700 3385 750 3415
rect 700 3365 715 3385
rect 735 3365 750 3385
rect 700 3335 750 3365
rect 700 3315 715 3335
rect 735 3315 750 3335
rect 700 3285 750 3315
rect 700 3265 715 3285
rect 735 3265 750 3285
rect 700 3235 750 3265
rect 700 3215 715 3235
rect 735 3215 750 3235
rect 700 3185 750 3215
rect 700 3165 715 3185
rect 735 3165 750 3185
rect 700 3150 750 3165
rect 850 3435 900 3450
rect 850 3415 865 3435
rect 885 3415 900 3435
rect 850 3385 900 3415
rect 850 3365 865 3385
rect 885 3365 900 3385
rect 850 3335 900 3365
rect 850 3315 865 3335
rect 885 3315 900 3335
rect 850 3285 900 3315
rect 850 3265 865 3285
rect 885 3265 900 3285
rect 850 3235 900 3265
rect 850 3215 865 3235
rect 885 3215 900 3235
rect 850 3185 900 3215
rect 850 3165 865 3185
rect 885 3165 900 3185
rect 550 3115 565 3135
rect 585 3115 600 3135
rect 550 3100 600 3115
rect 850 3135 900 3165
rect 1000 3435 1050 3465
rect 1300 3485 1350 3500
rect 1300 3465 1315 3485
rect 1335 3465 1350 3485
rect 1000 3415 1015 3435
rect 1035 3415 1050 3435
rect 1000 3385 1050 3415
rect 1000 3365 1015 3385
rect 1035 3365 1050 3385
rect 1000 3335 1050 3365
rect 1000 3315 1015 3335
rect 1035 3315 1050 3335
rect 1000 3285 1050 3315
rect 1000 3265 1015 3285
rect 1035 3265 1050 3285
rect 1000 3235 1050 3265
rect 1000 3215 1015 3235
rect 1035 3215 1050 3235
rect 1000 3185 1050 3215
rect 1000 3165 1015 3185
rect 1035 3165 1050 3185
rect 1000 3150 1050 3165
rect 1150 3435 1200 3450
rect 1150 3415 1165 3435
rect 1185 3415 1200 3435
rect 1150 3385 1200 3415
rect 1150 3365 1165 3385
rect 1185 3365 1200 3385
rect 1150 3335 1200 3365
rect 1150 3315 1165 3335
rect 1185 3315 1200 3335
rect 1150 3285 1200 3315
rect 1150 3265 1165 3285
rect 1185 3265 1200 3285
rect 1150 3235 1200 3265
rect 1150 3215 1165 3235
rect 1185 3215 1200 3235
rect 1150 3185 1200 3215
rect 1150 3165 1165 3185
rect 1185 3165 1200 3185
rect 850 3115 865 3135
rect 885 3115 900 3135
rect 850 3100 900 3115
rect 1150 3135 1200 3165
rect 1300 3435 1350 3465
rect 1600 3485 1650 3500
rect 1600 3465 1615 3485
rect 1635 3465 1650 3485
rect 1300 3415 1315 3435
rect 1335 3415 1350 3435
rect 1300 3385 1350 3415
rect 1300 3365 1315 3385
rect 1335 3365 1350 3385
rect 1300 3335 1350 3365
rect 1300 3315 1315 3335
rect 1335 3315 1350 3335
rect 1300 3285 1350 3315
rect 1300 3265 1315 3285
rect 1335 3265 1350 3285
rect 1300 3235 1350 3265
rect 1300 3215 1315 3235
rect 1335 3215 1350 3235
rect 1300 3185 1350 3215
rect 1300 3165 1315 3185
rect 1335 3165 1350 3185
rect 1300 3150 1350 3165
rect 1450 3435 1500 3450
rect 1450 3415 1465 3435
rect 1485 3415 1500 3435
rect 1450 3385 1500 3415
rect 1450 3365 1465 3385
rect 1485 3365 1500 3385
rect 1450 3335 1500 3365
rect 1450 3315 1465 3335
rect 1485 3315 1500 3335
rect 1450 3285 1500 3315
rect 1450 3265 1465 3285
rect 1485 3265 1500 3285
rect 1450 3235 1500 3265
rect 1450 3215 1465 3235
rect 1485 3215 1500 3235
rect 1450 3185 1500 3215
rect 1450 3165 1465 3185
rect 1485 3165 1500 3185
rect 1150 3115 1165 3135
rect 1185 3115 1200 3135
rect 1150 3100 1200 3115
rect 1450 3135 1500 3165
rect 1600 3435 1650 3465
rect 1600 3415 1615 3435
rect 1635 3415 1650 3435
rect 1600 3385 1650 3415
rect 1600 3365 1615 3385
rect 1635 3365 1650 3385
rect 1600 3335 1650 3365
rect 1600 3315 1615 3335
rect 1635 3315 1650 3335
rect 1600 3285 1650 3315
rect 1600 3265 1615 3285
rect 1635 3265 1650 3285
rect 1600 3235 1650 3265
rect 1600 3215 1615 3235
rect 1635 3215 1650 3235
rect 1600 3185 1650 3215
rect 1600 3165 1615 3185
rect 1635 3165 1650 3185
rect 1600 3150 1650 3165
rect 1750 3535 1800 3715
rect 1900 4085 1950 4100
rect 1900 4065 1915 4085
rect 1935 4065 1950 4085
rect 1900 4035 1950 4065
rect 1900 4015 1915 4035
rect 1935 4015 1950 4035
rect 1900 3985 1950 4015
rect 1900 3965 1915 3985
rect 1935 3965 1950 3985
rect 1900 3935 1950 3965
rect 1900 3915 1915 3935
rect 1935 3915 1950 3935
rect 1900 3885 1950 3915
rect 1900 3865 1915 3885
rect 1935 3865 1950 3885
rect 1900 3835 1950 3865
rect 1900 3815 1915 3835
rect 1935 3815 1950 3835
rect 1900 3785 1950 3815
rect 2050 4085 2100 4115
rect 2350 4135 2400 4150
rect 2350 4115 2365 4135
rect 2385 4115 2400 4135
rect 2050 4065 2065 4085
rect 2085 4065 2100 4085
rect 2050 4035 2100 4065
rect 2050 4015 2065 4035
rect 2085 4015 2100 4035
rect 2050 3985 2100 4015
rect 2050 3965 2065 3985
rect 2085 3965 2100 3985
rect 2050 3935 2100 3965
rect 2050 3915 2065 3935
rect 2085 3915 2100 3935
rect 2050 3885 2100 3915
rect 2050 3865 2065 3885
rect 2085 3865 2100 3885
rect 2050 3835 2100 3865
rect 2050 3815 2065 3835
rect 2085 3815 2100 3835
rect 2050 3800 2100 3815
rect 2200 4085 2250 4100
rect 2200 4065 2215 4085
rect 2235 4065 2250 4085
rect 2200 4035 2250 4065
rect 2200 4015 2215 4035
rect 2235 4015 2250 4035
rect 2200 3985 2250 4015
rect 2200 3965 2215 3985
rect 2235 3965 2250 3985
rect 2200 3935 2250 3965
rect 2200 3915 2215 3935
rect 2235 3915 2250 3935
rect 2200 3885 2250 3915
rect 2200 3865 2215 3885
rect 2235 3865 2250 3885
rect 2200 3835 2250 3865
rect 2200 3815 2215 3835
rect 2235 3815 2250 3835
rect 1900 3765 1915 3785
rect 1935 3765 1950 3785
rect 1900 3750 1950 3765
rect 2200 3785 2250 3815
rect 2200 3765 2215 3785
rect 2235 3765 2250 3785
rect 2200 3750 2250 3765
rect 1900 3735 2250 3750
rect 1900 3715 1915 3735
rect 1935 3715 2215 3735
rect 2235 3715 2250 3735
rect 1900 3700 2250 3715
rect 2350 4085 2400 4115
rect 2650 4135 2700 4150
rect 2650 4115 2665 4135
rect 2685 4115 2700 4135
rect 2350 4065 2365 4085
rect 2385 4065 2400 4085
rect 2350 4035 2400 4065
rect 2350 4015 2365 4035
rect 2385 4015 2400 4035
rect 2350 3985 2400 4015
rect 2350 3965 2365 3985
rect 2385 3965 2400 3985
rect 2350 3935 2400 3965
rect 2350 3915 2365 3935
rect 2385 3915 2400 3935
rect 2350 3885 2400 3915
rect 2350 3865 2365 3885
rect 2385 3865 2400 3885
rect 2350 3835 2400 3865
rect 2350 3815 2365 3835
rect 2385 3815 2400 3835
rect 2350 3785 2400 3815
rect 2350 3765 2365 3785
rect 2385 3765 2400 3785
rect 2350 3735 2400 3765
rect 2350 3715 2365 3735
rect 2385 3715 2400 3735
rect 1900 3640 1950 3650
rect 1900 3610 1910 3640
rect 1940 3610 1950 3640
rect 1900 3600 1950 3610
rect 2050 3640 2100 3700
rect 2050 3610 2060 3640
rect 2090 3610 2100 3640
rect 2050 3550 2100 3610
rect 2200 3640 2250 3650
rect 2200 3610 2210 3640
rect 2240 3610 2250 3640
rect 2200 3600 2250 3610
rect 1750 3515 1765 3535
rect 1785 3515 1800 3535
rect 1750 3485 1800 3515
rect 1750 3465 1765 3485
rect 1785 3465 1800 3485
rect 1750 3435 1800 3465
rect 1750 3415 1765 3435
rect 1785 3415 1800 3435
rect 1750 3385 1800 3415
rect 1750 3365 1765 3385
rect 1785 3365 1800 3385
rect 1750 3335 1800 3365
rect 1750 3315 1765 3335
rect 1785 3315 1800 3335
rect 1750 3285 1800 3315
rect 1750 3265 1765 3285
rect 1785 3265 1800 3285
rect 1750 3235 1800 3265
rect 1750 3215 1765 3235
rect 1785 3215 1800 3235
rect 1750 3185 1800 3215
rect 1750 3165 1765 3185
rect 1785 3165 1800 3185
rect 1450 3115 1465 3135
rect 1485 3115 1500 3135
rect 1450 3100 1500 3115
rect 1750 3135 1800 3165
rect 1900 3535 2250 3550
rect 1900 3515 1915 3535
rect 1935 3515 2215 3535
rect 2235 3515 2250 3535
rect 1900 3500 2250 3515
rect 1900 3485 1950 3500
rect 1900 3465 1915 3485
rect 1935 3465 1950 3485
rect 1900 3435 1950 3465
rect 2200 3485 2250 3500
rect 2200 3465 2215 3485
rect 2235 3465 2250 3485
rect 1900 3415 1915 3435
rect 1935 3415 1950 3435
rect 1900 3385 1950 3415
rect 1900 3365 1915 3385
rect 1935 3365 1950 3385
rect 1900 3335 1950 3365
rect 1900 3315 1915 3335
rect 1935 3315 1950 3335
rect 1900 3285 1950 3315
rect 1900 3265 1915 3285
rect 1935 3265 1950 3285
rect 1900 3235 1950 3265
rect 1900 3215 1915 3235
rect 1935 3215 1950 3235
rect 1900 3185 1950 3215
rect 1900 3165 1915 3185
rect 1935 3165 1950 3185
rect 1900 3150 1950 3165
rect 2050 3435 2100 3450
rect 2050 3415 2065 3435
rect 2085 3415 2100 3435
rect 2050 3385 2100 3415
rect 2050 3365 2065 3385
rect 2085 3365 2100 3385
rect 2050 3335 2100 3365
rect 2050 3315 2065 3335
rect 2085 3315 2100 3335
rect 2050 3285 2100 3315
rect 2050 3265 2065 3285
rect 2085 3265 2100 3285
rect 2050 3235 2100 3265
rect 2050 3215 2065 3235
rect 2085 3215 2100 3235
rect 2050 3185 2100 3215
rect 2050 3165 2065 3185
rect 2085 3165 2100 3185
rect 1750 3115 1765 3135
rect 1785 3115 1800 3135
rect 1750 3100 1800 3115
rect 2050 3135 2100 3165
rect 2200 3435 2250 3465
rect 2200 3415 2215 3435
rect 2235 3415 2250 3435
rect 2200 3385 2250 3415
rect 2200 3365 2215 3385
rect 2235 3365 2250 3385
rect 2200 3335 2250 3365
rect 2200 3315 2215 3335
rect 2235 3315 2250 3335
rect 2200 3285 2250 3315
rect 2200 3265 2215 3285
rect 2235 3265 2250 3285
rect 2200 3235 2250 3265
rect 2200 3215 2215 3235
rect 2235 3215 2250 3235
rect 2200 3185 2250 3215
rect 2200 3165 2215 3185
rect 2235 3165 2250 3185
rect 2200 3150 2250 3165
rect 2350 3535 2400 3715
rect 2500 4085 2550 4100
rect 2500 4065 2515 4085
rect 2535 4065 2550 4085
rect 2500 4035 2550 4065
rect 2500 4015 2515 4035
rect 2535 4015 2550 4035
rect 2500 3985 2550 4015
rect 2500 3965 2515 3985
rect 2535 3965 2550 3985
rect 2500 3935 2550 3965
rect 2500 3915 2515 3935
rect 2535 3915 2550 3935
rect 2500 3885 2550 3915
rect 2500 3865 2515 3885
rect 2535 3865 2550 3885
rect 2500 3835 2550 3865
rect 2500 3815 2515 3835
rect 2535 3815 2550 3835
rect 2500 3785 2550 3815
rect 2650 4085 2700 4115
rect 2950 4135 3000 4150
rect 2950 4115 2965 4135
rect 2985 4115 3000 4135
rect 2650 4065 2665 4085
rect 2685 4065 2700 4085
rect 2650 4035 2700 4065
rect 2650 4015 2665 4035
rect 2685 4015 2700 4035
rect 2650 3985 2700 4015
rect 2650 3965 2665 3985
rect 2685 3965 2700 3985
rect 2650 3935 2700 3965
rect 2650 3915 2665 3935
rect 2685 3915 2700 3935
rect 2650 3885 2700 3915
rect 2650 3865 2665 3885
rect 2685 3865 2700 3885
rect 2650 3835 2700 3865
rect 2650 3815 2665 3835
rect 2685 3815 2700 3835
rect 2650 3800 2700 3815
rect 2800 4085 2850 4100
rect 2800 4065 2815 4085
rect 2835 4065 2850 4085
rect 2800 4035 2850 4065
rect 2800 4015 2815 4035
rect 2835 4015 2850 4035
rect 2800 3985 2850 4015
rect 2800 3965 2815 3985
rect 2835 3965 2850 3985
rect 2800 3935 2850 3965
rect 2800 3915 2815 3935
rect 2835 3915 2850 3935
rect 2800 3885 2850 3915
rect 2800 3865 2815 3885
rect 2835 3865 2850 3885
rect 2800 3835 2850 3865
rect 2800 3815 2815 3835
rect 2835 3815 2850 3835
rect 2500 3765 2515 3785
rect 2535 3765 2550 3785
rect 2500 3750 2550 3765
rect 2800 3785 2850 3815
rect 2950 4085 3000 4115
rect 3250 4135 3300 4150
rect 3250 4115 3265 4135
rect 3285 4115 3300 4135
rect 2950 4065 2965 4085
rect 2985 4065 3000 4085
rect 2950 4035 3000 4065
rect 2950 4015 2965 4035
rect 2985 4015 3000 4035
rect 2950 3985 3000 4015
rect 2950 3965 2965 3985
rect 2985 3965 3000 3985
rect 2950 3935 3000 3965
rect 2950 3915 2965 3935
rect 2985 3915 3000 3935
rect 2950 3885 3000 3915
rect 2950 3865 2965 3885
rect 2985 3865 3000 3885
rect 2950 3835 3000 3865
rect 2950 3815 2965 3835
rect 2985 3815 3000 3835
rect 2950 3800 3000 3815
rect 3100 4085 3150 4100
rect 3100 4065 3115 4085
rect 3135 4065 3150 4085
rect 3100 4035 3150 4065
rect 3100 4015 3115 4035
rect 3135 4015 3150 4035
rect 3100 3985 3150 4015
rect 3100 3965 3115 3985
rect 3135 3965 3150 3985
rect 3100 3935 3150 3965
rect 3100 3915 3115 3935
rect 3135 3915 3150 3935
rect 3100 3885 3150 3915
rect 3100 3865 3115 3885
rect 3135 3865 3150 3885
rect 3100 3835 3150 3865
rect 3100 3815 3115 3835
rect 3135 3815 3150 3835
rect 2800 3765 2815 3785
rect 2835 3765 2850 3785
rect 2800 3750 2850 3765
rect 3100 3785 3150 3815
rect 3250 4085 3300 4115
rect 3550 4135 3600 4150
rect 3550 4115 3565 4135
rect 3585 4115 3600 4135
rect 3250 4065 3265 4085
rect 3285 4065 3300 4085
rect 3250 4035 3300 4065
rect 3250 4015 3265 4035
rect 3285 4015 3300 4035
rect 3250 3985 3300 4015
rect 3250 3965 3265 3985
rect 3285 3965 3300 3985
rect 3250 3935 3300 3965
rect 3250 3915 3265 3935
rect 3285 3915 3300 3935
rect 3250 3885 3300 3915
rect 3250 3865 3265 3885
rect 3285 3865 3300 3885
rect 3250 3835 3300 3865
rect 3250 3815 3265 3835
rect 3285 3815 3300 3835
rect 3250 3800 3300 3815
rect 3400 4085 3450 4100
rect 3400 4065 3415 4085
rect 3435 4065 3450 4085
rect 3400 4035 3450 4065
rect 3400 4015 3415 4035
rect 3435 4015 3450 4035
rect 3400 3985 3450 4015
rect 3400 3965 3415 3985
rect 3435 3965 3450 3985
rect 3400 3935 3450 3965
rect 3400 3915 3415 3935
rect 3435 3915 3450 3935
rect 3400 3885 3450 3915
rect 3400 3865 3415 3885
rect 3435 3865 3450 3885
rect 3400 3835 3450 3865
rect 3400 3815 3415 3835
rect 3435 3815 3450 3835
rect 3100 3765 3115 3785
rect 3135 3765 3150 3785
rect 3100 3750 3150 3765
rect 3400 3785 3450 3815
rect 3400 3765 3415 3785
rect 3435 3765 3450 3785
rect 3400 3750 3450 3765
rect 2500 3735 3450 3750
rect 2500 3715 3415 3735
rect 3435 3715 3450 3735
rect 2500 3700 3450 3715
rect 3550 4085 3600 4115
rect 3550 4065 3565 4085
rect 3585 4065 3600 4085
rect 3550 4035 3600 4065
rect 3550 4015 3565 4035
rect 3585 4015 3600 4035
rect 3550 3985 3600 4015
rect 3550 3965 3565 3985
rect 3585 3965 3600 3985
rect 3550 3935 3600 3965
rect 3550 3915 3565 3935
rect 3585 3915 3600 3935
rect 3550 3885 3600 3915
rect 3550 3865 3565 3885
rect 3585 3865 3600 3885
rect 3550 3835 3600 3865
rect 3550 3815 3565 3835
rect 3585 3815 3600 3835
rect 3550 3785 3600 3815
rect 3550 3765 3565 3785
rect 3585 3765 3600 3785
rect 3550 3735 3600 3765
rect 3550 3715 3565 3735
rect 3585 3715 3600 3735
rect 2500 3640 2550 3650
rect 2500 3610 2510 3640
rect 2540 3610 2550 3640
rect 2500 3600 2550 3610
rect 2800 3640 2850 3650
rect 2800 3610 2810 3640
rect 2840 3610 2850 3640
rect 2800 3600 2850 3610
rect 2950 3640 3000 3700
rect 2950 3610 2960 3640
rect 2990 3610 3000 3640
rect 2950 3550 3000 3610
rect 3100 3640 3150 3650
rect 3100 3610 3110 3640
rect 3140 3610 3150 3640
rect 3100 3600 3150 3610
rect 3400 3640 3450 3650
rect 3400 3610 3410 3640
rect 3440 3610 3450 3640
rect 3400 3600 3450 3610
rect 2350 3515 2365 3535
rect 2385 3515 2400 3535
rect 2350 3485 2400 3515
rect 2350 3465 2365 3485
rect 2385 3465 2400 3485
rect 2350 3435 2400 3465
rect 2350 3415 2365 3435
rect 2385 3415 2400 3435
rect 2350 3385 2400 3415
rect 2350 3365 2365 3385
rect 2385 3365 2400 3385
rect 2350 3335 2400 3365
rect 2350 3315 2365 3335
rect 2385 3315 2400 3335
rect 2350 3285 2400 3315
rect 2350 3265 2365 3285
rect 2385 3265 2400 3285
rect 2350 3235 2400 3265
rect 2350 3215 2365 3235
rect 2385 3215 2400 3235
rect 2350 3185 2400 3215
rect 2350 3165 2365 3185
rect 2385 3165 2400 3185
rect 2050 3115 2065 3135
rect 2085 3115 2100 3135
rect 2050 3100 2100 3115
rect 2350 3135 2400 3165
rect 2500 3535 3450 3550
rect 2500 3515 2515 3535
rect 2535 3515 2815 3535
rect 2835 3515 3115 3535
rect 3135 3515 3415 3535
rect 3435 3515 3450 3535
rect 2500 3500 3450 3515
rect 2500 3485 2550 3500
rect 2500 3465 2515 3485
rect 2535 3465 2550 3485
rect 2500 3435 2550 3465
rect 2800 3485 2850 3500
rect 2800 3465 2815 3485
rect 2835 3465 2850 3485
rect 2500 3415 2515 3435
rect 2535 3415 2550 3435
rect 2500 3385 2550 3415
rect 2500 3365 2515 3385
rect 2535 3365 2550 3385
rect 2500 3335 2550 3365
rect 2500 3315 2515 3335
rect 2535 3315 2550 3335
rect 2500 3285 2550 3315
rect 2500 3265 2515 3285
rect 2535 3265 2550 3285
rect 2500 3235 2550 3265
rect 2500 3215 2515 3235
rect 2535 3215 2550 3235
rect 2500 3185 2550 3215
rect 2500 3165 2515 3185
rect 2535 3165 2550 3185
rect 2500 3150 2550 3165
rect 2650 3435 2700 3450
rect 2650 3415 2665 3435
rect 2685 3415 2700 3435
rect 2650 3385 2700 3415
rect 2650 3365 2665 3385
rect 2685 3365 2700 3385
rect 2650 3335 2700 3365
rect 2650 3315 2665 3335
rect 2685 3315 2700 3335
rect 2650 3285 2700 3315
rect 2650 3265 2665 3285
rect 2685 3265 2700 3285
rect 2650 3235 2700 3265
rect 2650 3215 2665 3235
rect 2685 3215 2700 3235
rect 2650 3185 2700 3215
rect 2650 3165 2665 3185
rect 2685 3165 2700 3185
rect 2350 3115 2365 3135
rect 2385 3115 2400 3135
rect 2350 3100 2400 3115
rect 2650 3135 2700 3165
rect 2800 3435 2850 3465
rect 3100 3485 3150 3500
rect 3100 3465 3115 3485
rect 3135 3465 3150 3485
rect 2800 3415 2815 3435
rect 2835 3415 2850 3435
rect 2800 3385 2850 3415
rect 2800 3365 2815 3385
rect 2835 3365 2850 3385
rect 2800 3335 2850 3365
rect 2800 3315 2815 3335
rect 2835 3315 2850 3335
rect 2800 3285 2850 3315
rect 2800 3265 2815 3285
rect 2835 3265 2850 3285
rect 2800 3235 2850 3265
rect 2800 3215 2815 3235
rect 2835 3215 2850 3235
rect 2800 3185 2850 3215
rect 2800 3165 2815 3185
rect 2835 3165 2850 3185
rect 2800 3150 2850 3165
rect 2950 3435 3000 3450
rect 2950 3415 2965 3435
rect 2985 3415 3000 3435
rect 2950 3385 3000 3415
rect 2950 3365 2965 3385
rect 2985 3365 3000 3385
rect 2950 3335 3000 3365
rect 2950 3315 2965 3335
rect 2985 3315 3000 3335
rect 2950 3285 3000 3315
rect 2950 3265 2965 3285
rect 2985 3265 3000 3285
rect 2950 3235 3000 3265
rect 2950 3215 2965 3235
rect 2985 3215 3000 3235
rect 2950 3185 3000 3215
rect 2950 3165 2965 3185
rect 2985 3165 3000 3185
rect 2650 3115 2665 3135
rect 2685 3115 2700 3135
rect 2650 3100 2700 3115
rect 2950 3135 3000 3165
rect 3100 3435 3150 3465
rect 3400 3485 3450 3500
rect 3400 3465 3415 3485
rect 3435 3465 3450 3485
rect 3100 3415 3115 3435
rect 3135 3415 3150 3435
rect 3100 3385 3150 3415
rect 3100 3365 3115 3385
rect 3135 3365 3150 3385
rect 3100 3335 3150 3365
rect 3100 3315 3115 3335
rect 3135 3315 3150 3335
rect 3100 3285 3150 3315
rect 3100 3265 3115 3285
rect 3135 3265 3150 3285
rect 3100 3235 3150 3265
rect 3100 3215 3115 3235
rect 3135 3215 3150 3235
rect 3100 3185 3150 3215
rect 3100 3165 3115 3185
rect 3135 3165 3150 3185
rect 3100 3150 3150 3165
rect 3250 3435 3300 3450
rect 3250 3415 3265 3435
rect 3285 3415 3300 3435
rect 3250 3385 3300 3415
rect 3250 3365 3265 3385
rect 3285 3365 3300 3385
rect 3250 3335 3300 3365
rect 3250 3315 3265 3335
rect 3285 3315 3300 3335
rect 3250 3285 3300 3315
rect 3250 3265 3265 3285
rect 3285 3265 3300 3285
rect 3250 3235 3300 3265
rect 3250 3215 3265 3235
rect 3285 3215 3300 3235
rect 3250 3185 3300 3215
rect 3250 3165 3265 3185
rect 3285 3165 3300 3185
rect 2950 3115 2965 3135
rect 2985 3115 3000 3135
rect 2950 3100 3000 3115
rect 3250 3135 3300 3165
rect 3400 3435 3450 3465
rect 3400 3415 3415 3435
rect 3435 3415 3450 3435
rect 3400 3385 3450 3415
rect 3400 3365 3415 3385
rect 3435 3365 3450 3385
rect 3400 3335 3450 3365
rect 3400 3315 3415 3335
rect 3435 3315 3450 3335
rect 3400 3285 3450 3315
rect 3400 3265 3415 3285
rect 3435 3265 3450 3285
rect 3400 3235 3450 3265
rect 3400 3215 3415 3235
rect 3435 3215 3450 3235
rect 3400 3185 3450 3215
rect 3400 3165 3415 3185
rect 3435 3165 3450 3185
rect 3400 3150 3450 3165
rect 3550 3535 3600 3715
rect 4150 4185 4200 4260
rect 8350 4290 8400 4365
rect 8500 4835 8550 4850
rect 8500 4815 8515 4835
rect 8535 4815 8550 4835
rect 8500 4785 8550 4815
rect 8500 4765 8515 4785
rect 8535 4765 8550 4785
rect 8500 4735 8550 4765
rect 8500 4715 8515 4735
rect 8535 4715 8550 4735
rect 8500 4685 8550 4715
rect 8500 4665 8515 4685
rect 8535 4665 8550 4685
rect 8500 4635 8550 4665
rect 8500 4615 8515 4635
rect 8535 4615 8550 4635
rect 8500 4585 8550 4615
rect 8500 4565 8515 4585
rect 8535 4565 8550 4585
rect 8500 4535 8550 4565
rect 8500 4515 8515 4535
rect 8535 4515 8550 4535
rect 8500 4485 8550 4515
rect 8500 4465 8515 4485
rect 8535 4465 8550 4485
rect 8500 4435 8550 4465
rect 8500 4415 8515 4435
rect 8535 4415 8550 4435
rect 8500 4385 8550 4415
rect 8500 4365 8515 4385
rect 8535 4365 8550 4385
rect 8500 4350 8550 4365
rect 8650 4840 8700 5010
rect 8800 5485 8850 5500
rect 8800 5465 8815 5485
rect 8835 5465 8850 5485
rect 8800 5435 8850 5465
rect 8800 5415 8815 5435
rect 8835 5415 8850 5435
rect 8800 5385 8850 5415
rect 8800 5365 8815 5385
rect 8835 5365 8850 5385
rect 8800 5335 8850 5365
rect 8800 5315 8815 5335
rect 8835 5315 8850 5335
rect 8800 5285 8850 5315
rect 8800 5265 8815 5285
rect 8835 5265 8850 5285
rect 8800 5235 8850 5265
rect 8800 5215 8815 5235
rect 8835 5215 8850 5235
rect 8800 5185 8850 5215
rect 8800 5165 8815 5185
rect 8835 5165 8850 5185
rect 8800 5135 8850 5165
rect 8800 5115 8815 5135
rect 8835 5115 8850 5135
rect 8800 5085 8850 5115
rect 8800 5065 8815 5085
rect 8835 5065 8850 5085
rect 8800 5035 8850 5065
rect 8800 5015 8815 5035
rect 8835 5015 8850 5035
rect 8800 5000 8850 5015
rect 8950 5485 9000 5560
rect 9250 5590 9300 5600
rect 9250 5560 9260 5590
rect 9290 5560 9300 5590
rect 8950 5465 8965 5485
rect 8985 5465 9000 5485
rect 8950 5440 9000 5465
rect 8950 5410 8960 5440
rect 8990 5410 9000 5440
rect 8950 5385 9000 5410
rect 8950 5365 8965 5385
rect 8985 5365 9000 5385
rect 8950 5340 9000 5365
rect 8950 5310 8960 5340
rect 8990 5310 9000 5340
rect 8950 5285 9000 5310
rect 8950 5265 8965 5285
rect 8985 5265 9000 5285
rect 8950 5240 9000 5265
rect 8950 5210 8960 5240
rect 8990 5210 9000 5240
rect 8950 5185 9000 5210
rect 8950 5165 8965 5185
rect 8985 5165 9000 5185
rect 8950 5140 9000 5165
rect 8950 5110 8960 5140
rect 8990 5110 9000 5140
rect 8950 5085 9000 5110
rect 8950 5065 8965 5085
rect 8985 5065 9000 5085
rect 8950 5040 9000 5065
rect 8950 5010 8960 5040
rect 8990 5010 9000 5040
rect 8800 4940 8850 4950
rect 8800 4910 8810 4940
rect 8840 4910 8850 4940
rect 8800 4900 8850 4910
rect 8650 4810 8660 4840
rect 8690 4810 8700 4840
rect 8650 4785 8700 4810
rect 8650 4765 8665 4785
rect 8685 4765 8700 4785
rect 8650 4740 8700 4765
rect 8650 4710 8660 4740
rect 8690 4710 8700 4740
rect 8650 4685 8700 4710
rect 8650 4665 8665 4685
rect 8685 4665 8700 4685
rect 8650 4640 8700 4665
rect 8650 4610 8660 4640
rect 8690 4610 8700 4640
rect 8650 4585 8700 4610
rect 8650 4565 8665 4585
rect 8685 4565 8700 4585
rect 8650 4540 8700 4565
rect 8650 4510 8660 4540
rect 8690 4510 8700 4540
rect 8650 4485 8700 4510
rect 8650 4465 8665 4485
rect 8685 4465 8700 4485
rect 8650 4440 8700 4465
rect 8650 4410 8660 4440
rect 8690 4410 8700 4440
rect 8650 4385 8700 4410
rect 8650 4365 8665 4385
rect 8685 4365 8700 4385
rect 8350 4260 8360 4290
rect 8390 4260 8400 4290
rect 4150 4165 4165 4185
rect 4185 4165 4200 4185
rect 4150 4135 4200 4165
rect 4150 4115 4165 4135
rect 4185 4115 4200 4135
rect 4150 4085 4200 4115
rect 4150 4065 4165 4085
rect 4185 4065 4200 4085
rect 4150 4035 4200 4065
rect 4150 4015 4165 4035
rect 4185 4015 4200 4035
rect 4150 3985 4200 4015
rect 4150 3965 4165 3985
rect 4185 3965 4200 3985
rect 4150 3935 4200 3965
rect 4150 3915 4165 3935
rect 4185 3915 4200 3935
rect 4150 3885 4200 3915
rect 4150 3865 4165 3885
rect 4185 3865 4200 3885
rect 4150 3835 4200 3865
rect 4150 3815 4165 3835
rect 4185 3815 4200 3835
rect 3700 3640 3750 3650
rect 3700 3610 3710 3640
rect 3740 3610 3750 3640
rect 3700 3600 3750 3610
rect 4000 3640 4050 3650
rect 4000 3610 4010 3640
rect 4040 3610 4050 3640
rect 4000 3600 4050 3610
rect 3550 3515 3565 3535
rect 3585 3515 3600 3535
rect 3550 3485 3600 3515
rect 3550 3465 3565 3485
rect 3585 3465 3600 3485
rect 3550 3435 3600 3465
rect 3550 3415 3565 3435
rect 3585 3415 3600 3435
rect 3550 3385 3600 3415
rect 3550 3365 3565 3385
rect 3585 3365 3600 3385
rect 3550 3335 3600 3365
rect 3550 3315 3565 3335
rect 3585 3315 3600 3335
rect 3550 3285 3600 3315
rect 3550 3265 3565 3285
rect 3585 3265 3600 3285
rect 3550 3235 3600 3265
rect 3550 3215 3565 3235
rect 3585 3215 3600 3235
rect 3550 3185 3600 3215
rect 3550 3165 3565 3185
rect 3585 3165 3600 3185
rect 3250 3115 3265 3135
rect 3285 3115 3300 3135
rect 3250 3100 3300 3115
rect 3550 3135 3600 3165
rect 3550 3115 3565 3135
rect 3585 3115 3600 3135
rect 3550 3100 3600 3115
rect 550 3085 3600 3100
rect 550 3065 565 3085
rect 585 3065 865 3085
rect 885 3065 1165 3085
rect 1185 3065 1465 3085
rect 1485 3065 1765 3085
rect 1785 3065 2065 3085
rect 2085 3065 2365 3085
rect 2385 3065 2665 3085
rect 2685 3065 2965 3085
rect 2985 3065 3265 3085
rect 3285 3065 3565 3085
rect 3585 3065 3600 3085
rect 550 3050 3600 3065
rect 4150 3540 4200 3815
rect 4750 4185 7800 4200
rect 4750 4165 4765 4185
rect 4785 4165 5065 4185
rect 5085 4165 5365 4185
rect 5385 4165 5665 4185
rect 5685 4165 5965 4185
rect 5985 4165 6265 4185
rect 6285 4165 6565 4185
rect 6585 4165 6865 4185
rect 6885 4165 7165 4185
rect 7185 4165 7465 4185
rect 7485 4165 7765 4185
rect 7785 4165 7800 4185
rect 4750 4150 7800 4165
rect 4750 4135 4800 4150
rect 4750 4115 4765 4135
rect 4785 4115 4800 4135
rect 4750 4085 4800 4115
rect 5050 4135 5100 4150
rect 5050 4115 5065 4135
rect 5085 4115 5100 4135
rect 4750 4065 4765 4085
rect 4785 4065 4800 4085
rect 4750 4035 4800 4065
rect 4750 4015 4765 4035
rect 4785 4015 4800 4035
rect 4750 3985 4800 4015
rect 4750 3965 4765 3985
rect 4785 3965 4800 3985
rect 4750 3935 4800 3965
rect 4750 3915 4765 3935
rect 4785 3915 4800 3935
rect 4750 3885 4800 3915
rect 4750 3865 4765 3885
rect 4785 3865 4800 3885
rect 4750 3835 4800 3865
rect 4750 3815 4765 3835
rect 4785 3815 4800 3835
rect 4750 3785 4800 3815
rect 4750 3765 4765 3785
rect 4785 3765 4800 3785
rect 4750 3735 4800 3765
rect 4750 3715 4765 3735
rect 4785 3715 4800 3735
rect 4300 3640 4350 3650
rect 4300 3610 4310 3640
rect 4340 3610 4350 3640
rect 4300 3600 4350 3610
rect 4600 3640 4650 3650
rect 4600 3610 4610 3640
rect 4640 3610 4650 3640
rect 4600 3600 4650 3610
rect 4150 3510 4160 3540
rect 4190 3510 4200 3540
rect 4150 3440 4200 3510
rect 4150 3410 4160 3440
rect 4190 3410 4200 3440
rect 4150 3385 4200 3410
rect 4150 3365 4165 3385
rect 4185 3365 4200 3385
rect 4150 3340 4200 3365
rect 4150 3310 4160 3340
rect 4190 3310 4200 3340
rect 4150 3285 4200 3310
rect 4150 3265 4165 3285
rect 4185 3265 4200 3285
rect 4150 3240 4200 3265
rect 4150 3210 4160 3240
rect 4190 3210 4200 3240
rect 4150 3185 4200 3210
rect 4150 3165 4165 3185
rect 4185 3165 4200 3185
rect 4150 3140 4200 3165
rect 4150 3110 4160 3140
rect 4190 3110 4200 3140
rect 4150 3085 4200 3110
rect 4150 3065 4165 3085
rect 4185 3065 4200 3085
rect -50 2960 -40 2990
rect -10 2960 0 2990
rect -50 2950 0 2960
rect 4150 2990 4200 3065
rect 4750 3535 4800 3715
rect 4900 4085 4950 4100
rect 4900 4065 4915 4085
rect 4935 4065 4950 4085
rect 4900 4035 4950 4065
rect 4900 4015 4915 4035
rect 4935 4015 4950 4035
rect 4900 3985 4950 4015
rect 4900 3965 4915 3985
rect 4935 3965 4950 3985
rect 4900 3935 4950 3965
rect 4900 3915 4915 3935
rect 4935 3915 4950 3935
rect 4900 3885 4950 3915
rect 4900 3865 4915 3885
rect 4935 3865 4950 3885
rect 4900 3835 4950 3865
rect 4900 3815 4915 3835
rect 4935 3815 4950 3835
rect 4900 3785 4950 3815
rect 5050 4085 5100 4115
rect 5350 4135 5400 4150
rect 5350 4115 5365 4135
rect 5385 4115 5400 4135
rect 5050 4065 5065 4085
rect 5085 4065 5100 4085
rect 5050 4035 5100 4065
rect 5050 4015 5065 4035
rect 5085 4015 5100 4035
rect 5050 3985 5100 4015
rect 5050 3965 5065 3985
rect 5085 3965 5100 3985
rect 5050 3935 5100 3965
rect 5050 3915 5065 3935
rect 5085 3915 5100 3935
rect 5050 3885 5100 3915
rect 5050 3865 5065 3885
rect 5085 3865 5100 3885
rect 5050 3835 5100 3865
rect 5050 3815 5065 3835
rect 5085 3815 5100 3835
rect 5050 3800 5100 3815
rect 5200 4085 5250 4100
rect 5200 4065 5215 4085
rect 5235 4065 5250 4085
rect 5200 4035 5250 4065
rect 5200 4015 5215 4035
rect 5235 4015 5250 4035
rect 5200 3985 5250 4015
rect 5200 3965 5215 3985
rect 5235 3965 5250 3985
rect 5200 3935 5250 3965
rect 5200 3915 5215 3935
rect 5235 3915 5250 3935
rect 5200 3885 5250 3915
rect 5200 3865 5215 3885
rect 5235 3865 5250 3885
rect 5200 3835 5250 3865
rect 5200 3815 5215 3835
rect 5235 3815 5250 3835
rect 4900 3765 4915 3785
rect 4935 3765 4950 3785
rect 4900 3750 4950 3765
rect 5200 3785 5250 3815
rect 5350 4085 5400 4115
rect 5650 4135 5700 4150
rect 5650 4115 5665 4135
rect 5685 4115 5700 4135
rect 5350 4065 5365 4085
rect 5385 4065 5400 4085
rect 5350 4035 5400 4065
rect 5350 4015 5365 4035
rect 5385 4015 5400 4035
rect 5350 3985 5400 4015
rect 5350 3965 5365 3985
rect 5385 3965 5400 3985
rect 5350 3935 5400 3965
rect 5350 3915 5365 3935
rect 5385 3915 5400 3935
rect 5350 3885 5400 3915
rect 5350 3865 5365 3885
rect 5385 3865 5400 3885
rect 5350 3835 5400 3865
rect 5350 3815 5365 3835
rect 5385 3815 5400 3835
rect 5350 3800 5400 3815
rect 5500 4085 5550 4100
rect 5500 4065 5515 4085
rect 5535 4065 5550 4085
rect 5500 4035 5550 4065
rect 5500 4015 5515 4035
rect 5535 4015 5550 4035
rect 5500 3985 5550 4015
rect 5500 3965 5515 3985
rect 5535 3965 5550 3985
rect 5500 3935 5550 3965
rect 5500 3915 5515 3935
rect 5535 3915 5550 3935
rect 5500 3885 5550 3915
rect 5500 3865 5515 3885
rect 5535 3865 5550 3885
rect 5500 3835 5550 3865
rect 5500 3815 5515 3835
rect 5535 3815 5550 3835
rect 5200 3765 5215 3785
rect 5235 3765 5250 3785
rect 5200 3750 5250 3765
rect 5500 3785 5550 3815
rect 5650 4085 5700 4115
rect 5950 4135 6000 4150
rect 5950 4115 5965 4135
rect 5985 4115 6000 4135
rect 5650 4065 5665 4085
rect 5685 4065 5700 4085
rect 5650 4035 5700 4065
rect 5650 4015 5665 4035
rect 5685 4015 5700 4035
rect 5650 3985 5700 4015
rect 5650 3965 5665 3985
rect 5685 3965 5700 3985
rect 5650 3935 5700 3965
rect 5650 3915 5665 3935
rect 5685 3915 5700 3935
rect 5650 3885 5700 3915
rect 5650 3865 5665 3885
rect 5685 3865 5700 3885
rect 5650 3835 5700 3865
rect 5650 3815 5665 3835
rect 5685 3815 5700 3835
rect 5650 3800 5700 3815
rect 5800 4085 5850 4100
rect 5800 4065 5815 4085
rect 5835 4065 5850 4085
rect 5800 4035 5850 4065
rect 5800 4015 5815 4035
rect 5835 4015 5850 4035
rect 5800 3985 5850 4015
rect 5800 3965 5815 3985
rect 5835 3965 5850 3985
rect 5800 3935 5850 3965
rect 5800 3915 5815 3935
rect 5835 3915 5850 3935
rect 5800 3885 5850 3915
rect 5800 3865 5815 3885
rect 5835 3865 5850 3885
rect 5800 3835 5850 3865
rect 5800 3815 5815 3835
rect 5835 3815 5850 3835
rect 5500 3765 5515 3785
rect 5535 3765 5550 3785
rect 5500 3750 5550 3765
rect 5800 3785 5850 3815
rect 5800 3765 5815 3785
rect 5835 3765 5850 3785
rect 5800 3750 5850 3765
rect 4900 3735 5850 3750
rect 4900 3715 4915 3735
rect 4935 3715 5850 3735
rect 4900 3700 5850 3715
rect 5950 4085 6000 4115
rect 6250 4135 6300 4150
rect 6250 4115 6265 4135
rect 6285 4115 6300 4135
rect 5950 4065 5965 4085
rect 5985 4065 6000 4085
rect 5950 4035 6000 4065
rect 5950 4015 5965 4035
rect 5985 4015 6000 4035
rect 5950 3985 6000 4015
rect 5950 3965 5965 3985
rect 5985 3965 6000 3985
rect 5950 3935 6000 3965
rect 5950 3915 5965 3935
rect 5985 3915 6000 3935
rect 5950 3885 6000 3915
rect 5950 3865 5965 3885
rect 5985 3865 6000 3885
rect 5950 3835 6000 3865
rect 5950 3815 5965 3835
rect 5985 3815 6000 3835
rect 5950 3785 6000 3815
rect 5950 3765 5965 3785
rect 5985 3765 6000 3785
rect 5950 3735 6000 3765
rect 5950 3715 5965 3735
rect 5985 3715 6000 3735
rect 4900 3640 4950 3650
rect 4900 3610 4910 3640
rect 4940 3610 4950 3640
rect 4900 3600 4950 3610
rect 5200 3640 5250 3650
rect 5200 3610 5210 3640
rect 5240 3610 5250 3640
rect 5200 3600 5250 3610
rect 5350 3640 5400 3700
rect 5350 3610 5360 3640
rect 5390 3610 5400 3640
rect 5350 3550 5400 3610
rect 5500 3640 5550 3650
rect 5500 3610 5510 3640
rect 5540 3610 5550 3640
rect 5500 3600 5550 3610
rect 5800 3640 5850 3650
rect 5800 3610 5810 3640
rect 5840 3610 5850 3640
rect 5800 3600 5850 3610
rect 4750 3515 4765 3535
rect 4785 3515 4800 3535
rect 4750 3485 4800 3515
rect 4750 3465 4765 3485
rect 4785 3465 4800 3485
rect 4750 3435 4800 3465
rect 4750 3415 4765 3435
rect 4785 3415 4800 3435
rect 4750 3385 4800 3415
rect 4750 3365 4765 3385
rect 4785 3365 4800 3385
rect 4750 3335 4800 3365
rect 4750 3315 4765 3335
rect 4785 3315 4800 3335
rect 4750 3285 4800 3315
rect 4750 3265 4765 3285
rect 4785 3265 4800 3285
rect 4750 3235 4800 3265
rect 4750 3215 4765 3235
rect 4785 3215 4800 3235
rect 4750 3185 4800 3215
rect 4750 3165 4765 3185
rect 4785 3165 4800 3185
rect 4750 3135 4800 3165
rect 4900 3535 5850 3550
rect 4900 3515 4915 3535
rect 4935 3515 5215 3535
rect 5235 3515 5515 3535
rect 5535 3515 5815 3535
rect 5835 3515 5850 3535
rect 4900 3500 5850 3515
rect 4900 3485 4950 3500
rect 4900 3465 4915 3485
rect 4935 3465 4950 3485
rect 4900 3435 4950 3465
rect 5200 3485 5250 3500
rect 5200 3465 5215 3485
rect 5235 3465 5250 3485
rect 4900 3415 4915 3435
rect 4935 3415 4950 3435
rect 4900 3385 4950 3415
rect 4900 3365 4915 3385
rect 4935 3365 4950 3385
rect 4900 3335 4950 3365
rect 4900 3315 4915 3335
rect 4935 3315 4950 3335
rect 4900 3285 4950 3315
rect 4900 3265 4915 3285
rect 4935 3265 4950 3285
rect 4900 3235 4950 3265
rect 4900 3215 4915 3235
rect 4935 3215 4950 3235
rect 4900 3185 4950 3215
rect 4900 3165 4915 3185
rect 4935 3165 4950 3185
rect 4900 3150 4950 3165
rect 5050 3435 5100 3450
rect 5050 3415 5065 3435
rect 5085 3415 5100 3435
rect 5050 3385 5100 3415
rect 5050 3365 5065 3385
rect 5085 3365 5100 3385
rect 5050 3335 5100 3365
rect 5050 3315 5065 3335
rect 5085 3315 5100 3335
rect 5050 3285 5100 3315
rect 5050 3265 5065 3285
rect 5085 3265 5100 3285
rect 5050 3235 5100 3265
rect 5050 3215 5065 3235
rect 5085 3215 5100 3235
rect 5050 3185 5100 3215
rect 5050 3165 5065 3185
rect 5085 3165 5100 3185
rect 4750 3115 4765 3135
rect 4785 3115 4800 3135
rect 4750 3100 4800 3115
rect 5050 3135 5100 3165
rect 5200 3435 5250 3465
rect 5500 3485 5550 3500
rect 5500 3465 5515 3485
rect 5535 3465 5550 3485
rect 5200 3415 5215 3435
rect 5235 3415 5250 3435
rect 5200 3385 5250 3415
rect 5200 3365 5215 3385
rect 5235 3365 5250 3385
rect 5200 3335 5250 3365
rect 5200 3315 5215 3335
rect 5235 3315 5250 3335
rect 5200 3285 5250 3315
rect 5200 3265 5215 3285
rect 5235 3265 5250 3285
rect 5200 3235 5250 3265
rect 5200 3215 5215 3235
rect 5235 3215 5250 3235
rect 5200 3185 5250 3215
rect 5200 3165 5215 3185
rect 5235 3165 5250 3185
rect 5200 3150 5250 3165
rect 5350 3435 5400 3450
rect 5350 3415 5365 3435
rect 5385 3415 5400 3435
rect 5350 3385 5400 3415
rect 5350 3365 5365 3385
rect 5385 3365 5400 3385
rect 5350 3335 5400 3365
rect 5350 3315 5365 3335
rect 5385 3315 5400 3335
rect 5350 3285 5400 3315
rect 5350 3265 5365 3285
rect 5385 3265 5400 3285
rect 5350 3235 5400 3265
rect 5350 3215 5365 3235
rect 5385 3215 5400 3235
rect 5350 3185 5400 3215
rect 5350 3165 5365 3185
rect 5385 3165 5400 3185
rect 5050 3115 5065 3135
rect 5085 3115 5100 3135
rect 5050 3100 5100 3115
rect 5350 3135 5400 3165
rect 5500 3435 5550 3465
rect 5800 3485 5850 3500
rect 5800 3465 5815 3485
rect 5835 3465 5850 3485
rect 5500 3415 5515 3435
rect 5535 3415 5550 3435
rect 5500 3385 5550 3415
rect 5500 3365 5515 3385
rect 5535 3365 5550 3385
rect 5500 3335 5550 3365
rect 5500 3315 5515 3335
rect 5535 3315 5550 3335
rect 5500 3285 5550 3315
rect 5500 3265 5515 3285
rect 5535 3265 5550 3285
rect 5500 3235 5550 3265
rect 5500 3215 5515 3235
rect 5535 3215 5550 3235
rect 5500 3185 5550 3215
rect 5500 3165 5515 3185
rect 5535 3165 5550 3185
rect 5500 3150 5550 3165
rect 5650 3435 5700 3450
rect 5650 3415 5665 3435
rect 5685 3415 5700 3435
rect 5650 3385 5700 3415
rect 5650 3365 5665 3385
rect 5685 3365 5700 3385
rect 5650 3335 5700 3365
rect 5650 3315 5665 3335
rect 5685 3315 5700 3335
rect 5650 3285 5700 3315
rect 5650 3265 5665 3285
rect 5685 3265 5700 3285
rect 5650 3235 5700 3265
rect 5650 3215 5665 3235
rect 5685 3215 5700 3235
rect 5650 3185 5700 3215
rect 5650 3165 5665 3185
rect 5685 3165 5700 3185
rect 5350 3115 5365 3135
rect 5385 3115 5400 3135
rect 5350 3100 5400 3115
rect 5650 3135 5700 3165
rect 5800 3435 5850 3465
rect 5800 3415 5815 3435
rect 5835 3415 5850 3435
rect 5800 3385 5850 3415
rect 5800 3365 5815 3385
rect 5835 3365 5850 3385
rect 5800 3335 5850 3365
rect 5800 3315 5815 3335
rect 5835 3315 5850 3335
rect 5800 3285 5850 3315
rect 5800 3265 5815 3285
rect 5835 3265 5850 3285
rect 5800 3235 5850 3265
rect 5800 3215 5815 3235
rect 5835 3215 5850 3235
rect 5800 3185 5850 3215
rect 5800 3165 5815 3185
rect 5835 3165 5850 3185
rect 5800 3150 5850 3165
rect 5950 3535 6000 3715
rect 6100 4085 6150 4100
rect 6100 4065 6115 4085
rect 6135 4065 6150 4085
rect 6100 4035 6150 4065
rect 6100 4015 6115 4035
rect 6135 4015 6150 4035
rect 6100 3985 6150 4015
rect 6100 3965 6115 3985
rect 6135 3965 6150 3985
rect 6100 3935 6150 3965
rect 6100 3915 6115 3935
rect 6135 3915 6150 3935
rect 6100 3885 6150 3915
rect 6100 3865 6115 3885
rect 6135 3865 6150 3885
rect 6100 3835 6150 3865
rect 6100 3815 6115 3835
rect 6135 3815 6150 3835
rect 6100 3785 6150 3815
rect 6250 4085 6300 4115
rect 6550 4135 6600 4150
rect 6550 4115 6565 4135
rect 6585 4115 6600 4135
rect 6250 4065 6265 4085
rect 6285 4065 6300 4085
rect 6250 4035 6300 4065
rect 6250 4015 6265 4035
rect 6285 4015 6300 4035
rect 6250 3985 6300 4015
rect 6250 3965 6265 3985
rect 6285 3965 6300 3985
rect 6250 3935 6300 3965
rect 6250 3915 6265 3935
rect 6285 3915 6300 3935
rect 6250 3885 6300 3915
rect 6250 3865 6265 3885
rect 6285 3865 6300 3885
rect 6250 3835 6300 3865
rect 6250 3815 6265 3835
rect 6285 3815 6300 3835
rect 6250 3800 6300 3815
rect 6400 4085 6450 4100
rect 6400 4065 6415 4085
rect 6435 4065 6450 4085
rect 6400 4035 6450 4065
rect 6400 4015 6415 4035
rect 6435 4015 6450 4035
rect 6400 3985 6450 4015
rect 6400 3965 6415 3985
rect 6435 3965 6450 3985
rect 6400 3935 6450 3965
rect 6400 3915 6415 3935
rect 6435 3915 6450 3935
rect 6400 3885 6450 3915
rect 6400 3865 6415 3885
rect 6435 3865 6450 3885
rect 6400 3835 6450 3865
rect 6400 3815 6415 3835
rect 6435 3815 6450 3835
rect 6100 3765 6115 3785
rect 6135 3765 6150 3785
rect 6100 3750 6150 3765
rect 6400 3785 6450 3815
rect 6400 3765 6415 3785
rect 6435 3765 6450 3785
rect 6400 3750 6450 3765
rect 6100 3735 6450 3750
rect 6100 3715 6115 3735
rect 6135 3715 6415 3735
rect 6435 3715 6450 3735
rect 6100 3700 6450 3715
rect 6550 4085 6600 4115
rect 6850 4135 6900 4150
rect 6850 4115 6865 4135
rect 6885 4115 6900 4135
rect 6550 4065 6565 4085
rect 6585 4065 6600 4085
rect 6550 4035 6600 4065
rect 6550 4015 6565 4035
rect 6585 4015 6600 4035
rect 6550 3985 6600 4015
rect 6550 3965 6565 3985
rect 6585 3965 6600 3985
rect 6550 3935 6600 3965
rect 6550 3915 6565 3935
rect 6585 3915 6600 3935
rect 6550 3885 6600 3915
rect 6550 3865 6565 3885
rect 6585 3865 6600 3885
rect 6550 3835 6600 3865
rect 6550 3815 6565 3835
rect 6585 3815 6600 3835
rect 6550 3785 6600 3815
rect 6550 3765 6565 3785
rect 6585 3765 6600 3785
rect 6550 3735 6600 3765
rect 6550 3715 6565 3735
rect 6585 3715 6600 3735
rect 6100 3640 6150 3650
rect 6100 3610 6110 3640
rect 6140 3610 6150 3640
rect 6100 3600 6150 3610
rect 6250 3640 6300 3700
rect 6250 3610 6260 3640
rect 6290 3610 6300 3640
rect 6250 3550 6300 3610
rect 6400 3640 6450 3650
rect 6400 3610 6410 3640
rect 6440 3610 6450 3640
rect 6400 3600 6450 3610
rect 5950 3515 5965 3535
rect 5985 3515 6000 3535
rect 5950 3485 6000 3515
rect 5950 3465 5965 3485
rect 5985 3465 6000 3485
rect 5950 3435 6000 3465
rect 5950 3415 5965 3435
rect 5985 3415 6000 3435
rect 5950 3385 6000 3415
rect 5950 3365 5965 3385
rect 5985 3365 6000 3385
rect 5950 3335 6000 3365
rect 5950 3315 5965 3335
rect 5985 3315 6000 3335
rect 5950 3285 6000 3315
rect 5950 3265 5965 3285
rect 5985 3265 6000 3285
rect 5950 3235 6000 3265
rect 5950 3215 5965 3235
rect 5985 3215 6000 3235
rect 5950 3185 6000 3215
rect 5950 3165 5965 3185
rect 5985 3165 6000 3185
rect 5650 3115 5665 3135
rect 5685 3115 5700 3135
rect 5650 3100 5700 3115
rect 5950 3135 6000 3165
rect 6100 3535 6450 3550
rect 6100 3515 6115 3535
rect 6135 3515 6415 3535
rect 6435 3515 6450 3535
rect 6100 3500 6450 3515
rect 6100 3485 6150 3500
rect 6100 3465 6115 3485
rect 6135 3465 6150 3485
rect 6100 3435 6150 3465
rect 6400 3485 6450 3500
rect 6400 3465 6415 3485
rect 6435 3465 6450 3485
rect 6100 3415 6115 3435
rect 6135 3415 6150 3435
rect 6100 3385 6150 3415
rect 6100 3365 6115 3385
rect 6135 3365 6150 3385
rect 6100 3335 6150 3365
rect 6100 3315 6115 3335
rect 6135 3315 6150 3335
rect 6100 3285 6150 3315
rect 6100 3265 6115 3285
rect 6135 3265 6150 3285
rect 6100 3235 6150 3265
rect 6100 3215 6115 3235
rect 6135 3215 6150 3235
rect 6100 3185 6150 3215
rect 6100 3165 6115 3185
rect 6135 3165 6150 3185
rect 6100 3150 6150 3165
rect 6250 3435 6300 3450
rect 6250 3415 6265 3435
rect 6285 3415 6300 3435
rect 6250 3385 6300 3415
rect 6250 3365 6265 3385
rect 6285 3365 6300 3385
rect 6250 3335 6300 3365
rect 6250 3315 6265 3335
rect 6285 3315 6300 3335
rect 6250 3285 6300 3315
rect 6250 3265 6265 3285
rect 6285 3265 6300 3285
rect 6250 3235 6300 3265
rect 6250 3215 6265 3235
rect 6285 3215 6300 3235
rect 6250 3185 6300 3215
rect 6250 3165 6265 3185
rect 6285 3165 6300 3185
rect 5950 3115 5965 3135
rect 5985 3115 6000 3135
rect 5950 3100 6000 3115
rect 6250 3135 6300 3165
rect 6400 3435 6450 3465
rect 6400 3415 6415 3435
rect 6435 3415 6450 3435
rect 6400 3385 6450 3415
rect 6400 3365 6415 3385
rect 6435 3365 6450 3385
rect 6400 3335 6450 3365
rect 6400 3315 6415 3335
rect 6435 3315 6450 3335
rect 6400 3285 6450 3315
rect 6400 3265 6415 3285
rect 6435 3265 6450 3285
rect 6400 3235 6450 3265
rect 6400 3215 6415 3235
rect 6435 3215 6450 3235
rect 6400 3185 6450 3215
rect 6400 3165 6415 3185
rect 6435 3165 6450 3185
rect 6400 3150 6450 3165
rect 6550 3535 6600 3715
rect 6700 4085 6750 4100
rect 6700 4065 6715 4085
rect 6735 4065 6750 4085
rect 6700 4035 6750 4065
rect 6700 4015 6715 4035
rect 6735 4015 6750 4035
rect 6700 3985 6750 4015
rect 6700 3965 6715 3985
rect 6735 3965 6750 3985
rect 6700 3935 6750 3965
rect 6700 3915 6715 3935
rect 6735 3915 6750 3935
rect 6700 3885 6750 3915
rect 6700 3865 6715 3885
rect 6735 3865 6750 3885
rect 6700 3835 6750 3865
rect 6700 3815 6715 3835
rect 6735 3815 6750 3835
rect 6700 3785 6750 3815
rect 6850 4085 6900 4115
rect 7150 4135 7200 4150
rect 7150 4115 7165 4135
rect 7185 4115 7200 4135
rect 6850 4065 6865 4085
rect 6885 4065 6900 4085
rect 6850 4035 6900 4065
rect 6850 4015 6865 4035
rect 6885 4015 6900 4035
rect 6850 3985 6900 4015
rect 6850 3965 6865 3985
rect 6885 3965 6900 3985
rect 6850 3935 6900 3965
rect 6850 3915 6865 3935
rect 6885 3915 6900 3935
rect 6850 3885 6900 3915
rect 6850 3865 6865 3885
rect 6885 3865 6900 3885
rect 6850 3835 6900 3865
rect 6850 3815 6865 3835
rect 6885 3815 6900 3835
rect 6850 3800 6900 3815
rect 7000 4085 7050 4100
rect 7000 4065 7015 4085
rect 7035 4065 7050 4085
rect 7000 4035 7050 4065
rect 7000 4015 7015 4035
rect 7035 4015 7050 4035
rect 7000 3985 7050 4015
rect 7000 3965 7015 3985
rect 7035 3965 7050 3985
rect 7000 3935 7050 3965
rect 7000 3915 7015 3935
rect 7035 3915 7050 3935
rect 7000 3885 7050 3915
rect 7000 3865 7015 3885
rect 7035 3865 7050 3885
rect 7000 3835 7050 3865
rect 7000 3815 7015 3835
rect 7035 3815 7050 3835
rect 6700 3765 6715 3785
rect 6735 3765 6750 3785
rect 6700 3750 6750 3765
rect 7000 3785 7050 3815
rect 7150 4085 7200 4115
rect 7450 4135 7500 4150
rect 7450 4115 7465 4135
rect 7485 4115 7500 4135
rect 7150 4065 7165 4085
rect 7185 4065 7200 4085
rect 7150 4035 7200 4065
rect 7150 4015 7165 4035
rect 7185 4015 7200 4035
rect 7150 3985 7200 4015
rect 7150 3965 7165 3985
rect 7185 3965 7200 3985
rect 7150 3935 7200 3965
rect 7150 3915 7165 3935
rect 7185 3915 7200 3935
rect 7150 3885 7200 3915
rect 7150 3865 7165 3885
rect 7185 3865 7200 3885
rect 7150 3835 7200 3865
rect 7150 3815 7165 3835
rect 7185 3815 7200 3835
rect 7150 3800 7200 3815
rect 7300 4085 7350 4100
rect 7300 4065 7315 4085
rect 7335 4065 7350 4085
rect 7300 4035 7350 4065
rect 7300 4015 7315 4035
rect 7335 4015 7350 4035
rect 7300 3985 7350 4015
rect 7300 3965 7315 3985
rect 7335 3965 7350 3985
rect 7300 3935 7350 3965
rect 7300 3915 7315 3935
rect 7335 3915 7350 3935
rect 7300 3885 7350 3915
rect 7300 3865 7315 3885
rect 7335 3865 7350 3885
rect 7300 3835 7350 3865
rect 7300 3815 7315 3835
rect 7335 3815 7350 3835
rect 7000 3765 7015 3785
rect 7035 3765 7050 3785
rect 7000 3750 7050 3765
rect 7300 3785 7350 3815
rect 7450 4085 7500 4115
rect 7750 4135 7800 4150
rect 7750 4115 7765 4135
rect 7785 4115 7800 4135
rect 7450 4065 7465 4085
rect 7485 4065 7500 4085
rect 7450 4035 7500 4065
rect 7450 4015 7465 4035
rect 7485 4015 7500 4035
rect 7450 3985 7500 4015
rect 7450 3965 7465 3985
rect 7485 3965 7500 3985
rect 7450 3935 7500 3965
rect 7450 3915 7465 3935
rect 7485 3915 7500 3935
rect 7450 3885 7500 3915
rect 7450 3865 7465 3885
rect 7485 3865 7500 3885
rect 7450 3835 7500 3865
rect 7450 3815 7465 3835
rect 7485 3815 7500 3835
rect 7450 3800 7500 3815
rect 7600 4085 7650 4100
rect 7600 4065 7615 4085
rect 7635 4065 7650 4085
rect 7600 4035 7650 4065
rect 7600 4015 7615 4035
rect 7635 4015 7650 4035
rect 7600 3985 7650 4015
rect 7600 3965 7615 3985
rect 7635 3965 7650 3985
rect 7600 3935 7650 3965
rect 7600 3915 7615 3935
rect 7635 3915 7650 3935
rect 7600 3885 7650 3915
rect 7600 3865 7615 3885
rect 7635 3865 7650 3885
rect 7600 3835 7650 3865
rect 7600 3815 7615 3835
rect 7635 3815 7650 3835
rect 7300 3765 7315 3785
rect 7335 3765 7350 3785
rect 7300 3750 7350 3765
rect 7600 3785 7650 3815
rect 7600 3765 7615 3785
rect 7635 3765 7650 3785
rect 7600 3750 7650 3765
rect 6700 3735 7650 3750
rect 6700 3715 7615 3735
rect 7635 3715 7650 3735
rect 6700 3700 7650 3715
rect 7750 4085 7800 4115
rect 7750 4065 7765 4085
rect 7785 4065 7800 4085
rect 7750 4035 7800 4065
rect 7750 4015 7765 4035
rect 7785 4015 7800 4035
rect 7750 3985 7800 4015
rect 7750 3965 7765 3985
rect 7785 3965 7800 3985
rect 7750 3935 7800 3965
rect 7750 3915 7765 3935
rect 7785 3915 7800 3935
rect 7750 3885 7800 3915
rect 7750 3865 7765 3885
rect 7785 3865 7800 3885
rect 7750 3835 7800 3865
rect 7750 3815 7765 3835
rect 7785 3815 7800 3835
rect 7750 3785 7800 3815
rect 7750 3765 7765 3785
rect 7785 3765 7800 3785
rect 7750 3735 7800 3765
rect 7750 3715 7765 3735
rect 7785 3715 7800 3735
rect 6700 3640 6750 3650
rect 6700 3610 6710 3640
rect 6740 3610 6750 3640
rect 6700 3600 6750 3610
rect 7000 3640 7050 3650
rect 7000 3610 7010 3640
rect 7040 3610 7050 3640
rect 7000 3600 7050 3610
rect 7150 3640 7200 3700
rect 7150 3610 7160 3640
rect 7190 3610 7200 3640
rect 7150 3550 7200 3610
rect 7300 3640 7350 3650
rect 7300 3610 7310 3640
rect 7340 3610 7350 3640
rect 7300 3600 7350 3610
rect 7600 3640 7650 3650
rect 7600 3610 7610 3640
rect 7640 3610 7650 3640
rect 7600 3600 7650 3610
rect 6550 3515 6565 3535
rect 6585 3515 6600 3535
rect 6550 3485 6600 3515
rect 6550 3465 6565 3485
rect 6585 3465 6600 3485
rect 6550 3435 6600 3465
rect 6550 3415 6565 3435
rect 6585 3415 6600 3435
rect 6550 3385 6600 3415
rect 6550 3365 6565 3385
rect 6585 3365 6600 3385
rect 6550 3335 6600 3365
rect 6550 3315 6565 3335
rect 6585 3315 6600 3335
rect 6550 3285 6600 3315
rect 6550 3265 6565 3285
rect 6585 3265 6600 3285
rect 6550 3235 6600 3265
rect 6550 3215 6565 3235
rect 6585 3215 6600 3235
rect 6550 3185 6600 3215
rect 6550 3165 6565 3185
rect 6585 3165 6600 3185
rect 6250 3115 6265 3135
rect 6285 3115 6300 3135
rect 6250 3100 6300 3115
rect 6550 3135 6600 3165
rect 6700 3535 7650 3550
rect 6700 3515 6715 3535
rect 6735 3515 7015 3535
rect 7035 3515 7315 3535
rect 7335 3515 7615 3535
rect 7635 3515 7650 3535
rect 6700 3500 7650 3515
rect 6700 3485 6750 3500
rect 6700 3465 6715 3485
rect 6735 3465 6750 3485
rect 6700 3435 6750 3465
rect 7000 3485 7050 3500
rect 7000 3465 7015 3485
rect 7035 3465 7050 3485
rect 6700 3415 6715 3435
rect 6735 3415 6750 3435
rect 6700 3385 6750 3415
rect 6700 3365 6715 3385
rect 6735 3365 6750 3385
rect 6700 3335 6750 3365
rect 6700 3315 6715 3335
rect 6735 3315 6750 3335
rect 6700 3285 6750 3315
rect 6700 3265 6715 3285
rect 6735 3265 6750 3285
rect 6700 3235 6750 3265
rect 6700 3215 6715 3235
rect 6735 3215 6750 3235
rect 6700 3185 6750 3215
rect 6700 3165 6715 3185
rect 6735 3165 6750 3185
rect 6700 3150 6750 3165
rect 6850 3435 6900 3450
rect 6850 3415 6865 3435
rect 6885 3415 6900 3435
rect 6850 3385 6900 3415
rect 6850 3365 6865 3385
rect 6885 3365 6900 3385
rect 6850 3335 6900 3365
rect 6850 3315 6865 3335
rect 6885 3315 6900 3335
rect 6850 3285 6900 3315
rect 6850 3265 6865 3285
rect 6885 3265 6900 3285
rect 6850 3235 6900 3265
rect 6850 3215 6865 3235
rect 6885 3215 6900 3235
rect 6850 3185 6900 3215
rect 6850 3165 6865 3185
rect 6885 3165 6900 3185
rect 6550 3115 6565 3135
rect 6585 3115 6600 3135
rect 6550 3100 6600 3115
rect 6850 3135 6900 3165
rect 7000 3435 7050 3465
rect 7300 3485 7350 3500
rect 7300 3465 7315 3485
rect 7335 3465 7350 3485
rect 7000 3415 7015 3435
rect 7035 3415 7050 3435
rect 7000 3385 7050 3415
rect 7000 3365 7015 3385
rect 7035 3365 7050 3385
rect 7000 3335 7050 3365
rect 7000 3315 7015 3335
rect 7035 3315 7050 3335
rect 7000 3285 7050 3315
rect 7000 3265 7015 3285
rect 7035 3265 7050 3285
rect 7000 3235 7050 3265
rect 7000 3215 7015 3235
rect 7035 3215 7050 3235
rect 7000 3185 7050 3215
rect 7000 3165 7015 3185
rect 7035 3165 7050 3185
rect 7000 3150 7050 3165
rect 7150 3435 7200 3450
rect 7150 3415 7165 3435
rect 7185 3415 7200 3435
rect 7150 3385 7200 3415
rect 7150 3365 7165 3385
rect 7185 3365 7200 3385
rect 7150 3335 7200 3365
rect 7150 3315 7165 3335
rect 7185 3315 7200 3335
rect 7150 3285 7200 3315
rect 7150 3265 7165 3285
rect 7185 3265 7200 3285
rect 7150 3235 7200 3265
rect 7150 3215 7165 3235
rect 7185 3215 7200 3235
rect 7150 3185 7200 3215
rect 7150 3165 7165 3185
rect 7185 3165 7200 3185
rect 6850 3115 6865 3135
rect 6885 3115 6900 3135
rect 6850 3100 6900 3115
rect 7150 3135 7200 3165
rect 7300 3435 7350 3465
rect 7600 3485 7650 3500
rect 7600 3465 7615 3485
rect 7635 3465 7650 3485
rect 7300 3415 7315 3435
rect 7335 3415 7350 3435
rect 7300 3385 7350 3415
rect 7300 3365 7315 3385
rect 7335 3365 7350 3385
rect 7300 3335 7350 3365
rect 7300 3315 7315 3335
rect 7335 3315 7350 3335
rect 7300 3285 7350 3315
rect 7300 3265 7315 3285
rect 7335 3265 7350 3285
rect 7300 3235 7350 3265
rect 7300 3215 7315 3235
rect 7335 3215 7350 3235
rect 7300 3185 7350 3215
rect 7300 3165 7315 3185
rect 7335 3165 7350 3185
rect 7300 3150 7350 3165
rect 7450 3435 7500 3450
rect 7450 3415 7465 3435
rect 7485 3415 7500 3435
rect 7450 3385 7500 3415
rect 7450 3365 7465 3385
rect 7485 3365 7500 3385
rect 7450 3335 7500 3365
rect 7450 3315 7465 3335
rect 7485 3315 7500 3335
rect 7450 3285 7500 3315
rect 7450 3265 7465 3285
rect 7485 3265 7500 3285
rect 7450 3235 7500 3265
rect 7450 3215 7465 3235
rect 7485 3215 7500 3235
rect 7450 3185 7500 3215
rect 7450 3165 7465 3185
rect 7485 3165 7500 3185
rect 7150 3115 7165 3135
rect 7185 3115 7200 3135
rect 7150 3100 7200 3115
rect 7450 3135 7500 3165
rect 7600 3435 7650 3465
rect 7600 3415 7615 3435
rect 7635 3415 7650 3435
rect 7600 3385 7650 3415
rect 7600 3365 7615 3385
rect 7635 3365 7650 3385
rect 7600 3335 7650 3365
rect 7600 3315 7615 3335
rect 7635 3315 7650 3335
rect 7600 3285 7650 3315
rect 7600 3265 7615 3285
rect 7635 3265 7650 3285
rect 7600 3235 7650 3265
rect 7600 3215 7615 3235
rect 7635 3215 7650 3235
rect 7600 3185 7650 3215
rect 7600 3165 7615 3185
rect 7635 3165 7650 3185
rect 7600 3150 7650 3165
rect 7750 3535 7800 3715
rect 8350 4185 8400 4260
rect 8650 4290 8700 4365
rect 8800 4835 8850 4850
rect 8800 4815 8815 4835
rect 8835 4815 8850 4835
rect 8800 4785 8850 4815
rect 8800 4765 8815 4785
rect 8835 4765 8850 4785
rect 8800 4735 8850 4765
rect 8800 4715 8815 4735
rect 8835 4715 8850 4735
rect 8800 4685 8850 4715
rect 8800 4665 8815 4685
rect 8835 4665 8850 4685
rect 8800 4635 8850 4665
rect 8800 4615 8815 4635
rect 8835 4615 8850 4635
rect 8800 4585 8850 4615
rect 8800 4565 8815 4585
rect 8835 4565 8850 4585
rect 8800 4535 8850 4565
rect 8800 4515 8815 4535
rect 8835 4515 8850 4535
rect 8800 4485 8850 4515
rect 8800 4465 8815 4485
rect 8835 4465 8850 4485
rect 8800 4435 8850 4465
rect 8800 4415 8815 4435
rect 8835 4415 8850 4435
rect 8800 4385 8850 4415
rect 8800 4365 8815 4385
rect 8835 4365 8850 4385
rect 8800 4350 8850 4365
rect 8950 4840 9000 5010
rect 9100 5485 9150 5500
rect 9100 5465 9115 5485
rect 9135 5465 9150 5485
rect 9100 5435 9150 5465
rect 9100 5415 9115 5435
rect 9135 5415 9150 5435
rect 9100 5385 9150 5415
rect 9100 5365 9115 5385
rect 9135 5365 9150 5385
rect 9100 5335 9150 5365
rect 9100 5315 9115 5335
rect 9135 5315 9150 5335
rect 9100 5285 9150 5315
rect 9100 5265 9115 5285
rect 9135 5265 9150 5285
rect 9100 5235 9150 5265
rect 9100 5215 9115 5235
rect 9135 5215 9150 5235
rect 9100 5185 9150 5215
rect 9100 5165 9115 5185
rect 9135 5165 9150 5185
rect 9100 5135 9150 5165
rect 9100 5115 9115 5135
rect 9135 5115 9150 5135
rect 9100 5085 9150 5115
rect 9100 5065 9115 5085
rect 9135 5065 9150 5085
rect 9100 5035 9150 5065
rect 9100 5015 9115 5035
rect 9135 5015 9150 5035
rect 9100 5000 9150 5015
rect 9250 5485 9300 5560
rect 9550 5590 9600 5600
rect 9550 5560 9560 5590
rect 9590 5560 9600 5590
rect 9250 5465 9265 5485
rect 9285 5465 9300 5485
rect 9250 5440 9300 5465
rect 9250 5410 9260 5440
rect 9290 5410 9300 5440
rect 9250 5385 9300 5410
rect 9250 5365 9265 5385
rect 9285 5365 9300 5385
rect 9250 5340 9300 5365
rect 9250 5310 9260 5340
rect 9290 5310 9300 5340
rect 9250 5285 9300 5310
rect 9250 5265 9265 5285
rect 9285 5265 9300 5285
rect 9250 5240 9300 5265
rect 9250 5210 9260 5240
rect 9290 5210 9300 5240
rect 9250 5185 9300 5210
rect 9250 5165 9265 5185
rect 9285 5165 9300 5185
rect 9250 5140 9300 5165
rect 9250 5110 9260 5140
rect 9290 5110 9300 5140
rect 9250 5085 9300 5110
rect 9250 5065 9265 5085
rect 9285 5065 9300 5085
rect 9250 5040 9300 5065
rect 9250 5010 9260 5040
rect 9290 5010 9300 5040
rect 9100 4940 9150 4950
rect 9100 4910 9110 4940
rect 9140 4910 9150 4940
rect 9100 4900 9150 4910
rect 8950 4810 8960 4840
rect 8990 4810 9000 4840
rect 8950 4785 9000 4810
rect 8950 4765 8965 4785
rect 8985 4765 9000 4785
rect 8950 4740 9000 4765
rect 8950 4710 8960 4740
rect 8990 4710 9000 4740
rect 8950 4685 9000 4710
rect 8950 4665 8965 4685
rect 8985 4665 9000 4685
rect 8950 4640 9000 4665
rect 8950 4610 8960 4640
rect 8990 4610 9000 4640
rect 8950 4585 9000 4610
rect 8950 4565 8965 4585
rect 8985 4565 9000 4585
rect 8950 4540 9000 4565
rect 8950 4510 8960 4540
rect 8990 4510 9000 4540
rect 8950 4485 9000 4510
rect 8950 4465 8965 4485
rect 8985 4465 9000 4485
rect 8950 4440 9000 4465
rect 8950 4410 8960 4440
rect 8990 4410 9000 4440
rect 8950 4385 9000 4410
rect 8950 4365 8965 4385
rect 8985 4365 9000 4385
rect 8650 4260 8660 4290
rect 8690 4260 8700 4290
rect 8350 4165 8365 4185
rect 8385 4165 8400 4185
rect 8350 4140 8400 4165
rect 8350 4110 8360 4140
rect 8390 4110 8400 4140
rect 8350 4085 8400 4110
rect 8350 4065 8365 4085
rect 8385 4065 8400 4085
rect 8350 4040 8400 4065
rect 8350 4010 8360 4040
rect 8390 4010 8400 4040
rect 8350 3985 8400 4010
rect 8350 3965 8365 3985
rect 8385 3965 8400 3985
rect 8350 3940 8400 3965
rect 8350 3910 8360 3940
rect 8390 3910 8400 3940
rect 8350 3885 8400 3910
rect 8350 3865 8365 3885
rect 8385 3865 8400 3885
rect 8350 3840 8400 3865
rect 8350 3810 8360 3840
rect 8390 3810 8400 3840
rect 8350 3785 8400 3810
rect 8350 3765 8365 3785
rect 8385 3765 8400 3785
rect 8350 3740 8400 3765
rect 8350 3710 8360 3740
rect 8390 3710 8400 3740
rect 7900 3640 7950 3650
rect 7900 3610 7910 3640
rect 7940 3610 7950 3640
rect 7900 3600 7950 3610
rect 8200 3640 8250 3650
rect 8200 3610 8210 3640
rect 8240 3610 8250 3640
rect 8200 3600 8250 3610
rect 7750 3515 7765 3535
rect 7785 3515 7800 3535
rect 7750 3485 7800 3515
rect 7750 3465 7765 3485
rect 7785 3465 7800 3485
rect 7750 3435 7800 3465
rect 7750 3415 7765 3435
rect 7785 3415 7800 3435
rect 7750 3385 7800 3415
rect 7750 3365 7765 3385
rect 7785 3365 7800 3385
rect 7750 3335 7800 3365
rect 7750 3315 7765 3335
rect 7785 3315 7800 3335
rect 7750 3285 7800 3315
rect 7750 3265 7765 3285
rect 7785 3265 7800 3285
rect 7750 3235 7800 3265
rect 7750 3215 7765 3235
rect 7785 3215 7800 3235
rect 7750 3185 7800 3215
rect 7750 3165 7765 3185
rect 7785 3165 7800 3185
rect 7450 3115 7465 3135
rect 7485 3115 7500 3135
rect 7450 3100 7500 3115
rect 7750 3135 7800 3165
rect 7750 3115 7765 3135
rect 7785 3115 7800 3135
rect 7750 3100 7800 3115
rect 4750 3085 7800 3100
rect 4750 3065 4765 3085
rect 4785 3065 5065 3085
rect 5085 3065 5365 3085
rect 5385 3065 5665 3085
rect 5685 3065 5965 3085
rect 5985 3065 6265 3085
rect 6285 3065 6565 3085
rect 6585 3065 6865 3085
rect 6885 3065 7165 3085
rect 7185 3065 7465 3085
rect 7485 3065 7765 3085
rect 7785 3065 7800 3085
rect 4750 3050 7800 3065
rect 8350 3540 8400 3710
rect 8500 4185 8550 4200
rect 8500 4165 8515 4185
rect 8535 4165 8550 4185
rect 8500 4135 8550 4165
rect 8500 4115 8515 4135
rect 8535 4115 8550 4135
rect 8500 4085 8550 4115
rect 8500 4065 8515 4085
rect 8535 4065 8550 4085
rect 8500 4035 8550 4065
rect 8500 4015 8515 4035
rect 8535 4015 8550 4035
rect 8500 3985 8550 4015
rect 8500 3965 8515 3985
rect 8535 3965 8550 3985
rect 8500 3935 8550 3965
rect 8500 3915 8515 3935
rect 8535 3915 8550 3935
rect 8500 3885 8550 3915
rect 8500 3865 8515 3885
rect 8535 3865 8550 3885
rect 8500 3835 8550 3865
rect 8500 3815 8515 3835
rect 8535 3815 8550 3835
rect 8500 3785 8550 3815
rect 8500 3765 8515 3785
rect 8535 3765 8550 3785
rect 8500 3735 8550 3765
rect 8500 3715 8515 3735
rect 8535 3715 8550 3735
rect 8500 3700 8550 3715
rect 8650 4185 8700 4260
rect 8950 4290 9000 4365
rect 9100 4835 9150 4850
rect 9100 4815 9115 4835
rect 9135 4815 9150 4835
rect 9100 4785 9150 4815
rect 9100 4765 9115 4785
rect 9135 4765 9150 4785
rect 9100 4735 9150 4765
rect 9100 4715 9115 4735
rect 9135 4715 9150 4735
rect 9100 4685 9150 4715
rect 9100 4665 9115 4685
rect 9135 4665 9150 4685
rect 9100 4635 9150 4665
rect 9100 4615 9115 4635
rect 9135 4615 9150 4635
rect 9100 4585 9150 4615
rect 9100 4565 9115 4585
rect 9135 4565 9150 4585
rect 9100 4535 9150 4565
rect 9100 4515 9115 4535
rect 9135 4515 9150 4535
rect 9100 4485 9150 4515
rect 9100 4465 9115 4485
rect 9135 4465 9150 4485
rect 9100 4435 9150 4465
rect 9100 4415 9115 4435
rect 9135 4415 9150 4435
rect 9100 4385 9150 4415
rect 9100 4365 9115 4385
rect 9135 4365 9150 4385
rect 9100 4350 9150 4365
rect 9250 4840 9300 5010
rect 9400 5485 9450 5500
rect 9400 5465 9415 5485
rect 9435 5465 9450 5485
rect 9400 5435 9450 5465
rect 9400 5415 9415 5435
rect 9435 5415 9450 5435
rect 9400 5385 9450 5415
rect 9400 5365 9415 5385
rect 9435 5365 9450 5385
rect 9400 5335 9450 5365
rect 9400 5315 9415 5335
rect 9435 5315 9450 5335
rect 9400 5285 9450 5315
rect 9400 5265 9415 5285
rect 9435 5265 9450 5285
rect 9400 5235 9450 5265
rect 9400 5215 9415 5235
rect 9435 5215 9450 5235
rect 9400 5185 9450 5215
rect 9400 5165 9415 5185
rect 9435 5165 9450 5185
rect 9400 5135 9450 5165
rect 9400 5115 9415 5135
rect 9435 5115 9450 5135
rect 9400 5085 9450 5115
rect 9400 5065 9415 5085
rect 9435 5065 9450 5085
rect 9400 5035 9450 5065
rect 9400 5015 9415 5035
rect 9435 5015 9450 5035
rect 9400 5000 9450 5015
rect 9550 5485 9600 5560
rect 9850 5590 9900 5600
rect 9850 5560 9860 5590
rect 9890 5560 9900 5590
rect 9550 5465 9565 5485
rect 9585 5465 9600 5485
rect 9550 5440 9600 5465
rect 9550 5410 9560 5440
rect 9590 5410 9600 5440
rect 9550 5385 9600 5410
rect 9550 5365 9565 5385
rect 9585 5365 9600 5385
rect 9550 5340 9600 5365
rect 9550 5310 9560 5340
rect 9590 5310 9600 5340
rect 9550 5285 9600 5310
rect 9550 5265 9565 5285
rect 9585 5265 9600 5285
rect 9550 5240 9600 5265
rect 9550 5210 9560 5240
rect 9590 5210 9600 5240
rect 9550 5185 9600 5210
rect 9550 5165 9565 5185
rect 9585 5165 9600 5185
rect 9550 5140 9600 5165
rect 9550 5110 9560 5140
rect 9590 5110 9600 5140
rect 9550 5085 9600 5110
rect 9550 5065 9565 5085
rect 9585 5065 9600 5085
rect 9550 5040 9600 5065
rect 9550 5010 9560 5040
rect 9590 5010 9600 5040
rect 9400 4940 9450 4950
rect 9400 4910 9410 4940
rect 9440 4910 9450 4940
rect 9400 4900 9450 4910
rect 9250 4810 9260 4840
rect 9290 4810 9300 4840
rect 9250 4785 9300 4810
rect 9250 4765 9265 4785
rect 9285 4765 9300 4785
rect 9250 4740 9300 4765
rect 9250 4710 9260 4740
rect 9290 4710 9300 4740
rect 9250 4685 9300 4710
rect 9250 4665 9265 4685
rect 9285 4665 9300 4685
rect 9250 4640 9300 4665
rect 9250 4610 9260 4640
rect 9290 4610 9300 4640
rect 9250 4585 9300 4610
rect 9250 4565 9265 4585
rect 9285 4565 9300 4585
rect 9250 4540 9300 4565
rect 9250 4510 9260 4540
rect 9290 4510 9300 4540
rect 9250 4485 9300 4510
rect 9250 4465 9265 4485
rect 9285 4465 9300 4485
rect 9250 4440 9300 4465
rect 9250 4410 9260 4440
rect 9290 4410 9300 4440
rect 9250 4385 9300 4410
rect 9250 4365 9265 4385
rect 9285 4365 9300 4385
rect 8950 4260 8960 4290
rect 8990 4260 9000 4290
rect 8650 4165 8665 4185
rect 8685 4165 8700 4185
rect 8650 4140 8700 4165
rect 8650 4110 8660 4140
rect 8690 4110 8700 4140
rect 8650 4085 8700 4110
rect 8650 4065 8665 4085
rect 8685 4065 8700 4085
rect 8650 4040 8700 4065
rect 8650 4010 8660 4040
rect 8690 4010 8700 4040
rect 8650 3985 8700 4010
rect 8650 3965 8665 3985
rect 8685 3965 8700 3985
rect 8650 3940 8700 3965
rect 8650 3910 8660 3940
rect 8690 3910 8700 3940
rect 8650 3885 8700 3910
rect 8650 3865 8665 3885
rect 8685 3865 8700 3885
rect 8650 3840 8700 3865
rect 8650 3810 8660 3840
rect 8690 3810 8700 3840
rect 8650 3785 8700 3810
rect 8650 3765 8665 3785
rect 8685 3765 8700 3785
rect 8650 3740 8700 3765
rect 8650 3710 8660 3740
rect 8690 3710 8700 3740
rect 8500 3640 8550 3650
rect 8500 3610 8510 3640
rect 8540 3610 8550 3640
rect 8500 3600 8550 3610
rect 8350 3510 8360 3540
rect 8390 3510 8400 3540
rect 8350 3485 8400 3510
rect 8350 3465 8365 3485
rect 8385 3465 8400 3485
rect 8350 3440 8400 3465
rect 8350 3410 8360 3440
rect 8390 3410 8400 3440
rect 8350 3385 8400 3410
rect 8350 3365 8365 3385
rect 8385 3365 8400 3385
rect 8350 3340 8400 3365
rect 8350 3310 8360 3340
rect 8390 3310 8400 3340
rect 8350 3285 8400 3310
rect 8350 3265 8365 3285
rect 8385 3265 8400 3285
rect 8350 3240 8400 3265
rect 8350 3210 8360 3240
rect 8390 3210 8400 3240
rect 8350 3185 8400 3210
rect 8350 3165 8365 3185
rect 8385 3165 8400 3185
rect 8350 3140 8400 3165
rect 8350 3110 8360 3140
rect 8390 3110 8400 3140
rect 8350 3085 8400 3110
rect 8350 3065 8365 3085
rect 8385 3065 8400 3085
rect 4150 2960 4160 2990
rect 4190 2960 4200 2990
rect 4150 2950 4200 2960
rect 8350 2990 8400 3065
rect 8500 3535 8550 3550
rect 8500 3515 8515 3535
rect 8535 3515 8550 3535
rect 8500 3485 8550 3515
rect 8500 3465 8515 3485
rect 8535 3465 8550 3485
rect 8500 3435 8550 3465
rect 8500 3415 8515 3435
rect 8535 3415 8550 3435
rect 8500 3385 8550 3415
rect 8500 3365 8515 3385
rect 8535 3365 8550 3385
rect 8500 3335 8550 3365
rect 8500 3315 8515 3335
rect 8535 3315 8550 3335
rect 8500 3285 8550 3315
rect 8500 3265 8515 3285
rect 8535 3265 8550 3285
rect 8500 3235 8550 3265
rect 8500 3215 8515 3235
rect 8535 3215 8550 3235
rect 8500 3185 8550 3215
rect 8500 3165 8515 3185
rect 8535 3165 8550 3185
rect 8500 3135 8550 3165
rect 8500 3115 8515 3135
rect 8535 3115 8550 3135
rect 8500 3085 8550 3115
rect 8500 3065 8515 3085
rect 8535 3065 8550 3085
rect 8500 3050 8550 3065
rect 8650 3540 8700 3710
rect 8800 4185 8850 4200
rect 8800 4165 8815 4185
rect 8835 4165 8850 4185
rect 8800 4135 8850 4165
rect 8800 4115 8815 4135
rect 8835 4115 8850 4135
rect 8800 4085 8850 4115
rect 8800 4065 8815 4085
rect 8835 4065 8850 4085
rect 8800 4035 8850 4065
rect 8800 4015 8815 4035
rect 8835 4015 8850 4035
rect 8800 3985 8850 4015
rect 8800 3965 8815 3985
rect 8835 3965 8850 3985
rect 8800 3935 8850 3965
rect 8800 3915 8815 3935
rect 8835 3915 8850 3935
rect 8800 3885 8850 3915
rect 8800 3865 8815 3885
rect 8835 3865 8850 3885
rect 8800 3835 8850 3865
rect 8800 3815 8815 3835
rect 8835 3815 8850 3835
rect 8800 3785 8850 3815
rect 8800 3765 8815 3785
rect 8835 3765 8850 3785
rect 8800 3735 8850 3765
rect 8800 3715 8815 3735
rect 8835 3715 8850 3735
rect 8800 3700 8850 3715
rect 8950 4185 9000 4260
rect 9250 4290 9300 4365
rect 9400 4835 9450 4850
rect 9400 4815 9415 4835
rect 9435 4815 9450 4835
rect 9400 4785 9450 4815
rect 9400 4765 9415 4785
rect 9435 4765 9450 4785
rect 9400 4735 9450 4765
rect 9400 4715 9415 4735
rect 9435 4715 9450 4735
rect 9400 4685 9450 4715
rect 9400 4665 9415 4685
rect 9435 4665 9450 4685
rect 9400 4635 9450 4665
rect 9400 4615 9415 4635
rect 9435 4615 9450 4635
rect 9400 4585 9450 4615
rect 9400 4565 9415 4585
rect 9435 4565 9450 4585
rect 9400 4535 9450 4565
rect 9400 4515 9415 4535
rect 9435 4515 9450 4535
rect 9400 4485 9450 4515
rect 9400 4465 9415 4485
rect 9435 4465 9450 4485
rect 9400 4435 9450 4465
rect 9400 4415 9415 4435
rect 9435 4415 9450 4435
rect 9400 4385 9450 4415
rect 9400 4365 9415 4385
rect 9435 4365 9450 4385
rect 9400 4350 9450 4365
rect 9550 4840 9600 5010
rect 9700 5485 9750 5500
rect 9700 5465 9715 5485
rect 9735 5465 9750 5485
rect 9700 5435 9750 5465
rect 9700 5415 9715 5435
rect 9735 5415 9750 5435
rect 9700 5385 9750 5415
rect 9700 5365 9715 5385
rect 9735 5365 9750 5385
rect 9700 5335 9750 5365
rect 9700 5315 9715 5335
rect 9735 5315 9750 5335
rect 9700 5285 9750 5315
rect 9700 5265 9715 5285
rect 9735 5265 9750 5285
rect 9700 5235 9750 5265
rect 9700 5215 9715 5235
rect 9735 5215 9750 5235
rect 9700 5185 9750 5215
rect 9700 5165 9715 5185
rect 9735 5165 9750 5185
rect 9700 5135 9750 5165
rect 9700 5115 9715 5135
rect 9735 5115 9750 5135
rect 9700 5085 9750 5115
rect 9700 5065 9715 5085
rect 9735 5065 9750 5085
rect 9700 5035 9750 5065
rect 9700 5015 9715 5035
rect 9735 5015 9750 5035
rect 9700 5000 9750 5015
rect 9850 5485 9900 5560
rect 10150 5590 10200 5600
rect 10150 5560 10160 5590
rect 10190 5560 10200 5590
rect 9850 5465 9865 5485
rect 9885 5465 9900 5485
rect 9850 5440 9900 5465
rect 9850 5410 9860 5440
rect 9890 5410 9900 5440
rect 9850 5385 9900 5410
rect 9850 5365 9865 5385
rect 9885 5365 9900 5385
rect 9850 5340 9900 5365
rect 9850 5310 9860 5340
rect 9890 5310 9900 5340
rect 9850 5285 9900 5310
rect 9850 5265 9865 5285
rect 9885 5265 9900 5285
rect 9850 5240 9900 5265
rect 9850 5210 9860 5240
rect 9890 5210 9900 5240
rect 9850 5185 9900 5210
rect 9850 5165 9865 5185
rect 9885 5165 9900 5185
rect 9850 5140 9900 5165
rect 9850 5110 9860 5140
rect 9890 5110 9900 5140
rect 9850 5085 9900 5110
rect 9850 5065 9865 5085
rect 9885 5065 9900 5085
rect 9850 5040 9900 5065
rect 9850 5010 9860 5040
rect 9890 5010 9900 5040
rect 9700 4940 9750 4950
rect 9700 4910 9710 4940
rect 9740 4910 9750 4940
rect 9700 4900 9750 4910
rect 9550 4810 9560 4840
rect 9590 4810 9600 4840
rect 9550 4785 9600 4810
rect 9550 4765 9565 4785
rect 9585 4765 9600 4785
rect 9550 4740 9600 4765
rect 9550 4710 9560 4740
rect 9590 4710 9600 4740
rect 9550 4685 9600 4710
rect 9550 4665 9565 4685
rect 9585 4665 9600 4685
rect 9550 4640 9600 4665
rect 9550 4610 9560 4640
rect 9590 4610 9600 4640
rect 9550 4585 9600 4610
rect 9550 4565 9565 4585
rect 9585 4565 9600 4585
rect 9550 4540 9600 4565
rect 9550 4510 9560 4540
rect 9590 4510 9600 4540
rect 9550 4485 9600 4510
rect 9550 4465 9565 4485
rect 9585 4465 9600 4485
rect 9550 4440 9600 4465
rect 9550 4410 9560 4440
rect 9590 4410 9600 4440
rect 9550 4385 9600 4410
rect 9550 4365 9565 4385
rect 9585 4365 9600 4385
rect 9250 4260 9260 4290
rect 9290 4260 9300 4290
rect 8950 4165 8965 4185
rect 8985 4165 9000 4185
rect 8950 4140 9000 4165
rect 8950 4110 8960 4140
rect 8990 4110 9000 4140
rect 8950 4085 9000 4110
rect 8950 4065 8965 4085
rect 8985 4065 9000 4085
rect 8950 4040 9000 4065
rect 8950 4010 8960 4040
rect 8990 4010 9000 4040
rect 8950 3985 9000 4010
rect 8950 3965 8965 3985
rect 8985 3965 9000 3985
rect 8950 3940 9000 3965
rect 8950 3910 8960 3940
rect 8990 3910 9000 3940
rect 8950 3885 9000 3910
rect 8950 3865 8965 3885
rect 8985 3865 9000 3885
rect 8950 3840 9000 3865
rect 8950 3810 8960 3840
rect 8990 3810 9000 3840
rect 8950 3785 9000 3810
rect 8950 3765 8965 3785
rect 8985 3765 9000 3785
rect 8950 3740 9000 3765
rect 8950 3710 8960 3740
rect 8990 3710 9000 3740
rect 8800 3640 8850 3650
rect 8800 3610 8810 3640
rect 8840 3610 8850 3640
rect 8800 3600 8850 3610
rect 8650 3510 8660 3540
rect 8690 3510 8700 3540
rect 8650 3485 8700 3510
rect 8650 3465 8665 3485
rect 8685 3465 8700 3485
rect 8650 3440 8700 3465
rect 8650 3410 8660 3440
rect 8690 3410 8700 3440
rect 8650 3385 8700 3410
rect 8650 3365 8665 3385
rect 8685 3365 8700 3385
rect 8650 3340 8700 3365
rect 8650 3310 8660 3340
rect 8690 3310 8700 3340
rect 8650 3285 8700 3310
rect 8650 3265 8665 3285
rect 8685 3265 8700 3285
rect 8650 3240 8700 3265
rect 8650 3210 8660 3240
rect 8690 3210 8700 3240
rect 8650 3185 8700 3210
rect 8650 3165 8665 3185
rect 8685 3165 8700 3185
rect 8650 3140 8700 3165
rect 8650 3110 8660 3140
rect 8690 3110 8700 3140
rect 8650 3085 8700 3110
rect 8650 3065 8665 3085
rect 8685 3065 8700 3085
rect 8350 2960 8360 2990
rect 8390 2960 8400 2990
rect 8350 2950 8400 2960
rect 8650 2990 8700 3065
rect 8800 3535 8850 3550
rect 8800 3515 8815 3535
rect 8835 3515 8850 3535
rect 8800 3485 8850 3515
rect 8800 3465 8815 3485
rect 8835 3465 8850 3485
rect 8800 3435 8850 3465
rect 8800 3415 8815 3435
rect 8835 3415 8850 3435
rect 8800 3385 8850 3415
rect 8800 3365 8815 3385
rect 8835 3365 8850 3385
rect 8800 3335 8850 3365
rect 8800 3315 8815 3335
rect 8835 3315 8850 3335
rect 8800 3285 8850 3315
rect 8800 3265 8815 3285
rect 8835 3265 8850 3285
rect 8800 3235 8850 3265
rect 8800 3215 8815 3235
rect 8835 3215 8850 3235
rect 8800 3185 8850 3215
rect 8800 3165 8815 3185
rect 8835 3165 8850 3185
rect 8800 3135 8850 3165
rect 8800 3115 8815 3135
rect 8835 3115 8850 3135
rect 8800 3085 8850 3115
rect 8800 3065 8815 3085
rect 8835 3065 8850 3085
rect 8800 3050 8850 3065
rect 8950 3540 9000 3710
rect 9100 4185 9150 4200
rect 9100 4165 9115 4185
rect 9135 4165 9150 4185
rect 9100 4135 9150 4165
rect 9100 4115 9115 4135
rect 9135 4115 9150 4135
rect 9100 4085 9150 4115
rect 9100 4065 9115 4085
rect 9135 4065 9150 4085
rect 9100 4035 9150 4065
rect 9100 4015 9115 4035
rect 9135 4015 9150 4035
rect 9100 3985 9150 4015
rect 9100 3965 9115 3985
rect 9135 3965 9150 3985
rect 9100 3935 9150 3965
rect 9100 3915 9115 3935
rect 9135 3915 9150 3935
rect 9100 3885 9150 3915
rect 9100 3865 9115 3885
rect 9135 3865 9150 3885
rect 9100 3835 9150 3865
rect 9100 3815 9115 3835
rect 9135 3815 9150 3835
rect 9100 3785 9150 3815
rect 9100 3765 9115 3785
rect 9135 3765 9150 3785
rect 9100 3735 9150 3765
rect 9100 3715 9115 3735
rect 9135 3715 9150 3735
rect 9100 3700 9150 3715
rect 9250 4185 9300 4260
rect 9550 4290 9600 4365
rect 9700 4835 9750 4850
rect 9700 4815 9715 4835
rect 9735 4815 9750 4835
rect 9700 4785 9750 4815
rect 9700 4765 9715 4785
rect 9735 4765 9750 4785
rect 9700 4735 9750 4765
rect 9700 4715 9715 4735
rect 9735 4715 9750 4735
rect 9700 4685 9750 4715
rect 9700 4665 9715 4685
rect 9735 4665 9750 4685
rect 9700 4635 9750 4665
rect 9700 4615 9715 4635
rect 9735 4615 9750 4635
rect 9700 4585 9750 4615
rect 9700 4565 9715 4585
rect 9735 4565 9750 4585
rect 9700 4535 9750 4565
rect 9700 4515 9715 4535
rect 9735 4515 9750 4535
rect 9700 4485 9750 4515
rect 9700 4465 9715 4485
rect 9735 4465 9750 4485
rect 9700 4435 9750 4465
rect 9700 4415 9715 4435
rect 9735 4415 9750 4435
rect 9700 4385 9750 4415
rect 9700 4365 9715 4385
rect 9735 4365 9750 4385
rect 9700 4350 9750 4365
rect 9850 4840 9900 5010
rect 10000 5485 10050 5500
rect 10000 5465 10015 5485
rect 10035 5465 10050 5485
rect 10000 5435 10050 5465
rect 10000 5415 10015 5435
rect 10035 5415 10050 5435
rect 10000 5385 10050 5415
rect 10000 5365 10015 5385
rect 10035 5365 10050 5385
rect 10000 5335 10050 5365
rect 10000 5315 10015 5335
rect 10035 5315 10050 5335
rect 10000 5285 10050 5315
rect 10000 5265 10015 5285
rect 10035 5265 10050 5285
rect 10000 5235 10050 5265
rect 10000 5215 10015 5235
rect 10035 5215 10050 5235
rect 10000 5185 10050 5215
rect 10000 5165 10015 5185
rect 10035 5165 10050 5185
rect 10000 5135 10050 5165
rect 10000 5115 10015 5135
rect 10035 5115 10050 5135
rect 10000 5085 10050 5115
rect 10000 5065 10015 5085
rect 10035 5065 10050 5085
rect 10000 5035 10050 5065
rect 10000 5015 10015 5035
rect 10035 5015 10050 5035
rect 10000 5000 10050 5015
rect 10150 5485 10200 5560
rect 10450 5590 10500 5600
rect 10450 5560 10460 5590
rect 10490 5560 10500 5590
rect 10150 5465 10165 5485
rect 10185 5465 10200 5485
rect 10150 5440 10200 5465
rect 10150 5410 10160 5440
rect 10190 5410 10200 5440
rect 10150 5385 10200 5410
rect 10150 5365 10165 5385
rect 10185 5365 10200 5385
rect 10150 5340 10200 5365
rect 10150 5310 10160 5340
rect 10190 5310 10200 5340
rect 10150 5285 10200 5310
rect 10150 5265 10165 5285
rect 10185 5265 10200 5285
rect 10150 5240 10200 5265
rect 10150 5210 10160 5240
rect 10190 5210 10200 5240
rect 10150 5185 10200 5210
rect 10150 5165 10165 5185
rect 10185 5165 10200 5185
rect 10150 5140 10200 5165
rect 10150 5110 10160 5140
rect 10190 5110 10200 5140
rect 10150 5085 10200 5110
rect 10150 5065 10165 5085
rect 10185 5065 10200 5085
rect 10150 5040 10200 5065
rect 10150 5010 10160 5040
rect 10190 5010 10200 5040
rect 10000 4940 10050 4950
rect 10000 4910 10010 4940
rect 10040 4910 10050 4940
rect 10000 4900 10050 4910
rect 9850 4810 9860 4840
rect 9890 4810 9900 4840
rect 9850 4785 9900 4810
rect 9850 4765 9865 4785
rect 9885 4765 9900 4785
rect 9850 4740 9900 4765
rect 9850 4710 9860 4740
rect 9890 4710 9900 4740
rect 9850 4685 9900 4710
rect 9850 4665 9865 4685
rect 9885 4665 9900 4685
rect 9850 4640 9900 4665
rect 9850 4610 9860 4640
rect 9890 4610 9900 4640
rect 9850 4585 9900 4610
rect 9850 4565 9865 4585
rect 9885 4565 9900 4585
rect 9850 4540 9900 4565
rect 9850 4510 9860 4540
rect 9890 4510 9900 4540
rect 9850 4485 9900 4510
rect 9850 4465 9865 4485
rect 9885 4465 9900 4485
rect 9850 4440 9900 4465
rect 9850 4410 9860 4440
rect 9890 4410 9900 4440
rect 9850 4385 9900 4410
rect 9850 4365 9865 4385
rect 9885 4365 9900 4385
rect 9550 4260 9560 4290
rect 9590 4260 9600 4290
rect 9250 4165 9265 4185
rect 9285 4165 9300 4185
rect 9250 4140 9300 4165
rect 9250 4110 9260 4140
rect 9290 4110 9300 4140
rect 9250 4085 9300 4110
rect 9250 4065 9265 4085
rect 9285 4065 9300 4085
rect 9250 4040 9300 4065
rect 9250 4010 9260 4040
rect 9290 4010 9300 4040
rect 9250 3985 9300 4010
rect 9250 3965 9265 3985
rect 9285 3965 9300 3985
rect 9250 3940 9300 3965
rect 9250 3910 9260 3940
rect 9290 3910 9300 3940
rect 9250 3885 9300 3910
rect 9250 3865 9265 3885
rect 9285 3865 9300 3885
rect 9250 3840 9300 3865
rect 9250 3810 9260 3840
rect 9290 3810 9300 3840
rect 9250 3785 9300 3810
rect 9250 3765 9265 3785
rect 9285 3765 9300 3785
rect 9250 3740 9300 3765
rect 9250 3710 9260 3740
rect 9290 3710 9300 3740
rect 9100 3640 9150 3650
rect 9100 3610 9110 3640
rect 9140 3610 9150 3640
rect 9100 3600 9150 3610
rect 8950 3510 8960 3540
rect 8990 3510 9000 3540
rect 8950 3485 9000 3510
rect 8950 3465 8965 3485
rect 8985 3465 9000 3485
rect 8950 3440 9000 3465
rect 8950 3410 8960 3440
rect 8990 3410 9000 3440
rect 8950 3385 9000 3410
rect 8950 3365 8965 3385
rect 8985 3365 9000 3385
rect 8950 3340 9000 3365
rect 8950 3310 8960 3340
rect 8990 3310 9000 3340
rect 8950 3285 9000 3310
rect 8950 3265 8965 3285
rect 8985 3265 9000 3285
rect 8950 3240 9000 3265
rect 8950 3210 8960 3240
rect 8990 3210 9000 3240
rect 8950 3185 9000 3210
rect 8950 3165 8965 3185
rect 8985 3165 9000 3185
rect 8950 3140 9000 3165
rect 8950 3110 8960 3140
rect 8990 3110 9000 3140
rect 8950 3085 9000 3110
rect 8950 3065 8965 3085
rect 8985 3065 9000 3085
rect 8650 2960 8660 2990
rect 8690 2960 8700 2990
rect 8650 2950 8700 2960
rect 8950 2990 9000 3065
rect 9100 3535 9150 3550
rect 9100 3515 9115 3535
rect 9135 3515 9150 3535
rect 9100 3485 9150 3515
rect 9100 3465 9115 3485
rect 9135 3465 9150 3485
rect 9100 3435 9150 3465
rect 9100 3415 9115 3435
rect 9135 3415 9150 3435
rect 9100 3385 9150 3415
rect 9100 3365 9115 3385
rect 9135 3365 9150 3385
rect 9100 3335 9150 3365
rect 9100 3315 9115 3335
rect 9135 3315 9150 3335
rect 9100 3285 9150 3315
rect 9100 3265 9115 3285
rect 9135 3265 9150 3285
rect 9100 3235 9150 3265
rect 9100 3215 9115 3235
rect 9135 3215 9150 3235
rect 9100 3185 9150 3215
rect 9100 3165 9115 3185
rect 9135 3165 9150 3185
rect 9100 3135 9150 3165
rect 9100 3115 9115 3135
rect 9135 3115 9150 3135
rect 9100 3085 9150 3115
rect 9100 3065 9115 3085
rect 9135 3065 9150 3085
rect 9100 3050 9150 3065
rect 9250 3540 9300 3710
rect 9400 4185 9450 4200
rect 9400 4165 9415 4185
rect 9435 4165 9450 4185
rect 9400 4135 9450 4165
rect 9400 4115 9415 4135
rect 9435 4115 9450 4135
rect 9400 4085 9450 4115
rect 9400 4065 9415 4085
rect 9435 4065 9450 4085
rect 9400 4035 9450 4065
rect 9400 4015 9415 4035
rect 9435 4015 9450 4035
rect 9400 3985 9450 4015
rect 9400 3965 9415 3985
rect 9435 3965 9450 3985
rect 9400 3935 9450 3965
rect 9400 3915 9415 3935
rect 9435 3915 9450 3935
rect 9400 3885 9450 3915
rect 9400 3865 9415 3885
rect 9435 3865 9450 3885
rect 9400 3835 9450 3865
rect 9400 3815 9415 3835
rect 9435 3815 9450 3835
rect 9400 3785 9450 3815
rect 9400 3765 9415 3785
rect 9435 3765 9450 3785
rect 9400 3735 9450 3765
rect 9400 3715 9415 3735
rect 9435 3715 9450 3735
rect 9400 3700 9450 3715
rect 9550 4185 9600 4260
rect 9850 4290 9900 4365
rect 10000 4835 10050 4850
rect 10000 4815 10015 4835
rect 10035 4815 10050 4835
rect 10000 4785 10050 4815
rect 10000 4765 10015 4785
rect 10035 4765 10050 4785
rect 10000 4735 10050 4765
rect 10000 4715 10015 4735
rect 10035 4715 10050 4735
rect 10000 4685 10050 4715
rect 10000 4665 10015 4685
rect 10035 4665 10050 4685
rect 10000 4635 10050 4665
rect 10000 4615 10015 4635
rect 10035 4615 10050 4635
rect 10000 4585 10050 4615
rect 10000 4565 10015 4585
rect 10035 4565 10050 4585
rect 10000 4535 10050 4565
rect 10000 4515 10015 4535
rect 10035 4515 10050 4535
rect 10000 4485 10050 4515
rect 10000 4465 10015 4485
rect 10035 4465 10050 4485
rect 10000 4435 10050 4465
rect 10000 4415 10015 4435
rect 10035 4415 10050 4435
rect 10000 4385 10050 4415
rect 10000 4365 10015 4385
rect 10035 4365 10050 4385
rect 10000 4350 10050 4365
rect 10150 4840 10200 5010
rect 10300 5485 10350 5500
rect 10300 5465 10315 5485
rect 10335 5465 10350 5485
rect 10300 5435 10350 5465
rect 10300 5415 10315 5435
rect 10335 5415 10350 5435
rect 10300 5385 10350 5415
rect 10300 5365 10315 5385
rect 10335 5365 10350 5385
rect 10300 5335 10350 5365
rect 10300 5315 10315 5335
rect 10335 5315 10350 5335
rect 10300 5285 10350 5315
rect 10300 5265 10315 5285
rect 10335 5265 10350 5285
rect 10300 5235 10350 5265
rect 10300 5215 10315 5235
rect 10335 5215 10350 5235
rect 10300 5185 10350 5215
rect 10300 5165 10315 5185
rect 10335 5165 10350 5185
rect 10300 5135 10350 5165
rect 10300 5115 10315 5135
rect 10335 5115 10350 5135
rect 10300 5085 10350 5115
rect 10300 5065 10315 5085
rect 10335 5065 10350 5085
rect 10300 5035 10350 5065
rect 10300 5015 10315 5035
rect 10335 5015 10350 5035
rect 10300 5000 10350 5015
rect 10450 5485 10500 5560
rect 10750 5590 10800 5600
rect 10750 5560 10760 5590
rect 10790 5560 10800 5590
rect 10450 5465 10465 5485
rect 10485 5465 10500 5485
rect 10450 5440 10500 5465
rect 10450 5410 10460 5440
rect 10490 5410 10500 5440
rect 10450 5385 10500 5410
rect 10450 5365 10465 5385
rect 10485 5365 10500 5385
rect 10450 5340 10500 5365
rect 10450 5310 10460 5340
rect 10490 5310 10500 5340
rect 10450 5285 10500 5310
rect 10450 5265 10465 5285
rect 10485 5265 10500 5285
rect 10450 5240 10500 5265
rect 10450 5210 10460 5240
rect 10490 5210 10500 5240
rect 10450 5185 10500 5210
rect 10450 5165 10465 5185
rect 10485 5165 10500 5185
rect 10450 5140 10500 5165
rect 10450 5110 10460 5140
rect 10490 5110 10500 5140
rect 10450 5085 10500 5110
rect 10450 5065 10465 5085
rect 10485 5065 10500 5085
rect 10450 5040 10500 5065
rect 10450 5010 10460 5040
rect 10490 5010 10500 5040
rect 10300 4940 10350 4950
rect 10300 4910 10310 4940
rect 10340 4910 10350 4940
rect 10300 4900 10350 4910
rect 10150 4810 10160 4840
rect 10190 4810 10200 4840
rect 10150 4785 10200 4810
rect 10150 4765 10165 4785
rect 10185 4765 10200 4785
rect 10150 4740 10200 4765
rect 10150 4710 10160 4740
rect 10190 4710 10200 4740
rect 10150 4685 10200 4710
rect 10150 4665 10165 4685
rect 10185 4665 10200 4685
rect 10150 4640 10200 4665
rect 10150 4610 10160 4640
rect 10190 4610 10200 4640
rect 10150 4585 10200 4610
rect 10150 4565 10165 4585
rect 10185 4565 10200 4585
rect 10150 4540 10200 4565
rect 10150 4510 10160 4540
rect 10190 4510 10200 4540
rect 10150 4485 10200 4510
rect 10150 4465 10165 4485
rect 10185 4465 10200 4485
rect 10150 4440 10200 4465
rect 10150 4410 10160 4440
rect 10190 4410 10200 4440
rect 10150 4385 10200 4410
rect 10150 4365 10165 4385
rect 10185 4365 10200 4385
rect 9850 4260 9860 4290
rect 9890 4260 9900 4290
rect 9550 4165 9565 4185
rect 9585 4165 9600 4185
rect 9550 4140 9600 4165
rect 9550 4110 9560 4140
rect 9590 4110 9600 4140
rect 9550 4085 9600 4110
rect 9550 4065 9565 4085
rect 9585 4065 9600 4085
rect 9550 4040 9600 4065
rect 9550 4010 9560 4040
rect 9590 4010 9600 4040
rect 9550 3985 9600 4010
rect 9550 3965 9565 3985
rect 9585 3965 9600 3985
rect 9550 3940 9600 3965
rect 9550 3910 9560 3940
rect 9590 3910 9600 3940
rect 9550 3885 9600 3910
rect 9550 3865 9565 3885
rect 9585 3865 9600 3885
rect 9550 3840 9600 3865
rect 9550 3810 9560 3840
rect 9590 3810 9600 3840
rect 9550 3785 9600 3810
rect 9550 3765 9565 3785
rect 9585 3765 9600 3785
rect 9550 3740 9600 3765
rect 9550 3710 9560 3740
rect 9590 3710 9600 3740
rect 9400 3640 9450 3650
rect 9400 3610 9410 3640
rect 9440 3610 9450 3640
rect 9400 3600 9450 3610
rect 9250 3510 9260 3540
rect 9290 3510 9300 3540
rect 9250 3485 9300 3510
rect 9250 3465 9265 3485
rect 9285 3465 9300 3485
rect 9250 3440 9300 3465
rect 9250 3410 9260 3440
rect 9290 3410 9300 3440
rect 9250 3385 9300 3410
rect 9250 3365 9265 3385
rect 9285 3365 9300 3385
rect 9250 3340 9300 3365
rect 9250 3310 9260 3340
rect 9290 3310 9300 3340
rect 9250 3285 9300 3310
rect 9250 3265 9265 3285
rect 9285 3265 9300 3285
rect 9250 3240 9300 3265
rect 9250 3210 9260 3240
rect 9290 3210 9300 3240
rect 9250 3185 9300 3210
rect 9250 3165 9265 3185
rect 9285 3165 9300 3185
rect 9250 3140 9300 3165
rect 9250 3110 9260 3140
rect 9290 3110 9300 3140
rect 9250 3085 9300 3110
rect 9250 3065 9265 3085
rect 9285 3065 9300 3085
rect 8950 2960 8960 2990
rect 8990 2960 9000 2990
rect 8950 2950 9000 2960
rect 9250 2990 9300 3065
rect 9400 3535 9450 3550
rect 9400 3515 9415 3535
rect 9435 3515 9450 3535
rect 9400 3485 9450 3515
rect 9400 3465 9415 3485
rect 9435 3465 9450 3485
rect 9400 3435 9450 3465
rect 9400 3415 9415 3435
rect 9435 3415 9450 3435
rect 9400 3385 9450 3415
rect 9400 3365 9415 3385
rect 9435 3365 9450 3385
rect 9400 3335 9450 3365
rect 9400 3315 9415 3335
rect 9435 3315 9450 3335
rect 9400 3285 9450 3315
rect 9400 3265 9415 3285
rect 9435 3265 9450 3285
rect 9400 3235 9450 3265
rect 9400 3215 9415 3235
rect 9435 3215 9450 3235
rect 9400 3185 9450 3215
rect 9400 3165 9415 3185
rect 9435 3165 9450 3185
rect 9400 3135 9450 3165
rect 9400 3115 9415 3135
rect 9435 3115 9450 3135
rect 9400 3085 9450 3115
rect 9400 3065 9415 3085
rect 9435 3065 9450 3085
rect 9400 3050 9450 3065
rect 9550 3540 9600 3710
rect 9700 4185 9750 4200
rect 9700 4165 9715 4185
rect 9735 4165 9750 4185
rect 9700 4135 9750 4165
rect 9700 4115 9715 4135
rect 9735 4115 9750 4135
rect 9700 4085 9750 4115
rect 9700 4065 9715 4085
rect 9735 4065 9750 4085
rect 9700 4035 9750 4065
rect 9700 4015 9715 4035
rect 9735 4015 9750 4035
rect 9700 3985 9750 4015
rect 9700 3965 9715 3985
rect 9735 3965 9750 3985
rect 9700 3935 9750 3965
rect 9700 3915 9715 3935
rect 9735 3915 9750 3935
rect 9700 3885 9750 3915
rect 9700 3865 9715 3885
rect 9735 3865 9750 3885
rect 9700 3835 9750 3865
rect 9700 3815 9715 3835
rect 9735 3815 9750 3835
rect 9700 3785 9750 3815
rect 9700 3765 9715 3785
rect 9735 3765 9750 3785
rect 9700 3735 9750 3765
rect 9700 3715 9715 3735
rect 9735 3715 9750 3735
rect 9700 3700 9750 3715
rect 9850 4185 9900 4260
rect 10150 4290 10200 4365
rect 10300 4835 10350 4850
rect 10300 4815 10315 4835
rect 10335 4815 10350 4835
rect 10300 4785 10350 4815
rect 10300 4765 10315 4785
rect 10335 4765 10350 4785
rect 10300 4735 10350 4765
rect 10300 4715 10315 4735
rect 10335 4715 10350 4735
rect 10300 4685 10350 4715
rect 10300 4665 10315 4685
rect 10335 4665 10350 4685
rect 10300 4635 10350 4665
rect 10300 4615 10315 4635
rect 10335 4615 10350 4635
rect 10300 4585 10350 4615
rect 10300 4565 10315 4585
rect 10335 4565 10350 4585
rect 10300 4535 10350 4565
rect 10300 4515 10315 4535
rect 10335 4515 10350 4535
rect 10300 4485 10350 4515
rect 10300 4465 10315 4485
rect 10335 4465 10350 4485
rect 10300 4435 10350 4465
rect 10300 4415 10315 4435
rect 10335 4415 10350 4435
rect 10300 4385 10350 4415
rect 10300 4365 10315 4385
rect 10335 4365 10350 4385
rect 10300 4350 10350 4365
rect 10450 4840 10500 5010
rect 10600 5485 10650 5500
rect 10600 5465 10615 5485
rect 10635 5465 10650 5485
rect 10600 5435 10650 5465
rect 10600 5415 10615 5435
rect 10635 5415 10650 5435
rect 10600 5385 10650 5415
rect 10600 5365 10615 5385
rect 10635 5365 10650 5385
rect 10600 5335 10650 5365
rect 10600 5315 10615 5335
rect 10635 5315 10650 5335
rect 10600 5285 10650 5315
rect 10600 5265 10615 5285
rect 10635 5265 10650 5285
rect 10600 5235 10650 5265
rect 10600 5215 10615 5235
rect 10635 5215 10650 5235
rect 10600 5185 10650 5215
rect 10600 5165 10615 5185
rect 10635 5165 10650 5185
rect 10600 5135 10650 5165
rect 10600 5115 10615 5135
rect 10635 5115 10650 5135
rect 10600 5085 10650 5115
rect 10600 5065 10615 5085
rect 10635 5065 10650 5085
rect 10600 5035 10650 5065
rect 10600 5015 10615 5035
rect 10635 5015 10650 5035
rect 10600 5000 10650 5015
rect 10750 5485 10800 5560
rect 11950 5590 12000 5600
rect 11950 5560 11960 5590
rect 11990 5560 12000 5590
rect 10750 5465 10765 5485
rect 10785 5465 10800 5485
rect 10750 5440 10800 5465
rect 10750 5410 10760 5440
rect 10790 5410 10800 5440
rect 10750 5385 10800 5410
rect 10750 5365 10765 5385
rect 10785 5365 10800 5385
rect 10750 5340 10800 5365
rect 10750 5310 10760 5340
rect 10790 5310 10800 5340
rect 10750 5285 10800 5310
rect 10750 5265 10765 5285
rect 10785 5265 10800 5285
rect 10750 5240 10800 5265
rect 10750 5210 10760 5240
rect 10790 5210 10800 5240
rect 10750 5185 10800 5210
rect 10750 5165 10765 5185
rect 10785 5165 10800 5185
rect 10750 5140 10800 5165
rect 10750 5110 10760 5140
rect 10790 5110 10800 5140
rect 10750 5085 10800 5110
rect 10750 5065 10765 5085
rect 10785 5065 10800 5085
rect 10750 5040 10800 5065
rect 10750 5010 10760 5040
rect 10790 5010 10800 5040
rect 10600 4940 10650 4950
rect 10600 4910 10610 4940
rect 10640 4910 10650 4940
rect 10600 4900 10650 4910
rect 10450 4810 10460 4840
rect 10490 4810 10500 4840
rect 10450 4785 10500 4810
rect 10450 4765 10465 4785
rect 10485 4765 10500 4785
rect 10450 4740 10500 4765
rect 10450 4710 10460 4740
rect 10490 4710 10500 4740
rect 10450 4685 10500 4710
rect 10450 4665 10465 4685
rect 10485 4665 10500 4685
rect 10450 4640 10500 4665
rect 10450 4610 10460 4640
rect 10490 4610 10500 4640
rect 10450 4585 10500 4610
rect 10450 4565 10465 4585
rect 10485 4565 10500 4585
rect 10450 4540 10500 4565
rect 10450 4510 10460 4540
rect 10490 4510 10500 4540
rect 10450 4485 10500 4510
rect 10450 4465 10465 4485
rect 10485 4465 10500 4485
rect 10450 4440 10500 4465
rect 10450 4410 10460 4440
rect 10490 4410 10500 4440
rect 10450 4385 10500 4410
rect 10450 4365 10465 4385
rect 10485 4365 10500 4385
rect 10150 4260 10160 4290
rect 10190 4260 10200 4290
rect 9850 4165 9865 4185
rect 9885 4165 9900 4185
rect 9850 4140 9900 4165
rect 9850 4110 9860 4140
rect 9890 4110 9900 4140
rect 9850 4085 9900 4110
rect 9850 4065 9865 4085
rect 9885 4065 9900 4085
rect 9850 4040 9900 4065
rect 9850 4010 9860 4040
rect 9890 4010 9900 4040
rect 9850 3985 9900 4010
rect 9850 3965 9865 3985
rect 9885 3965 9900 3985
rect 9850 3940 9900 3965
rect 9850 3910 9860 3940
rect 9890 3910 9900 3940
rect 9850 3885 9900 3910
rect 9850 3865 9865 3885
rect 9885 3865 9900 3885
rect 9850 3840 9900 3865
rect 9850 3810 9860 3840
rect 9890 3810 9900 3840
rect 9850 3785 9900 3810
rect 9850 3765 9865 3785
rect 9885 3765 9900 3785
rect 9850 3740 9900 3765
rect 9850 3710 9860 3740
rect 9890 3710 9900 3740
rect 9700 3640 9750 3650
rect 9700 3610 9710 3640
rect 9740 3610 9750 3640
rect 9700 3600 9750 3610
rect 9550 3510 9560 3540
rect 9590 3510 9600 3540
rect 9550 3485 9600 3510
rect 9550 3465 9565 3485
rect 9585 3465 9600 3485
rect 9550 3440 9600 3465
rect 9550 3410 9560 3440
rect 9590 3410 9600 3440
rect 9550 3385 9600 3410
rect 9550 3365 9565 3385
rect 9585 3365 9600 3385
rect 9550 3340 9600 3365
rect 9550 3310 9560 3340
rect 9590 3310 9600 3340
rect 9550 3285 9600 3310
rect 9550 3265 9565 3285
rect 9585 3265 9600 3285
rect 9550 3240 9600 3265
rect 9550 3210 9560 3240
rect 9590 3210 9600 3240
rect 9550 3185 9600 3210
rect 9550 3165 9565 3185
rect 9585 3165 9600 3185
rect 9550 3140 9600 3165
rect 9550 3110 9560 3140
rect 9590 3110 9600 3140
rect 9550 3085 9600 3110
rect 9550 3065 9565 3085
rect 9585 3065 9600 3085
rect 9250 2960 9260 2990
rect 9290 2960 9300 2990
rect 9250 2950 9300 2960
rect 9550 2990 9600 3065
rect 9700 3535 9750 3550
rect 9700 3515 9715 3535
rect 9735 3515 9750 3535
rect 9700 3485 9750 3515
rect 9700 3465 9715 3485
rect 9735 3465 9750 3485
rect 9700 3435 9750 3465
rect 9700 3415 9715 3435
rect 9735 3415 9750 3435
rect 9700 3385 9750 3415
rect 9700 3365 9715 3385
rect 9735 3365 9750 3385
rect 9700 3335 9750 3365
rect 9700 3315 9715 3335
rect 9735 3315 9750 3335
rect 9700 3285 9750 3315
rect 9700 3265 9715 3285
rect 9735 3265 9750 3285
rect 9700 3235 9750 3265
rect 9700 3215 9715 3235
rect 9735 3215 9750 3235
rect 9700 3185 9750 3215
rect 9700 3165 9715 3185
rect 9735 3165 9750 3185
rect 9700 3135 9750 3165
rect 9700 3115 9715 3135
rect 9735 3115 9750 3135
rect 9700 3085 9750 3115
rect 9700 3065 9715 3085
rect 9735 3065 9750 3085
rect 9700 3050 9750 3065
rect 9850 3540 9900 3710
rect 10000 4185 10050 4200
rect 10000 4165 10015 4185
rect 10035 4165 10050 4185
rect 10000 4135 10050 4165
rect 10000 4115 10015 4135
rect 10035 4115 10050 4135
rect 10000 4085 10050 4115
rect 10000 4065 10015 4085
rect 10035 4065 10050 4085
rect 10000 4035 10050 4065
rect 10000 4015 10015 4035
rect 10035 4015 10050 4035
rect 10000 3985 10050 4015
rect 10000 3965 10015 3985
rect 10035 3965 10050 3985
rect 10000 3935 10050 3965
rect 10000 3915 10015 3935
rect 10035 3915 10050 3935
rect 10000 3885 10050 3915
rect 10000 3865 10015 3885
rect 10035 3865 10050 3885
rect 10000 3835 10050 3865
rect 10000 3815 10015 3835
rect 10035 3815 10050 3835
rect 10000 3785 10050 3815
rect 10000 3765 10015 3785
rect 10035 3765 10050 3785
rect 10000 3735 10050 3765
rect 10000 3715 10015 3735
rect 10035 3715 10050 3735
rect 10000 3700 10050 3715
rect 10150 4185 10200 4260
rect 10450 4290 10500 4365
rect 10600 4835 10650 4850
rect 10600 4815 10615 4835
rect 10635 4815 10650 4835
rect 10600 4785 10650 4815
rect 10600 4765 10615 4785
rect 10635 4765 10650 4785
rect 10600 4735 10650 4765
rect 10600 4715 10615 4735
rect 10635 4715 10650 4735
rect 10600 4685 10650 4715
rect 10600 4665 10615 4685
rect 10635 4665 10650 4685
rect 10600 4635 10650 4665
rect 10600 4615 10615 4635
rect 10635 4615 10650 4635
rect 10600 4585 10650 4615
rect 10600 4565 10615 4585
rect 10635 4565 10650 4585
rect 10600 4535 10650 4565
rect 10600 4515 10615 4535
rect 10635 4515 10650 4535
rect 10600 4485 10650 4515
rect 10600 4465 10615 4485
rect 10635 4465 10650 4485
rect 10600 4435 10650 4465
rect 10600 4415 10615 4435
rect 10635 4415 10650 4435
rect 10600 4385 10650 4415
rect 10600 4365 10615 4385
rect 10635 4365 10650 4385
rect 10600 4350 10650 4365
rect 10750 4840 10800 5010
rect 11350 5485 11400 5500
rect 11350 5465 11365 5485
rect 11385 5465 11400 5485
rect 11350 5435 11400 5465
rect 11350 5415 11365 5435
rect 11385 5415 11400 5435
rect 11350 5385 11400 5415
rect 11350 5365 11365 5385
rect 11385 5365 11400 5385
rect 11350 5335 11400 5365
rect 11350 5315 11365 5335
rect 11385 5315 11400 5335
rect 11350 5285 11400 5315
rect 11350 5265 11365 5285
rect 11385 5265 11400 5285
rect 11350 5235 11400 5265
rect 11350 5215 11365 5235
rect 11385 5215 11400 5235
rect 11350 5185 11400 5215
rect 11350 5165 11365 5185
rect 11385 5165 11400 5185
rect 11350 5135 11400 5165
rect 11350 5115 11365 5135
rect 11385 5115 11400 5135
rect 11350 5085 11400 5115
rect 11350 5065 11365 5085
rect 11385 5065 11400 5085
rect 11350 5035 11400 5065
rect 11350 5015 11365 5035
rect 11385 5015 11400 5035
rect 10900 4940 10950 4950
rect 10900 4910 10910 4940
rect 10940 4910 10950 4940
rect 10900 4900 10950 4910
rect 11200 4940 11250 4950
rect 11200 4910 11210 4940
rect 11240 4910 11250 4940
rect 11200 4900 11250 4910
rect 11350 4940 11400 5015
rect 11950 5485 12000 5560
rect 13150 5590 13200 5600
rect 13150 5560 13160 5590
rect 13190 5560 13200 5590
rect 11950 5465 11965 5485
rect 11985 5465 12000 5485
rect 11950 5440 12000 5465
rect 11950 5410 11960 5440
rect 11990 5410 12000 5440
rect 11950 5385 12000 5410
rect 11950 5365 11965 5385
rect 11985 5365 12000 5385
rect 11950 5340 12000 5365
rect 11950 5310 11960 5340
rect 11990 5310 12000 5340
rect 11950 5285 12000 5310
rect 11950 5265 11965 5285
rect 11985 5265 12000 5285
rect 11950 5240 12000 5265
rect 11950 5210 11960 5240
rect 11990 5210 12000 5240
rect 11950 5185 12000 5210
rect 11950 5165 11965 5185
rect 11985 5165 12000 5185
rect 11950 5140 12000 5165
rect 11950 5110 11960 5140
rect 11990 5110 12000 5140
rect 11950 5085 12000 5110
rect 11950 5065 11965 5085
rect 11985 5065 12000 5085
rect 11950 5040 12000 5065
rect 11950 5010 11960 5040
rect 11990 5010 12000 5040
rect 11350 4910 11360 4940
rect 11390 4910 11400 4940
rect 10750 4810 10760 4840
rect 10790 4810 10800 4840
rect 10750 4785 10800 4810
rect 10750 4765 10765 4785
rect 10785 4765 10800 4785
rect 10750 4740 10800 4765
rect 10750 4710 10760 4740
rect 10790 4710 10800 4740
rect 10750 4685 10800 4710
rect 10750 4665 10765 4685
rect 10785 4665 10800 4685
rect 10750 4640 10800 4665
rect 10750 4610 10760 4640
rect 10790 4610 10800 4640
rect 10750 4585 10800 4610
rect 10750 4565 10765 4585
rect 10785 4565 10800 4585
rect 10750 4540 10800 4565
rect 10750 4510 10760 4540
rect 10790 4510 10800 4540
rect 10750 4485 10800 4510
rect 10750 4465 10765 4485
rect 10785 4465 10800 4485
rect 10750 4440 10800 4465
rect 10750 4410 10760 4440
rect 10790 4410 10800 4440
rect 10750 4385 10800 4410
rect 10750 4365 10765 4385
rect 10785 4365 10800 4385
rect 10450 4260 10460 4290
rect 10490 4260 10500 4290
rect 10150 4165 10165 4185
rect 10185 4165 10200 4185
rect 10150 4140 10200 4165
rect 10150 4110 10160 4140
rect 10190 4110 10200 4140
rect 10150 4085 10200 4110
rect 10150 4065 10165 4085
rect 10185 4065 10200 4085
rect 10150 4040 10200 4065
rect 10150 4010 10160 4040
rect 10190 4010 10200 4040
rect 10150 3985 10200 4010
rect 10150 3965 10165 3985
rect 10185 3965 10200 3985
rect 10150 3940 10200 3965
rect 10150 3910 10160 3940
rect 10190 3910 10200 3940
rect 10150 3885 10200 3910
rect 10150 3865 10165 3885
rect 10185 3865 10200 3885
rect 10150 3840 10200 3865
rect 10150 3810 10160 3840
rect 10190 3810 10200 3840
rect 10150 3785 10200 3810
rect 10150 3765 10165 3785
rect 10185 3765 10200 3785
rect 10150 3740 10200 3765
rect 10150 3710 10160 3740
rect 10190 3710 10200 3740
rect 10000 3640 10050 3650
rect 10000 3610 10010 3640
rect 10040 3610 10050 3640
rect 10000 3600 10050 3610
rect 9850 3510 9860 3540
rect 9890 3510 9900 3540
rect 9850 3485 9900 3510
rect 9850 3465 9865 3485
rect 9885 3465 9900 3485
rect 9850 3440 9900 3465
rect 9850 3410 9860 3440
rect 9890 3410 9900 3440
rect 9850 3385 9900 3410
rect 9850 3365 9865 3385
rect 9885 3365 9900 3385
rect 9850 3340 9900 3365
rect 9850 3310 9860 3340
rect 9890 3310 9900 3340
rect 9850 3285 9900 3310
rect 9850 3265 9865 3285
rect 9885 3265 9900 3285
rect 9850 3240 9900 3265
rect 9850 3210 9860 3240
rect 9890 3210 9900 3240
rect 9850 3185 9900 3210
rect 9850 3165 9865 3185
rect 9885 3165 9900 3185
rect 9850 3140 9900 3165
rect 9850 3110 9860 3140
rect 9890 3110 9900 3140
rect 9850 3085 9900 3110
rect 9850 3065 9865 3085
rect 9885 3065 9900 3085
rect 9550 2960 9560 2990
rect 9590 2960 9600 2990
rect 9550 2950 9600 2960
rect 9850 2990 9900 3065
rect 10000 3535 10050 3550
rect 10000 3515 10015 3535
rect 10035 3515 10050 3535
rect 10000 3485 10050 3515
rect 10000 3465 10015 3485
rect 10035 3465 10050 3485
rect 10000 3435 10050 3465
rect 10000 3415 10015 3435
rect 10035 3415 10050 3435
rect 10000 3385 10050 3415
rect 10000 3365 10015 3385
rect 10035 3365 10050 3385
rect 10000 3335 10050 3365
rect 10000 3315 10015 3335
rect 10035 3315 10050 3335
rect 10000 3285 10050 3315
rect 10000 3265 10015 3285
rect 10035 3265 10050 3285
rect 10000 3235 10050 3265
rect 10000 3215 10015 3235
rect 10035 3215 10050 3235
rect 10000 3185 10050 3215
rect 10000 3165 10015 3185
rect 10035 3165 10050 3185
rect 10000 3135 10050 3165
rect 10000 3115 10015 3135
rect 10035 3115 10050 3135
rect 10000 3085 10050 3115
rect 10000 3065 10015 3085
rect 10035 3065 10050 3085
rect 10000 3050 10050 3065
rect 10150 3540 10200 3710
rect 10300 4185 10350 4200
rect 10300 4165 10315 4185
rect 10335 4165 10350 4185
rect 10300 4135 10350 4165
rect 10300 4115 10315 4135
rect 10335 4115 10350 4135
rect 10300 4085 10350 4115
rect 10300 4065 10315 4085
rect 10335 4065 10350 4085
rect 10300 4035 10350 4065
rect 10300 4015 10315 4035
rect 10335 4015 10350 4035
rect 10300 3985 10350 4015
rect 10300 3965 10315 3985
rect 10335 3965 10350 3985
rect 10300 3935 10350 3965
rect 10300 3915 10315 3935
rect 10335 3915 10350 3935
rect 10300 3885 10350 3915
rect 10300 3865 10315 3885
rect 10335 3865 10350 3885
rect 10300 3835 10350 3865
rect 10300 3815 10315 3835
rect 10335 3815 10350 3835
rect 10300 3785 10350 3815
rect 10300 3765 10315 3785
rect 10335 3765 10350 3785
rect 10300 3735 10350 3765
rect 10300 3715 10315 3735
rect 10335 3715 10350 3735
rect 10300 3700 10350 3715
rect 10450 4185 10500 4260
rect 10750 4290 10800 4365
rect 10750 4260 10760 4290
rect 10790 4260 10800 4290
rect 10450 4165 10465 4185
rect 10485 4165 10500 4185
rect 10450 4140 10500 4165
rect 10450 4110 10460 4140
rect 10490 4110 10500 4140
rect 10450 4085 10500 4110
rect 10450 4065 10465 4085
rect 10485 4065 10500 4085
rect 10450 4040 10500 4065
rect 10450 4010 10460 4040
rect 10490 4010 10500 4040
rect 10450 3985 10500 4010
rect 10450 3965 10465 3985
rect 10485 3965 10500 3985
rect 10450 3940 10500 3965
rect 10450 3910 10460 3940
rect 10490 3910 10500 3940
rect 10450 3885 10500 3910
rect 10450 3865 10465 3885
rect 10485 3865 10500 3885
rect 10450 3840 10500 3865
rect 10450 3810 10460 3840
rect 10490 3810 10500 3840
rect 10450 3785 10500 3810
rect 10450 3765 10465 3785
rect 10485 3765 10500 3785
rect 10450 3740 10500 3765
rect 10450 3710 10460 3740
rect 10490 3710 10500 3740
rect 10300 3640 10350 3650
rect 10300 3610 10310 3640
rect 10340 3610 10350 3640
rect 10300 3600 10350 3610
rect 10150 3510 10160 3540
rect 10190 3510 10200 3540
rect 10150 3485 10200 3510
rect 10150 3465 10165 3485
rect 10185 3465 10200 3485
rect 10150 3440 10200 3465
rect 10150 3410 10160 3440
rect 10190 3410 10200 3440
rect 10150 3385 10200 3410
rect 10150 3365 10165 3385
rect 10185 3365 10200 3385
rect 10150 3340 10200 3365
rect 10150 3310 10160 3340
rect 10190 3310 10200 3340
rect 10150 3285 10200 3310
rect 10150 3265 10165 3285
rect 10185 3265 10200 3285
rect 10150 3240 10200 3265
rect 10150 3210 10160 3240
rect 10190 3210 10200 3240
rect 10150 3185 10200 3210
rect 10150 3165 10165 3185
rect 10185 3165 10200 3185
rect 10150 3140 10200 3165
rect 10150 3110 10160 3140
rect 10190 3110 10200 3140
rect 10150 3085 10200 3110
rect 10150 3065 10165 3085
rect 10185 3065 10200 3085
rect 9850 2960 9860 2990
rect 9890 2960 9900 2990
rect 9850 2950 9900 2960
rect 10150 2990 10200 3065
rect 10300 3535 10350 3550
rect 10300 3515 10315 3535
rect 10335 3515 10350 3535
rect 10300 3485 10350 3515
rect 10300 3465 10315 3485
rect 10335 3465 10350 3485
rect 10300 3435 10350 3465
rect 10300 3415 10315 3435
rect 10335 3415 10350 3435
rect 10300 3385 10350 3415
rect 10300 3365 10315 3385
rect 10335 3365 10350 3385
rect 10300 3335 10350 3365
rect 10300 3315 10315 3335
rect 10335 3315 10350 3335
rect 10300 3285 10350 3315
rect 10300 3265 10315 3285
rect 10335 3265 10350 3285
rect 10300 3235 10350 3265
rect 10300 3215 10315 3235
rect 10335 3215 10350 3235
rect 10300 3185 10350 3215
rect 10300 3165 10315 3185
rect 10335 3165 10350 3185
rect 10300 3135 10350 3165
rect 10300 3115 10315 3135
rect 10335 3115 10350 3135
rect 10300 3085 10350 3115
rect 10300 3065 10315 3085
rect 10335 3065 10350 3085
rect 10300 3050 10350 3065
rect 10450 3540 10500 3710
rect 10600 4185 10650 4200
rect 10600 4165 10615 4185
rect 10635 4165 10650 4185
rect 10600 4135 10650 4165
rect 10600 4115 10615 4135
rect 10635 4115 10650 4135
rect 10600 4085 10650 4115
rect 10600 4065 10615 4085
rect 10635 4065 10650 4085
rect 10600 4035 10650 4065
rect 10600 4015 10615 4035
rect 10635 4015 10650 4035
rect 10600 3985 10650 4015
rect 10600 3965 10615 3985
rect 10635 3965 10650 3985
rect 10600 3935 10650 3965
rect 10600 3915 10615 3935
rect 10635 3915 10650 3935
rect 10600 3885 10650 3915
rect 10600 3865 10615 3885
rect 10635 3865 10650 3885
rect 10600 3835 10650 3865
rect 10600 3815 10615 3835
rect 10635 3815 10650 3835
rect 10600 3785 10650 3815
rect 10600 3765 10615 3785
rect 10635 3765 10650 3785
rect 10600 3735 10650 3765
rect 10600 3715 10615 3735
rect 10635 3715 10650 3735
rect 10600 3700 10650 3715
rect 10750 4185 10800 4260
rect 10750 4165 10765 4185
rect 10785 4165 10800 4185
rect 10750 4140 10800 4165
rect 10750 4110 10760 4140
rect 10790 4110 10800 4140
rect 10750 4085 10800 4110
rect 10750 4065 10765 4085
rect 10785 4065 10800 4085
rect 10750 4040 10800 4065
rect 10750 4010 10760 4040
rect 10790 4010 10800 4040
rect 10750 3985 10800 4010
rect 10750 3965 10765 3985
rect 10785 3965 10800 3985
rect 10750 3940 10800 3965
rect 10750 3910 10760 3940
rect 10790 3910 10800 3940
rect 10750 3885 10800 3910
rect 10750 3865 10765 3885
rect 10785 3865 10800 3885
rect 10750 3840 10800 3865
rect 10750 3810 10760 3840
rect 10790 3810 10800 3840
rect 10750 3785 10800 3810
rect 10750 3765 10765 3785
rect 10785 3765 10800 3785
rect 10750 3740 10800 3765
rect 10750 3710 10760 3740
rect 10790 3710 10800 3740
rect 10600 3640 10650 3650
rect 10600 3610 10610 3640
rect 10640 3610 10650 3640
rect 10600 3600 10650 3610
rect 10450 3510 10460 3540
rect 10490 3510 10500 3540
rect 10450 3485 10500 3510
rect 10450 3465 10465 3485
rect 10485 3465 10500 3485
rect 10450 3440 10500 3465
rect 10450 3410 10460 3440
rect 10490 3410 10500 3440
rect 10450 3385 10500 3410
rect 10450 3365 10465 3385
rect 10485 3365 10500 3385
rect 10450 3340 10500 3365
rect 10450 3310 10460 3340
rect 10490 3310 10500 3340
rect 10450 3285 10500 3310
rect 10450 3265 10465 3285
rect 10485 3265 10500 3285
rect 10450 3240 10500 3265
rect 10450 3210 10460 3240
rect 10490 3210 10500 3240
rect 10450 3185 10500 3210
rect 10450 3165 10465 3185
rect 10485 3165 10500 3185
rect 10450 3140 10500 3165
rect 10450 3110 10460 3140
rect 10490 3110 10500 3140
rect 10450 3085 10500 3110
rect 10450 3065 10465 3085
rect 10485 3065 10500 3085
rect 10150 2960 10160 2990
rect 10190 2960 10200 2990
rect 10150 2950 10200 2960
rect 10450 2990 10500 3065
rect 10600 3535 10650 3550
rect 10600 3515 10615 3535
rect 10635 3515 10650 3535
rect 10600 3485 10650 3515
rect 10600 3465 10615 3485
rect 10635 3465 10650 3485
rect 10600 3435 10650 3465
rect 10600 3415 10615 3435
rect 10635 3415 10650 3435
rect 10600 3385 10650 3415
rect 10600 3365 10615 3385
rect 10635 3365 10650 3385
rect 10600 3335 10650 3365
rect 10600 3315 10615 3335
rect 10635 3315 10650 3335
rect 10600 3285 10650 3315
rect 10600 3265 10615 3285
rect 10635 3265 10650 3285
rect 10600 3235 10650 3265
rect 10600 3215 10615 3235
rect 10635 3215 10650 3235
rect 10600 3185 10650 3215
rect 10600 3165 10615 3185
rect 10635 3165 10650 3185
rect 10600 3135 10650 3165
rect 10600 3115 10615 3135
rect 10635 3115 10650 3135
rect 10600 3085 10650 3115
rect 10600 3065 10615 3085
rect 10635 3065 10650 3085
rect 10600 3050 10650 3065
rect 10750 3540 10800 3710
rect 11350 4835 11400 4910
rect 11500 4940 11550 4950
rect 11500 4910 11510 4940
rect 11540 4910 11550 4940
rect 11500 4900 11550 4910
rect 11800 4940 11850 4950
rect 11800 4910 11810 4940
rect 11840 4910 11850 4940
rect 11800 4900 11850 4910
rect 11350 4815 11365 4835
rect 11385 4815 11400 4835
rect 11350 4785 11400 4815
rect 11350 4765 11365 4785
rect 11385 4765 11400 4785
rect 11350 4735 11400 4765
rect 11350 4715 11365 4735
rect 11385 4715 11400 4735
rect 11350 4685 11400 4715
rect 11350 4665 11365 4685
rect 11385 4665 11400 4685
rect 11350 4635 11400 4665
rect 11350 4615 11365 4635
rect 11385 4615 11400 4635
rect 11350 4585 11400 4615
rect 11350 4565 11365 4585
rect 11385 4565 11400 4585
rect 11350 4535 11400 4565
rect 11350 4515 11365 4535
rect 11385 4515 11400 4535
rect 11350 4485 11400 4515
rect 11350 4465 11365 4485
rect 11385 4465 11400 4485
rect 11350 4435 11400 4465
rect 11350 4415 11365 4435
rect 11385 4415 11400 4435
rect 11350 4385 11400 4415
rect 11350 4365 11365 4385
rect 11385 4365 11400 4385
rect 11350 4185 11400 4365
rect 11350 4165 11365 4185
rect 11385 4165 11400 4185
rect 11350 4135 11400 4165
rect 11350 4115 11365 4135
rect 11385 4115 11400 4135
rect 11350 4085 11400 4115
rect 11350 4065 11365 4085
rect 11385 4065 11400 4085
rect 11350 4035 11400 4065
rect 11350 4015 11365 4035
rect 11385 4015 11400 4035
rect 11350 3985 11400 4015
rect 11350 3965 11365 3985
rect 11385 3965 11400 3985
rect 11350 3935 11400 3965
rect 11350 3915 11365 3935
rect 11385 3915 11400 3935
rect 11350 3885 11400 3915
rect 11350 3865 11365 3885
rect 11385 3865 11400 3885
rect 11350 3835 11400 3865
rect 11350 3815 11365 3835
rect 11385 3815 11400 3835
rect 11350 3785 11400 3815
rect 11350 3765 11365 3785
rect 11385 3765 11400 3785
rect 11350 3735 11400 3765
rect 11350 3715 11365 3735
rect 11385 3715 11400 3735
rect 10900 3640 10950 3650
rect 10900 3610 10910 3640
rect 10940 3610 10950 3640
rect 10900 3600 10950 3610
rect 11200 3640 11250 3650
rect 11200 3610 11210 3640
rect 11240 3610 11250 3640
rect 11200 3600 11250 3610
rect 11350 3640 11400 3715
rect 11950 4840 12000 5010
rect 12550 5485 12600 5500
rect 12550 5465 12565 5485
rect 12585 5465 12600 5485
rect 12550 5435 12600 5465
rect 12550 5415 12565 5435
rect 12585 5415 12600 5435
rect 12550 5385 12600 5415
rect 12550 5365 12565 5385
rect 12585 5365 12600 5385
rect 12550 5335 12600 5365
rect 12550 5315 12565 5335
rect 12585 5315 12600 5335
rect 12550 5285 12600 5315
rect 12550 5265 12565 5285
rect 12585 5265 12600 5285
rect 12550 5235 12600 5265
rect 12550 5215 12565 5235
rect 12585 5215 12600 5235
rect 12550 5185 12600 5215
rect 12550 5165 12565 5185
rect 12585 5165 12600 5185
rect 12550 5135 12600 5165
rect 12550 5115 12565 5135
rect 12585 5115 12600 5135
rect 12550 5085 12600 5115
rect 12550 5065 12565 5085
rect 12585 5065 12600 5085
rect 12550 5035 12600 5065
rect 12550 5015 12565 5035
rect 12585 5015 12600 5035
rect 12100 4940 12150 4950
rect 12100 4910 12110 4940
rect 12140 4910 12150 4940
rect 12100 4900 12150 4910
rect 12400 4940 12450 4950
rect 12400 4910 12410 4940
rect 12440 4910 12450 4940
rect 12400 4900 12450 4910
rect 12550 4940 12600 5015
rect 13150 5485 13200 5560
rect 14350 5590 14400 5600
rect 14350 5560 14360 5590
rect 14390 5560 14400 5590
rect 13150 5465 13165 5485
rect 13185 5465 13200 5485
rect 13150 5440 13200 5465
rect 13150 5410 13160 5440
rect 13190 5410 13200 5440
rect 13150 5385 13200 5410
rect 13150 5365 13165 5385
rect 13185 5365 13200 5385
rect 13150 5340 13200 5365
rect 13150 5310 13160 5340
rect 13190 5310 13200 5340
rect 13150 5285 13200 5310
rect 13150 5265 13165 5285
rect 13185 5265 13200 5285
rect 13150 5240 13200 5265
rect 13150 5210 13160 5240
rect 13190 5210 13200 5240
rect 13150 5185 13200 5210
rect 13150 5165 13165 5185
rect 13185 5165 13200 5185
rect 13150 5140 13200 5165
rect 13150 5110 13160 5140
rect 13190 5110 13200 5140
rect 13150 5085 13200 5110
rect 13150 5065 13165 5085
rect 13185 5065 13200 5085
rect 13150 5040 13200 5065
rect 13150 5010 13160 5040
rect 13190 5010 13200 5040
rect 12550 4910 12560 4940
rect 12590 4910 12600 4940
rect 11950 4810 11960 4840
rect 11990 4810 12000 4840
rect 11950 4785 12000 4810
rect 11950 4765 11965 4785
rect 11985 4765 12000 4785
rect 11950 4740 12000 4765
rect 11950 4710 11960 4740
rect 11990 4710 12000 4740
rect 11950 4685 12000 4710
rect 11950 4665 11965 4685
rect 11985 4665 12000 4685
rect 11950 4640 12000 4665
rect 11950 4610 11960 4640
rect 11990 4610 12000 4640
rect 11950 4585 12000 4610
rect 11950 4565 11965 4585
rect 11985 4565 12000 4585
rect 11950 4540 12000 4565
rect 11950 4510 11960 4540
rect 11990 4510 12000 4540
rect 11950 4485 12000 4510
rect 11950 4465 11965 4485
rect 11985 4465 12000 4485
rect 11950 4440 12000 4465
rect 11950 4410 11960 4440
rect 11990 4410 12000 4440
rect 11950 4385 12000 4410
rect 11950 4365 11965 4385
rect 11985 4365 12000 4385
rect 11950 4290 12000 4365
rect 11950 4260 11960 4290
rect 11990 4260 12000 4290
rect 11950 4185 12000 4260
rect 11950 4165 11965 4185
rect 11985 4165 12000 4185
rect 11950 4140 12000 4165
rect 11950 4110 11960 4140
rect 11990 4110 12000 4140
rect 11950 4085 12000 4110
rect 11950 4065 11965 4085
rect 11985 4065 12000 4085
rect 11950 4040 12000 4065
rect 11950 4010 11960 4040
rect 11990 4010 12000 4040
rect 11950 3985 12000 4010
rect 11950 3965 11965 3985
rect 11985 3965 12000 3985
rect 11950 3940 12000 3965
rect 11950 3910 11960 3940
rect 11990 3910 12000 3940
rect 11950 3885 12000 3910
rect 11950 3865 11965 3885
rect 11985 3865 12000 3885
rect 11950 3840 12000 3865
rect 11950 3810 11960 3840
rect 11990 3810 12000 3840
rect 11950 3785 12000 3810
rect 11950 3765 11965 3785
rect 11985 3765 12000 3785
rect 11950 3740 12000 3765
rect 11950 3710 11960 3740
rect 11990 3710 12000 3740
rect 11350 3610 11360 3640
rect 11390 3610 11400 3640
rect 10750 3510 10760 3540
rect 10790 3510 10800 3540
rect 10750 3485 10800 3510
rect 10750 3465 10765 3485
rect 10785 3465 10800 3485
rect 10750 3440 10800 3465
rect 10750 3410 10760 3440
rect 10790 3410 10800 3440
rect 10750 3385 10800 3410
rect 10750 3365 10765 3385
rect 10785 3365 10800 3385
rect 10750 3340 10800 3365
rect 10750 3310 10760 3340
rect 10790 3310 10800 3340
rect 10750 3285 10800 3310
rect 10750 3265 10765 3285
rect 10785 3265 10800 3285
rect 10750 3240 10800 3265
rect 10750 3210 10760 3240
rect 10790 3210 10800 3240
rect 10750 3185 10800 3210
rect 10750 3165 10765 3185
rect 10785 3165 10800 3185
rect 10750 3140 10800 3165
rect 10750 3110 10760 3140
rect 10790 3110 10800 3140
rect 10750 3085 10800 3110
rect 10750 3065 10765 3085
rect 10785 3065 10800 3085
rect 10450 2960 10460 2990
rect 10490 2960 10500 2990
rect 10450 2950 10500 2960
rect 10750 2990 10800 3065
rect 11350 3535 11400 3610
rect 11500 3640 11550 3650
rect 11500 3610 11510 3640
rect 11540 3610 11550 3640
rect 11500 3600 11550 3610
rect 11800 3640 11850 3650
rect 11800 3610 11810 3640
rect 11840 3610 11850 3640
rect 11800 3600 11850 3610
rect 11350 3515 11365 3535
rect 11385 3515 11400 3535
rect 11350 3485 11400 3515
rect 11350 3465 11365 3485
rect 11385 3465 11400 3485
rect 11350 3435 11400 3465
rect 11350 3415 11365 3435
rect 11385 3415 11400 3435
rect 11350 3385 11400 3415
rect 11350 3365 11365 3385
rect 11385 3365 11400 3385
rect 11350 3335 11400 3365
rect 11350 3315 11365 3335
rect 11385 3315 11400 3335
rect 11350 3285 11400 3315
rect 11350 3265 11365 3285
rect 11385 3265 11400 3285
rect 11350 3235 11400 3265
rect 11350 3215 11365 3235
rect 11385 3215 11400 3235
rect 11350 3185 11400 3215
rect 11350 3165 11365 3185
rect 11385 3165 11400 3185
rect 11350 3135 11400 3165
rect 11350 3115 11365 3135
rect 11385 3115 11400 3135
rect 11350 3085 11400 3115
rect 11350 3065 11365 3085
rect 11385 3065 11400 3085
rect 11350 3050 11400 3065
rect 11950 3540 12000 3710
rect 12550 4835 12600 4910
rect 12700 4940 12750 4950
rect 12700 4910 12710 4940
rect 12740 4910 12750 4940
rect 12700 4900 12750 4910
rect 13000 4940 13050 4950
rect 13000 4910 13010 4940
rect 13040 4910 13050 4940
rect 13000 4900 13050 4910
rect 12550 4815 12565 4835
rect 12585 4815 12600 4835
rect 12550 4785 12600 4815
rect 12550 4765 12565 4785
rect 12585 4765 12600 4785
rect 12550 4735 12600 4765
rect 12550 4715 12565 4735
rect 12585 4715 12600 4735
rect 12550 4685 12600 4715
rect 12550 4665 12565 4685
rect 12585 4665 12600 4685
rect 12550 4635 12600 4665
rect 12550 4615 12565 4635
rect 12585 4615 12600 4635
rect 12550 4585 12600 4615
rect 12550 4565 12565 4585
rect 12585 4565 12600 4585
rect 12550 4535 12600 4565
rect 12550 4515 12565 4535
rect 12585 4515 12600 4535
rect 12550 4485 12600 4515
rect 12550 4465 12565 4485
rect 12585 4465 12600 4485
rect 12550 4435 12600 4465
rect 12550 4415 12565 4435
rect 12585 4415 12600 4435
rect 12550 4385 12600 4415
rect 12550 4365 12565 4385
rect 12585 4365 12600 4385
rect 12550 4185 12600 4365
rect 12550 4165 12565 4185
rect 12585 4165 12600 4185
rect 12550 4135 12600 4165
rect 12550 4115 12565 4135
rect 12585 4115 12600 4135
rect 12550 4085 12600 4115
rect 12550 4065 12565 4085
rect 12585 4065 12600 4085
rect 12550 4035 12600 4065
rect 12550 4015 12565 4035
rect 12585 4015 12600 4035
rect 12550 3985 12600 4015
rect 12550 3965 12565 3985
rect 12585 3965 12600 3985
rect 12550 3935 12600 3965
rect 12550 3915 12565 3935
rect 12585 3915 12600 3935
rect 12550 3885 12600 3915
rect 12550 3865 12565 3885
rect 12585 3865 12600 3885
rect 12550 3835 12600 3865
rect 12550 3815 12565 3835
rect 12585 3815 12600 3835
rect 12550 3785 12600 3815
rect 12550 3765 12565 3785
rect 12585 3765 12600 3785
rect 12550 3735 12600 3765
rect 12550 3715 12565 3735
rect 12585 3715 12600 3735
rect 12100 3640 12150 3650
rect 12100 3610 12110 3640
rect 12140 3610 12150 3640
rect 12100 3600 12150 3610
rect 12400 3640 12450 3650
rect 12400 3610 12410 3640
rect 12440 3610 12450 3640
rect 12400 3600 12450 3610
rect 12550 3640 12600 3715
rect 13150 4840 13200 5010
rect 13750 5485 13800 5500
rect 13750 5465 13765 5485
rect 13785 5465 13800 5485
rect 13750 5435 13800 5465
rect 13750 5415 13765 5435
rect 13785 5415 13800 5435
rect 13750 5385 13800 5415
rect 13750 5365 13765 5385
rect 13785 5365 13800 5385
rect 13750 5335 13800 5365
rect 13750 5315 13765 5335
rect 13785 5315 13800 5335
rect 13750 5285 13800 5315
rect 13750 5265 13765 5285
rect 13785 5265 13800 5285
rect 13750 5235 13800 5265
rect 13750 5215 13765 5235
rect 13785 5215 13800 5235
rect 13750 5185 13800 5215
rect 13750 5165 13765 5185
rect 13785 5165 13800 5185
rect 13750 5135 13800 5165
rect 13750 5115 13765 5135
rect 13785 5115 13800 5135
rect 13750 5085 13800 5115
rect 13750 5065 13765 5085
rect 13785 5065 13800 5085
rect 13750 5035 13800 5065
rect 13750 5015 13765 5035
rect 13785 5015 13800 5035
rect 13300 4940 13350 4950
rect 13300 4910 13310 4940
rect 13340 4910 13350 4940
rect 13300 4900 13350 4910
rect 13600 4940 13650 4950
rect 13600 4910 13610 4940
rect 13640 4910 13650 4940
rect 13600 4900 13650 4910
rect 13750 4940 13800 5015
rect 14350 5485 14400 5560
rect 15550 5590 15600 5600
rect 15550 5560 15560 5590
rect 15590 5560 15600 5590
rect 14350 5465 14365 5485
rect 14385 5465 14400 5485
rect 14350 5440 14400 5465
rect 14350 5410 14360 5440
rect 14390 5410 14400 5440
rect 14350 5385 14400 5410
rect 14350 5365 14365 5385
rect 14385 5365 14400 5385
rect 14350 5340 14400 5365
rect 14350 5310 14360 5340
rect 14390 5310 14400 5340
rect 14350 5285 14400 5310
rect 14350 5265 14365 5285
rect 14385 5265 14400 5285
rect 14350 5240 14400 5265
rect 14350 5210 14360 5240
rect 14390 5210 14400 5240
rect 14350 5185 14400 5210
rect 14350 5165 14365 5185
rect 14385 5165 14400 5185
rect 14350 5140 14400 5165
rect 14350 5110 14360 5140
rect 14390 5110 14400 5140
rect 14350 5085 14400 5110
rect 14350 5065 14365 5085
rect 14385 5065 14400 5085
rect 14350 5040 14400 5065
rect 14350 5010 14360 5040
rect 14390 5010 14400 5040
rect 13750 4910 13760 4940
rect 13790 4910 13800 4940
rect 13150 4810 13160 4840
rect 13190 4810 13200 4840
rect 13150 4785 13200 4810
rect 13150 4765 13165 4785
rect 13185 4765 13200 4785
rect 13150 4740 13200 4765
rect 13150 4710 13160 4740
rect 13190 4710 13200 4740
rect 13150 4685 13200 4710
rect 13150 4665 13165 4685
rect 13185 4665 13200 4685
rect 13150 4640 13200 4665
rect 13150 4610 13160 4640
rect 13190 4610 13200 4640
rect 13150 4585 13200 4610
rect 13150 4565 13165 4585
rect 13185 4565 13200 4585
rect 13150 4540 13200 4565
rect 13150 4510 13160 4540
rect 13190 4510 13200 4540
rect 13150 4485 13200 4510
rect 13150 4465 13165 4485
rect 13185 4465 13200 4485
rect 13150 4440 13200 4465
rect 13150 4410 13160 4440
rect 13190 4410 13200 4440
rect 13150 4385 13200 4410
rect 13150 4365 13165 4385
rect 13185 4365 13200 4385
rect 13150 4290 13200 4365
rect 13150 4260 13160 4290
rect 13190 4260 13200 4290
rect 13150 4185 13200 4260
rect 13150 4165 13165 4185
rect 13185 4165 13200 4185
rect 13150 4140 13200 4165
rect 13150 4110 13160 4140
rect 13190 4110 13200 4140
rect 13150 4085 13200 4110
rect 13150 4065 13165 4085
rect 13185 4065 13200 4085
rect 13150 4040 13200 4065
rect 13150 4010 13160 4040
rect 13190 4010 13200 4040
rect 13150 3985 13200 4010
rect 13150 3965 13165 3985
rect 13185 3965 13200 3985
rect 13150 3940 13200 3965
rect 13150 3910 13160 3940
rect 13190 3910 13200 3940
rect 13150 3885 13200 3910
rect 13150 3865 13165 3885
rect 13185 3865 13200 3885
rect 13150 3840 13200 3865
rect 13150 3810 13160 3840
rect 13190 3810 13200 3840
rect 13150 3785 13200 3810
rect 13150 3765 13165 3785
rect 13185 3765 13200 3785
rect 13150 3740 13200 3765
rect 13150 3710 13160 3740
rect 13190 3710 13200 3740
rect 12550 3610 12560 3640
rect 12590 3610 12600 3640
rect 11950 3510 11960 3540
rect 11990 3510 12000 3540
rect 11950 3485 12000 3510
rect 11950 3465 11965 3485
rect 11985 3465 12000 3485
rect 11950 3440 12000 3465
rect 11950 3410 11960 3440
rect 11990 3410 12000 3440
rect 11950 3385 12000 3410
rect 11950 3365 11965 3385
rect 11985 3365 12000 3385
rect 11950 3340 12000 3365
rect 11950 3310 11960 3340
rect 11990 3310 12000 3340
rect 11950 3285 12000 3310
rect 11950 3265 11965 3285
rect 11985 3265 12000 3285
rect 11950 3240 12000 3265
rect 11950 3210 11960 3240
rect 11990 3210 12000 3240
rect 11950 3185 12000 3210
rect 11950 3165 11965 3185
rect 11985 3165 12000 3185
rect 11950 3140 12000 3165
rect 11950 3110 11960 3140
rect 11990 3110 12000 3140
rect 11950 3085 12000 3110
rect 11950 3065 11965 3085
rect 11985 3065 12000 3085
rect 10750 2960 10760 2990
rect 10790 2960 10800 2990
rect 10750 2950 10800 2960
rect 11950 2990 12000 3065
rect 12550 3535 12600 3610
rect 12700 3640 12750 3650
rect 12700 3610 12710 3640
rect 12740 3610 12750 3640
rect 12700 3600 12750 3610
rect 13000 3640 13050 3650
rect 13000 3610 13010 3640
rect 13040 3610 13050 3640
rect 13000 3600 13050 3610
rect 12550 3515 12565 3535
rect 12585 3515 12600 3535
rect 12550 3485 12600 3515
rect 12550 3465 12565 3485
rect 12585 3465 12600 3485
rect 12550 3435 12600 3465
rect 12550 3415 12565 3435
rect 12585 3415 12600 3435
rect 12550 3385 12600 3415
rect 12550 3365 12565 3385
rect 12585 3365 12600 3385
rect 12550 3335 12600 3365
rect 12550 3315 12565 3335
rect 12585 3315 12600 3335
rect 12550 3285 12600 3315
rect 12550 3265 12565 3285
rect 12585 3265 12600 3285
rect 12550 3235 12600 3265
rect 12550 3215 12565 3235
rect 12585 3215 12600 3235
rect 12550 3185 12600 3215
rect 12550 3165 12565 3185
rect 12585 3165 12600 3185
rect 12550 3135 12600 3165
rect 12550 3115 12565 3135
rect 12585 3115 12600 3135
rect 12550 3085 12600 3115
rect 12550 3065 12565 3085
rect 12585 3065 12600 3085
rect 12550 3050 12600 3065
rect 13150 3540 13200 3710
rect 13750 4835 13800 4910
rect 13900 4940 13950 4950
rect 13900 4910 13910 4940
rect 13940 4910 13950 4940
rect 13900 4900 13950 4910
rect 14200 4940 14250 4950
rect 14200 4910 14210 4940
rect 14240 4910 14250 4940
rect 14200 4900 14250 4910
rect 13750 4815 13765 4835
rect 13785 4815 13800 4835
rect 13750 4785 13800 4815
rect 13750 4765 13765 4785
rect 13785 4765 13800 4785
rect 13750 4735 13800 4765
rect 13750 4715 13765 4735
rect 13785 4715 13800 4735
rect 13750 4685 13800 4715
rect 13750 4665 13765 4685
rect 13785 4665 13800 4685
rect 13750 4635 13800 4665
rect 13750 4615 13765 4635
rect 13785 4615 13800 4635
rect 13750 4585 13800 4615
rect 13750 4565 13765 4585
rect 13785 4565 13800 4585
rect 13750 4535 13800 4565
rect 13750 4515 13765 4535
rect 13785 4515 13800 4535
rect 13750 4485 13800 4515
rect 13750 4465 13765 4485
rect 13785 4465 13800 4485
rect 13750 4435 13800 4465
rect 13750 4415 13765 4435
rect 13785 4415 13800 4435
rect 13750 4385 13800 4415
rect 13750 4365 13765 4385
rect 13785 4365 13800 4385
rect 13750 4185 13800 4365
rect 13750 4165 13765 4185
rect 13785 4165 13800 4185
rect 13750 4135 13800 4165
rect 13750 4115 13765 4135
rect 13785 4115 13800 4135
rect 13750 4085 13800 4115
rect 13750 4065 13765 4085
rect 13785 4065 13800 4085
rect 13750 4035 13800 4065
rect 13750 4015 13765 4035
rect 13785 4015 13800 4035
rect 13750 3985 13800 4015
rect 13750 3965 13765 3985
rect 13785 3965 13800 3985
rect 13750 3935 13800 3965
rect 13750 3915 13765 3935
rect 13785 3915 13800 3935
rect 13750 3885 13800 3915
rect 13750 3865 13765 3885
rect 13785 3865 13800 3885
rect 13750 3835 13800 3865
rect 13750 3815 13765 3835
rect 13785 3815 13800 3835
rect 13750 3785 13800 3815
rect 13750 3765 13765 3785
rect 13785 3765 13800 3785
rect 13750 3735 13800 3765
rect 13750 3715 13765 3735
rect 13785 3715 13800 3735
rect 13300 3640 13350 3650
rect 13300 3610 13310 3640
rect 13340 3610 13350 3640
rect 13300 3600 13350 3610
rect 13600 3640 13650 3650
rect 13600 3610 13610 3640
rect 13640 3610 13650 3640
rect 13600 3600 13650 3610
rect 13750 3640 13800 3715
rect 14350 4840 14400 5010
rect 14950 5485 15000 5500
rect 14950 5465 14965 5485
rect 14985 5465 15000 5485
rect 14950 5435 15000 5465
rect 14950 5415 14965 5435
rect 14985 5415 15000 5435
rect 14950 5385 15000 5415
rect 14950 5365 14965 5385
rect 14985 5365 15000 5385
rect 14950 5335 15000 5365
rect 14950 5315 14965 5335
rect 14985 5315 15000 5335
rect 14950 5285 15000 5315
rect 14950 5265 14965 5285
rect 14985 5265 15000 5285
rect 14950 5235 15000 5265
rect 14950 5215 14965 5235
rect 14985 5215 15000 5235
rect 14950 5185 15000 5215
rect 14950 5165 14965 5185
rect 14985 5165 15000 5185
rect 14950 5135 15000 5165
rect 14950 5115 14965 5135
rect 14985 5115 15000 5135
rect 14950 5085 15000 5115
rect 14950 5065 14965 5085
rect 14985 5065 15000 5085
rect 14950 5035 15000 5065
rect 14950 5015 14965 5035
rect 14985 5015 15000 5035
rect 14500 4940 14550 4950
rect 14500 4910 14510 4940
rect 14540 4910 14550 4940
rect 14500 4900 14550 4910
rect 14800 4940 14850 4950
rect 14800 4910 14810 4940
rect 14840 4910 14850 4940
rect 14800 4900 14850 4910
rect 14950 4940 15000 5015
rect 15550 5485 15600 5560
rect 20350 5590 20400 5600
rect 20350 5560 20360 5590
rect 20390 5560 20400 5590
rect 15550 5465 15565 5485
rect 15585 5465 15600 5485
rect 15550 5440 15600 5465
rect 15550 5410 15560 5440
rect 15590 5410 15600 5440
rect 15550 5385 15600 5410
rect 15550 5365 15565 5385
rect 15585 5365 15600 5385
rect 15550 5340 15600 5365
rect 15550 5310 15560 5340
rect 15590 5310 15600 5340
rect 15550 5285 15600 5310
rect 15550 5265 15565 5285
rect 15585 5265 15600 5285
rect 15550 5240 15600 5265
rect 15550 5210 15560 5240
rect 15590 5210 15600 5240
rect 15550 5185 15600 5210
rect 15550 5165 15565 5185
rect 15585 5165 15600 5185
rect 15550 5140 15600 5165
rect 15550 5110 15560 5140
rect 15590 5110 15600 5140
rect 15550 5085 15600 5110
rect 15550 5065 15565 5085
rect 15585 5065 15600 5085
rect 15550 5040 15600 5065
rect 15550 5010 15560 5040
rect 15590 5010 15600 5040
rect 14950 4910 14960 4940
rect 14990 4910 15000 4940
rect 14350 4810 14360 4840
rect 14390 4810 14400 4840
rect 14350 4785 14400 4810
rect 14350 4765 14365 4785
rect 14385 4765 14400 4785
rect 14350 4740 14400 4765
rect 14350 4710 14360 4740
rect 14390 4710 14400 4740
rect 14350 4685 14400 4710
rect 14350 4665 14365 4685
rect 14385 4665 14400 4685
rect 14350 4640 14400 4665
rect 14350 4610 14360 4640
rect 14390 4610 14400 4640
rect 14350 4585 14400 4610
rect 14350 4565 14365 4585
rect 14385 4565 14400 4585
rect 14350 4540 14400 4565
rect 14350 4510 14360 4540
rect 14390 4510 14400 4540
rect 14350 4485 14400 4510
rect 14350 4465 14365 4485
rect 14385 4465 14400 4485
rect 14350 4440 14400 4465
rect 14350 4410 14360 4440
rect 14390 4410 14400 4440
rect 14350 4385 14400 4410
rect 14350 4365 14365 4385
rect 14385 4365 14400 4385
rect 14350 4290 14400 4365
rect 14350 4260 14360 4290
rect 14390 4260 14400 4290
rect 14350 4185 14400 4260
rect 14350 4165 14365 4185
rect 14385 4165 14400 4185
rect 14350 4140 14400 4165
rect 14350 4110 14360 4140
rect 14390 4110 14400 4140
rect 14350 4085 14400 4110
rect 14350 4065 14365 4085
rect 14385 4065 14400 4085
rect 14350 4040 14400 4065
rect 14350 4010 14360 4040
rect 14390 4010 14400 4040
rect 14350 3985 14400 4010
rect 14350 3965 14365 3985
rect 14385 3965 14400 3985
rect 14350 3940 14400 3965
rect 14350 3910 14360 3940
rect 14390 3910 14400 3940
rect 14350 3885 14400 3910
rect 14350 3865 14365 3885
rect 14385 3865 14400 3885
rect 14350 3840 14400 3865
rect 14350 3810 14360 3840
rect 14390 3810 14400 3840
rect 14350 3785 14400 3810
rect 14350 3765 14365 3785
rect 14385 3765 14400 3785
rect 14350 3740 14400 3765
rect 14350 3710 14360 3740
rect 14390 3710 14400 3740
rect 13750 3610 13760 3640
rect 13790 3610 13800 3640
rect 13150 3510 13160 3540
rect 13190 3510 13200 3540
rect 13150 3485 13200 3510
rect 13150 3465 13165 3485
rect 13185 3465 13200 3485
rect 13150 3440 13200 3465
rect 13150 3410 13160 3440
rect 13190 3410 13200 3440
rect 13150 3385 13200 3410
rect 13150 3365 13165 3385
rect 13185 3365 13200 3385
rect 13150 3340 13200 3365
rect 13150 3310 13160 3340
rect 13190 3310 13200 3340
rect 13150 3285 13200 3310
rect 13150 3265 13165 3285
rect 13185 3265 13200 3285
rect 13150 3240 13200 3265
rect 13150 3210 13160 3240
rect 13190 3210 13200 3240
rect 13150 3185 13200 3210
rect 13150 3165 13165 3185
rect 13185 3165 13200 3185
rect 13150 3140 13200 3165
rect 13150 3110 13160 3140
rect 13190 3110 13200 3140
rect 13150 3085 13200 3110
rect 13150 3065 13165 3085
rect 13185 3065 13200 3085
rect 11950 2960 11960 2990
rect 11990 2960 12000 2990
rect 11950 2950 12000 2960
rect 13150 2990 13200 3065
rect 13750 3535 13800 3610
rect 13900 3640 13950 3650
rect 13900 3610 13910 3640
rect 13940 3610 13950 3640
rect 13900 3600 13950 3610
rect 14200 3640 14250 3650
rect 14200 3610 14210 3640
rect 14240 3610 14250 3640
rect 14200 3600 14250 3610
rect 13750 3515 13765 3535
rect 13785 3515 13800 3535
rect 13750 3485 13800 3515
rect 13750 3465 13765 3485
rect 13785 3465 13800 3485
rect 13750 3435 13800 3465
rect 13750 3415 13765 3435
rect 13785 3415 13800 3435
rect 13750 3385 13800 3415
rect 13750 3365 13765 3385
rect 13785 3365 13800 3385
rect 13750 3335 13800 3365
rect 13750 3315 13765 3335
rect 13785 3315 13800 3335
rect 13750 3285 13800 3315
rect 13750 3265 13765 3285
rect 13785 3265 13800 3285
rect 13750 3235 13800 3265
rect 13750 3215 13765 3235
rect 13785 3215 13800 3235
rect 13750 3185 13800 3215
rect 13750 3165 13765 3185
rect 13785 3165 13800 3185
rect 13750 3135 13800 3165
rect 13750 3115 13765 3135
rect 13785 3115 13800 3135
rect 13750 3085 13800 3115
rect 13750 3065 13765 3085
rect 13785 3065 13800 3085
rect 13750 3050 13800 3065
rect 14350 3540 14400 3710
rect 14950 4835 15000 4910
rect 15100 4940 15150 4950
rect 15100 4910 15110 4940
rect 15140 4910 15150 4940
rect 15100 4900 15150 4910
rect 15400 4940 15450 4950
rect 15400 4910 15410 4940
rect 15440 4910 15450 4940
rect 15400 4900 15450 4910
rect 14950 4815 14965 4835
rect 14985 4815 15000 4835
rect 14950 4785 15000 4815
rect 14950 4765 14965 4785
rect 14985 4765 15000 4785
rect 14950 4735 15000 4765
rect 14950 4715 14965 4735
rect 14985 4715 15000 4735
rect 14950 4685 15000 4715
rect 14950 4665 14965 4685
rect 14985 4665 15000 4685
rect 14950 4635 15000 4665
rect 14950 4615 14965 4635
rect 14985 4615 15000 4635
rect 14950 4585 15000 4615
rect 14950 4565 14965 4585
rect 14985 4565 15000 4585
rect 14950 4535 15000 4565
rect 14950 4515 14965 4535
rect 14985 4515 15000 4535
rect 14950 4485 15000 4515
rect 14950 4465 14965 4485
rect 14985 4465 15000 4485
rect 14950 4435 15000 4465
rect 14950 4415 14965 4435
rect 14985 4415 15000 4435
rect 14950 4385 15000 4415
rect 14950 4365 14965 4385
rect 14985 4365 15000 4385
rect 14950 4185 15000 4365
rect 14950 4165 14965 4185
rect 14985 4165 15000 4185
rect 14950 4135 15000 4165
rect 14950 4115 14965 4135
rect 14985 4115 15000 4135
rect 14950 4085 15000 4115
rect 14950 4065 14965 4085
rect 14985 4065 15000 4085
rect 14950 4035 15000 4065
rect 14950 4015 14965 4035
rect 14985 4015 15000 4035
rect 14950 3985 15000 4015
rect 14950 3965 14965 3985
rect 14985 3965 15000 3985
rect 14950 3935 15000 3965
rect 14950 3915 14965 3935
rect 14985 3915 15000 3935
rect 14950 3885 15000 3915
rect 14950 3865 14965 3885
rect 14985 3865 15000 3885
rect 14950 3835 15000 3865
rect 14950 3815 14965 3835
rect 14985 3815 15000 3835
rect 14950 3785 15000 3815
rect 14950 3765 14965 3785
rect 14985 3765 15000 3785
rect 14950 3735 15000 3765
rect 14950 3715 14965 3735
rect 14985 3715 15000 3735
rect 14500 3640 14550 3650
rect 14500 3610 14510 3640
rect 14540 3610 14550 3640
rect 14500 3600 14550 3610
rect 14800 3640 14850 3650
rect 14800 3610 14810 3640
rect 14840 3610 14850 3640
rect 14800 3600 14850 3610
rect 14950 3640 15000 3715
rect 15550 4840 15600 5010
rect 16150 5485 19800 5500
rect 16150 5465 16165 5485
rect 16185 5465 16465 5485
rect 16485 5465 16765 5485
rect 16785 5465 17065 5485
rect 17085 5465 17365 5485
rect 17385 5465 18565 5485
rect 18585 5465 18865 5485
rect 18885 5465 19165 5485
rect 19185 5465 19465 5485
rect 19485 5465 19765 5485
rect 19785 5465 19800 5485
rect 16150 5450 19800 5465
rect 16150 5435 16200 5450
rect 16150 5415 16165 5435
rect 16185 5415 16200 5435
rect 16150 5385 16200 5415
rect 16450 5435 16500 5450
rect 16450 5415 16465 5435
rect 16485 5415 16500 5435
rect 16150 5365 16165 5385
rect 16185 5365 16200 5385
rect 16150 5335 16200 5365
rect 16150 5315 16165 5335
rect 16185 5315 16200 5335
rect 16150 5285 16200 5315
rect 16150 5265 16165 5285
rect 16185 5265 16200 5285
rect 16150 5235 16200 5265
rect 16150 5215 16165 5235
rect 16185 5215 16200 5235
rect 16150 5185 16200 5215
rect 16150 5165 16165 5185
rect 16185 5165 16200 5185
rect 16150 5135 16200 5165
rect 16150 5115 16165 5135
rect 16185 5115 16200 5135
rect 16150 5085 16200 5115
rect 16150 5065 16165 5085
rect 16185 5065 16200 5085
rect 16150 5035 16200 5065
rect 16150 5015 16165 5035
rect 16185 5015 16200 5035
rect 15700 4940 15750 4950
rect 15700 4910 15710 4940
rect 15740 4910 15750 4940
rect 15700 4900 15750 4910
rect 16000 4940 16050 4950
rect 16000 4910 16010 4940
rect 16040 4910 16050 4940
rect 16000 4900 16050 4910
rect 15550 4810 15560 4840
rect 15590 4810 15600 4840
rect 15550 4785 15600 4810
rect 15550 4765 15565 4785
rect 15585 4765 15600 4785
rect 15550 4740 15600 4765
rect 15550 4710 15560 4740
rect 15590 4710 15600 4740
rect 15550 4685 15600 4710
rect 15550 4665 15565 4685
rect 15585 4665 15600 4685
rect 15550 4640 15600 4665
rect 15550 4610 15560 4640
rect 15590 4610 15600 4640
rect 15550 4585 15600 4610
rect 15550 4565 15565 4585
rect 15585 4565 15600 4585
rect 15550 4540 15600 4565
rect 15550 4510 15560 4540
rect 15590 4510 15600 4540
rect 15550 4485 15600 4510
rect 15550 4465 15565 4485
rect 15585 4465 15600 4485
rect 15550 4440 15600 4465
rect 15550 4410 15560 4440
rect 15590 4410 15600 4440
rect 15550 4385 15600 4410
rect 15550 4365 15565 4385
rect 15585 4365 15600 4385
rect 15550 4290 15600 4365
rect 16150 4835 16200 5015
rect 16300 5385 16350 5400
rect 16300 5365 16315 5385
rect 16335 5365 16350 5385
rect 16300 5335 16350 5365
rect 16300 5315 16315 5335
rect 16335 5315 16350 5335
rect 16300 5285 16350 5315
rect 16300 5265 16315 5285
rect 16335 5265 16350 5285
rect 16300 5235 16350 5265
rect 16300 5215 16315 5235
rect 16335 5215 16350 5235
rect 16300 5185 16350 5215
rect 16300 5165 16315 5185
rect 16335 5165 16350 5185
rect 16300 5135 16350 5165
rect 16300 5115 16315 5135
rect 16335 5115 16350 5135
rect 16300 5085 16350 5115
rect 16450 5385 16500 5415
rect 16750 5435 16800 5450
rect 16750 5415 16765 5435
rect 16785 5415 16800 5435
rect 16450 5365 16465 5385
rect 16485 5365 16500 5385
rect 16450 5335 16500 5365
rect 16450 5315 16465 5335
rect 16485 5315 16500 5335
rect 16450 5285 16500 5315
rect 16450 5265 16465 5285
rect 16485 5265 16500 5285
rect 16450 5235 16500 5265
rect 16450 5215 16465 5235
rect 16485 5215 16500 5235
rect 16450 5185 16500 5215
rect 16450 5165 16465 5185
rect 16485 5165 16500 5185
rect 16450 5135 16500 5165
rect 16450 5115 16465 5135
rect 16485 5115 16500 5135
rect 16450 5100 16500 5115
rect 16600 5385 16650 5400
rect 16600 5365 16615 5385
rect 16635 5365 16650 5385
rect 16600 5335 16650 5365
rect 16600 5315 16615 5335
rect 16635 5315 16650 5335
rect 16600 5285 16650 5315
rect 16600 5265 16615 5285
rect 16635 5265 16650 5285
rect 16600 5235 16650 5265
rect 16600 5215 16615 5235
rect 16635 5215 16650 5235
rect 16600 5185 16650 5215
rect 16600 5165 16615 5185
rect 16635 5165 16650 5185
rect 16600 5135 16650 5165
rect 16600 5115 16615 5135
rect 16635 5115 16650 5135
rect 16300 5065 16315 5085
rect 16335 5065 16350 5085
rect 16300 5050 16350 5065
rect 16600 5085 16650 5115
rect 16750 5385 16800 5415
rect 17050 5435 17100 5450
rect 17050 5415 17065 5435
rect 17085 5415 17100 5435
rect 16750 5365 16765 5385
rect 16785 5365 16800 5385
rect 16750 5335 16800 5365
rect 16750 5315 16765 5335
rect 16785 5315 16800 5335
rect 16750 5285 16800 5315
rect 16750 5265 16765 5285
rect 16785 5265 16800 5285
rect 16750 5235 16800 5265
rect 16750 5215 16765 5235
rect 16785 5215 16800 5235
rect 16750 5185 16800 5215
rect 16750 5165 16765 5185
rect 16785 5165 16800 5185
rect 16750 5135 16800 5165
rect 16750 5115 16765 5135
rect 16785 5115 16800 5135
rect 16750 5100 16800 5115
rect 16900 5385 16950 5400
rect 16900 5365 16915 5385
rect 16935 5365 16950 5385
rect 16900 5335 16950 5365
rect 16900 5315 16915 5335
rect 16935 5315 16950 5335
rect 16900 5285 16950 5315
rect 16900 5265 16915 5285
rect 16935 5265 16950 5285
rect 16900 5235 16950 5265
rect 16900 5215 16915 5235
rect 16935 5215 16950 5235
rect 16900 5185 16950 5215
rect 16900 5165 16915 5185
rect 16935 5165 16950 5185
rect 16900 5135 16950 5165
rect 16900 5115 16915 5135
rect 16935 5115 16950 5135
rect 16600 5065 16615 5085
rect 16635 5065 16650 5085
rect 16600 5050 16650 5065
rect 16900 5085 16950 5115
rect 17050 5385 17100 5415
rect 17350 5435 17400 5450
rect 17350 5415 17365 5435
rect 17385 5415 17400 5435
rect 17050 5365 17065 5385
rect 17085 5365 17100 5385
rect 17050 5335 17100 5365
rect 17050 5315 17065 5335
rect 17085 5315 17100 5335
rect 17050 5285 17100 5315
rect 17050 5265 17065 5285
rect 17085 5265 17100 5285
rect 17050 5235 17100 5265
rect 17050 5215 17065 5235
rect 17085 5215 17100 5235
rect 17050 5185 17100 5215
rect 17050 5165 17065 5185
rect 17085 5165 17100 5185
rect 17050 5135 17100 5165
rect 17050 5115 17065 5135
rect 17085 5115 17100 5135
rect 17050 5100 17100 5115
rect 17200 5385 17250 5400
rect 17200 5365 17215 5385
rect 17235 5365 17250 5385
rect 17200 5335 17250 5365
rect 17200 5315 17215 5335
rect 17235 5315 17250 5335
rect 17200 5285 17250 5315
rect 17200 5265 17215 5285
rect 17235 5265 17250 5285
rect 17200 5235 17250 5265
rect 17200 5215 17215 5235
rect 17235 5215 17250 5235
rect 17200 5185 17250 5215
rect 17200 5165 17215 5185
rect 17235 5165 17250 5185
rect 17200 5135 17250 5165
rect 17200 5115 17215 5135
rect 17235 5115 17250 5135
rect 16900 5065 16915 5085
rect 16935 5065 16950 5085
rect 16900 5050 16950 5065
rect 17200 5085 17250 5115
rect 17200 5065 17215 5085
rect 17235 5065 17250 5085
rect 17200 5050 17250 5065
rect 16300 5035 17250 5050
rect 16300 5015 16315 5035
rect 16335 5015 16615 5035
rect 16635 5015 16915 5035
rect 16935 5015 17215 5035
rect 17235 5015 17250 5035
rect 16300 5000 17250 5015
rect 17350 5385 17400 5415
rect 18550 5435 18600 5450
rect 18550 5415 18565 5435
rect 18585 5415 18600 5435
rect 17350 5365 17365 5385
rect 17385 5365 17400 5385
rect 17350 5335 17400 5365
rect 17350 5315 17365 5335
rect 17385 5315 17400 5335
rect 17350 5285 17400 5315
rect 17350 5265 17365 5285
rect 17385 5265 17400 5285
rect 17350 5235 17400 5265
rect 17350 5215 17365 5235
rect 17385 5215 17400 5235
rect 17350 5185 17400 5215
rect 17350 5165 17365 5185
rect 17385 5165 17400 5185
rect 17350 5135 17400 5165
rect 17350 5115 17365 5135
rect 17385 5115 17400 5135
rect 17350 5085 17400 5115
rect 17350 5065 17365 5085
rect 17385 5065 17400 5085
rect 17350 5035 17400 5065
rect 17350 5015 17365 5035
rect 17385 5015 17400 5035
rect 16300 4940 16350 4950
rect 16300 4910 16310 4940
rect 16340 4910 16350 4940
rect 16300 4900 16350 4910
rect 16450 4850 16500 5000
rect 16600 4940 16650 4950
rect 16600 4910 16610 4940
rect 16640 4910 16650 4940
rect 16600 4900 16650 4910
rect 16750 4940 16800 5000
rect 16750 4910 16760 4940
rect 16790 4910 16800 4940
rect 16750 4850 16800 4910
rect 16900 4940 16950 4950
rect 16900 4910 16910 4940
rect 16940 4910 16950 4940
rect 16900 4900 16950 4910
rect 17050 4850 17100 5000
rect 17200 4940 17250 4950
rect 17200 4910 17210 4940
rect 17240 4910 17250 4940
rect 17200 4900 17250 4910
rect 16150 4815 16165 4835
rect 16185 4815 16200 4835
rect 16150 4785 16200 4815
rect 16150 4765 16165 4785
rect 16185 4765 16200 4785
rect 16150 4735 16200 4765
rect 16150 4715 16165 4735
rect 16185 4715 16200 4735
rect 16150 4685 16200 4715
rect 16150 4665 16165 4685
rect 16185 4665 16200 4685
rect 16150 4635 16200 4665
rect 16150 4615 16165 4635
rect 16185 4615 16200 4635
rect 16150 4585 16200 4615
rect 16150 4565 16165 4585
rect 16185 4565 16200 4585
rect 16150 4535 16200 4565
rect 16150 4515 16165 4535
rect 16185 4515 16200 4535
rect 16150 4485 16200 4515
rect 16150 4465 16165 4485
rect 16185 4465 16200 4485
rect 16150 4435 16200 4465
rect 16300 4835 17250 4850
rect 16300 4815 16315 4835
rect 16335 4815 16615 4835
rect 16635 4815 16915 4835
rect 16935 4815 17215 4835
rect 17235 4815 17250 4835
rect 16300 4800 17250 4815
rect 16300 4785 16350 4800
rect 16300 4765 16315 4785
rect 16335 4765 16350 4785
rect 16300 4735 16350 4765
rect 16600 4785 16650 4800
rect 16600 4765 16615 4785
rect 16635 4765 16650 4785
rect 16300 4715 16315 4735
rect 16335 4715 16350 4735
rect 16300 4685 16350 4715
rect 16300 4665 16315 4685
rect 16335 4665 16350 4685
rect 16300 4635 16350 4665
rect 16300 4615 16315 4635
rect 16335 4615 16350 4635
rect 16300 4585 16350 4615
rect 16300 4565 16315 4585
rect 16335 4565 16350 4585
rect 16300 4535 16350 4565
rect 16300 4515 16315 4535
rect 16335 4515 16350 4535
rect 16300 4485 16350 4515
rect 16300 4465 16315 4485
rect 16335 4465 16350 4485
rect 16300 4450 16350 4465
rect 16450 4735 16500 4750
rect 16450 4715 16465 4735
rect 16485 4715 16500 4735
rect 16450 4685 16500 4715
rect 16450 4665 16465 4685
rect 16485 4665 16500 4685
rect 16450 4635 16500 4665
rect 16450 4615 16465 4635
rect 16485 4615 16500 4635
rect 16450 4585 16500 4615
rect 16450 4565 16465 4585
rect 16485 4565 16500 4585
rect 16450 4535 16500 4565
rect 16450 4515 16465 4535
rect 16485 4515 16500 4535
rect 16450 4485 16500 4515
rect 16450 4465 16465 4485
rect 16485 4465 16500 4485
rect 16150 4415 16165 4435
rect 16185 4415 16200 4435
rect 16150 4400 16200 4415
rect 16450 4435 16500 4465
rect 16600 4735 16650 4765
rect 16900 4785 16950 4800
rect 16900 4765 16915 4785
rect 16935 4765 16950 4785
rect 16600 4715 16615 4735
rect 16635 4715 16650 4735
rect 16600 4685 16650 4715
rect 16600 4665 16615 4685
rect 16635 4665 16650 4685
rect 16600 4635 16650 4665
rect 16600 4615 16615 4635
rect 16635 4615 16650 4635
rect 16600 4585 16650 4615
rect 16600 4565 16615 4585
rect 16635 4565 16650 4585
rect 16600 4535 16650 4565
rect 16600 4515 16615 4535
rect 16635 4515 16650 4535
rect 16600 4485 16650 4515
rect 16600 4465 16615 4485
rect 16635 4465 16650 4485
rect 16600 4450 16650 4465
rect 16750 4735 16800 4750
rect 16750 4715 16765 4735
rect 16785 4715 16800 4735
rect 16750 4685 16800 4715
rect 16750 4665 16765 4685
rect 16785 4665 16800 4685
rect 16750 4635 16800 4665
rect 16750 4615 16765 4635
rect 16785 4615 16800 4635
rect 16750 4585 16800 4615
rect 16750 4565 16765 4585
rect 16785 4565 16800 4585
rect 16750 4535 16800 4565
rect 16750 4515 16765 4535
rect 16785 4515 16800 4535
rect 16750 4485 16800 4515
rect 16750 4465 16765 4485
rect 16785 4465 16800 4485
rect 16450 4415 16465 4435
rect 16485 4415 16500 4435
rect 16450 4400 16500 4415
rect 16750 4435 16800 4465
rect 16900 4735 16950 4765
rect 17200 4785 17250 4800
rect 17200 4765 17215 4785
rect 17235 4765 17250 4785
rect 16900 4715 16915 4735
rect 16935 4715 16950 4735
rect 16900 4685 16950 4715
rect 16900 4665 16915 4685
rect 16935 4665 16950 4685
rect 16900 4635 16950 4665
rect 16900 4615 16915 4635
rect 16935 4615 16950 4635
rect 16900 4585 16950 4615
rect 16900 4565 16915 4585
rect 16935 4565 16950 4585
rect 16900 4535 16950 4565
rect 16900 4515 16915 4535
rect 16935 4515 16950 4535
rect 16900 4485 16950 4515
rect 16900 4465 16915 4485
rect 16935 4465 16950 4485
rect 16900 4450 16950 4465
rect 17050 4735 17100 4750
rect 17050 4715 17065 4735
rect 17085 4715 17100 4735
rect 17050 4685 17100 4715
rect 17050 4665 17065 4685
rect 17085 4665 17100 4685
rect 17050 4635 17100 4665
rect 17050 4615 17065 4635
rect 17085 4615 17100 4635
rect 17050 4585 17100 4615
rect 17050 4565 17065 4585
rect 17085 4565 17100 4585
rect 17050 4535 17100 4565
rect 17050 4515 17065 4535
rect 17085 4515 17100 4535
rect 17050 4485 17100 4515
rect 17050 4465 17065 4485
rect 17085 4465 17100 4485
rect 16750 4415 16765 4435
rect 16785 4415 16800 4435
rect 16750 4400 16800 4415
rect 17050 4435 17100 4465
rect 17200 4735 17250 4765
rect 17200 4715 17215 4735
rect 17235 4715 17250 4735
rect 17200 4685 17250 4715
rect 17200 4665 17215 4685
rect 17235 4665 17250 4685
rect 17200 4635 17250 4665
rect 17200 4615 17215 4635
rect 17235 4615 17250 4635
rect 17200 4585 17250 4615
rect 17200 4565 17215 4585
rect 17235 4565 17250 4585
rect 17200 4535 17250 4565
rect 17200 4515 17215 4535
rect 17235 4515 17250 4535
rect 17200 4485 17250 4515
rect 17200 4465 17215 4485
rect 17235 4465 17250 4485
rect 17200 4450 17250 4465
rect 17350 4835 17400 5015
rect 17950 5385 18000 5400
rect 17950 5365 17965 5385
rect 17985 5365 18000 5385
rect 17950 5340 18000 5365
rect 17950 5310 17960 5340
rect 17990 5310 18000 5340
rect 17950 5285 18000 5310
rect 17950 5265 17965 5285
rect 17985 5265 18000 5285
rect 17950 5240 18000 5265
rect 17950 5210 17960 5240
rect 17990 5210 18000 5240
rect 17950 5185 18000 5210
rect 17950 5165 17965 5185
rect 17985 5165 18000 5185
rect 17950 5140 18000 5165
rect 17950 5110 17960 5140
rect 17990 5110 18000 5140
rect 17950 5085 18000 5110
rect 17950 5065 17965 5085
rect 17985 5065 18000 5085
rect 17950 5040 18000 5065
rect 17950 5010 17960 5040
rect 17990 5010 18000 5040
rect 17500 4940 17550 4950
rect 17500 4910 17510 4940
rect 17540 4910 17550 4940
rect 17500 4900 17550 4910
rect 17800 4940 17850 4950
rect 17800 4910 17810 4940
rect 17840 4910 17850 4940
rect 17800 4900 17850 4910
rect 17350 4815 17365 4835
rect 17385 4815 17400 4835
rect 17350 4785 17400 4815
rect 17350 4765 17365 4785
rect 17385 4765 17400 4785
rect 17350 4735 17400 4765
rect 17350 4715 17365 4735
rect 17385 4715 17400 4735
rect 17350 4685 17400 4715
rect 17350 4665 17365 4685
rect 17385 4665 17400 4685
rect 17350 4635 17400 4665
rect 17350 4615 17365 4635
rect 17385 4615 17400 4635
rect 17350 4585 17400 4615
rect 17350 4565 17365 4585
rect 17385 4565 17400 4585
rect 17350 4535 17400 4565
rect 17350 4515 17365 4535
rect 17385 4515 17400 4535
rect 17350 4485 17400 4515
rect 17350 4465 17365 4485
rect 17385 4465 17400 4485
rect 17050 4415 17065 4435
rect 17085 4415 17100 4435
rect 17050 4400 17100 4415
rect 17350 4435 17400 4465
rect 17950 4840 18000 5010
rect 18550 5385 18600 5415
rect 18850 5435 18900 5450
rect 18850 5415 18865 5435
rect 18885 5415 18900 5435
rect 18550 5365 18565 5385
rect 18585 5365 18600 5385
rect 18550 5335 18600 5365
rect 18550 5315 18565 5335
rect 18585 5315 18600 5335
rect 18550 5285 18600 5315
rect 18550 5265 18565 5285
rect 18585 5265 18600 5285
rect 18550 5235 18600 5265
rect 18550 5215 18565 5235
rect 18585 5215 18600 5235
rect 18550 5185 18600 5215
rect 18550 5165 18565 5185
rect 18585 5165 18600 5185
rect 18550 5135 18600 5165
rect 18550 5115 18565 5135
rect 18585 5115 18600 5135
rect 18550 5085 18600 5115
rect 18550 5065 18565 5085
rect 18585 5065 18600 5085
rect 18550 5035 18600 5065
rect 18550 5015 18565 5035
rect 18585 5015 18600 5035
rect 18100 4940 18150 4950
rect 18100 4910 18110 4940
rect 18140 4910 18150 4940
rect 18100 4900 18150 4910
rect 18400 4940 18450 4950
rect 18400 4910 18410 4940
rect 18440 4910 18450 4940
rect 18400 4900 18450 4910
rect 17950 4810 17960 4840
rect 17990 4810 18000 4840
rect 17950 4785 18000 4810
rect 17950 4765 17965 4785
rect 17985 4765 18000 4785
rect 17950 4740 18000 4765
rect 17950 4710 17960 4740
rect 17990 4710 18000 4740
rect 17950 4685 18000 4710
rect 17950 4665 17965 4685
rect 17985 4665 18000 4685
rect 17950 4640 18000 4665
rect 17950 4610 17960 4640
rect 17990 4610 18000 4640
rect 17950 4585 18000 4610
rect 17950 4565 17965 4585
rect 17985 4565 18000 4585
rect 17950 4540 18000 4565
rect 17950 4510 17960 4540
rect 17990 4510 18000 4540
rect 17950 4485 18000 4510
rect 17950 4465 17965 4485
rect 17985 4465 18000 4485
rect 17950 4450 18000 4465
rect 18550 4835 18600 5015
rect 18700 5385 18750 5400
rect 18700 5365 18715 5385
rect 18735 5365 18750 5385
rect 18700 5335 18750 5365
rect 18700 5315 18715 5335
rect 18735 5315 18750 5335
rect 18700 5285 18750 5315
rect 18700 5265 18715 5285
rect 18735 5265 18750 5285
rect 18700 5235 18750 5265
rect 18700 5215 18715 5235
rect 18735 5215 18750 5235
rect 18700 5185 18750 5215
rect 18700 5165 18715 5185
rect 18735 5165 18750 5185
rect 18700 5135 18750 5165
rect 18700 5115 18715 5135
rect 18735 5115 18750 5135
rect 18700 5085 18750 5115
rect 18850 5385 18900 5415
rect 19150 5435 19200 5450
rect 19150 5415 19165 5435
rect 19185 5415 19200 5435
rect 18850 5365 18865 5385
rect 18885 5365 18900 5385
rect 18850 5335 18900 5365
rect 18850 5315 18865 5335
rect 18885 5315 18900 5335
rect 18850 5285 18900 5315
rect 18850 5265 18865 5285
rect 18885 5265 18900 5285
rect 18850 5235 18900 5265
rect 18850 5215 18865 5235
rect 18885 5215 18900 5235
rect 18850 5185 18900 5215
rect 18850 5165 18865 5185
rect 18885 5165 18900 5185
rect 18850 5135 18900 5165
rect 18850 5115 18865 5135
rect 18885 5115 18900 5135
rect 18850 5100 18900 5115
rect 19000 5385 19050 5400
rect 19000 5365 19015 5385
rect 19035 5365 19050 5385
rect 19000 5335 19050 5365
rect 19000 5315 19015 5335
rect 19035 5315 19050 5335
rect 19000 5285 19050 5315
rect 19000 5265 19015 5285
rect 19035 5265 19050 5285
rect 19000 5235 19050 5265
rect 19000 5215 19015 5235
rect 19035 5215 19050 5235
rect 19000 5185 19050 5215
rect 19000 5165 19015 5185
rect 19035 5165 19050 5185
rect 19000 5135 19050 5165
rect 19000 5115 19015 5135
rect 19035 5115 19050 5135
rect 18700 5065 18715 5085
rect 18735 5065 18750 5085
rect 18700 5050 18750 5065
rect 19000 5085 19050 5115
rect 19150 5385 19200 5415
rect 19450 5435 19500 5450
rect 19450 5415 19465 5435
rect 19485 5415 19500 5435
rect 19150 5365 19165 5385
rect 19185 5365 19200 5385
rect 19150 5335 19200 5365
rect 19150 5315 19165 5335
rect 19185 5315 19200 5335
rect 19150 5285 19200 5315
rect 19150 5265 19165 5285
rect 19185 5265 19200 5285
rect 19150 5235 19200 5265
rect 19150 5215 19165 5235
rect 19185 5215 19200 5235
rect 19150 5185 19200 5215
rect 19150 5165 19165 5185
rect 19185 5165 19200 5185
rect 19150 5135 19200 5165
rect 19150 5115 19165 5135
rect 19185 5115 19200 5135
rect 19150 5100 19200 5115
rect 19300 5385 19350 5400
rect 19300 5365 19315 5385
rect 19335 5365 19350 5385
rect 19300 5335 19350 5365
rect 19300 5315 19315 5335
rect 19335 5315 19350 5335
rect 19300 5285 19350 5315
rect 19300 5265 19315 5285
rect 19335 5265 19350 5285
rect 19300 5235 19350 5265
rect 19300 5215 19315 5235
rect 19335 5215 19350 5235
rect 19300 5185 19350 5215
rect 19300 5165 19315 5185
rect 19335 5165 19350 5185
rect 19300 5135 19350 5165
rect 19300 5115 19315 5135
rect 19335 5115 19350 5135
rect 19000 5065 19015 5085
rect 19035 5065 19050 5085
rect 19000 5050 19050 5065
rect 19300 5085 19350 5115
rect 19450 5385 19500 5415
rect 19750 5435 19800 5450
rect 19750 5415 19765 5435
rect 19785 5415 19800 5435
rect 19450 5365 19465 5385
rect 19485 5365 19500 5385
rect 19450 5335 19500 5365
rect 19450 5315 19465 5335
rect 19485 5315 19500 5335
rect 19450 5285 19500 5315
rect 19450 5265 19465 5285
rect 19485 5265 19500 5285
rect 19450 5235 19500 5265
rect 19450 5215 19465 5235
rect 19485 5215 19500 5235
rect 19450 5185 19500 5215
rect 19450 5165 19465 5185
rect 19485 5165 19500 5185
rect 19450 5135 19500 5165
rect 19450 5115 19465 5135
rect 19485 5115 19500 5135
rect 19450 5100 19500 5115
rect 19600 5385 19650 5400
rect 19600 5365 19615 5385
rect 19635 5365 19650 5385
rect 19600 5335 19650 5365
rect 19600 5315 19615 5335
rect 19635 5315 19650 5335
rect 19600 5285 19650 5315
rect 19600 5265 19615 5285
rect 19635 5265 19650 5285
rect 19600 5235 19650 5265
rect 19600 5215 19615 5235
rect 19635 5215 19650 5235
rect 19600 5185 19650 5215
rect 19600 5165 19615 5185
rect 19635 5165 19650 5185
rect 19600 5135 19650 5165
rect 19600 5115 19615 5135
rect 19635 5115 19650 5135
rect 19300 5065 19315 5085
rect 19335 5065 19350 5085
rect 19300 5050 19350 5065
rect 19600 5085 19650 5115
rect 19600 5065 19615 5085
rect 19635 5065 19650 5085
rect 19600 5050 19650 5065
rect 18700 5035 19650 5050
rect 18700 5015 18715 5035
rect 18735 5015 19015 5035
rect 19035 5015 19315 5035
rect 19335 5015 19615 5035
rect 19635 5015 19650 5035
rect 18700 5000 19650 5015
rect 19750 5385 19800 5415
rect 19750 5365 19765 5385
rect 19785 5365 19800 5385
rect 19750 5335 19800 5365
rect 19750 5315 19765 5335
rect 19785 5315 19800 5335
rect 19750 5285 19800 5315
rect 19750 5265 19765 5285
rect 19785 5265 19800 5285
rect 19750 5235 19800 5265
rect 19750 5215 19765 5235
rect 19785 5215 19800 5235
rect 19750 5185 19800 5215
rect 19750 5165 19765 5185
rect 19785 5165 19800 5185
rect 19750 5135 19800 5165
rect 19750 5115 19765 5135
rect 19785 5115 19800 5135
rect 19750 5085 19800 5115
rect 19750 5065 19765 5085
rect 19785 5065 19800 5085
rect 19750 5035 19800 5065
rect 19750 5015 19765 5035
rect 19785 5015 19800 5035
rect 18700 4940 18750 4950
rect 18700 4910 18710 4940
rect 18740 4910 18750 4940
rect 18700 4900 18750 4910
rect 19000 4940 19050 4950
rect 19000 4910 19010 4940
rect 19040 4910 19050 4940
rect 19000 4900 19050 4910
rect 19150 4940 19200 5000
rect 19150 4910 19160 4940
rect 19190 4910 19200 4940
rect 19150 4850 19200 4910
rect 19300 4940 19350 4950
rect 19300 4910 19310 4940
rect 19340 4910 19350 4940
rect 19300 4900 19350 4910
rect 19600 4940 19650 4950
rect 19600 4910 19610 4940
rect 19640 4910 19650 4940
rect 19600 4900 19650 4910
rect 18550 4815 18565 4835
rect 18585 4815 18600 4835
rect 18550 4785 18600 4815
rect 18550 4765 18565 4785
rect 18585 4765 18600 4785
rect 18550 4735 18600 4765
rect 18550 4715 18565 4735
rect 18585 4715 18600 4735
rect 18550 4685 18600 4715
rect 18550 4665 18565 4685
rect 18585 4665 18600 4685
rect 18550 4635 18600 4665
rect 18550 4615 18565 4635
rect 18585 4615 18600 4635
rect 18550 4585 18600 4615
rect 18550 4565 18565 4585
rect 18585 4565 18600 4585
rect 18550 4535 18600 4565
rect 18550 4515 18565 4535
rect 18585 4515 18600 4535
rect 18550 4485 18600 4515
rect 18550 4465 18565 4485
rect 18585 4465 18600 4485
rect 17350 4415 17365 4435
rect 17385 4415 17400 4435
rect 17350 4400 17400 4415
rect 18550 4435 18600 4465
rect 18700 4835 19650 4850
rect 18700 4815 18715 4835
rect 18735 4815 19015 4835
rect 19035 4815 19315 4835
rect 19335 4815 19615 4835
rect 19635 4815 19650 4835
rect 18700 4800 19650 4815
rect 18700 4785 18750 4800
rect 18700 4765 18715 4785
rect 18735 4765 18750 4785
rect 18700 4735 18750 4765
rect 19000 4785 19050 4800
rect 19000 4765 19015 4785
rect 19035 4765 19050 4785
rect 18700 4715 18715 4735
rect 18735 4715 18750 4735
rect 18700 4685 18750 4715
rect 18700 4665 18715 4685
rect 18735 4665 18750 4685
rect 18700 4635 18750 4665
rect 18700 4615 18715 4635
rect 18735 4615 18750 4635
rect 18700 4585 18750 4615
rect 18700 4565 18715 4585
rect 18735 4565 18750 4585
rect 18700 4535 18750 4565
rect 18700 4515 18715 4535
rect 18735 4515 18750 4535
rect 18700 4485 18750 4515
rect 18700 4465 18715 4485
rect 18735 4465 18750 4485
rect 18700 4450 18750 4465
rect 18850 4735 18900 4750
rect 18850 4715 18865 4735
rect 18885 4715 18900 4735
rect 18850 4685 18900 4715
rect 18850 4665 18865 4685
rect 18885 4665 18900 4685
rect 18850 4635 18900 4665
rect 18850 4615 18865 4635
rect 18885 4615 18900 4635
rect 18850 4585 18900 4615
rect 18850 4565 18865 4585
rect 18885 4565 18900 4585
rect 18850 4535 18900 4565
rect 18850 4515 18865 4535
rect 18885 4515 18900 4535
rect 18850 4485 18900 4515
rect 18850 4465 18865 4485
rect 18885 4465 18900 4485
rect 18550 4415 18565 4435
rect 18585 4415 18600 4435
rect 18550 4400 18600 4415
rect 18850 4435 18900 4465
rect 19000 4735 19050 4765
rect 19300 4785 19350 4800
rect 19300 4765 19315 4785
rect 19335 4765 19350 4785
rect 19000 4715 19015 4735
rect 19035 4715 19050 4735
rect 19000 4685 19050 4715
rect 19000 4665 19015 4685
rect 19035 4665 19050 4685
rect 19000 4635 19050 4665
rect 19000 4615 19015 4635
rect 19035 4615 19050 4635
rect 19000 4585 19050 4615
rect 19000 4565 19015 4585
rect 19035 4565 19050 4585
rect 19000 4535 19050 4565
rect 19000 4515 19015 4535
rect 19035 4515 19050 4535
rect 19000 4485 19050 4515
rect 19000 4465 19015 4485
rect 19035 4465 19050 4485
rect 19000 4450 19050 4465
rect 19150 4735 19200 4750
rect 19150 4715 19165 4735
rect 19185 4715 19200 4735
rect 19150 4685 19200 4715
rect 19150 4665 19165 4685
rect 19185 4665 19200 4685
rect 19150 4635 19200 4665
rect 19150 4615 19165 4635
rect 19185 4615 19200 4635
rect 19150 4585 19200 4615
rect 19150 4565 19165 4585
rect 19185 4565 19200 4585
rect 19150 4535 19200 4565
rect 19150 4515 19165 4535
rect 19185 4515 19200 4535
rect 19150 4485 19200 4515
rect 19150 4465 19165 4485
rect 19185 4465 19200 4485
rect 18850 4415 18865 4435
rect 18885 4415 18900 4435
rect 18850 4400 18900 4415
rect 19150 4435 19200 4465
rect 19300 4735 19350 4765
rect 19600 4785 19650 4800
rect 19600 4765 19615 4785
rect 19635 4765 19650 4785
rect 19300 4715 19315 4735
rect 19335 4715 19350 4735
rect 19300 4685 19350 4715
rect 19300 4665 19315 4685
rect 19335 4665 19350 4685
rect 19300 4635 19350 4665
rect 19300 4615 19315 4635
rect 19335 4615 19350 4635
rect 19300 4585 19350 4615
rect 19300 4565 19315 4585
rect 19335 4565 19350 4585
rect 19300 4535 19350 4565
rect 19300 4515 19315 4535
rect 19335 4515 19350 4535
rect 19300 4485 19350 4515
rect 19300 4465 19315 4485
rect 19335 4465 19350 4485
rect 19300 4450 19350 4465
rect 19450 4735 19500 4750
rect 19450 4715 19465 4735
rect 19485 4715 19500 4735
rect 19450 4685 19500 4715
rect 19450 4665 19465 4685
rect 19485 4665 19500 4685
rect 19450 4635 19500 4665
rect 19450 4615 19465 4635
rect 19485 4615 19500 4635
rect 19450 4585 19500 4615
rect 19450 4565 19465 4585
rect 19485 4565 19500 4585
rect 19450 4535 19500 4565
rect 19450 4515 19465 4535
rect 19485 4515 19500 4535
rect 19450 4485 19500 4515
rect 19450 4465 19465 4485
rect 19485 4465 19500 4485
rect 19150 4415 19165 4435
rect 19185 4415 19200 4435
rect 19150 4400 19200 4415
rect 19450 4435 19500 4465
rect 19600 4735 19650 4765
rect 19600 4715 19615 4735
rect 19635 4715 19650 4735
rect 19600 4685 19650 4715
rect 19600 4665 19615 4685
rect 19635 4665 19650 4685
rect 19600 4635 19650 4665
rect 19600 4615 19615 4635
rect 19635 4615 19650 4635
rect 19600 4585 19650 4615
rect 19600 4565 19615 4585
rect 19635 4565 19650 4585
rect 19600 4535 19650 4565
rect 19600 4515 19615 4535
rect 19635 4515 19650 4535
rect 19600 4485 19650 4515
rect 19600 4465 19615 4485
rect 19635 4465 19650 4485
rect 19600 4450 19650 4465
rect 19750 4835 19800 5015
rect 20350 5485 20400 5560
rect 22450 5590 22500 5600
rect 22450 5560 22460 5590
rect 22490 5560 22500 5590
rect 20350 5465 20365 5485
rect 20385 5465 20400 5485
rect 20350 5440 20400 5465
rect 20350 5410 20360 5440
rect 20390 5410 20400 5440
rect 20350 5385 20400 5410
rect 20350 5365 20365 5385
rect 20385 5365 20400 5385
rect 20350 5340 20400 5365
rect 20350 5310 20360 5340
rect 20390 5310 20400 5340
rect 20350 5285 20400 5310
rect 20350 5265 20365 5285
rect 20385 5265 20400 5285
rect 20350 5240 20400 5265
rect 20350 5210 20360 5240
rect 20390 5210 20400 5240
rect 20350 5185 20400 5210
rect 20350 5165 20365 5185
rect 20385 5165 20400 5185
rect 20350 5140 20400 5165
rect 20350 5110 20360 5140
rect 20390 5110 20400 5140
rect 20350 5085 20400 5110
rect 20350 5065 20365 5085
rect 20385 5065 20400 5085
rect 20350 5040 20400 5065
rect 20350 5010 20360 5040
rect 20390 5010 20400 5040
rect 19900 4940 19950 4950
rect 19900 4910 19910 4940
rect 19940 4910 19950 4940
rect 19900 4900 19950 4910
rect 20200 4940 20250 4950
rect 20200 4910 20210 4940
rect 20240 4910 20250 4940
rect 20200 4900 20250 4910
rect 19750 4815 19765 4835
rect 19785 4815 19800 4835
rect 19750 4785 19800 4815
rect 19750 4765 19765 4785
rect 19785 4765 19800 4785
rect 19750 4735 19800 4765
rect 19750 4715 19765 4735
rect 19785 4715 19800 4735
rect 19750 4685 19800 4715
rect 19750 4665 19765 4685
rect 19785 4665 19800 4685
rect 19750 4635 19800 4665
rect 19750 4615 19765 4635
rect 19785 4615 19800 4635
rect 19750 4585 19800 4615
rect 19750 4565 19765 4585
rect 19785 4565 19800 4585
rect 19750 4535 19800 4565
rect 19750 4515 19765 4535
rect 19785 4515 19800 4535
rect 19750 4485 19800 4515
rect 19750 4465 19765 4485
rect 19785 4465 19800 4485
rect 19450 4415 19465 4435
rect 19485 4415 19500 4435
rect 19450 4400 19500 4415
rect 19750 4435 19800 4465
rect 19750 4415 19765 4435
rect 19785 4415 19800 4435
rect 19750 4400 19800 4415
rect 16150 4385 19800 4400
rect 16150 4365 16165 4385
rect 16185 4365 16465 4385
rect 16485 4365 16765 4385
rect 16785 4365 17065 4385
rect 17085 4365 17365 4385
rect 17385 4365 18565 4385
rect 18585 4365 18865 4385
rect 18885 4365 19165 4385
rect 19185 4365 19465 4385
rect 19485 4365 19765 4385
rect 19785 4365 19800 4385
rect 16150 4350 19800 4365
rect 20350 4840 20400 5010
rect 20950 5485 21000 5500
rect 20950 5465 20965 5485
rect 20985 5465 21000 5485
rect 20950 5435 21000 5465
rect 20950 5415 20965 5435
rect 20985 5415 21000 5435
rect 20950 5385 21000 5415
rect 20950 5365 20965 5385
rect 20985 5365 21000 5385
rect 20950 5335 21000 5365
rect 20950 5315 20965 5335
rect 20985 5315 21000 5335
rect 20950 5285 21000 5315
rect 20950 5265 20965 5285
rect 20985 5265 21000 5285
rect 20950 5235 21000 5265
rect 20950 5215 20965 5235
rect 20985 5215 21000 5235
rect 20950 5185 21000 5215
rect 20950 5165 20965 5185
rect 20985 5165 21000 5185
rect 20950 5135 21000 5165
rect 20950 5115 20965 5135
rect 20985 5115 21000 5135
rect 20950 5085 21000 5115
rect 20950 5065 20965 5085
rect 20985 5065 21000 5085
rect 20950 5035 21000 5065
rect 20950 5015 20965 5035
rect 20985 5015 21000 5035
rect 20500 4940 20550 4950
rect 20500 4910 20510 4940
rect 20540 4910 20550 4940
rect 20500 4900 20550 4910
rect 20800 4940 20850 4950
rect 20800 4910 20810 4940
rect 20840 4910 20850 4940
rect 20800 4900 20850 4910
rect 20950 4940 21000 5015
rect 21400 5485 21450 5500
rect 21400 5465 21415 5485
rect 21435 5465 21450 5485
rect 21400 5435 21450 5465
rect 21400 5415 21415 5435
rect 21435 5415 21450 5435
rect 21400 5385 21450 5415
rect 21400 5365 21415 5385
rect 21435 5365 21450 5385
rect 21400 5335 21450 5365
rect 21400 5315 21415 5335
rect 21435 5315 21450 5335
rect 21400 5285 21450 5315
rect 21400 5265 21415 5285
rect 21435 5265 21450 5285
rect 21400 5235 21450 5265
rect 21400 5215 21415 5235
rect 21435 5215 21450 5235
rect 21400 5185 21450 5215
rect 21400 5165 21415 5185
rect 21435 5165 21450 5185
rect 21400 5135 21450 5165
rect 21400 5115 21415 5135
rect 21435 5115 21450 5135
rect 21400 5085 21450 5115
rect 21400 5065 21415 5085
rect 21435 5065 21450 5085
rect 21400 5035 21450 5065
rect 21400 5015 21415 5035
rect 21435 5015 21450 5035
rect 20950 4910 20960 4940
rect 20990 4910 21000 4940
rect 20350 4810 20360 4840
rect 20390 4810 20400 4840
rect 20350 4785 20400 4810
rect 20350 4765 20365 4785
rect 20385 4765 20400 4785
rect 20350 4740 20400 4765
rect 20350 4710 20360 4740
rect 20390 4710 20400 4740
rect 20350 4685 20400 4710
rect 20350 4665 20365 4685
rect 20385 4665 20400 4685
rect 20350 4640 20400 4665
rect 20350 4610 20360 4640
rect 20390 4610 20400 4640
rect 20350 4585 20400 4610
rect 20350 4565 20365 4585
rect 20385 4565 20400 4585
rect 20350 4540 20400 4565
rect 20350 4510 20360 4540
rect 20390 4510 20400 4540
rect 20350 4485 20400 4510
rect 20350 4465 20365 4485
rect 20385 4465 20400 4485
rect 20350 4440 20400 4465
rect 20350 4410 20360 4440
rect 20390 4410 20400 4440
rect 20350 4385 20400 4410
rect 20350 4365 20365 4385
rect 20385 4365 20400 4385
rect 15550 4260 15560 4290
rect 15590 4260 15600 4290
rect 15550 4185 15600 4260
rect 17950 4200 18000 4350
rect 20350 4290 20400 4365
rect 20350 4260 20360 4290
rect 20390 4260 20400 4290
rect 15550 4165 15565 4185
rect 15585 4165 15600 4185
rect 15550 4140 15600 4165
rect 15550 4110 15560 4140
rect 15590 4110 15600 4140
rect 15550 4085 15600 4110
rect 15550 4065 15565 4085
rect 15585 4065 15600 4085
rect 15550 4040 15600 4065
rect 15550 4010 15560 4040
rect 15590 4010 15600 4040
rect 15550 3985 15600 4010
rect 15550 3965 15565 3985
rect 15585 3965 15600 3985
rect 15550 3940 15600 3965
rect 15550 3910 15560 3940
rect 15590 3910 15600 3940
rect 15550 3885 15600 3910
rect 15550 3865 15565 3885
rect 15585 3865 15600 3885
rect 15550 3840 15600 3865
rect 15550 3810 15560 3840
rect 15590 3810 15600 3840
rect 15550 3785 15600 3810
rect 15550 3765 15565 3785
rect 15585 3765 15600 3785
rect 15550 3740 15600 3765
rect 15550 3710 15560 3740
rect 15590 3710 15600 3740
rect 14950 3610 14960 3640
rect 14990 3610 15000 3640
rect 14350 3510 14360 3540
rect 14390 3510 14400 3540
rect 14350 3485 14400 3510
rect 14350 3465 14365 3485
rect 14385 3465 14400 3485
rect 14350 3440 14400 3465
rect 14350 3410 14360 3440
rect 14390 3410 14400 3440
rect 14350 3385 14400 3410
rect 14350 3365 14365 3385
rect 14385 3365 14400 3385
rect 14350 3340 14400 3365
rect 14350 3310 14360 3340
rect 14390 3310 14400 3340
rect 14350 3285 14400 3310
rect 14350 3265 14365 3285
rect 14385 3265 14400 3285
rect 14350 3240 14400 3265
rect 14350 3210 14360 3240
rect 14390 3210 14400 3240
rect 14350 3185 14400 3210
rect 14350 3165 14365 3185
rect 14385 3165 14400 3185
rect 14350 3140 14400 3165
rect 14350 3110 14360 3140
rect 14390 3110 14400 3140
rect 14350 3085 14400 3110
rect 14350 3065 14365 3085
rect 14385 3065 14400 3085
rect 13150 2960 13160 2990
rect 13190 2960 13200 2990
rect 13150 2950 13200 2960
rect 14350 2990 14400 3065
rect 14950 3535 15000 3610
rect 15100 3640 15150 3650
rect 15100 3610 15110 3640
rect 15140 3610 15150 3640
rect 15100 3600 15150 3610
rect 15400 3640 15450 3650
rect 15400 3610 15410 3640
rect 15440 3610 15450 3640
rect 15400 3600 15450 3610
rect 14950 3515 14965 3535
rect 14985 3515 15000 3535
rect 14950 3485 15000 3515
rect 14950 3465 14965 3485
rect 14985 3465 15000 3485
rect 14950 3435 15000 3465
rect 14950 3415 14965 3435
rect 14985 3415 15000 3435
rect 14950 3385 15000 3415
rect 14950 3365 14965 3385
rect 14985 3365 15000 3385
rect 14950 3335 15000 3365
rect 14950 3315 14965 3335
rect 14985 3315 15000 3335
rect 14950 3285 15000 3315
rect 14950 3265 14965 3285
rect 14985 3265 15000 3285
rect 14950 3235 15000 3265
rect 14950 3215 14965 3235
rect 14985 3215 15000 3235
rect 14950 3185 15000 3215
rect 14950 3165 14965 3185
rect 14985 3165 15000 3185
rect 14950 3135 15000 3165
rect 14950 3115 14965 3135
rect 14985 3115 15000 3135
rect 14950 3085 15000 3115
rect 14950 3065 14965 3085
rect 14985 3065 15000 3085
rect 14950 3050 15000 3065
rect 15550 3540 15600 3710
rect 16150 4185 19800 4200
rect 16150 4165 16165 4185
rect 16185 4165 16465 4185
rect 16485 4165 16765 4185
rect 16785 4165 17065 4185
rect 17085 4165 17365 4185
rect 17385 4165 18565 4185
rect 18585 4165 18865 4185
rect 18885 4165 19165 4185
rect 19185 4165 19465 4185
rect 19485 4165 19765 4185
rect 19785 4165 19800 4185
rect 16150 4150 19800 4165
rect 16150 4135 16200 4150
rect 16150 4115 16165 4135
rect 16185 4115 16200 4135
rect 16150 4085 16200 4115
rect 16450 4135 16500 4150
rect 16450 4115 16465 4135
rect 16485 4115 16500 4135
rect 16150 4065 16165 4085
rect 16185 4065 16200 4085
rect 16150 4035 16200 4065
rect 16150 4015 16165 4035
rect 16185 4015 16200 4035
rect 16150 3985 16200 4015
rect 16150 3965 16165 3985
rect 16185 3965 16200 3985
rect 16150 3935 16200 3965
rect 16150 3915 16165 3935
rect 16185 3915 16200 3935
rect 16150 3885 16200 3915
rect 16150 3865 16165 3885
rect 16185 3865 16200 3885
rect 16150 3835 16200 3865
rect 16150 3815 16165 3835
rect 16185 3815 16200 3835
rect 16150 3785 16200 3815
rect 16150 3765 16165 3785
rect 16185 3765 16200 3785
rect 16150 3735 16200 3765
rect 16150 3715 16165 3735
rect 16185 3715 16200 3735
rect 15700 3640 15750 3650
rect 15700 3610 15710 3640
rect 15740 3610 15750 3640
rect 15700 3600 15750 3610
rect 16000 3640 16050 3650
rect 16000 3610 16010 3640
rect 16040 3610 16050 3640
rect 16000 3600 16050 3610
rect 15550 3510 15560 3540
rect 15590 3510 15600 3540
rect 15550 3485 15600 3510
rect 15550 3465 15565 3485
rect 15585 3465 15600 3485
rect 15550 3440 15600 3465
rect 15550 3410 15560 3440
rect 15590 3410 15600 3440
rect 15550 3385 15600 3410
rect 15550 3365 15565 3385
rect 15585 3365 15600 3385
rect 15550 3340 15600 3365
rect 15550 3310 15560 3340
rect 15590 3310 15600 3340
rect 15550 3285 15600 3310
rect 15550 3265 15565 3285
rect 15585 3265 15600 3285
rect 15550 3240 15600 3265
rect 15550 3210 15560 3240
rect 15590 3210 15600 3240
rect 15550 3185 15600 3210
rect 15550 3165 15565 3185
rect 15585 3165 15600 3185
rect 15550 3140 15600 3165
rect 15550 3110 15560 3140
rect 15590 3110 15600 3140
rect 15550 3085 15600 3110
rect 15550 3065 15565 3085
rect 15585 3065 15600 3085
rect 14350 2960 14360 2990
rect 14390 2960 14400 2990
rect 14350 2950 14400 2960
rect 15550 2990 15600 3065
rect 16150 3535 16200 3715
rect 16300 4085 16350 4100
rect 16300 4065 16315 4085
rect 16335 4065 16350 4085
rect 16300 4035 16350 4065
rect 16300 4015 16315 4035
rect 16335 4015 16350 4035
rect 16300 3985 16350 4015
rect 16300 3965 16315 3985
rect 16335 3965 16350 3985
rect 16300 3935 16350 3965
rect 16300 3915 16315 3935
rect 16335 3915 16350 3935
rect 16300 3885 16350 3915
rect 16300 3865 16315 3885
rect 16335 3865 16350 3885
rect 16300 3835 16350 3865
rect 16300 3815 16315 3835
rect 16335 3815 16350 3835
rect 16300 3785 16350 3815
rect 16450 4085 16500 4115
rect 16750 4135 16800 4150
rect 16750 4115 16765 4135
rect 16785 4115 16800 4135
rect 16450 4065 16465 4085
rect 16485 4065 16500 4085
rect 16450 4035 16500 4065
rect 16450 4015 16465 4035
rect 16485 4015 16500 4035
rect 16450 3985 16500 4015
rect 16450 3965 16465 3985
rect 16485 3965 16500 3985
rect 16450 3935 16500 3965
rect 16450 3915 16465 3935
rect 16485 3915 16500 3935
rect 16450 3885 16500 3915
rect 16450 3865 16465 3885
rect 16485 3865 16500 3885
rect 16450 3835 16500 3865
rect 16450 3815 16465 3835
rect 16485 3815 16500 3835
rect 16450 3800 16500 3815
rect 16600 4085 16650 4100
rect 16600 4065 16615 4085
rect 16635 4065 16650 4085
rect 16600 4035 16650 4065
rect 16600 4015 16615 4035
rect 16635 4015 16650 4035
rect 16600 3985 16650 4015
rect 16600 3965 16615 3985
rect 16635 3965 16650 3985
rect 16600 3935 16650 3965
rect 16600 3915 16615 3935
rect 16635 3915 16650 3935
rect 16600 3885 16650 3915
rect 16600 3865 16615 3885
rect 16635 3865 16650 3885
rect 16600 3835 16650 3865
rect 16600 3815 16615 3835
rect 16635 3815 16650 3835
rect 16300 3765 16315 3785
rect 16335 3765 16350 3785
rect 16300 3750 16350 3765
rect 16600 3785 16650 3815
rect 16750 4085 16800 4115
rect 17050 4135 17100 4150
rect 17050 4115 17065 4135
rect 17085 4115 17100 4135
rect 16750 4065 16765 4085
rect 16785 4065 16800 4085
rect 16750 4035 16800 4065
rect 16750 4015 16765 4035
rect 16785 4015 16800 4035
rect 16750 3985 16800 4015
rect 16750 3965 16765 3985
rect 16785 3965 16800 3985
rect 16750 3935 16800 3965
rect 16750 3915 16765 3935
rect 16785 3915 16800 3935
rect 16750 3885 16800 3915
rect 16750 3865 16765 3885
rect 16785 3865 16800 3885
rect 16750 3835 16800 3865
rect 16750 3815 16765 3835
rect 16785 3815 16800 3835
rect 16750 3800 16800 3815
rect 16900 4085 16950 4100
rect 16900 4065 16915 4085
rect 16935 4065 16950 4085
rect 16900 4035 16950 4065
rect 16900 4015 16915 4035
rect 16935 4015 16950 4035
rect 16900 3985 16950 4015
rect 16900 3965 16915 3985
rect 16935 3965 16950 3985
rect 16900 3935 16950 3965
rect 16900 3915 16915 3935
rect 16935 3915 16950 3935
rect 16900 3885 16950 3915
rect 16900 3865 16915 3885
rect 16935 3865 16950 3885
rect 16900 3835 16950 3865
rect 16900 3815 16915 3835
rect 16935 3815 16950 3835
rect 16600 3765 16615 3785
rect 16635 3765 16650 3785
rect 16600 3750 16650 3765
rect 16900 3785 16950 3815
rect 17050 4085 17100 4115
rect 17350 4135 17400 4150
rect 17350 4115 17365 4135
rect 17385 4115 17400 4135
rect 17050 4065 17065 4085
rect 17085 4065 17100 4085
rect 17050 4035 17100 4065
rect 17050 4015 17065 4035
rect 17085 4015 17100 4035
rect 17050 3985 17100 4015
rect 17050 3965 17065 3985
rect 17085 3965 17100 3985
rect 17050 3935 17100 3965
rect 17050 3915 17065 3935
rect 17085 3915 17100 3935
rect 17050 3885 17100 3915
rect 17050 3865 17065 3885
rect 17085 3865 17100 3885
rect 17050 3835 17100 3865
rect 17050 3815 17065 3835
rect 17085 3815 17100 3835
rect 17050 3800 17100 3815
rect 17200 4085 17250 4100
rect 17200 4065 17215 4085
rect 17235 4065 17250 4085
rect 17200 4035 17250 4065
rect 17200 4015 17215 4035
rect 17235 4015 17250 4035
rect 17200 3985 17250 4015
rect 17200 3965 17215 3985
rect 17235 3965 17250 3985
rect 17200 3935 17250 3965
rect 17200 3915 17215 3935
rect 17235 3915 17250 3935
rect 17200 3885 17250 3915
rect 17200 3865 17215 3885
rect 17235 3865 17250 3885
rect 17200 3835 17250 3865
rect 17200 3815 17215 3835
rect 17235 3815 17250 3835
rect 16900 3765 16915 3785
rect 16935 3765 16950 3785
rect 16900 3750 16950 3765
rect 17200 3785 17250 3815
rect 17200 3765 17215 3785
rect 17235 3765 17250 3785
rect 17200 3750 17250 3765
rect 16300 3735 17250 3750
rect 16300 3715 16315 3735
rect 16335 3715 16615 3735
rect 16635 3715 16915 3735
rect 16935 3715 17215 3735
rect 17235 3715 17250 3735
rect 16300 3700 17250 3715
rect 17350 4085 17400 4115
rect 18550 4135 18600 4150
rect 18550 4115 18565 4135
rect 18585 4115 18600 4135
rect 17350 4065 17365 4085
rect 17385 4065 17400 4085
rect 17350 4035 17400 4065
rect 17350 4015 17365 4035
rect 17385 4015 17400 4035
rect 17350 3985 17400 4015
rect 17350 3965 17365 3985
rect 17385 3965 17400 3985
rect 17350 3935 17400 3965
rect 17350 3915 17365 3935
rect 17385 3915 17400 3935
rect 17350 3885 17400 3915
rect 17350 3865 17365 3885
rect 17385 3865 17400 3885
rect 17350 3835 17400 3865
rect 17350 3815 17365 3835
rect 17385 3815 17400 3835
rect 17350 3785 17400 3815
rect 17350 3765 17365 3785
rect 17385 3765 17400 3785
rect 17350 3735 17400 3765
rect 17350 3715 17365 3735
rect 17385 3715 17400 3735
rect 16300 3640 16350 3650
rect 16300 3610 16310 3640
rect 16340 3610 16350 3640
rect 16300 3600 16350 3610
rect 16600 3640 16650 3650
rect 16600 3610 16610 3640
rect 16640 3610 16650 3640
rect 16600 3600 16650 3610
rect 16750 3640 16800 3700
rect 16750 3610 16760 3640
rect 16790 3610 16800 3640
rect 16750 3550 16800 3610
rect 16900 3640 16950 3650
rect 16900 3610 16910 3640
rect 16940 3610 16950 3640
rect 16900 3600 16950 3610
rect 17200 3640 17250 3650
rect 17200 3610 17210 3640
rect 17240 3610 17250 3640
rect 17200 3600 17250 3610
rect 16150 3515 16165 3535
rect 16185 3515 16200 3535
rect 16150 3485 16200 3515
rect 16150 3465 16165 3485
rect 16185 3465 16200 3485
rect 16150 3435 16200 3465
rect 16150 3415 16165 3435
rect 16185 3415 16200 3435
rect 16150 3385 16200 3415
rect 16150 3365 16165 3385
rect 16185 3365 16200 3385
rect 16150 3335 16200 3365
rect 16150 3315 16165 3335
rect 16185 3315 16200 3335
rect 16150 3285 16200 3315
rect 16150 3265 16165 3285
rect 16185 3265 16200 3285
rect 16150 3235 16200 3265
rect 16150 3215 16165 3235
rect 16185 3215 16200 3235
rect 16150 3185 16200 3215
rect 16150 3165 16165 3185
rect 16185 3165 16200 3185
rect 16150 3135 16200 3165
rect 16300 3535 17250 3550
rect 16300 3515 16315 3535
rect 16335 3515 16615 3535
rect 16635 3515 16915 3535
rect 16935 3515 17215 3535
rect 17235 3515 17250 3535
rect 16300 3500 17250 3515
rect 16300 3485 16350 3500
rect 16300 3465 16315 3485
rect 16335 3465 16350 3485
rect 16300 3435 16350 3465
rect 16600 3485 16650 3500
rect 16600 3465 16615 3485
rect 16635 3465 16650 3485
rect 16300 3415 16315 3435
rect 16335 3415 16350 3435
rect 16300 3385 16350 3415
rect 16300 3365 16315 3385
rect 16335 3365 16350 3385
rect 16300 3335 16350 3365
rect 16300 3315 16315 3335
rect 16335 3315 16350 3335
rect 16300 3285 16350 3315
rect 16300 3265 16315 3285
rect 16335 3265 16350 3285
rect 16300 3235 16350 3265
rect 16300 3215 16315 3235
rect 16335 3215 16350 3235
rect 16300 3185 16350 3215
rect 16300 3165 16315 3185
rect 16335 3165 16350 3185
rect 16300 3150 16350 3165
rect 16450 3435 16500 3450
rect 16450 3415 16465 3435
rect 16485 3415 16500 3435
rect 16450 3385 16500 3415
rect 16450 3365 16465 3385
rect 16485 3365 16500 3385
rect 16450 3335 16500 3365
rect 16450 3315 16465 3335
rect 16485 3315 16500 3335
rect 16450 3285 16500 3315
rect 16450 3265 16465 3285
rect 16485 3265 16500 3285
rect 16450 3235 16500 3265
rect 16450 3215 16465 3235
rect 16485 3215 16500 3235
rect 16450 3185 16500 3215
rect 16450 3165 16465 3185
rect 16485 3165 16500 3185
rect 16150 3115 16165 3135
rect 16185 3115 16200 3135
rect 16150 3100 16200 3115
rect 16450 3135 16500 3165
rect 16600 3435 16650 3465
rect 16900 3485 16950 3500
rect 16900 3465 16915 3485
rect 16935 3465 16950 3485
rect 16600 3415 16615 3435
rect 16635 3415 16650 3435
rect 16600 3385 16650 3415
rect 16600 3365 16615 3385
rect 16635 3365 16650 3385
rect 16600 3335 16650 3365
rect 16600 3315 16615 3335
rect 16635 3315 16650 3335
rect 16600 3285 16650 3315
rect 16600 3265 16615 3285
rect 16635 3265 16650 3285
rect 16600 3235 16650 3265
rect 16600 3215 16615 3235
rect 16635 3215 16650 3235
rect 16600 3185 16650 3215
rect 16600 3165 16615 3185
rect 16635 3165 16650 3185
rect 16600 3150 16650 3165
rect 16750 3435 16800 3450
rect 16750 3415 16765 3435
rect 16785 3415 16800 3435
rect 16750 3385 16800 3415
rect 16750 3365 16765 3385
rect 16785 3365 16800 3385
rect 16750 3335 16800 3365
rect 16750 3315 16765 3335
rect 16785 3315 16800 3335
rect 16750 3285 16800 3315
rect 16750 3265 16765 3285
rect 16785 3265 16800 3285
rect 16750 3235 16800 3265
rect 16750 3215 16765 3235
rect 16785 3215 16800 3235
rect 16750 3185 16800 3215
rect 16750 3165 16765 3185
rect 16785 3165 16800 3185
rect 16450 3115 16465 3135
rect 16485 3115 16500 3135
rect 16450 3100 16500 3115
rect 16750 3135 16800 3165
rect 16900 3435 16950 3465
rect 17200 3485 17250 3500
rect 17200 3465 17215 3485
rect 17235 3465 17250 3485
rect 16900 3415 16915 3435
rect 16935 3415 16950 3435
rect 16900 3385 16950 3415
rect 16900 3365 16915 3385
rect 16935 3365 16950 3385
rect 16900 3335 16950 3365
rect 16900 3315 16915 3335
rect 16935 3315 16950 3335
rect 16900 3285 16950 3315
rect 16900 3265 16915 3285
rect 16935 3265 16950 3285
rect 16900 3235 16950 3265
rect 16900 3215 16915 3235
rect 16935 3215 16950 3235
rect 16900 3185 16950 3215
rect 16900 3165 16915 3185
rect 16935 3165 16950 3185
rect 16900 3150 16950 3165
rect 17050 3435 17100 3450
rect 17050 3415 17065 3435
rect 17085 3415 17100 3435
rect 17050 3385 17100 3415
rect 17050 3365 17065 3385
rect 17085 3365 17100 3385
rect 17050 3335 17100 3365
rect 17050 3315 17065 3335
rect 17085 3315 17100 3335
rect 17050 3285 17100 3315
rect 17050 3265 17065 3285
rect 17085 3265 17100 3285
rect 17050 3235 17100 3265
rect 17050 3215 17065 3235
rect 17085 3215 17100 3235
rect 17050 3185 17100 3215
rect 17050 3165 17065 3185
rect 17085 3165 17100 3185
rect 16750 3115 16765 3135
rect 16785 3115 16800 3135
rect 16750 3100 16800 3115
rect 17050 3135 17100 3165
rect 17200 3435 17250 3465
rect 17200 3415 17215 3435
rect 17235 3415 17250 3435
rect 17200 3385 17250 3415
rect 17200 3365 17215 3385
rect 17235 3365 17250 3385
rect 17200 3335 17250 3365
rect 17200 3315 17215 3335
rect 17235 3315 17250 3335
rect 17200 3285 17250 3315
rect 17200 3265 17215 3285
rect 17235 3265 17250 3285
rect 17200 3235 17250 3265
rect 17200 3215 17215 3235
rect 17235 3215 17250 3235
rect 17200 3185 17250 3215
rect 17200 3165 17215 3185
rect 17235 3165 17250 3185
rect 17200 3150 17250 3165
rect 17350 3535 17400 3715
rect 17950 4085 18000 4100
rect 17950 4065 17965 4085
rect 17985 4065 18000 4085
rect 17950 4040 18000 4065
rect 17950 4010 17960 4040
rect 17990 4010 18000 4040
rect 17950 3985 18000 4010
rect 17950 3965 17965 3985
rect 17985 3965 18000 3985
rect 17950 3940 18000 3965
rect 17950 3910 17960 3940
rect 17990 3910 18000 3940
rect 17950 3885 18000 3910
rect 17950 3865 17965 3885
rect 17985 3865 18000 3885
rect 17950 3840 18000 3865
rect 17950 3810 17960 3840
rect 17990 3810 18000 3840
rect 17950 3785 18000 3810
rect 17950 3765 17965 3785
rect 17985 3765 18000 3785
rect 17950 3740 18000 3765
rect 17950 3710 17960 3740
rect 17990 3710 18000 3740
rect 17500 3640 17550 3650
rect 17500 3610 17510 3640
rect 17540 3610 17550 3640
rect 17500 3600 17550 3610
rect 17800 3640 17850 3650
rect 17800 3610 17810 3640
rect 17840 3610 17850 3640
rect 17800 3600 17850 3610
rect 17350 3515 17365 3535
rect 17385 3515 17400 3535
rect 17350 3485 17400 3515
rect 17350 3465 17365 3485
rect 17385 3465 17400 3485
rect 17350 3435 17400 3465
rect 17350 3415 17365 3435
rect 17385 3415 17400 3435
rect 17350 3385 17400 3415
rect 17350 3365 17365 3385
rect 17385 3365 17400 3385
rect 17350 3335 17400 3365
rect 17350 3315 17365 3335
rect 17385 3315 17400 3335
rect 17350 3285 17400 3315
rect 17350 3265 17365 3285
rect 17385 3265 17400 3285
rect 17350 3235 17400 3265
rect 17350 3215 17365 3235
rect 17385 3215 17400 3235
rect 17350 3185 17400 3215
rect 17350 3165 17365 3185
rect 17385 3165 17400 3185
rect 17050 3115 17065 3135
rect 17085 3115 17100 3135
rect 17050 3100 17100 3115
rect 17350 3135 17400 3165
rect 17950 3540 18000 3710
rect 18550 4085 18600 4115
rect 18850 4135 18900 4150
rect 18850 4115 18865 4135
rect 18885 4115 18900 4135
rect 18550 4065 18565 4085
rect 18585 4065 18600 4085
rect 18550 4035 18600 4065
rect 18550 4015 18565 4035
rect 18585 4015 18600 4035
rect 18550 3985 18600 4015
rect 18550 3965 18565 3985
rect 18585 3965 18600 3985
rect 18550 3935 18600 3965
rect 18550 3915 18565 3935
rect 18585 3915 18600 3935
rect 18550 3885 18600 3915
rect 18550 3865 18565 3885
rect 18585 3865 18600 3885
rect 18550 3835 18600 3865
rect 18550 3815 18565 3835
rect 18585 3815 18600 3835
rect 18550 3785 18600 3815
rect 18550 3765 18565 3785
rect 18585 3765 18600 3785
rect 18550 3735 18600 3765
rect 18550 3715 18565 3735
rect 18585 3715 18600 3735
rect 18100 3640 18150 3650
rect 18100 3610 18110 3640
rect 18140 3610 18150 3640
rect 18100 3600 18150 3610
rect 18400 3640 18450 3650
rect 18400 3610 18410 3640
rect 18440 3610 18450 3640
rect 18400 3600 18450 3610
rect 17950 3510 17960 3540
rect 17990 3510 18000 3540
rect 17950 3485 18000 3510
rect 17950 3465 17965 3485
rect 17985 3465 18000 3485
rect 17950 3440 18000 3465
rect 17950 3410 17960 3440
rect 17990 3410 18000 3440
rect 17950 3385 18000 3410
rect 17950 3365 17965 3385
rect 17985 3365 18000 3385
rect 17950 3340 18000 3365
rect 17950 3310 17960 3340
rect 17990 3310 18000 3340
rect 17950 3285 18000 3310
rect 17950 3265 17965 3285
rect 17985 3265 18000 3285
rect 17950 3240 18000 3265
rect 17950 3210 17960 3240
rect 17990 3210 18000 3240
rect 17950 3185 18000 3210
rect 17950 3165 17965 3185
rect 17985 3165 18000 3185
rect 17950 3150 18000 3165
rect 18550 3535 18600 3715
rect 18700 4085 18750 4100
rect 18700 4065 18715 4085
rect 18735 4065 18750 4085
rect 18700 4035 18750 4065
rect 18700 4015 18715 4035
rect 18735 4015 18750 4035
rect 18700 3985 18750 4015
rect 18700 3965 18715 3985
rect 18735 3965 18750 3985
rect 18700 3935 18750 3965
rect 18700 3915 18715 3935
rect 18735 3915 18750 3935
rect 18700 3885 18750 3915
rect 18700 3865 18715 3885
rect 18735 3865 18750 3885
rect 18700 3835 18750 3865
rect 18700 3815 18715 3835
rect 18735 3815 18750 3835
rect 18700 3785 18750 3815
rect 18850 4085 18900 4115
rect 19150 4135 19200 4150
rect 19150 4115 19165 4135
rect 19185 4115 19200 4135
rect 18850 4065 18865 4085
rect 18885 4065 18900 4085
rect 18850 4035 18900 4065
rect 18850 4015 18865 4035
rect 18885 4015 18900 4035
rect 18850 3985 18900 4015
rect 18850 3965 18865 3985
rect 18885 3965 18900 3985
rect 18850 3935 18900 3965
rect 18850 3915 18865 3935
rect 18885 3915 18900 3935
rect 18850 3885 18900 3915
rect 18850 3865 18865 3885
rect 18885 3865 18900 3885
rect 18850 3835 18900 3865
rect 18850 3815 18865 3835
rect 18885 3815 18900 3835
rect 18850 3800 18900 3815
rect 19000 4085 19050 4100
rect 19000 4065 19015 4085
rect 19035 4065 19050 4085
rect 19000 4035 19050 4065
rect 19000 4015 19015 4035
rect 19035 4015 19050 4035
rect 19000 3985 19050 4015
rect 19000 3965 19015 3985
rect 19035 3965 19050 3985
rect 19000 3935 19050 3965
rect 19000 3915 19015 3935
rect 19035 3915 19050 3935
rect 19000 3885 19050 3915
rect 19000 3865 19015 3885
rect 19035 3865 19050 3885
rect 19000 3835 19050 3865
rect 19000 3815 19015 3835
rect 19035 3815 19050 3835
rect 18700 3765 18715 3785
rect 18735 3765 18750 3785
rect 18700 3750 18750 3765
rect 19000 3785 19050 3815
rect 19150 4085 19200 4115
rect 19450 4135 19500 4150
rect 19450 4115 19465 4135
rect 19485 4115 19500 4135
rect 19150 4065 19165 4085
rect 19185 4065 19200 4085
rect 19150 4035 19200 4065
rect 19150 4015 19165 4035
rect 19185 4015 19200 4035
rect 19150 3985 19200 4015
rect 19150 3965 19165 3985
rect 19185 3965 19200 3985
rect 19150 3935 19200 3965
rect 19150 3915 19165 3935
rect 19185 3915 19200 3935
rect 19150 3885 19200 3915
rect 19150 3865 19165 3885
rect 19185 3865 19200 3885
rect 19150 3835 19200 3865
rect 19150 3815 19165 3835
rect 19185 3815 19200 3835
rect 19150 3800 19200 3815
rect 19300 4085 19350 4100
rect 19300 4065 19315 4085
rect 19335 4065 19350 4085
rect 19300 4035 19350 4065
rect 19300 4015 19315 4035
rect 19335 4015 19350 4035
rect 19300 3985 19350 4015
rect 19300 3965 19315 3985
rect 19335 3965 19350 3985
rect 19300 3935 19350 3965
rect 19300 3915 19315 3935
rect 19335 3915 19350 3935
rect 19300 3885 19350 3915
rect 19300 3865 19315 3885
rect 19335 3865 19350 3885
rect 19300 3835 19350 3865
rect 19300 3815 19315 3835
rect 19335 3815 19350 3835
rect 19000 3765 19015 3785
rect 19035 3765 19050 3785
rect 19000 3750 19050 3765
rect 19300 3785 19350 3815
rect 19450 4085 19500 4115
rect 19750 4135 19800 4150
rect 19750 4115 19765 4135
rect 19785 4115 19800 4135
rect 19450 4065 19465 4085
rect 19485 4065 19500 4085
rect 19450 4035 19500 4065
rect 19450 4015 19465 4035
rect 19485 4015 19500 4035
rect 19450 3985 19500 4015
rect 19450 3965 19465 3985
rect 19485 3965 19500 3985
rect 19450 3935 19500 3965
rect 19450 3915 19465 3935
rect 19485 3915 19500 3935
rect 19450 3885 19500 3915
rect 19450 3865 19465 3885
rect 19485 3865 19500 3885
rect 19450 3835 19500 3865
rect 19450 3815 19465 3835
rect 19485 3815 19500 3835
rect 19450 3800 19500 3815
rect 19600 4085 19650 4100
rect 19600 4065 19615 4085
rect 19635 4065 19650 4085
rect 19600 4035 19650 4065
rect 19600 4015 19615 4035
rect 19635 4015 19650 4035
rect 19600 3985 19650 4015
rect 19600 3965 19615 3985
rect 19635 3965 19650 3985
rect 19600 3935 19650 3965
rect 19600 3915 19615 3935
rect 19635 3915 19650 3935
rect 19600 3885 19650 3915
rect 19600 3865 19615 3885
rect 19635 3865 19650 3885
rect 19600 3835 19650 3865
rect 19600 3815 19615 3835
rect 19635 3815 19650 3835
rect 19300 3765 19315 3785
rect 19335 3765 19350 3785
rect 19300 3750 19350 3765
rect 19600 3785 19650 3815
rect 19600 3765 19615 3785
rect 19635 3765 19650 3785
rect 19600 3750 19650 3765
rect 18700 3735 19650 3750
rect 18700 3715 18715 3735
rect 18735 3715 19015 3735
rect 19035 3715 19315 3735
rect 19335 3715 19615 3735
rect 19635 3715 19650 3735
rect 18700 3700 19650 3715
rect 19750 4085 19800 4115
rect 19750 4065 19765 4085
rect 19785 4065 19800 4085
rect 19750 4035 19800 4065
rect 19750 4015 19765 4035
rect 19785 4015 19800 4035
rect 19750 3985 19800 4015
rect 19750 3965 19765 3985
rect 19785 3965 19800 3985
rect 19750 3935 19800 3965
rect 19750 3915 19765 3935
rect 19785 3915 19800 3935
rect 19750 3885 19800 3915
rect 19750 3865 19765 3885
rect 19785 3865 19800 3885
rect 19750 3835 19800 3865
rect 19750 3815 19765 3835
rect 19785 3815 19800 3835
rect 19750 3785 19800 3815
rect 19750 3765 19765 3785
rect 19785 3765 19800 3785
rect 19750 3735 19800 3765
rect 19750 3715 19765 3735
rect 19785 3715 19800 3735
rect 18700 3640 18750 3650
rect 18700 3610 18710 3640
rect 18740 3610 18750 3640
rect 18700 3600 18750 3610
rect 19000 3640 19050 3650
rect 19000 3610 19010 3640
rect 19040 3610 19050 3640
rect 19000 3600 19050 3610
rect 19150 3640 19200 3700
rect 19150 3610 19160 3640
rect 19190 3610 19200 3640
rect 19150 3550 19200 3610
rect 19300 3640 19350 3650
rect 19300 3610 19310 3640
rect 19340 3610 19350 3640
rect 19300 3600 19350 3610
rect 19600 3640 19650 3650
rect 19600 3610 19610 3640
rect 19640 3610 19650 3640
rect 19600 3600 19650 3610
rect 18550 3515 18565 3535
rect 18585 3515 18600 3535
rect 18550 3485 18600 3515
rect 18550 3465 18565 3485
rect 18585 3465 18600 3485
rect 18550 3435 18600 3465
rect 18550 3415 18565 3435
rect 18585 3415 18600 3435
rect 18550 3385 18600 3415
rect 18550 3365 18565 3385
rect 18585 3365 18600 3385
rect 18550 3335 18600 3365
rect 18550 3315 18565 3335
rect 18585 3315 18600 3335
rect 18550 3285 18600 3315
rect 18550 3265 18565 3285
rect 18585 3265 18600 3285
rect 18550 3235 18600 3265
rect 18550 3215 18565 3235
rect 18585 3215 18600 3235
rect 18550 3185 18600 3215
rect 18550 3165 18565 3185
rect 18585 3165 18600 3185
rect 17350 3115 17365 3135
rect 17385 3115 17400 3135
rect 17350 3100 17400 3115
rect 18550 3135 18600 3165
rect 18700 3535 19650 3550
rect 18700 3515 18715 3535
rect 18735 3515 19015 3535
rect 19035 3515 19315 3535
rect 19335 3515 19615 3535
rect 19635 3515 19650 3535
rect 18700 3500 19650 3515
rect 18700 3485 18750 3500
rect 18700 3465 18715 3485
rect 18735 3465 18750 3485
rect 18700 3435 18750 3465
rect 19000 3485 19050 3500
rect 19000 3465 19015 3485
rect 19035 3465 19050 3485
rect 18700 3415 18715 3435
rect 18735 3415 18750 3435
rect 18700 3385 18750 3415
rect 18700 3365 18715 3385
rect 18735 3365 18750 3385
rect 18700 3335 18750 3365
rect 18700 3315 18715 3335
rect 18735 3315 18750 3335
rect 18700 3285 18750 3315
rect 18700 3265 18715 3285
rect 18735 3265 18750 3285
rect 18700 3235 18750 3265
rect 18700 3215 18715 3235
rect 18735 3215 18750 3235
rect 18700 3185 18750 3215
rect 18700 3165 18715 3185
rect 18735 3165 18750 3185
rect 18700 3150 18750 3165
rect 18850 3435 18900 3450
rect 18850 3415 18865 3435
rect 18885 3415 18900 3435
rect 18850 3385 18900 3415
rect 18850 3365 18865 3385
rect 18885 3365 18900 3385
rect 18850 3335 18900 3365
rect 18850 3315 18865 3335
rect 18885 3315 18900 3335
rect 18850 3285 18900 3315
rect 18850 3265 18865 3285
rect 18885 3265 18900 3285
rect 18850 3235 18900 3265
rect 18850 3215 18865 3235
rect 18885 3215 18900 3235
rect 18850 3185 18900 3215
rect 18850 3165 18865 3185
rect 18885 3165 18900 3185
rect 18550 3115 18565 3135
rect 18585 3115 18600 3135
rect 18550 3100 18600 3115
rect 18850 3135 18900 3165
rect 19000 3435 19050 3465
rect 19300 3485 19350 3500
rect 19300 3465 19315 3485
rect 19335 3465 19350 3485
rect 19000 3415 19015 3435
rect 19035 3415 19050 3435
rect 19000 3385 19050 3415
rect 19000 3365 19015 3385
rect 19035 3365 19050 3385
rect 19000 3335 19050 3365
rect 19000 3315 19015 3335
rect 19035 3315 19050 3335
rect 19000 3285 19050 3315
rect 19000 3265 19015 3285
rect 19035 3265 19050 3285
rect 19000 3235 19050 3265
rect 19000 3215 19015 3235
rect 19035 3215 19050 3235
rect 19000 3185 19050 3215
rect 19000 3165 19015 3185
rect 19035 3165 19050 3185
rect 19000 3150 19050 3165
rect 19150 3435 19200 3450
rect 19150 3415 19165 3435
rect 19185 3415 19200 3435
rect 19150 3385 19200 3415
rect 19150 3365 19165 3385
rect 19185 3365 19200 3385
rect 19150 3335 19200 3365
rect 19150 3315 19165 3335
rect 19185 3315 19200 3335
rect 19150 3285 19200 3315
rect 19150 3265 19165 3285
rect 19185 3265 19200 3285
rect 19150 3235 19200 3265
rect 19150 3215 19165 3235
rect 19185 3215 19200 3235
rect 19150 3185 19200 3215
rect 19150 3165 19165 3185
rect 19185 3165 19200 3185
rect 18850 3115 18865 3135
rect 18885 3115 18900 3135
rect 18850 3100 18900 3115
rect 19150 3135 19200 3165
rect 19300 3435 19350 3465
rect 19600 3485 19650 3500
rect 19600 3465 19615 3485
rect 19635 3465 19650 3485
rect 19300 3415 19315 3435
rect 19335 3415 19350 3435
rect 19300 3385 19350 3415
rect 19300 3365 19315 3385
rect 19335 3365 19350 3385
rect 19300 3335 19350 3365
rect 19300 3315 19315 3335
rect 19335 3315 19350 3335
rect 19300 3285 19350 3315
rect 19300 3265 19315 3285
rect 19335 3265 19350 3285
rect 19300 3235 19350 3265
rect 19300 3215 19315 3235
rect 19335 3215 19350 3235
rect 19300 3185 19350 3215
rect 19300 3165 19315 3185
rect 19335 3165 19350 3185
rect 19300 3150 19350 3165
rect 19450 3435 19500 3450
rect 19450 3415 19465 3435
rect 19485 3415 19500 3435
rect 19450 3385 19500 3415
rect 19450 3365 19465 3385
rect 19485 3365 19500 3385
rect 19450 3335 19500 3365
rect 19450 3315 19465 3335
rect 19485 3315 19500 3335
rect 19450 3285 19500 3315
rect 19450 3265 19465 3285
rect 19485 3265 19500 3285
rect 19450 3235 19500 3265
rect 19450 3215 19465 3235
rect 19485 3215 19500 3235
rect 19450 3185 19500 3215
rect 19450 3165 19465 3185
rect 19485 3165 19500 3185
rect 19150 3115 19165 3135
rect 19185 3115 19200 3135
rect 19150 3100 19200 3115
rect 19450 3135 19500 3165
rect 19600 3435 19650 3465
rect 19600 3415 19615 3435
rect 19635 3415 19650 3435
rect 19600 3385 19650 3415
rect 19600 3365 19615 3385
rect 19635 3365 19650 3385
rect 19600 3335 19650 3365
rect 19600 3315 19615 3335
rect 19635 3315 19650 3335
rect 19600 3285 19650 3315
rect 19600 3265 19615 3285
rect 19635 3265 19650 3285
rect 19600 3235 19650 3265
rect 19600 3215 19615 3235
rect 19635 3215 19650 3235
rect 19600 3185 19650 3215
rect 19600 3165 19615 3185
rect 19635 3165 19650 3185
rect 19600 3150 19650 3165
rect 19750 3535 19800 3715
rect 20350 4185 20400 4260
rect 20350 4165 20365 4185
rect 20385 4165 20400 4185
rect 20350 4140 20400 4165
rect 20350 4110 20360 4140
rect 20390 4110 20400 4140
rect 20350 4085 20400 4110
rect 20350 4065 20365 4085
rect 20385 4065 20400 4085
rect 20350 4040 20400 4065
rect 20350 4010 20360 4040
rect 20390 4010 20400 4040
rect 20350 3985 20400 4010
rect 20350 3965 20365 3985
rect 20385 3965 20400 3985
rect 20350 3940 20400 3965
rect 20350 3910 20360 3940
rect 20390 3910 20400 3940
rect 20350 3885 20400 3910
rect 20350 3865 20365 3885
rect 20385 3865 20400 3885
rect 20350 3840 20400 3865
rect 20350 3810 20360 3840
rect 20390 3810 20400 3840
rect 20350 3785 20400 3810
rect 20350 3765 20365 3785
rect 20385 3765 20400 3785
rect 20350 3740 20400 3765
rect 20350 3710 20360 3740
rect 20390 3710 20400 3740
rect 19900 3640 19950 3650
rect 19900 3610 19910 3640
rect 19940 3610 19950 3640
rect 19900 3600 19950 3610
rect 20200 3640 20250 3650
rect 20200 3610 20210 3640
rect 20240 3610 20250 3640
rect 20200 3600 20250 3610
rect 19750 3515 19765 3535
rect 19785 3515 19800 3535
rect 19750 3485 19800 3515
rect 19750 3465 19765 3485
rect 19785 3465 19800 3485
rect 19750 3435 19800 3465
rect 19750 3415 19765 3435
rect 19785 3415 19800 3435
rect 19750 3385 19800 3415
rect 19750 3365 19765 3385
rect 19785 3365 19800 3385
rect 19750 3335 19800 3365
rect 19750 3315 19765 3335
rect 19785 3315 19800 3335
rect 19750 3285 19800 3315
rect 19750 3265 19765 3285
rect 19785 3265 19800 3285
rect 19750 3235 19800 3265
rect 19750 3215 19765 3235
rect 19785 3215 19800 3235
rect 19750 3185 19800 3215
rect 19750 3165 19765 3185
rect 19785 3165 19800 3185
rect 19450 3115 19465 3135
rect 19485 3115 19500 3135
rect 19450 3100 19500 3115
rect 19750 3135 19800 3165
rect 19750 3115 19765 3135
rect 19785 3115 19800 3135
rect 19750 3100 19800 3115
rect 16150 3085 19800 3100
rect 16150 3065 16165 3085
rect 16185 3065 16465 3085
rect 16485 3065 16765 3085
rect 16785 3065 17065 3085
rect 17085 3065 17365 3085
rect 17385 3065 18565 3085
rect 18585 3065 18865 3085
rect 18885 3065 19165 3085
rect 19185 3065 19465 3085
rect 19485 3065 19765 3085
rect 19785 3065 19800 3085
rect 16150 3050 19800 3065
rect 20350 3540 20400 3710
rect 20950 4835 21000 4910
rect 21100 4940 21150 4950
rect 21100 4910 21110 4940
rect 21140 4910 21150 4940
rect 21100 4900 21150 4910
rect 21400 4940 21450 5015
rect 21850 5485 21900 5500
rect 21850 5465 21865 5485
rect 21885 5465 21900 5485
rect 21850 5435 21900 5465
rect 21850 5415 21865 5435
rect 21885 5415 21900 5435
rect 21850 5385 21900 5415
rect 21850 5365 21865 5385
rect 21885 5365 21900 5385
rect 21850 5335 21900 5365
rect 21850 5315 21865 5335
rect 21885 5315 21900 5335
rect 21850 5285 21900 5315
rect 21850 5265 21865 5285
rect 21885 5265 21900 5285
rect 21850 5235 21900 5265
rect 21850 5215 21865 5235
rect 21885 5215 21900 5235
rect 21850 5185 21900 5215
rect 21850 5165 21865 5185
rect 21885 5165 21900 5185
rect 21850 5135 21900 5165
rect 21850 5115 21865 5135
rect 21885 5115 21900 5135
rect 21850 5085 21900 5115
rect 21850 5065 21865 5085
rect 21885 5065 21900 5085
rect 21850 5035 21900 5065
rect 21850 5015 21865 5035
rect 21885 5015 21900 5035
rect 21400 4910 21410 4940
rect 21440 4910 21450 4940
rect 20950 4815 20965 4835
rect 20985 4815 21000 4835
rect 20950 4785 21000 4815
rect 20950 4765 20965 4785
rect 20985 4765 21000 4785
rect 20950 4735 21000 4765
rect 20950 4715 20965 4735
rect 20985 4715 21000 4735
rect 20950 4685 21000 4715
rect 20950 4665 20965 4685
rect 20985 4665 21000 4685
rect 20950 4635 21000 4665
rect 20950 4615 20965 4635
rect 20985 4615 21000 4635
rect 20950 4585 21000 4615
rect 20950 4565 20965 4585
rect 20985 4565 21000 4585
rect 20950 4535 21000 4565
rect 20950 4515 20965 4535
rect 20985 4515 21000 4535
rect 20950 4485 21000 4515
rect 20950 4465 20965 4485
rect 20985 4465 21000 4485
rect 20950 4435 21000 4465
rect 20950 4415 20965 4435
rect 20985 4415 21000 4435
rect 20950 4385 21000 4415
rect 20950 4365 20965 4385
rect 20985 4365 21000 4385
rect 20950 4185 21000 4365
rect 20950 4165 20965 4185
rect 20985 4165 21000 4185
rect 20950 4135 21000 4165
rect 20950 4115 20965 4135
rect 20985 4115 21000 4135
rect 20950 4085 21000 4115
rect 20950 4065 20965 4085
rect 20985 4065 21000 4085
rect 20950 4035 21000 4065
rect 20950 4015 20965 4035
rect 20985 4015 21000 4035
rect 20950 3985 21000 4015
rect 20950 3965 20965 3985
rect 20985 3965 21000 3985
rect 20950 3935 21000 3965
rect 20950 3915 20965 3935
rect 20985 3915 21000 3935
rect 20950 3885 21000 3915
rect 20950 3865 20965 3885
rect 20985 3865 21000 3885
rect 20950 3835 21000 3865
rect 20950 3815 20965 3835
rect 20985 3815 21000 3835
rect 20950 3785 21000 3815
rect 20950 3765 20965 3785
rect 20985 3765 21000 3785
rect 20950 3735 21000 3765
rect 20950 3715 20965 3735
rect 20985 3715 21000 3735
rect 20500 3640 20550 3650
rect 20500 3610 20510 3640
rect 20540 3610 20550 3640
rect 20500 3600 20550 3610
rect 20800 3640 20850 3650
rect 20800 3610 20810 3640
rect 20840 3610 20850 3640
rect 20800 3600 20850 3610
rect 20950 3640 21000 3715
rect 21400 4835 21450 4910
rect 21700 4940 21750 4950
rect 21700 4910 21710 4940
rect 21740 4910 21750 4940
rect 21700 4900 21750 4910
rect 21850 4940 21900 5015
rect 22450 5485 22500 5560
rect 24550 5590 24600 5600
rect 24550 5560 24560 5590
rect 24590 5560 24600 5590
rect 22450 5465 22465 5485
rect 22485 5465 22500 5485
rect 22450 5440 22500 5465
rect 22450 5410 22460 5440
rect 22490 5410 22500 5440
rect 22450 5385 22500 5410
rect 22450 5365 22465 5385
rect 22485 5365 22500 5385
rect 22450 5340 22500 5365
rect 22450 5310 22460 5340
rect 22490 5310 22500 5340
rect 22450 5285 22500 5310
rect 22450 5265 22465 5285
rect 22485 5265 22500 5285
rect 22450 5240 22500 5265
rect 22450 5210 22460 5240
rect 22490 5210 22500 5240
rect 22450 5185 22500 5210
rect 22450 5165 22465 5185
rect 22485 5165 22500 5185
rect 22450 5140 22500 5165
rect 22450 5110 22460 5140
rect 22490 5110 22500 5140
rect 22450 5085 22500 5110
rect 22450 5065 22465 5085
rect 22485 5065 22500 5085
rect 22450 5040 22500 5065
rect 22450 5010 22460 5040
rect 22490 5010 22500 5040
rect 21850 4910 21860 4940
rect 21890 4910 21900 4940
rect 21400 4815 21415 4835
rect 21435 4815 21450 4835
rect 21400 4785 21450 4815
rect 21400 4765 21415 4785
rect 21435 4765 21450 4785
rect 21400 4735 21450 4765
rect 21400 4715 21415 4735
rect 21435 4715 21450 4735
rect 21400 4685 21450 4715
rect 21400 4665 21415 4685
rect 21435 4665 21450 4685
rect 21400 4635 21450 4665
rect 21400 4615 21415 4635
rect 21435 4615 21450 4635
rect 21400 4585 21450 4615
rect 21400 4565 21415 4585
rect 21435 4565 21450 4585
rect 21400 4535 21450 4565
rect 21400 4515 21415 4535
rect 21435 4515 21450 4535
rect 21400 4485 21450 4515
rect 21400 4465 21415 4485
rect 21435 4465 21450 4485
rect 21400 4435 21450 4465
rect 21400 4415 21415 4435
rect 21435 4415 21450 4435
rect 21400 4385 21450 4415
rect 21400 4365 21415 4385
rect 21435 4365 21450 4385
rect 21400 4185 21450 4365
rect 21400 4165 21415 4185
rect 21435 4165 21450 4185
rect 21400 4135 21450 4165
rect 21400 4115 21415 4135
rect 21435 4115 21450 4135
rect 21400 4085 21450 4115
rect 21400 4065 21415 4085
rect 21435 4065 21450 4085
rect 21400 4035 21450 4065
rect 21400 4015 21415 4035
rect 21435 4015 21450 4035
rect 21400 3985 21450 4015
rect 21400 3965 21415 3985
rect 21435 3965 21450 3985
rect 21400 3935 21450 3965
rect 21400 3915 21415 3935
rect 21435 3915 21450 3935
rect 21400 3885 21450 3915
rect 21400 3865 21415 3885
rect 21435 3865 21450 3885
rect 21400 3835 21450 3865
rect 21400 3815 21415 3835
rect 21435 3815 21450 3835
rect 21400 3785 21450 3815
rect 21400 3765 21415 3785
rect 21435 3765 21450 3785
rect 21400 3735 21450 3765
rect 21400 3715 21415 3735
rect 21435 3715 21450 3735
rect 20950 3610 20960 3640
rect 20990 3610 21000 3640
rect 20350 3510 20360 3540
rect 20390 3510 20400 3540
rect 20350 3485 20400 3510
rect 20350 3465 20365 3485
rect 20385 3465 20400 3485
rect 20350 3440 20400 3465
rect 20350 3410 20360 3440
rect 20390 3410 20400 3440
rect 20350 3385 20400 3410
rect 20350 3365 20365 3385
rect 20385 3365 20400 3385
rect 20350 3340 20400 3365
rect 20350 3310 20360 3340
rect 20390 3310 20400 3340
rect 20350 3285 20400 3310
rect 20350 3265 20365 3285
rect 20385 3265 20400 3285
rect 20350 3240 20400 3265
rect 20350 3210 20360 3240
rect 20390 3210 20400 3240
rect 20350 3185 20400 3210
rect 20350 3165 20365 3185
rect 20385 3165 20400 3185
rect 20350 3140 20400 3165
rect 20350 3110 20360 3140
rect 20390 3110 20400 3140
rect 20350 3085 20400 3110
rect 20350 3065 20365 3085
rect 20385 3065 20400 3085
rect 15550 2960 15560 2990
rect 15590 2960 15600 2990
rect 15550 2950 15600 2960
rect 20350 2990 20400 3065
rect 20950 3535 21000 3610
rect 21100 3640 21150 3650
rect 21100 3610 21110 3640
rect 21140 3610 21150 3640
rect 21100 3600 21150 3610
rect 21400 3640 21450 3715
rect 21850 4835 21900 4910
rect 22000 4940 22050 4950
rect 22000 4910 22010 4940
rect 22040 4910 22050 4940
rect 22000 4900 22050 4910
rect 22300 4940 22350 4950
rect 22300 4910 22310 4940
rect 22340 4910 22350 4940
rect 22300 4900 22350 4910
rect 21850 4815 21865 4835
rect 21885 4815 21900 4835
rect 21850 4785 21900 4815
rect 21850 4765 21865 4785
rect 21885 4765 21900 4785
rect 21850 4735 21900 4765
rect 21850 4715 21865 4735
rect 21885 4715 21900 4735
rect 21850 4685 21900 4715
rect 21850 4665 21865 4685
rect 21885 4665 21900 4685
rect 21850 4635 21900 4665
rect 21850 4615 21865 4635
rect 21885 4615 21900 4635
rect 21850 4585 21900 4615
rect 21850 4565 21865 4585
rect 21885 4565 21900 4585
rect 21850 4535 21900 4565
rect 21850 4515 21865 4535
rect 21885 4515 21900 4535
rect 21850 4485 21900 4515
rect 21850 4465 21865 4485
rect 21885 4465 21900 4485
rect 21850 4435 21900 4465
rect 21850 4415 21865 4435
rect 21885 4415 21900 4435
rect 21850 4385 21900 4415
rect 21850 4365 21865 4385
rect 21885 4365 21900 4385
rect 21850 4185 21900 4365
rect 21850 4165 21865 4185
rect 21885 4165 21900 4185
rect 21850 4135 21900 4165
rect 21850 4115 21865 4135
rect 21885 4115 21900 4135
rect 21850 4085 21900 4115
rect 21850 4065 21865 4085
rect 21885 4065 21900 4085
rect 21850 4035 21900 4065
rect 21850 4015 21865 4035
rect 21885 4015 21900 4035
rect 21850 3985 21900 4015
rect 21850 3965 21865 3985
rect 21885 3965 21900 3985
rect 21850 3935 21900 3965
rect 21850 3915 21865 3935
rect 21885 3915 21900 3935
rect 21850 3885 21900 3915
rect 21850 3865 21865 3885
rect 21885 3865 21900 3885
rect 21850 3835 21900 3865
rect 21850 3815 21865 3835
rect 21885 3815 21900 3835
rect 21850 3785 21900 3815
rect 21850 3765 21865 3785
rect 21885 3765 21900 3785
rect 21850 3735 21900 3765
rect 21850 3715 21865 3735
rect 21885 3715 21900 3735
rect 21400 3610 21410 3640
rect 21440 3610 21450 3640
rect 20950 3515 20965 3535
rect 20985 3515 21000 3535
rect 20950 3485 21000 3515
rect 20950 3465 20965 3485
rect 20985 3465 21000 3485
rect 20950 3435 21000 3465
rect 20950 3415 20965 3435
rect 20985 3415 21000 3435
rect 20950 3385 21000 3415
rect 20950 3365 20965 3385
rect 20985 3365 21000 3385
rect 20950 3335 21000 3365
rect 20950 3315 20965 3335
rect 20985 3315 21000 3335
rect 20950 3285 21000 3315
rect 20950 3265 20965 3285
rect 20985 3265 21000 3285
rect 20950 3235 21000 3265
rect 20950 3215 20965 3235
rect 20985 3215 21000 3235
rect 20950 3185 21000 3215
rect 20950 3165 20965 3185
rect 20985 3165 21000 3185
rect 20950 3135 21000 3165
rect 20950 3115 20965 3135
rect 20985 3115 21000 3135
rect 20950 3085 21000 3115
rect 20950 3065 20965 3085
rect 20985 3065 21000 3085
rect 20950 3050 21000 3065
rect 21400 3535 21450 3610
rect 21700 3640 21750 3650
rect 21700 3610 21710 3640
rect 21740 3610 21750 3640
rect 21700 3600 21750 3610
rect 21850 3640 21900 3715
rect 22450 4840 22500 5010
rect 23050 5485 23100 5500
rect 23050 5465 23065 5485
rect 23085 5465 23100 5485
rect 23050 5435 23100 5465
rect 23050 5415 23065 5435
rect 23085 5415 23100 5435
rect 23050 5385 23100 5415
rect 23050 5365 23065 5385
rect 23085 5365 23100 5385
rect 23050 5335 23100 5365
rect 23050 5315 23065 5335
rect 23085 5315 23100 5335
rect 23050 5285 23100 5315
rect 23050 5265 23065 5285
rect 23085 5265 23100 5285
rect 23050 5235 23100 5265
rect 23050 5215 23065 5235
rect 23085 5215 23100 5235
rect 23050 5185 23100 5215
rect 23050 5165 23065 5185
rect 23085 5165 23100 5185
rect 23050 5135 23100 5165
rect 23050 5115 23065 5135
rect 23085 5115 23100 5135
rect 23050 5085 23100 5115
rect 23050 5065 23065 5085
rect 23085 5065 23100 5085
rect 23050 5035 23100 5065
rect 23050 5015 23065 5035
rect 23085 5015 23100 5035
rect 22600 4940 22650 4950
rect 22600 4910 22610 4940
rect 22640 4910 22650 4940
rect 22600 4900 22650 4910
rect 22900 4940 22950 4950
rect 22900 4910 22910 4940
rect 22940 4910 22950 4940
rect 22900 4900 22950 4910
rect 23050 4940 23100 5015
rect 23500 5485 23550 5500
rect 23500 5465 23515 5485
rect 23535 5465 23550 5485
rect 23500 5435 23550 5465
rect 23500 5415 23515 5435
rect 23535 5415 23550 5435
rect 23500 5385 23550 5415
rect 23500 5365 23515 5385
rect 23535 5365 23550 5385
rect 23500 5335 23550 5365
rect 23500 5315 23515 5335
rect 23535 5315 23550 5335
rect 23500 5285 23550 5315
rect 23500 5265 23515 5285
rect 23535 5265 23550 5285
rect 23500 5235 23550 5265
rect 23500 5215 23515 5235
rect 23535 5215 23550 5235
rect 23500 5185 23550 5215
rect 23500 5165 23515 5185
rect 23535 5165 23550 5185
rect 23500 5135 23550 5165
rect 23500 5115 23515 5135
rect 23535 5115 23550 5135
rect 23500 5085 23550 5115
rect 23500 5065 23515 5085
rect 23535 5065 23550 5085
rect 23500 5035 23550 5065
rect 23500 5015 23515 5035
rect 23535 5015 23550 5035
rect 23050 4910 23060 4940
rect 23090 4910 23100 4940
rect 22450 4810 22460 4840
rect 22490 4810 22500 4840
rect 22450 4785 22500 4810
rect 22450 4765 22465 4785
rect 22485 4765 22500 4785
rect 22450 4740 22500 4765
rect 22450 4710 22460 4740
rect 22490 4710 22500 4740
rect 22450 4685 22500 4710
rect 22450 4665 22465 4685
rect 22485 4665 22500 4685
rect 22450 4640 22500 4665
rect 22450 4610 22460 4640
rect 22490 4610 22500 4640
rect 22450 4585 22500 4610
rect 22450 4565 22465 4585
rect 22485 4565 22500 4585
rect 22450 4540 22500 4565
rect 22450 4510 22460 4540
rect 22490 4510 22500 4540
rect 22450 4485 22500 4510
rect 22450 4465 22465 4485
rect 22485 4465 22500 4485
rect 22450 4440 22500 4465
rect 22450 4410 22460 4440
rect 22490 4410 22500 4440
rect 22450 4385 22500 4410
rect 22450 4365 22465 4385
rect 22485 4365 22500 4385
rect 22450 4290 22500 4365
rect 22450 4260 22460 4290
rect 22490 4260 22500 4290
rect 22450 4185 22500 4260
rect 22450 4165 22465 4185
rect 22485 4165 22500 4185
rect 22450 4140 22500 4165
rect 22450 4110 22460 4140
rect 22490 4110 22500 4140
rect 22450 4085 22500 4110
rect 22450 4065 22465 4085
rect 22485 4065 22500 4085
rect 22450 4040 22500 4065
rect 22450 4010 22460 4040
rect 22490 4010 22500 4040
rect 22450 3985 22500 4010
rect 22450 3965 22465 3985
rect 22485 3965 22500 3985
rect 22450 3940 22500 3965
rect 22450 3910 22460 3940
rect 22490 3910 22500 3940
rect 22450 3885 22500 3910
rect 22450 3865 22465 3885
rect 22485 3865 22500 3885
rect 22450 3840 22500 3865
rect 22450 3810 22460 3840
rect 22490 3810 22500 3840
rect 22450 3785 22500 3810
rect 22450 3765 22465 3785
rect 22485 3765 22500 3785
rect 22450 3740 22500 3765
rect 22450 3710 22460 3740
rect 22490 3710 22500 3740
rect 21850 3610 21860 3640
rect 21890 3610 21900 3640
rect 21400 3515 21415 3535
rect 21435 3515 21450 3535
rect 21400 3485 21450 3515
rect 21400 3465 21415 3485
rect 21435 3465 21450 3485
rect 21400 3435 21450 3465
rect 21400 3415 21415 3435
rect 21435 3415 21450 3435
rect 21400 3385 21450 3415
rect 21400 3365 21415 3385
rect 21435 3365 21450 3385
rect 21400 3335 21450 3365
rect 21400 3315 21415 3335
rect 21435 3315 21450 3335
rect 21400 3285 21450 3315
rect 21400 3265 21415 3285
rect 21435 3265 21450 3285
rect 21400 3235 21450 3265
rect 21400 3215 21415 3235
rect 21435 3215 21450 3235
rect 21400 3185 21450 3215
rect 21400 3165 21415 3185
rect 21435 3165 21450 3185
rect 21400 3135 21450 3165
rect 21400 3115 21415 3135
rect 21435 3115 21450 3135
rect 21400 3085 21450 3115
rect 21400 3065 21415 3085
rect 21435 3065 21450 3085
rect 21400 3050 21450 3065
rect 21850 3535 21900 3610
rect 22000 3640 22050 3650
rect 22000 3610 22010 3640
rect 22040 3610 22050 3640
rect 22000 3600 22050 3610
rect 22300 3640 22350 3650
rect 22300 3610 22310 3640
rect 22340 3610 22350 3640
rect 22300 3600 22350 3610
rect 21850 3515 21865 3535
rect 21885 3515 21900 3535
rect 21850 3485 21900 3515
rect 21850 3465 21865 3485
rect 21885 3465 21900 3485
rect 21850 3435 21900 3465
rect 21850 3415 21865 3435
rect 21885 3415 21900 3435
rect 21850 3385 21900 3415
rect 21850 3365 21865 3385
rect 21885 3365 21900 3385
rect 21850 3335 21900 3365
rect 21850 3315 21865 3335
rect 21885 3315 21900 3335
rect 21850 3285 21900 3315
rect 21850 3265 21865 3285
rect 21885 3265 21900 3285
rect 21850 3235 21900 3265
rect 21850 3215 21865 3235
rect 21885 3215 21900 3235
rect 21850 3185 21900 3215
rect 21850 3165 21865 3185
rect 21885 3165 21900 3185
rect 21850 3135 21900 3165
rect 21850 3115 21865 3135
rect 21885 3115 21900 3135
rect 21850 3085 21900 3115
rect 21850 3065 21865 3085
rect 21885 3065 21900 3085
rect 21850 3050 21900 3065
rect 22450 3540 22500 3710
rect 23050 4835 23100 4910
rect 23200 4940 23250 4950
rect 23200 4910 23210 4940
rect 23240 4910 23250 4940
rect 23200 4900 23250 4910
rect 23350 4940 23400 4950
rect 23350 4910 23360 4940
rect 23390 4910 23400 4940
rect 23350 4900 23400 4910
rect 23500 4940 23550 5015
rect 23950 5485 24000 5500
rect 23950 5465 23965 5485
rect 23985 5465 24000 5485
rect 23950 5435 24000 5465
rect 23950 5415 23965 5435
rect 23985 5415 24000 5435
rect 23950 5385 24000 5415
rect 23950 5365 23965 5385
rect 23985 5365 24000 5385
rect 23950 5335 24000 5365
rect 23950 5315 23965 5335
rect 23985 5315 24000 5335
rect 23950 5285 24000 5315
rect 23950 5265 23965 5285
rect 23985 5265 24000 5285
rect 23950 5235 24000 5265
rect 23950 5215 23965 5235
rect 23985 5215 24000 5235
rect 23950 5185 24000 5215
rect 23950 5165 23965 5185
rect 23985 5165 24000 5185
rect 23950 5135 24000 5165
rect 23950 5115 23965 5135
rect 23985 5115 24000 5135
rect 23950 5085 24000 5115
rect 23950 5065 23965 5085
rect 23985 5065 24000 5085
rect 23950 5035 24000 5065
rect 23950 5015 23965 5035
rect 23985 5015 24000 5035
rect 23500 4910 23510 4940
rect 23540 4910 23550 4940
rect 23050 4815 23065 4835
rect 23085 4815 23100 4835
rect 23050 4785 23100 4815
rect 23050 4765 23065 4785
rect 23085 4765 23100 4785
rect 23050 4735 23100 4765
rect 23050 4715 23065 4735
rect 23085 4715 23100 4735
rect 23050 4685 23100 4715
rect 23050 4665 23065 4685
rect 23085 4665 23100 4685
rect 23050 4635 23100 4665
rect 23050 4615 23065 4635
rect 23085 4615 23100 4635
rect 23050 4585 23100 4615
rect 23050 4565 23065 4585
rect 23085 4565 23100 4585
rect 23050 4535 23100 4565
rect 23050 4515 23065 4535
rect 23085 4515 23100 4535
rect 23050 4485 23100 4515
rect 23050 4465 23065 4485
rect 23085 4465 23100 4485
rect 23050 4435 23100 4465
rect 23050 4415 23065 4435
rect 23085 4415 23100 4435
rect 23050 4385 23100 4415
rect 23050 4365 23065 4385
rect 23085 4365 23100 4385
rect 23050 4185 23100 4365
rect 23050 4165 23065 4185
rect 23085 4165 23100 4185
rect 23050 4135 23100 4165
rect 23050 4115 23065 4135
rect 23085 4115 23100 4135
rect 23050 4085 23100 4115
rect 23050 4065 23065 4085
rect 23085 4065 23100 4085
rect 23050 4035 23100 4065
rect 23050 4015 23065 4035
rect 23085 4015 23100 4035
rect 23050 3985 23100 4015
rect 23050 3965 23065 3985
rect 23085 3965 23100 3985
rect 23050 3935 23100 3965
rect 23050 3915 23065 3935
rect 23085 3915 23100 3935
rect 23050 3885 23100 3915
rect 23050 3865 23065 3885
rect 23085 3865 23100 3885
rect 23050 3835 23100 3865
rect 23050 3815 23065 3835
rect 23085 3815 23100 3835
rect 23050 3785 23100 3815
rect 23050 3765 23065 3785
rect 23085 3765 23100 3785
rect 23050 3735 23100 3765
rect 23050 3715 23065 3735
rect 23085 3715 23100 3735
rect 22600 3640 22650 3650
rect 22600 3610 22610 3640
rect 22640 3610 22650 3640
rect 22600 3600 22650 3610
rect 22900 3640 22950 3650
rect 22900 3610 22910 3640
rect 22940 3610 22950 3640
rect 22900 3600 22950 3610
rect 23050 3640 23100 3715
rect 23500 4835 23550 4910
rect 23650 4940 23700 4950
rect 23650 4910 23660 4940
rect 23690 4910 23700 4940
rect 23650 4900 23700 4910
rect 23800 4940 23850 4950
rect 23800 4910 23810 4940
rect 23840 4910 23850 4940
rect 23800 4900 23850 4910
rect 23950 4940 24000 5015
rect 24550 5485 24600 5560
rect 26650 5590 26700 5600
rect 26650 5560 26660 5590
rect 26690 5560 26700 5590
rect 24550 5465 24565 5485
rect 24585 5465 24600 5485
rect 24550 5440 24600 5465
rect 24550 5410 24560 5440
rect 24590 5410 24600 5440
rect 24550 5385 24600 5410
rect 24550 5365 24565 5385
rect 24585 5365 24600 5385
rect 24550 5340 24600 5365
rect 24550 5310 24560 5340
rect 24590 5310 24600 5340
rect 24550 5285 24600 5310
rect 24550 5265 24565 5285
rect 24585 5265 24600 5285
rect 24550 5240 24600 5265
rect 24550 5210 24560 5240
rect 24590 5210 24600 5240
rect 24550 5185 24600 5210
rect 24550 5165 24565 5185
rect 24585 5165 24600 5185
rect 24550 5140 24600 5165
rect 24550 5110 24560 5140
rect 24590 5110 24600 5140
rect 24550 5085 24600 5110
rect 24550 5065 24565 5085
rect 24585 5065 24600 5085
rect 24550 5040 24600 5065
rect 24550 5010 24560 5040
rect 24590 5010 24600 5040
rect 23950 4910 23960 4940
rect 23990 4910 24000 4940
rect 23500 4815 23515 4835
rect 23535 4815 23550 4835
rect 23500 4785 23550 4815
rect 23500 4765 23515 4785
rect 23535 4765 23550 4785
rect 23500 4735 23550 4765
rect 23500 4715 23515 4735
rect 23535 4715 23550 4735
rect 23500 4685 23550 4715
rect 23500 4665 23515 4685
rect 23535 4665 23550 4685
rect 23500 4635 23550 4665
rect 23500 4615 23515 4635
rect 23535 4615 23550 4635
rect 23500 4585 23550 4615
rect 23500 4565 23515 4585
rect 23535 4565 23550 4585
rect 23500 4535 23550 4565
rect 23500 4515 23515 4535
rect 23535 4515 23550 4535
rect 23500 4485 23550 4515
rect 23500 4465 23515 4485
rect 23535 4465 23550 4485
rect 23500 4435 23550 4465
rect 23500 4415 23515 4435
rect 23535 4415 23550 4435
rect 23500 4385 23550 4415
rect 23500 4365 23515 4385
rect 23535 4365 23550 4385
rect 23500 4185 23550 4365
rect 23500 4165 23515 4185
rect 23535 4165 23550 4185
rect 23500 4135 23550 4165
rect 23500 4115 23515 4135
rect 23535 4115 23550 4135
rect 23500 4085 23550 4115
rect 23500 4065 23515 4085
rect 23535 4065 23550 4085
rect 23500 4035 23550 4065
rect 23500 4015 23515 4035
rect 23535 4015 23550 4035
rect 23500 3985 23550 4015
rect 23500 3965 23515 3985
rect 23535 3965 23550 3985
rect 23500 3935 23550 3965
rect 23500 3915 23515 3935
rect 23535 3915 23550 3935
rect 23500 3885 23550 3915
rect 23500 3865 23515 3885
rect 23535 3865 23550 3885
rect 23500 3835 23550 3865
rect 23500 3815 23515 3835
rect 23535 3815 23550 3835
rect 23500 3785 23550 3815
rect 23500 3765 23515 3785
rect 23535 3765 23550 3785
rect 23500 3735 23550 3765
rect 23500 3715 23515 3735
rect 23535 3715 23550 3735
rect 23050 3610 23060 3640
rect 23090 3610 23100 3640
rect 22450 3510 22460 3540
rect 22490 3510 22500 3540
rect 22450 3485 22500 3510
rect 22450 3465 22465 3485
rect 22485 3465 22500 3485
rect 22450 3440 22500 3465
rect 22450 3410 22460 3440
rect 22490 3410 22500 3440
rect 22450 3385 22500 3410
rect 22450 3365 22465 3385
rect 22485 3365 22500 3385
rect 22450 3340 22500 3365
rect 22450 3310 22460 3340
rect 22490 3310 22500 3340
rect 22450 3285 22500 3310
rect 22450 3265 22465 3285
rect 22485 3265 22500 3285
rect 22450 3240 22500 3265
rect 22450 3210 22460 3240
rect 22490 3210 22500 3240
rect 22450 3185 22500 3210
rect 22450 3165 22465 3185
rect 22485 3165 22500 3185
rect 22450 3140 22500 3165
rect 22450 3110 22460 3140
rect 22490 3110 22500 3140
rect 22450 3085 22500 3110
rect 22450 3065 22465 3085
rect 22485 3065 22500 3085
rect 22450 3000 22500 3065
rect 23050 3535 23100 3610
rect 23200 3640 23250 3650
rect 23200 3610 23210 3640
rect 23240 3610 23250 3640
rect 23200 3600 23250 3610
rect 23350 3640 23400 3650
rect 23350 3610 23360 3640
rect 23390 3610 23400 3640
rect 23350 3600 23400 3610
rect 23500 3640 23550 3715
rect 23950 4835 24000 4910
rect 24100 4940 24150 4950
rect 24100 4910 24110 4940
rect 24140 4910 24150 4940
rect 24100 4900 24150 4910
rect 24400 4940 24450 4950
rect 24400 4910 24410 4940
rect 24440 4910 24450 4940
rect 24400 4900 24450 4910
rect 23950 4815 23965 4835
rect 23985 4815 24000 4835
rect 23950 4785 24000 4815
rect 23950 4765 23965 4785
rect 23985 4765 24000 4785
rect 23950 4735 24000 4765
rect 23950 4715 23965 4735
rect 23985 4715 24000 4735
rect 23950 4685 24000 4715
rect 23950 4665 23965 4685
rect 23985 4665 24000 4685
rect 23950 4635 24000 4665
rect 23950 4615 23965 4635
rect 23985 4615 24000 4635
rect 23950 4585 24000 4615
rect 23950 4565 23965 4585
rect 23985 4565 24000 4585
rect 23950 4535 24000 4565
rect 23950 4515 23965 4535
rect 23985 4515 24000 4535
rect 23950 4485 24000 4515
rect 23950 4465 23965 4485
rect 23985 4465 24000 4485
rect 23950 4435 24000 4465
rect 23950 4415 23965 4435
rect 23985 4415 24000 4435
rect 23950 4385 24000 4415
rect 23950 4365 23965 4385
rect 23985 4365 24000 4385
rect 23950 4185 24000 4365
rect 23950 4165 23965 4185
rect 23985 4165 24000 4185
rect 23950 4135 24000 4165
rect 23950 4115 23965 4135
rect 23985 4115 24000 4135
rect 23950 4085 24000 4115
rect 23950 4065 23965 4085
rect 23985 4065 24000 4085
rect 23950 4035 24000 4065
rect 23950 4015 23965 4035
rect 23985 4015 24000 4035
rect 23950 3985 24000 4015
rect 23950 3965 23965 3985
rect 23985 3965 24000 3985
rect 23950 3935 24000 3965
rect 23950 3915 23965 3935
rect 23985 3915 24000 3935
rect 23950 3885 24000 3915
rect 23950 3865 23965 3885
rect 23985 3865 24000 3885
rect 23950 3835 24000 3865
rect 23950 3815 23965 3835
rect 23985 3815 24000 3835
rect 23950 3785 24000 3815
rect 23950 3765 23965 3785
rect 23985 3765 24000 3785
rect 23950 3735 24000 3765
rect 23950 3715 23965 3735
rect 23985 3715 24000 3735
rect 23500 3610 23510 3640
rect 23540 3610 23550 3640
rect 23050 3515 23065 3535
rect 23085 3515 23100 3535
rect 23050 3485 23100 3515
rect 23050 3465 23065 3485
rect 23085 3465 23100 3485
rect 23050 3435 23100 3465
rect 23050 3415 23065 3435
rect 23085 3415 23100 3435
rect 23050 3385 23100 3415
rect 23050 3365 23065 3385
rect 23085 3365 23100 3385
rect 23050 3335 23100 3365
rect 23050 3315 23065 3335
rect 23085 3315 23100 3335
rect 23050 3285 23100 3315
rect 23050 3265 23065 3285
rect 23085 3265 23100 3285
rect 23050 3235 23100 3265
rect 23050 3215 23065 3235
rect 23085 3215 23100 3235
rect 23050 3185 23100 3215
rect 23050 3165 23065 3185
rect 23085 3165 23100 3185
rect 23050 3135 23100 3165
rect 23050 3115 23065 3135
rect 23085 3115 23100 3135
rect 23050 3085 23100 3115
rect 23050 3065 23065 3085
rect 23085 3065 23100 3085
rect 23050 3050 23100 3065
rect 23500 3535 23550 3610
rect 23650 3640 23700 3650
rect 23650 3610 23660 3640
rect 23690 3610 23700 3640
rect 23650 3600 23700 3610
rect 23800 3640 23850 3650
rect 23800 3610 23810 3640
rect 23840 3610 23850 3640
rect 23800 3600 23850 3610
rect 23950 3640 24000 3715
rect 24550 4840 24600 5010
rect 25150 5485 25200 5500
rect 25150 5465 25165 5485
rect 25185 5465 25200 5485
rect 25150 5435 25200 5465
rect 25150 5415 25165 5435
rect 25185 5415 25200 5435
rect 25150 5385 25200 5415
rect 25150 5365 25165 5385
rect 25185 5365 25200 5385
rect 25150 5335 25200 5365
rect 25150 5315 25165 5335
rect 25185 5315 25200 5335
rect 25150 5285 25200 5315
rect 25150 5265 25165 5285
rect 25185 5265 25200 5285
rect 25150 5235 25200 5265
rect 25150 5215 25165 5235
rect 25185 5215 25200 5235
rect 25150 5185 25200 5215
rect 25150 5165 25165 5185
rect 25185 5165 25200 5185
rect 25150 5135 25200 5165
rect 25150 5115 25165 5135
rect 25185 5115 25200 5135
rect 25150 5085 25200 5115
rect 25150 5065 25165 5085
rect 25185 5065 25200 5085
rect 25150 5035 25200 5065
rect 25150 5015 25165 5035
rect 25185 5015 25200 5035
rect 24700 4940 24750 4950
rect 24700 4910 24710 4940
rect 24740 4910 24750 4940
rect 24700 4900 24750 4910
rect 25000 4940 25050 4950
rect 25000 4910 25010 4940
rect 25040 4910 25050 4940
rect 25000 4900 25050 4910
rect 24550 4810 24560 4840
rect 24590 4810 24600 4840
rect 24550 4785 24600 4810
rect 24550 4765 24565 4785
rect 24585 4765 24600 4785
rect 24550 4740 24600 4765
rect 24550 4710 24560 4740
rect 24590 4710 24600 4740
rect 24550 4685 24600 4710
rect 24550 4665 24565 4685
rect 24585 4665 24600 4685
rect 24550 4640 24600 4665
rect 24550 4610 24560 4640
rect 24590 4610 24600 4640
rect 24550 4585 24600 4610
rect 24550 4565 24565 4585
rect 24585 4565 24600 4585
rect 24550 4540 24600 4565
rect 24550 4510 24560 4540
rect 24590 4510 24600 4540
rect 24550 4485 24600 4510
rect 24550 4465 24565 4485
rect 24585 4465 24600 4485
rect 24550 4440 24600 4465
rect 24550 4410 24560 4440
rect 24590 4410 24600 4440
rect 24550 4385 24600 4410
rect 24550 4365 24565 4385
rect 24585 4365 24600 4385
rect 24550 4290 24600 4365
rect 25150 4835 25200 5015
rect 25600 5485 25650 5500
rect 25600 5465 25615 5485
rect 25635 5465 25650 5485
rect 25600 5435 25650 5465
rect 25600 5415 25615 5435
rect 25635 5415 25650 5435
rect 25600 5385 25650 5415
rect 25600 5365 25615 5385
rect 25635 5365 25650 5385
rect 25600 5335 25650 5365
rect 25600 5315 25615 5335
rect 25635 5315 25650 5335
rect 25600 5285 25650 5315
rect 25600 5265 25615 5285
rect 25635 5265 25650 5285
rect 25600 5235 25650 5265
rect 25600 5215 25615 5235
rect 25635 5215 25650 5235
rect 25600 5185 25650 5215
rect 25600 5165 25615 5185
rect 25635 5165 25650 5185
rect 25600 5135 25650 5165
rect 25600 5115 25615 5135
rect 25635 5115 25650 5135
rect 25600 5085 25650 5115
rect 25600 5065 25615 5085
rect 25635 5065 25650 5085
rect 25600 5035 25650 5065
rect 25600 5015 25615 5035
rect 25635 5015 25650 5035
rect 25450 4940 25500 4950
rect 25450 4910 25460 4940
rect 25490 4910 25500 4940
rect 25450 4900 25500 4910
rect 25600 4940 25650 5015
rect 26050 5485 26100 5500
rect 26050 5465 26065 5485
rect 26085 5465 26100 5485
rect 26050 5435 26100 5465
rect 26050 5415 26065 5435
rect 26085 5415 26100 5435
rect 26050 5385 26100 5415
rect 26050 5365 26065 5385
rect 26085 5365 26100 5385
rect 26050 5335 26100 5365
rect 26050 5315 26065 5335
rect 26085 5315 26100 5335
rect 26050 5285 26100 5315
rect 26050 5265 26065 5285
rect 26085 5265 26100 5285
rect 26050 5235 26100 5265
rect 26050 5215 26065 5235
rect 26085 5215 26100 5235
rect 26050 5185 26100 5215
rect 26050 5165 26065 5185
rect 26085 5165 26100 5185
rect 26050 5135 26100 5165
rect 26050 5115 26065 5135
rect 26085 5115 26100 5135
rect 26050 5085 26100 5115
rect 26050 5065 26065 5085
rect 26085 5065 26100 5085
rect 26050 5035 26100 5065
rect 26050 5015 26065 5035
rect 26085 5015 26100 5035
rect 25600 4910 25610 4940
rect 25640 4910 25650 4940
rect 25150 4815 25165 4835
rect 25185 4815 25200 4835
rect 25150 4785 25200 4815
rect 25150 4765 25165 4785
rect 25185 4765 25200 4785
rect 25150 4735 25200 4765
rect 25150 4715 25165 4735
rect 25185 4715 25200 4735
rect 25150 4685 25200 4715
rect 25150 4665 25165 4685
rect 25185 4665 25200 4685
rect 25150 4635 25200 4665
rect 25150 4615 25165 4635
rect 25185 4615 25200 4635
rect 25150 4585 25200 4615
rect 25150 4565 25165 4585
rect 25185 4565 25200 4585
rect 25150 4535 25200 4565
rect 25150 4515 25165 4535
rect 25185 4515 25200 4535
rect 25150 4485 25200 4515
rect 25150 4465 25165 4485
rect 25185 4465 25200 4485
rect 25150 4435 25200 4465
rect 25150 4415 25165 4435
rect 25185 4415 25200 4435
rect 25150 4385 25200 4415
rect 25150 4365 25165 4385
rect 25185 4365 25200 4385
rect 25150 4350 25200 4365
rect 25600 4835 25650 4910
rect 25750 4940 25800 4950
rect 25750 4910 25760 4940
rect 25790 4910 25800 4940
rect 25750 4900 25800 4910
rect 25600 4815 25615 4835
rect 25635 4815 25650 4835
rect 25600 4785 25650 4815
rect 25600 4765 25615 4785
rect 25635 4765 25650 4785
rect 25600 4735 25650 4765
rect 25600 4715 25615 4735
rect 25635 4715 25650 4735
rect 25600 4685 25650 4715
rect 25600 4665 25615 4685
rect 25635 4665 25650 4685
rect 25600 4635 25650 4665
rect 25600 4615 25615 4635
rect 25635 4615 25650 4635
rect 25600 4585 25650 4615
rect 25600 4565 25615 4585
rect 25635 4565 25650 4585
rect 25600 4535 25650 4565
rect 25600 4515 25615 4535
rect 25635 4515 25650 4535
rect 25600 4485 25650 4515
rect 25600 4465 25615 4485
rect 25635 4465 25650 4485
rect 25600 4435 25650 4465
rect 25600 4415 25615 4435
rect 25635 4415 25650 4435
rect 25600 4385 25650 4415
rect 25600 4365 25615 4385
rect 25635 4365 25650 4385
rect 24550 4260 24560 4290
rect 24590 4260 24600 4290
rect 24550 4185 24600 4260
rect 24550 4165 24565 4185
rect 24585 4165 24600 4185
rect 24550 4140 24600 4165
rect 24550 4110 24560 4140
rect 24590 4110 24600 4140
rect 24550 4085 24600 4110
rect 24550 4065 24565 4085
rect 24585 4065 24600 4085
rect 24550 4040 24600 4065
rect 24550 4010 24560 4040
rect 24590 4010 24600 4040
rect 24550 3985 24600 4010
rect 24550 3965 24565 3985
rect 24585 3965 24600 3985
rect 24550 3940 24600 3965
rect 24550 3910 24560 3940
rect 24590 3910 24600 3940
rect 24550 3885 24600 3910
rect 24550 3865 24565 3885
rect 24585 3865 24600 3885
rect 24550 3840 24600 3865
rect 24550 3810 24560 3840
rect 24590 3810 24600 3840
rect 24550 3785 24600 3810
rect 24550 3765 24565 3785
rect 24585 3765 24600 3785
rect 24550 3740 24600 3765
rect 24550 3710 24560 3740
rect 24590 3710 24600 3740
rect 23950 3610 23960 3640
rect 23990 3610 24000 3640
rect 23500 3515 23515 3535
rect 23535 3515 23550 3535
rect 23500 3485 23550 3515
rect 23500 3465 23515 3485
rect 23535 3465 23550 3485
rect 23500 3435 23550 3465
rect 23500 3415 23515 3435
rect 23535 3415 23550 3435
rect 23500 3385 23550 3415
rect 23500 3365 23515 3385
rect 23535 3365 23550 3385
rect 23500 3335 23550 3365
rect 23500 3315 23515 3335
rect 23535 3315 23550 3335
rect 23500 3285 23550 3315
rect 23500 3265 23515 3285
rect 23535 3265 23550 3285
rect 23500 3235 23550 3265
rect 23500 3215 23515 3235
rect 23535 3215 23550 3235
rect 23500 3185 23550 3215
rect 23500 3165 23515 3185
rect 23535 3165 23550 3185
rect 23500 3135 23550 3165
rect 23500 3115 23515 3135
rect 23535 3115 23550 3135
rect 23500 3085 23550 3115
rect 23500 3065 23515 3085
rect 23535 3065 23550 3085
rect 23500 3050 23550 3065
rect 23950 3535 24000 3610
rect 24100 3640 24150 3650
rect 24100 3610 24110 3640
rect 24140 3610 24150 3640
rect 24100 3600 24150 3610
rect 24400 3640 24450 3650
rect 24400 3610 24410 3640
rect 24440 3610 24450 3640
rect 24400 3600 24450 3610
rect 23950 3515 23965 3535
rect 23985 3515 24000 3535
rect 23950 3485 24000 3515
rect 23950 3465 23965 3485
rect 23985 3465 24000 3485
rect 23950 3435 24000 3465
rect 23950 3415 23965 3435
rect 23985 3415 24000 3435
rect 23950 3385 24000 3415
rect 23950 3365 23965 3385
rect 23985 3365 24000 3385
rect 23950 3335 24000 3365
rect 23950 3315 23965 3335
rect 23985 3315 24000 3335
rect 23950 3285 24000 3315
rect 23950 3265 23965 3285
rect 23985 3265 24000 3285
rect 23950 3235 24000 3265
rect 23950 3215 23965 3235
rect 23985 3215 24000 3235
rect 23950 3185 24000 3215
rect 23950 3165 23965 3185
rect 23985 3165 24000 3185
rect 23950 3135 24000 3165
rect 23950 3115 23965 3135
rect 23985 3115 24000 3135
rect 23950 3085 24000 3115
rect 23950 3065 23965 3085
rect 23985 3065 24000 3085
rect 23950 3050 24000 3065
rect 24550 3540 24600 3710
rect 25150 4185 25200 4200
rect 25150 4165 25165 4185
rect 25185 4165 25200 4185
rect 25150 4135 25200 4165
rect 25150 4115 25165 4135
rect 25185 4115 25200 4135
rect 25150 4085 25200 4115
rect 25150 4065 25165 4085
rect 25185 4065 25200 4085
rect 25150 4035 25200 4065
rect 25150 4015 25165 4035
rect 25185 4015 25200 4035
rect 25150 3985 25200 4015
rect 25150 3965 25165 3985
rect 25185 3965 25200 3985
rect 25150 3935 25200 3965
rect 25150 3915 25165 3935
rect 25185 3915 25200 3935
rect 25150 3885 25200 3915
rect 25150 3865 25165 3885
rect 25185 3865 25200 3885
rect 25150 3835 25200 3865
rect 25150 3815 25165 3835
rect 25185 3815 25200 3835
rect 25150 3785 25200 3815
rect 25150 3765 25165 3785
rect 25185 3765 25200 3785
rect 25150 3735 25200 3765
rect 25150 3715 25165 3735
rect 25185 3715 25200 3735
rect 24700 3640 24750 3650
rect 24700 3610 24710 3640
rect 24740 3610 24750 3640
rect 24700 3600 24750 3610
rect 25000 3640 25050 3650
rect 25000 3610 25010 3640
rect 25040 3610 25050 3640
rect 25000 3600 25050 3610
rect 24550 3510 24560 3540
rect 24590 3510 24600 3540
rect 24550 3485 24600 3510
rect 24550 3465 24565 3485
rect 24585 3465 24600 3485
rect 24550 3440 24600 3465
rect 24550 3410 24560 3440
rect 24590 3410 24600 3440
rect 24550 3385 24600 3410
rect 24550 3365 24565 3385
rect 24585 3365 24600 3385
rect 24550 3340 24600 3365
rect 24550 3310 24560 3340
rect 24590 3310 24600 3340
rect 24550 3285 24600 3310
rect 24550 3265 24565 3285
rect 24585 3265 24600 3285
rect 24550 3240 24600 3265
rect 24550 3210 24560 3240
rect 24590 3210 24600 3240
rect 24550 3185 24600 3210
rect 24550 3165 24565 3185
rect 24585 3165 24600 3185
rect 24550 3140 24600 3165
rect 24550 3110 24560 3140
rect 24590 3110 24600 3140
rect 24550 3085 24600 3110
rect 24550 3065 24565 3085
rect 24585 3065 24600 3085
rect 20350 2960 20360 2990
rect 20390 2960 20400 2990
rect 20350 2950 20400 2960
rect 24550 2990 24600 3065
rect 25150 3535 25200 3715
rect 25600 4185 25650 4365
rect 26050 4835 26100 5015
rect 26650 5485 26700 5560
rect 28150 5590 28200 5600
rect 28150 5560 28160 5590
rect 28190 5560 28200 5590
rect 26650 5465 26665 5485
rect 26685 5465 26700 5485
rect 26650 5440 26700 5465
rect 26650 5410 26660 5440
rect 26690 5410 26700 5440
rect 26650 5385 26700 5410
rect 26650 5365 26665 5385
rect 26685 5365 26700 5385
rect 26650 5340 26700 5365
rect 26650 5310 26660 5340
rect 26690 5310 26700 5340
rect 26650 5285 26700 5310
rect 26650 5265 26665 5285
rect 26685 5265 26700 5285
rect 26650 5240 26700 5265
rect 26650 5210 26660 5240
rect 26690 5210 26700 5240
rect 26650 5185 26700 5210
rect 26650 5165 26665 5185
rect 26685 5165 26700 5185
rect 26650 5140 26700 5165
rect 26650 5110 26660 5140
rect 26690 5110 26700 5140
rect 26650 5085 26700 5110
rect 26650 5065 26665 5085
rect 26685 5065 26700 5085
rect 26650 5040 26700 5065
rect 26650 5010 26660 5040
rect 26690 5010 26700 5040
rect 26200 4940 26250 4950
rect 26200 4910 26210 4940
rect 26240 4910 26250 4940
rect 26200 4900 26250 4910
rect 26500 4940 26550 4950
rect 26500 4910 26510 4940
rect 26540 4910 26550 4940
rect 26500 4900 26550 4910
rect 26050 4815 26065 4835
rect 26085 4815 26100 4835
rect 26050 4785 26100 4815
rect 26050 4765 26065 4785
rect 26085 4765 26100 4785
rect 26050 4735 26100 4765
rect 26050 4715 26065 4735
rect 26085 4715 26100 4735
rect 26050 4685 26100 4715
rect 26050 4665 26065 4685
rect 26085 4665 26100 4685
rect 26050 4635 26100 4665
rect 26050 4615 26065 4635
rect 26085 4615 26100 4635
rect 26050 4585 26100 4615
rect 26050 4565 26065 4585
rect 26085 4565 26100 4585
rect 26050 4535 26100 4565
rect 26050 4515 26065 4535
rect 26085 4515 26100 4535
rect 26050 4485 26100 4515
rect 26050 4465 26065 4485
rect 26085 4465 26100 4485
rect 26050 4435 26100 4465
rect 26050 4415 26065 4435
rect 26085 4415 26100 4435
rect 26050 4385 26100 4415
rect 26050 4365 26065 4385
rect 26085 4365 26100 4385
rect 26050 4350 26100 4365
rect 26650 4840 26700 5010
rect 27250 5485 27300 5500
rect 27250 5465 27265 5485
rect 27285 5465 27300 5485
rect 27250 5435 27300 5465
rect 27250 5415 27265 5435
rect 27285 5415 27300 5435
rect 27250 5385 27300 5415
rect 27250 5365 27265 5385
rect 27285 5365 27300 5385
rect 27250 5335 27300 5365
rect 27250 5315 27265 5335
rect 27285 5315 27300 5335
rect 27250 5285 27300 5315
rect 27250 5265 27265 5285
rect 27285 5265 27300 5285
rect 27250 5235 27300 5265
rect 27250 5215 27265 5235
rect 27285 5215 27300 5235
rect 27250 5185 27300 5215
rect 27250 5165 27265 5185
rect 27285 5165 27300 5185
rect 27250 5135 27300 5165
rect 27250 5115 27265 5135
rect 27285 5115 27300 5135
rect 27250 5085 27300 5115
rect 27250 5065 27265 5085
rect 27285 5065 27300 5085
rect 27250 5035 27300 5065
rect 27250 5015 27265 5035
rect 27285 5015 27300 5035
rect 26800 4940 26850 4950
rect 26800 4910 26810 4940
rect 26840 4910 26850 4940
rect 26800 4900 26850 4910
rect 27100 4940 27150 4950
rect 27100 4910 27110 4940
rect 27140 4910 27150 4940
rect 27100 4900 27150 4910
rect 26650 4810 26660 4840
rect 26690 4810 26700 4840
rect 26650 4785 26700 4810
rect 26650 4765 26665 4785
rect 26685 4765 26700 4785
rect 26650 4740 26700 4765
rect 26650 4710 26660 4740
rect 26690 4710 26700 4740
rect 26650 4685 26700 4710
rect 26650 4665 26665 4685
rect 26685 4665 26700 4685
rect 26650 4640 26700 4665
rect 26650 4610 26660 4640
rect 26690 4610 26700 4640
rect 26650 4585 26700 4610
rect 26650 4565 26665 4585
rect 26685 4565 26700 4585
rect 26650 4540 26700 4565
rect 26650 4510 26660 4540
rect 26690 4510 26700 4540
rect 26650 4485 26700 4510
rect 26650 4465 26665 4485
rect 26685 4465 26700 4485
rect 26650 4440 26700 4465
rect 26650 4410 26660 4440
rect 26690 4410 26700 4440
rect 26650 4385 26700 4410
rect 26650 4365 26665 4385
rect 26685 4365 26700 4385
rect 26650 4290 26700 4365
rect 27250 4835 27300 5015
rect 27700 5485 27750 5500
rect 27700 5465 27715 5485
rect 27735 5465 27750 5485
rect 27700 5435 27750 5465
rect 27700 5415 27715 5435
rect 27735 5415 27750 5435
rect 27700 5385 27750 5415
rect 27700 5365 27715 5385
rect 27735 5365 27750 5385
rect 27700 5335 27750 5365
rect 27700 5315 27715 5335
rect 27735 5315 27750 5335
rect 27700 5285 27750 5315
rect 27700 5265 27715 5285
rect 27735 5265 27750 5285
rect 27700 5235 27750 5265
rect 27700 5215 27715 5235
rect 27735 5215 27750 5235
rect 27700 5185 27750 5215
rect 27700 5165 27715 5185
rect 27735 5165 27750 5185
rect 27700 5135 27750 5165
rect 27700 5115 27715 5135
rect 27735 5115 27750 5135
rect 27700 5085 27750 5115
rect 27700 5065 27715 5085
rect 27735 5065 27750 5085
rect 27700 5035 27750 5065
rect 27700 5015 27715 5035
rect 27735 5015 27750 5035
rect 27550 4940 27600 4950
rect 27550 4910 27560 4940
rect 27590 4910 27600 4940
rect 27550 4900 27600 4910
rect 27700 4940 27750 5015
rect 28150 5485 28200 5560
rect 28150 5465 28165 5485
rect 28185 5465 28200 5485
rect 28150 5440 28200 5465
rect 28150 5410 28160 5440
rect 28190 5410 28200 5440
rect 28150 5385 28200 5410
rect 28150 5365 28165 5385
rect 28185 5365 28200 5385
rect 28150 5340 28200 5365
rect 28150 5310 28160 5340
rect 28190 5310 28200 5340
rect 28150 5285 28200 5310
rect 28150 5265 28165 5285
rect 28185 5265 28200 5285
rect 28150 5240 28200 5265
rect 28150 5210 28160 5240
rect 28190 5210 28200 5240
rect 28150 5185 28200 5210
rect 28150 5165 28165 5185
rect 28185 5165 28200 5185
rect 28150 5140 28200 5165
rect 28150 5110 28160 5140
rect 28190 5110 28200 5140
rect 28150 5085 28200 5110
rect 28150 5065 28165 5085
rect 28185 5065 28200 5085
rect 28150 5040 28200 5065
rect 28150 5010 28160 5040
rect 28190 5010 28200 5040
rect 27700 4910 27710 4940
rect 27740 4910 27750 4940
rect 27250 4815 27265 4835
rect 27285 4815 27300 4835
rect 27250 4785 27300 4815
rect 27250 4765 27265 4785
rect 27285 4765 27300 4785
rect 27250 4735 27300 4765
rect 27250 4715 27265 4735
rect 27285 4715 27300 4735
rect 27250 4685 27300 4715
rect 27250 4665 27265 4685
rect 27285 4665 27300 4685
rect 27250 4635 27300 4665
rect 27250 4615 27265 4635
rect 27285 4615 27300 4635
rect 27250 4585 27300 4615
rect 27250 4565 27265 4585
rect 27285 4565 27300 4585
rect 27250 4535 27300 4565
rect 27250 4515 27265 4535
rect 27285 4515 27300 4535
rect 27250 4485 27300 4515
rect 27250 4465 27265 4485
rect 27285 4465 27300 4485
rect 27250 4435 27300 4465
rect 27250 4415 27265 4435
rect 27285 4415 27300 4435
rect 27250 4385 27300 4415
rect 27250 4365 27265 4385
rect 27285 4365 27300 4385
rect 27250 4350 27300 4365
rect 27700 4835 27750 4910
rect 27850 4940 27900 4950
rect 27850 4910 27860 4940
rect 27890 4910 27900 4940
rect 27850 4900 27900 4910
rect 27700 4815 27715 4835
rect 27735 4815 27750 4835
rect 27700 4785 27750 4815
rect 27700 4765 27715 4785
rect 27735 4765 27750 4785
rect 27700 4735 27750 4765
rect 27700 4715 27715 4735
rect 27735 4715 27750 4735
rect 27700 4685 27750 4715
rect 27700 4665 27715 4685
rect 27735 4665 27750 4685
rect 27700 4635 27750 4665
rect 27700 4615 27715 4635
rect 27735 4615 27750 4635
rect 27700 4585 27750 4615
rect 27700 4565 27715 4585
rect 27735 4565 27750 4585
rect 27700 4535 27750 4565
rect 27700 4515 27715 4535
rect 27735 4515 27750 4535
rect 27700 4485 27750 4515
rect 27700 4465 27715 4485
rect 27735 4465 27750 4485
rect 27700 4435 27750 4465
rect 27700 4415 27715 4435
rect 27735 4415 27750 4435
rect 27700 4385 27750 4415
rect 27700 4365 27715 4385
rect 27735 4365 27750 4385
rect 26650 4260 26660 4290
rect 26690 4260 26700 4290
rect 25600 4165 25615 4185
rect 25635 4165 25650 4185
rect 25600 4135 25650 4165
rect 25600 4115 25615 4135
rect 25635 4115 25650 4135
rect 25600 4085 25650 4115
rect 25600 4065 25615 4085
rect 25635 4065 25650 4085
rect 25600 4035 25650 4065
rect 25600 4015 25615 4035
rect 25635 4015 25650 4035
rect 25600 3985 25650 4015
rect 25600 3965 25615 3985
rect 25635 3965 25650 3985
rect 25600 3935 25650 3965
rect 25600 3915 25615 3935
rect 25635 3915 25650 3935
rect 25600 3885 25650 3915
rect 25600 3865 25615 3885
rect 25635 3865 25650 3885
rect 25600 3835 25650 3865
rect 25600 3815 25615 3835
rect 25635 3815 25650 3835
rect 25600 3785 25650 3815
rect 25600 3765 25615 3785
rect 25635 3765 25650 3785
rect 25600 3735 25650 3765
rect 25600 3715 25615 3735
rect 25635 3715 25650 3735
rect 25450 3640 25500 3650
rect 25450 3610 25460 3640
rect 25490 3610 25500 3640
rect 25450 3600 25500 3610
rect 25600 3640 25650 3715
rect 26050 4185 26100 4200
rect 26050 4165 26065 4185
rect 26085 4165 26100 4185
rect 26050 4135 26100 4165
rect 26050 4115 26065 4135
rect 26085 4115 26100 4135
rect 26050 4085 26100 4115
rect 26050 4065 26065 4085
rect 26085 4065 26100 4085
rect 26050 4035 26100 4065
rect 26050 4015 26065 4035
rect 26085 4015 26100 4035
rect 26050 3985 26100 4015
rect 26050 3965 26065 3985
rect 26085 3965 26100 3985
rect 26050 3935 26100 3965
rect 26050 3915 26065 3935
rect 26085 3915 26100 3935
rect 26050 3885 26100 3915
rect 26050 3865 26065 3885
rect 26085 3865 26100 3885
rect 26050 3835 26100 3865
rect 26050 3815 26065 3835
rect 26085 3815 26100 3835
rect 26050 3785 26100 3815
rect 26050 3765 26065 3785
rect 26085 3765 26100 3785
rect 26050 3735 26100 3765
rect 26050 3715 26065 3735
rect 26085 3715 26100 3735
rect 25600 3610 25610 3640
rect 25640 3610 25650 3640
rect 25150 3515 25165 3535
rect 25185 3515 25200 3535
rect 25150 3485 25200 3515
rect 25150 3465 25165 3485
rect 25185 3465 25200 3485
rect 25150 3435 25200 3465
rect 25150 3415 25165 3435
rect 25185 3415 25200 3435
rect 25150 3385 25200 3415
rect 25150 3365 25165 3385
rect 25185 3365 25200 3385
rect 25150 3335 25200 3365
rect 25150 3315 25165 3335
rect 25185 3315 25200 3335
rect 25150 3285 25200 3315
rect 25150 3265 25165 3285
rect 25185 3265 25200 3285
rect 25150 3235 25200 3265
rect 25150 3215 25165 3235
rect 25185 3215 25200 3235
rect 25150 3185 25200 3215
rect 25150 3165 25165 3185
rect 25185 3165 25200 3185
rect 25150 3135 25200 3165
rect 25150 3115 25165 3135
rect 25185 3115 25200 3135
rect 25150 3085 25200 3115
rect 25150 3065 25165 3085
rect 25185 3065 25200 3085
rect 25150 3050 25200 3065
rect 25600 3535 25650 3610
rect 25750 3640 25800 3650
rect 25750 3610 25760 3640
rect 25790 3610 25800 3640
rect 25750 3600 25800 3610
rect 25600 3515 25615 3535
rect 25635 3515 25650 3535
rect 25600 3485 25650 3515
rect 25600 3465 25615 3485
rect 25635 3465 25650 3485
rect 25600 3435 25650 3465
rect 25600 3415 25615 3435
rect 25635 3415 25650 3435
rect 25600 3385 25650 3415
rect 25600 3365 25615 3385
rect 25635 3365 25650 3385
rect 25600 3335 25650 3365
rect 25600 3315 25615 3335
rect 25635 3315 25650 3335
rect 25600 3285 25650 3315
rect 25600 3265 25615 3285
rect 25635 3265 25650 3285
rect 25600 3235 25650 3265
rect 25600 3215 25615 3235
rect 25635 3215 25650 3235
rect 25600 3185 25650 3215
rect 25600 3165 25615 3185
rect 25635 3165 25650 3185
rect 25600 3135 25650 3165
rect 25600 3115 25615 3135
rect 25635 3115 25650 3135
rect 25600 3085 25650 3115
rect 25600 3065 25615 3085
rect 25635 3065 25650 3085
rect 25600 3050 25650 3065
rect 26050 3535 26100 3715
rect 26650 4185 26700 4260
rect 26650 4165 26665 4185
rect 26685 4165 26700 4185
rect 26650 4140 26700 4165
rect 26650 4110 26660 4140
rect 26690 4110 26700 4140
rect 26650 4085 26700 4110
rect 26650 4065 26665 4085
rect 26685 4065 26700 4085
rect 26650 4040 26700 4065
rect 26650 4010 26660 4040
rect 26690 4010 26700 4040
rect 26650 3985 26700 4010
rect 26650 3965 26665 3985
rect 26685 3965 26700 3985
rect 26650 3940 26700 3965
rect 26650 3910 26660 3940
rect 26690 3910 26700 3940
rect 26650 3885 26700 3910
rect 26650 3865 26665 3885
rect 26685 3865 26700 3885
rect 26650 3840 26700 3865
rect 26650 3810 26660 3840
rect 26690 3810 26700 3840
rect 26650 3785 26700 3810
rect 26650 3765 26665 3785
rect 26685 3765 26700 3785
rect 26650 3740 26700 3765
rect 26650 3710 26660 3740
rect 26690 3710 26700 3740
rect 26200 3640 26250 3650
rect 26200 3610 26210 3640
rect 26240 3610 26250 3640
rect 26200 3600 26250 3610
rect 26500 3640 26550 3650
rect 26500 3610 26510 3640
rect 26540 3610 26550 3640
rect 26500 3600 26550 3610
rect 26050 3515 26065 3535
rect 26085 3515 26100 3535
rect 26050 3485 26100 3515
rect 26050 3465 26065 3485
rect 26085 3465 26100 3485
rect 26050 3435 26100 3465
rect 26050 3415 26065 3435
rect 26085 3415 26100 3435
rect 26050 3385 26100 3415
rect 26050 3365 26065 3385
rect 26085 3365 26100 3385
rect 26050 3335 26100 3365
rect 26050 3315 26065 3335
rect 26085 3315 26100 3335
rect 26050 3285 26100 3315
rect 26050 3265 26065 3285
rect 26085 3265 26100 3285
rect 26050 3235 26100 3265
rect 26050 3215 26065 3235
rect 26085 3215 26100 3235
rect 26050 3185 26100 3215
rect 26050 3165 26065 3185
rect 26085 3165 26100 3185
rect 26050 3135 26100 3165
rect 26050 3115 26065 3135
rect 26085 3115 26100 3135
rect 26050 3085 26100 3115
rect 26050 3065 26065 3085
rect 26085 3065 26100 3085
rect 26050 3050 26100 3065
rect 26650 3540 26700 3710
rect 27250 4185 27300 4200
rect 27250 4165 27265 4185
rect 27285 4165 27300 4185
rect 27250 4135 27300 4165
rect 27250 4115 27265 4135
rect 27285 4115 27300 4135
rect 27250 4085 27300 4115
rect 27250 4065 27265 4085
rect 27285 4065 27300 4085
rect 27250 4035 27300 4065
rect 27250 4015 27265 4035
rect 27285 4015 27300 4035
rect 27250 3985 27300 4015
rect 27250 3965 27265 3985
rect 27285 3965 27300 3985
rect 27250 3935 27300 3965
rect 27250 3915 27265 3935
rect 27285 3915 27300 3935
rect 27250 3885 27300 3915
rect 27250 3865 27265 3885
rect 27285 3865 27300 3885
rect 27250 3835 27300 3865
rect 27250 3815 27265 3835
rect 27285 3815 27300 3835
rect 27250 3785 27300 3815
rect 27250 3765 27265 3785
rect 27285 3765 27300 3785
rect 27250 3735 27300 3765
rect 27250 3715 27265 3735
rect 27285 3715 27300 3735
rect 26800 3640 26850 3650
rect 26800 3610 26810 3640
rect 26840 3610 26850 3640
rect 26800 3600 26850 3610
rect 27100 3640 27150 3650
rect 27100 3610 27110 3640
rect 27140 3610 27150 3640
rect 27100 3600 27150 3610
rect 26650 3510 26660 3540
rect 26690 3510 26700 3540
rect 26650 3485 26700 3510
rect 26650 3465 26665 3485
rect 26685 3465 26700 3485
rect 26650 3440 26700 3465
rect 26650 3410 26660 3440
rect 26690 3410 26700 3440
rect 26650 3385 26700 3410
rect 26650 3365 26665 3385
rect 26685 3365 26700 3385
rect 26650 3340 26700 3365
rect 26650 3310 26660 3340
rect 26690 3310 26700 3340
rect 26650 3285 26700 3310
rect 26650 3265 26665 3285
rect 26685 3265 26700 3285
rect 26650 3240 26700 3265
rect 26650 3210 26660 3240
rect 26690 3210 26700 3240
rect 26650 3185 26700 3210
rect 26650 3165 26665 3185
rect 26685 3165 26700 3185
rect 26650 3140 26700 3165
rect 26650 3110 26660 3140
rect 26690 3110 26700 3140
rect 26650 3085 26700 3110
rect 26650 3065 26665 3085
rect 26685 3065 26700 3085
rect 26650 3050 26700 3065
rect 27250 3535 27300 3715
rect 27700 4185 27750 4365
rect 27700 4165 27715 4185
rect 27735 4165 27750 4185
rect 27700 4135 27750 4165
rect 27700 4115 27715 4135
rect 27735 4115 27750 4135
rect 27700 4085 27750 4115
rect 27700 4065 27715 4085
rect 27735 4065 27750 4085
rect 27700 4035 27750 4065
rect 27700 4015 27715 4035
rect 27735 4015 27750 4035
rect 27700 3985 27750 4015
rect 27700 3965 27715 3985
rect 27735 3965 27750 3985
rect 27700 3935 27750 3965
rect 27700 3915 27715 3935
rect 27735 3915 27750 3935
rect 27700 3885 27750 3915
rect 27700 3865 27715 3885
rect 27735 3865 27750 3885
rect 27700 3835 27750 3865
rect 27700 3815 27715 3835
rect 27735 3815 27750 3835
rect 27700 3785 27750 3815
rect 27700 3765 27715 3785
rect 27735 3765 27750 3785
rect 27700 3735 27750 3765
rect 27700 3715 27715 3735
rect 27735 3715 27750 3735
rect 27550 3640 27600 3650
rect 27550 3610 27560 3640
rect 27590 3610 27600 3640
rect 27550 3600 27600 3610
rect 27700 3640 27750 3715
rect 28150 4840 28200 5010
rect 28750 5590 28800 5600
rect 28750 5560 28760 5590
rect 28790 5560 28800 5590
rect 28750 5485 28800 5560
rect 32050 5590 32100 5600
rect 32050 5560 32060 5590
rect 32090 5560 32100 5590
rect 28750 5465 28765 5485
rect 28785 5465 28800 5485
rect 28750 5440 28800 5465
rect 28750 5410 28760 5440
rect 28790 5410 28800 5440
rect 28750 5385 28800 5410
rect 28750 5365 28765 5385
rect 28785 5365 28800 5385
rect 28750 5340 28800 5365
rect 28750 5310 28760 5340
rect 28790 5310 28800 5340
rect 28750 5285 28800 5310
rect 28750 5265 28765 5285
rect 28785 5265 28800 5285
rect 28750 5240 28800 5265
rect 28750 5210 28760 5240
rect 28790 5210 28800 5240
rect 28750 5185 28800 5210
rect 28750 5165 28765 5185
rect 28785 5165 28800 5185
rect 28750 5140 28800 5165
rect 28750 5110 28760 5140
rect 28790 5110 28800 5140
rect 28750 5085 28800 5110
rect 28750 5065 28765 5085
rect 28785 5065 28800 5085
rect 28750 5040 28800 5065
rect 28750 5010 28760 5040
rect 28790 5010 28800 5040
rect 28300 4940 28350 4950
rect 28300 4910 28310 4940
rect 28340 4910 28350 4940
rect 28300 4900 28350 4910
rect 28600 4940 28650 4950
rect 28600 4910 28610 4940
rect 28640 4910 28650 4940
rect 28600 4900 28650 4910
rect 28750 4940 28800 5010
rect 29350 5485 29700 5500
rect 29350 5465 29365 5485
rect 29385 5465 29665 5485
rect 29685 5465 29700 5485
rect 29350 5450 29700 5465
rect 29350 5435 29400 5450
rect 29350 5415 29365 5435
rect 29385 5415 29400 5435
rect 29350 5385 29400 5415
rect 29650 5435 29700 5450
rect 29650 5415 29665 5435
rect 29685 5415 29700 5435
rect 29350 5365 29365 5385
rect 29385 5365 29400 5385
rect 29350 5335 29400 5365
rect 29350 5315 29365 5335
rect 29385 5315 29400 5335
rect 29350 5285 29400 5315
rect 29350 5265 29365 5285
rect 29385 5265 29400 5285
rect 29350 5235 29400 5265
rect 29350 5215 29365 5235
rect 29385 5215 29400 5235
rect 29350 5185 29400 5215
rect 29350 5165 29365 5185
rect 29385 5165 29400 5185
rect 29350 5135 29400 5165
rect 29350 5115 29365 5135
rect 29385 5115 29400 5135
rect 29350 5085 29400 5115
rect 29350 5065 29365 5085
rect 29385 5065 29400 5085
rect 29350 5035 29400 5065
rect 29350 5015 29365 5035
rect 29385 5015 29400 5035
rect 28750 4910 28760 4940
rect 28790 4910 28800 4940
rect 28150 4810 28160 4840
rect 28190 4810 28200 4840
rect 28150 4785 28200 4810
rect 28150 4765 28165 4785
rect 28185 4765 28200 4785
rect 28150 4740 28200 4765
rect 28150 4710 28160 4740
rect 28190 4710 28200 4740
rect 28150 4685 28200 4710
rect 28150 4665 28165 4685
rect 28185 4665 28200 4685
rect 28150 4640 28200 4665
rect 28150 4610 28160 4640
rect 28190 4610 28200 4640
rect 28150 4585 28200 4610
rect 28150 4565 28165 4585
rect 28185 4565 28200 4585
rect 28150 4540 28200 4565
rect 28150 4510 28160 4540
rect 28190 4510 28200 4540
rect 28150 4485 28200 4510
rect 28150 4465 28165 4485
rect 28185 4465 28200 4485
rect 28150 4440 28200 4465
rect 28150 4410 28160 4440
rect 28190 4410 28200 4440
rect 28150 4385 28200 4410
rect 28150 4365 28165 4385
rect 28185 4365 28200 4385
rect 28150 4290 28200 4365
rect 28150 4260 28160 4290
rect 28190 4260 28200 4290
rect 28150 4185 28200 4260
rect 28150 4165 28165 4185
rect 28185 4165 28200 4185
rect 28150 4140 28200 4165
rect 28150 4110 28160 4140
rect 28190 4110 28200 4140
rect 28150 4085 28200 4110
rect 28150 4065 28165 4085
rect 28185 4065 28200 4085
rect 28150 4040 28200 4065
rect 28150 4010 28160 4040
rect 28190 4010 28200 4040
rect 28150 3985 28200 4010
rect 28150 3965 28165 3985
rect 28185 3965 28200 3985
rect 28150 3940 28200 3965
rect 28150 3910 28160 3940
rect 28190 3910 28200 3940
rect 28150 3885 28200 3910
rect 28150 3865 28165 3885
rect 28185 3865 28200 3885
rect 28150 3840 28200 3865
rect 28150 3810 28160 3840
rect 28190 3810 28200 3840
rect 28150 3785 28200 3810
rect 28150 3765 28165 3785
rect 28185 3765 28200 3785
rect 28150 3740 28200 3765
rect 28150 3710 28160 3740
rect 28190 3710 28200 3740
rect 27700 3610 27710 3640
rect 27740 3610 27750 3640
rect 27250 3515 27265 3535
rect 27285 3515 27300 3535
rect 27250 3485 27300 3515
rect 27250 3465 27265 3485
rect 27285 3465 27300 3485
rect 27250 3435 27300 3465
rect 27250 3415 27265 3435
rect 27285 3415 27300 3435
rect 27250 3385 27300 3415
rect 27250 3365 27265 3385
rect 27285 3365 27300 3385
rect 27250 3335 27300 3365
rect 27250 3315 27265 3335
rect 27285 3315 27300 3335
rect 27250 3285 27300 3315
rect 27250 3265 27265 3285
rect 27285 3265 27300 3285
rect 27250 3235 27300 3265
rect 27250 3215 27265 3235
rect 27285 3215 27300 3235
rect 27250 3185 27300 3215
rect 27250 3165 27265 3185
rect 27285 3165 27300 3185
rect 27250 3135 27300 3165
rect 27250 3115 27265 3135
rect 27285 3115 27300 3135
rect 27250 3085 27300 3115
rect 27250 3065 27265 3085
rect 27285 3065 27300 3085
rect 27250 3050 27300 3065
rect 27700 3535 27750 3610
rect 27850 3640 27900 3650
rect 27850 3610 27860 3640
rect 27890 3610 27900 3640
rect 27850 3600 27900 3610
rect 27700 3515 27715 3535
rect 27735 3515 27750 3535
rect 27700 3485 27750 3515
rect 27700 3465 27715 3485
rect 27735 3465 27750 3485
rect 27700 3435 27750 3465
rect 27700 3415 27715 3435
rect 27735 3415 27750 3435
rect 27700 3385 27750 3415
rect 27700 3365 27715 3385
rect 27735 3365 27750 3385
rect 27700 3335 27750 3365
rect 27700 3315 27715 3335
rect 27735 3315 27750 3335
rect 27700 3285 27750 3315
rect 27700 3265 27715 3285
rect 27735 3265 27750 3285
rect 27700 3235 27750 3265
rect 27700 3215 27715 3235
rect 27735 3215 27750 3235
rect 27700 3185 27750 3215
rect 27700 3165 27715 3185
rect 27735 3165 27750 3185
rect 27700 3135 27750 3165
rect 27700 3115 27715 3135
rect 27735 3115 27750 3135
rect 27700 3085 27750 3115
rect 27700 3065 27715 3085
rect 27735 3065 27750 3085
rect 27700 3050 27750 3065
rect 28150 3540 28200 3710
rect 28750 4840 28800 4910
rect 28900 4940 28950 4950
rect 28900 4910 28910 4940
rect 28940 4910 28950 4940
rect 28900 4900 28950 4910
rect 29200 4940 29250 4950
rect 29200 4910 29210 4940
rect 29240 4910 29250 4940
rect 29200 4900 29250 4910
rect 29350 4940 29400 5015
rect 29500 5385 29550 5400
rect 29500 5365 29515 5385
rect 29535 5365 29550 5385
rect 29500 5335 29550 5365
rect 29500 5315 29515 5335
rect 29535 5315 29550 5335
rect 29500 5285 29550 5315
rect 29500 5265 29515 5285
rect 29535 5265 29550 5285
rect 29500 5235 29550 5265
rect 29500 5215 29515 5235
rect 29535 5215 29550 5235
rect 29500 5185 29550 5215
rect 29500 5165 29515 5185
rect 29535 5165 29550 5185
rect 29500 5135 29550 5165
rect 29500 5115 29515 5135
rect 29535 5115 29550 5135
rect 29500 5085 29550 5115
rect 29650 5385 29700 5415
rect 29650 5365 29665 5385
rect 29685 5365 29700 5385
rect 29650 5335 29700 5365
rect 29650 5315 29665 5335
rect 29685 5315 29700 5335
rect 29650 5285 29700 5315
rect 29650 5265 29665 5285
rect 29685 5265 29700 5285
rect 29650 5235 29700 5265
rect 29650 5215 29665 5235
rect 29685 5215 29700 5235
rect 29650 5185 29700 5215
rect 29650 5165 29665 5185
rect 29685 5165 29700 5185
rect 29650 5135 29700 5165
rect 29650 5115 29665 5135
rect 29685 5115 29700 5135
rect 29650 5100 29700 5115
rect 29800 5485 29850 5500
rect 29800 5465 29815 5485
rect 29835 5465 29850 5485
rect 29800 5435 29850 5465
rect 29800 5415 29815 5435
rect 29835 5415 29850 5435
rect 29800 5385 29850 5415
rect 29800 5365 29815 5385
rect 29835 5365 29850 5385
rect 29800 5335 29850 5365
rect 29800 5315 29815 5335
rect 29835 5315 29850 5335
rect 29800 5285 29850 5315
rect 29800 5265 29815 5285
rect 29835 5265 29850 5285
rect 29800 5235 29850 5265
rect 29800 5215 29815 5235
rect 29835 5215 29850 5235
rect 29800 5185 29850 5215
rect 29800 5165 29815 5185
rect 29835 5165 29850 5185
rect 29800 5135 29850 5165
rect 29800 5115 29815 5135
rect 29835 5115 29850 5135
rect 29500 5065 29515 5085
rect 29535 5065 29550 5085
rect 29500 5050 29550 5065
rect 29800 5085 29850 5115
rect 29950 5485 30900 5500
rect 29950 5465 29965 5485
rect 29985 5465 30265 5485
rect 30285 5465 30415 5485
rect 30435 5465 30565 5485
rect 30585 5465 30865 5485
rect 30885 5465 30900 5485
rect 29950 5450 30900 5465
rect 29950 5435 30000 5450
rect 29950 5415 29965 5435
rect 29985 5415 30000 5435
rect 29950 5385 30000 5415
rect 30250 5435 30300 5450
rect 30250 5415 30265 5435
rect 30285 5415 30300 5435
rect 29950 5365 29965 5385
rect 29985 5365 30000 5385
rect 29950 5335 30000 5365
rect 29950 5315 29965 5335
rect 29985 5315 30000 5335
rect 29950 5285 30000 5315
rect 29950 5265 29965 5285
rect 29985 5265 30000 5285
rect 29950 5235 30000 5265
rect 29950 5215 29965 5235
rect 29985 5215 30000 5235
rect 29950 5185 30000 5215
rect 29950 5165 29965 5185
rect 29985 5165 30000 5185
rect 29950 5135 30000 5165
rect 29950 5115 29965 5135
rect 29985 5115 30000 5135
rect 29950 5100 30000 5115
rect 30100 5385 30150 5400
rect 30100 5365 30115 5385
rect 30135 5365 30150 5385
rect 30100 5335 30150 5365
rect 30100 5315 30115 5335
rect 30135 5315 30150 5335
rect 30100 5285 30150 5315
rect 30100 5265 30115 5285
rect 30135 5265 30150 5285
rect 30100 5235 30150 5265
rect 30100 5215 30115 5235
rect 30135 5215 30150 5235
rect 30100 5185 30150 5215
rect 30100 5165 30115 5185
rect 30135 5165 30150 5185
rect 30100 5135 30150 5165
rect 30100 5115 30115 5135
rect 30135 5115 30150 5135
rect 29800 5065 29815 5085
rect 29835 5065 29850 5085
rect 29800 5050 29850 5065
rect 30100 5085 30150 5115
rect 30250 5385 30300 5415
rect 30250 5365 30265 5385
rect 30285 5365 30300 5385
rect 30250 5335 30300 5365
rect 30250 5315 30265 5335
rect 30285 5315 30300 5335
rect 30250 5285 30300 5315
rect 30250 5265 30265 5285
rect 30285 5265 30300 5285
rect 30250 5235 30300 5265
rect 30250 5215 30265 5235
rect 30285 5215 30300 5235
rect 30250 5185 30300 5215
rect 30250 5165 30265 5185
rect 30285 5165 30300 5185
rect 30250 5135 30300 5165
rect 30250 5115 30265 5135
rect 30285 5115 30300 5135
rect 30250 5100 30300 5115
rect 30400 5435 30450 5450
rect 30400 5415 30415 5435
rect 30435 5415 30450 5435
rect 30400 5385 30450 5415
rect 30400 5365 30415 5385
rect 30435 5365 30450 5385
rect 30400 5335 30450 5365
rect 30400 5315 30415 5335
rect 30435 5315 30450 5335
rect 30400 5285 30450 5315
rect 30400 5265 30415 5285
rect 30435 5265 30450 5285
rect 30400 5235 30450 5265
rect 30400 5215 30415 5235
rect 30435 5215 30450 5235
rect 30400 5185 30450 5215
rect 30400 5165 30415 5185
rect 30435 5165 30450 5185
rect 30400 5135 30450 5165
rect 30400 5115 30415 5135
rect 30435 5115 30450 5135
rect 30100 5065 30115 5085
rect 30135 5065 30150 5085
rect 30100 5050 30150 5065
rect 30400 5085 30450 5115
rect 30550 5435 30600 5450
rect 30550 5415 30565 5435
rect 30585 5415 30600 5435
rect 30550 5385 30600 5415
rect 30850 5435 30900 5450
rect 30850 5415 30865 5435
rect 30885 5415 30900 5435
rect 30550 5365 30565 5385
rect 30585 5365 30600 5385
rect 30550 5335 30600 5365
rect 30550 5315 30565 5335
rect 30585 5315 30600 5335
rect 30550 5285 30600 5315
rect 30550 5265 30565 5285
rect 30585 5265 30600 5285
rect 30550 5235 30600 5265
rect 30550 5215 30565 5235
rect 30585 5215 30600 5235
rect 30550 5185 30600 5215
rect 30550 5165 30565 5185
rect 30585 5165 30600 5185
rect 30550 5135 30600 5165
rect 30550 5115 30565 5135
rect 30585 5115 30600 5135
rect 30550 5100 30600 5115
rect 30700 5385 30750 5400
rect 30700 5365 30715 5385
rect 30735 5365 30750 5385
rect 30700 5335 30750 5365
rect 30700 5315 30715 5335
rect 30735 5315 30750 5335
rect 30700 5285 30750 5315
rect 30700 5265 30715 5285
rect 30735 5265 30750 5285
rect 30700 5235 30750 5265
rect 30700 5215 30715 5235
rect 30735 5215 30750 5235
rect 30700 5185 30750 5215
rect 30700 5165 30715 5185
rect 30735 5165 30750 5185
rect 30700 5135 30750 5165
rect 30700 5115 30715 5135
rect 30735 5115 30750 5135
rect 30400 5065 30415 5085
rect 30435 5065 30450 5085
rect 30400 5050 30450 5065
rect 30700 5085 30750 5115
rect 30850 5385 30900 5415
rect 30850 5365 30865 5385
rect 30885 5365 30900 5385
rect 30850 5335 30900 5365
rect 30850 5315 30865 5335
rect 30885 5315 30900 5335
rect 30850 5285 30900 5315
rect 30850 5265 30865 5285
rect 30885 5265 30900 5285
rect 30850 5235 30900 5265
rect 30850 5215 30865 5235
rect 30885 5215 30900 5235
rect 30850 5185 30900 5215
rect 30850 5165 30865 5185
rect 30885 5165 30900 5185
rect 30850 5135 30900 5165
rect 30850 5115 30865 5135
rect 30885 5115 30900 5135
rect 30850 5100 30900 5115
rect 31000 5485 31050 5500
rect 31000 5465 31015 5485
rect 31035 5465 31050 5485
rect 31000 5435 31050 5465
rect 31000 5415 31015 5435
rect 31035 5415 31050 5435
rect 31000 5385 31050 5415
rect 31000 5365 31015 5385
rect 31035 5365 31050 5385
rect 31000 5335 31050 5365
rect 31000 5315 31015 5335
rect 31035 5315 31050 5335
rect 31000 5285 31050 5315
rect 31000 5265 31015 5285
rect 31035 5265 31050 5285
rect 31000 5235 31050 5265
rect 31000 5215 31015 5235
rect 31035 5215 31050 5235
rect 31000 5185 31050 5215
rect 31000 5165 31015 5185
rect 31035 5165 31050 5185
rect 31000 5135 31050 5165
rect 31000 5115 31015 5135
rect 31035 5115 31050 5135
rect 30700 5065 30715 5085
rect 30735 5065 30750 5085
rect 30700 5050 30750 5065
rect 31000 5085 31050 5115
rect 31150 5485 31500 5500
rect 31150 5465 31165 5485
rect 31185 5465 31465 5485
rect 31485 5465 31500 5485
rect 31150 5450 31500 5465
rect 31150 5435 31200 5450
rect 31150 5415 31165 5435
rect 31185 5415 31200 5435
rect 31150 5385 31200 5415
rect 31450 5435 31500 5450
rect 31450 5415 31465 5435
rect 31485 5415 31500 5435
rect 31150 5365 31165 5385
rect 31185 5365 31200 5385
rect 31150 5335 31200 5365
rect 31150 5315 31165 5335
rect 31185 5315 31200 5335
rect 31150 5285 31200 5315
rect 31150 5265 31165 5285
rect 31185 5265 31200 5285
rect 31150 5235 31200 5265
rect 31150 5215 31165 5235
rect 31185 5215 31200 5235
rect 31150 5185 31200 5215
rect 31150 5165 31165 5185
rect 31185 5165 31200 5185
rect 31150 5135 31200 5165
rect 31150 5115 31165 5135
rect 31185 5115 31200 5135
rect 31150 5100 31200 5115
rect 31300 5385 31350 5400
rect 31300 5365 31315 5385
rect 31335 5365 31350 5385
rect 31300 5335 31350 5365
rect 31300 5315 31315 5335
rect 31335 5315 31350 5335
rect 31300 5285 31350 5315
rect 31300 5265 31315 5285
rect 31335 5265 31350 5285
rect 31300 5235 31350 5265
rect 31300 5215 31315 5235
rect 31335 5215 31350 5235
rect 31300 5185 31350 5215
rect 31300 5165 31315 5185
rect 31335 5165 31350 5185
rect 31300 5135 31350 5165
rect 31300 5115 31315 5135
rect 31335 5115 31350 5135
rect 31000 5065 31015 5085
rect 31035 5065 31050 5085
rect 31000 5050 31050 5065
rect 31300 5085 31350 5115
rect 31300 5065 31315 5085
rect 31335 5065 31350 5085
rect 31300 5050 31350 5065
rect 29500 5035 31350 5050
rect 29500 5015 29515 5035
rect 29535 5015 29815 5035
rect 29835 5015 30115 5035
rect 30135 5015 30415 5035
rect 30435 5015 30715 5035
rect 30735 5015 31015 5035
rect 31035 5015 31315 5035
rect 31335 5015 31350 5035
rect 29500 5000 31350 5015
rect 31450 5385 31500 5415
rect 31450 5365 31465 5385
rect 31485 5365 31500 5385
rect 31450 5335 31500 5365
rect 31450 5315 31465 5335
rect 31485 5315 31500 5335
rect 31450 5285 31500 5315
rect 31450 5265 31465 5285
rect 31485 5265 31500 5285
rect 31450 5235 31500 5265
rect 31450 5215 31465 5235
rect 31485 5215 31500 5235
rect 31450 5185 31500 5215
rect 31450 5165 31465 5185
rect 31485 5165 31500 5185
rect 31450 5135 31500 5165
rect 31450 5115 31465 5135
rect 31485 5115 31500 5135
rect 31450 5085 31500 5115
rect 31450 5065 31465 5085
rect 31485 5065 31500 5085
rect 31450 5035 31500 5065
rect 31450 5015 31465 5035
rect 31485 5015 31500 5035
rect 29350 4910 29360 4940
rect 29390 4910 29400 4940
rect 28750 4810 28760 4840
rect 28790 4810 28800 4840
rect 28750 4785 28800 4810
rect 28750 4765 28765 4785
rect 28785 4765 28800 4785
rect 28750 4740 28800 4765
rect 28750 4710 28760 4740
rect 28790 4710 28800 4740
rect 28750 4685 28800 4710
rect 28750 4665 28765 4685
rect 28785 4665 28800 4685
rect 28750 4640 28800 4665
rect 28750 4610 28760 4640
rect 28790 4610 28800 4640
rect 28750 4585 28800 4610
rect 28750 4565 28765 4585
rect 28785 4565 28800 4585
rect 28750 4540 28800 4565
rect 28750 4510 28760 4540
rect 28790 4510 28800 4540
rect 28750 4485 28800 4510
rect 28750 4465 28765 4485
rect 28785 4465 28800 4485
rect 28750 4440 28800 4465
rect 28750 4410 28760 4440
rect 28790 4410 28800 4440
rect 28750 4385 28800 4410
rect 28750 4365 28765 4385
rect 28785 4365 28800 4385
rect 28750 4290 28800 4365
rect 28750 4260 28760 4290
rect 28790 4260 28800 4290
rect 28750 4185 28800 4260
rect 28750 4165 28765 4185
rect 28785 4165 28800 4185
rect 28750 4140 28800 4165
rect 28750 4110 28760 4140
rect 28790 4110 28800 4140
rect 28750 4085 28800 4110
rect 28750 4065 28765 4085
rect 28785 4065 28800 4085
rect 28750 4040 28800 4065
rect 28750 4010 28760 4040
rect 28790 4010 28800 4040
rect 28750 3985 28800 4010
rect 28750 3965 28765 3985
rect 28785 3965 28800 3985
rect 28750 3940 28800 3965
rect 28750 3910 28760 3940
rect 28790 3910 28800 3940
rect 28750 3885 28800 3910
rect 28750 3865 28765 3885
rect 28785 3865 28800 3885
rect 28750 3840 28800 3865
rect 28750 3810 28760 3840
rect 28790 3810 28800 3840
rect 28750 3785 28800 3810
rect 28750 3765 28765 3785
rect 28785 3765 28800 3785
rect 28750 3740 28800 3765
rect 28750 3710 28760 3740
rect 28790 3710 28800 3740
rect 28300 3640 28350 3650
rect 28300 3610 28310 3640
rect 28340 3610 28350 3640
rect 28300 3600 28350 3610
rect 28600 3640 28650 3650
rect 28600 3610 28610 3640
rect 28640 3610 28650 3640
rect 28600 3600 28650 3610
rect 28750 3640 28800 3710
rect 29350 4835 29400 4910
rect 29650 4940 29700 4950
rect 29650 4910 29660 4940
rect 29690 4910 29700 4940
rect 29650 4900 29700 4910
rect 29950 4940 30000 4950
rect 29950 4910 29960 4940
rect 29990 4910 30000 4940
rect 29950 4900 30000 4910
rect 30250 4940 30300 4950
rect 30250 4910 30260 4940
rect 30290 4910 30300 4940
rect 30250 4900 30300 4910
rect 30550 4940 30600 4950
rect 30550 4910 30560 4940
rect 30590 4910 30600 4940
rect 30550 4900 30600 4910
rect 30850 4940 30900 4950
rect 30850 4910 30860 4940
rect 30890 4910 30900 4940
rect 30850 4900 30900 4910
rect 31150 4940 31200 4950
rect 31150 4910 31160 4940
rect 31190 4910 31200 4940
rect 31150 4900 31200 4910
rect 31450 4940 31500 5015
rect 32050 5485 32100 5560
rect 32050 5465 32065 5485
rect 32085 5465 32100 5485
rect 32050 5440 32100 5465
rect 32050 5410 32060 5440
rect 32090 5410 32100 5440
rect 32050 5385 32100 5410
rect 32050 5365 32065 5385
rect 32085 5365 32100 5385
rect 32050 5340 32100 5365
rect 32050 5310 32060 5340
rect 32090 5310 32100 5340
rect 32050 5285 32100 5310
rect 32050 5265 32065 5285
rect 32085 5265 32100 5285
rect 32050 5240 32100 5265
rect 32050 5210 32060 5240
rect 32090 5210 32100 5240
rect 32050 5185 32100 5210
rect 32050 5165 32065 5185
rect 32085 5165 32100 5185
rect 32050 5140 32100 5165
rect 32050 5110 32060 5140
rect 32090 5110 32100 5140
rect 32050 5085 32100 5110
rect 32050 5065 32065 5085
rect 32085 5065 32100 5085
rect 32050 5040 32100 5065
rect 32050 5010 32060 5040
rect 32090 5010 32100 5040
rect 31450 4910 31460 4940
rect 31490 4910 31500 4940
rect 29350 4815 29365 4835
rect 29385 4815 29400 4835
rect 29350 4785 29400 4815
rect 29350 4765 29365 4785
rect 29385 4765 29400 4785
rect 29350 4735 29400 4765
rect 29350 4715 29365 4735
rect 29385 4715 29400 4735
rect 29350 4685 29400 4715
rect 29350 4665 29365 4685
rect 29385 4665 29400 4685
rect 29350 4635 29400 4665
rect 29350 4615 29365 4635
rect 29385 4615 29400 4635
rect 29350 4585 29400 4615
rect 29350 4565 29365 4585
rect 29385 4565 29400 4585
rect 29350 4535 29400 4565
rect 29350 4515 29365 4535
rect 29385 4515 29400 4535
rect 29350 4485 29400 4515
rect 29350 4465 29365 4485
rect 29385 4465 29400 4485
rect 29350 4435 29400 4465
rect 29500 4835 31350 4850
rect 29500 4815 29515 4835
rect 29535 4815 29815 4835
rect 29835 4815 30115 4835
rect 30135 4815 30415 4835
rect 30435 4815 30715 4835
rect 30735 4815 31015 4835
rect 31035 4815 31315 4835
rect 31335 4815 31350 4835
rect 29500 4800 31350 4815
rect 29500 4785 29550 4800
rect 29500 4765 29515 4785
rect 29535 4765 29550 4785
rect 29500 4735 29550 4765
rect 29800 4785 29850 4800
rect 29800 4765 29815 4785
rect 29835 4765 29850 4785
rect 29500 4715 29515 4735
rect 29535 4715 29550 4735
rect 29500 4685 29550 4715
rect 29500 4665 29515 4685
rect 29535 4665 29550 4685
rect 29500 4635 29550 4665
rect 29500 4615 29515 4635
rect 29535 4615 29550 4635
rect 29500 4585 29550 4615
rect 29500 4565 29515 4585
rect 29535 4565 29550 4585
rect 29500 4535 29550 4565
rect 29500 4515 29515 4535
rect 29535 4515 29550 4535
rect 29500 4485 29550 4515
rect 29500 4465 29515 4485
rect 29535 4465 29550 4485
rect 29500 4450 29550 4465
rect 29650 4735 29700 4750
rect 29650 4715 29665 4735
rect 29685 4715 29700 4735
rect 29650 4685 29700 4715
rect 29650 4665 29665 4685
rect 29685 4665 29700 4685
rect 29650 4635 29700 4665
rect 29650 4615 29665 4635
rect 29685 4615 29700 4635
rect 29650 4585 29700 4615
rect 29650 4565 29665 4585
rect 29685 4565 29700 4585
rect 29650 4535 29700 4565
rect 29650 4515 29665 4535
rect 29685 4515 29700 4535
rect 29650 4485 29700 4515
rect 29650 4465 29665 4485
rect 29685 4465 29700 4485
rect 29350 4415 29365 4435
rect 29385 4415 29400 4435
rect 29350 4400 29400 4415
rect 29650 4435 29700 4465
rect 29650 4415 29665 4435
rect 29685 4415 29700 4435
rect 29650 4400 29700 4415
rect 29350 4385 29700 4400
rect 29350 4365 29365 4385
rect 29385 4365 29665 4385
rect 29685 4365 29700 4385
rect 29350 4350 29700 4365
rect 29800 4735 29850 4765
rect 30100 4785 30150 4800
rect 30100 4765 30115 4785
rect 30135 4765 30150 4785
rect 29800 4715 29815 4735
rect 29835 4715 29850 4735
rect 29800 4685 29850 4715
rect 29800 4665 29815 4685
rect 29835 4665 29850 4685
rect 29800 4635 29850 4665
rect 29800 4615 29815 4635
rect 29835 4615 29850 4635
rect 29800 4585 29850 4615
rect 29800 4565 29815 4585
rect 29835 4565 29850 4585
rect 29800 4535 29850 4565
rect 29800 4515 29815 4535
rect 29835 4515 29850 4535
rect 29800 4485 29850 4515
rect 29800 4465 29815 4485
rect 29835 4465 29850 4485
rect 29800 4435 29850 4465
rect 29800 4415 29815 4435
rect 29835 4415 29850 4435
rect 29800 4385 29850 4415
rect 29800 4365 29815 4385
rect 29835 4365 29850 4385
rect 29800 4350 29850 4365
rect 29950 4735 30000 4750
rect 29950 4715 29965 4735
rect 29985 4715 30000 4735
rect 29950 4685 30000 4715
rect 29950 4665 29965 4685
rect 29985 4665 30000 4685
rect 29950 4635 30000 4665
rect 29950 4615 29965 4635
rect 29985 4615 30000 4635
rect 29950 4585 30000 4615
rect 29950 4565 29965 4585
rect 29985 4565 30000 4585
rect 29950 4535 30000 4565
rect 29950 4515 29965 4535
rect 29985 4515 30000 4535
rect 29950 4485 30000 4515
rect 29950 4465 29965 4485
rect 29985 4465 30000 4485
rect 29950 4435 30000 4465
rect 30100 4735 30150 4765
rect 30400 4785 30450 4800
rect 30400 4765 30415 4785
rect 30435 4765 30450 4785
rect 30100 4715 30115 4735
rect 30135 4715 30150 4735
rect 30100 4685 30150 4715
rect 30100 4665 30115 4685
rect 30135 4665 30150 4685
rect 30100 4635 30150 4665
rect 30100 4615 30115 4635
rect 30135 4615 30150 4635
rect 30100 4585 30150 4615
rect 30100 4565 30115 4585
rect 30135 4565 30150 4585
rect 30100 4535 30150 4565
rect 30100 4515 30115 4535
rect 30135 4515 30150 4535
rect 30100 4485 30150 4515
rect 30100 4465 30115 4485
rect 30135 4465 30150 4485
rect 30100 4450 30150 4465
rect 30250 4735 30300 4750
rect 30250 4715 30265 4735
rect 30285 4715 30300 4735
rect 30250 4685 30300 4715
rect 30250 4665 30265 4685
rect 30285 4665 30300 4685
rect 30250 4635 30300 4665
rect 30250 4615 30265 4635
rect 30285 4615 30300 4635
rect 30250 4585 30300 4615
rect 30250 4565 30265 4585
rect 30285 4565 30300 4585
rect 30250 4535 30300 4565
rect 30250 4515 30265 4535
rect 30285 4515 30300 4535
rect 30250 4485 30300 4515
rect 30250 4465 30265 4485
rect 30285 4465 30300 4485
rect 29950 4415 29965 4435
rect 29985 4415 30000 4435
rect 29950 4400 30000 4415
rect 30250 4435 30300 4465
rect 30250 4415 30265 4435
rect 30285 4415 30300 4435
rect 30250 4400 30300 4415
rect 30400 4735 30450 4765
rect 30700 4785 30750 4800
rect 30700 4765 30715 4785
rect 30735 4765 30750 4785
rect 30400 4715 30415 4735
rect 30435 4715 30450 4735
rect 30400 4685 30450 4715
rect 30400 4665 30415 4685
rect 30435 4665 30450 4685
rect 30400 4635 30450 4665
rect 30400 4615 30415 4635
rect 30435 4615 30450 4635
rect 30400 4585 30450 4615
rect 30400 4565 30415 4585
rect 30435 4565 30450 4585
rect 30400 4535 30450 4565
rect 30400 4515 30415 4535
rect 30435 4515 30450 4535
rect 30400 4485 30450 4515
rect 30400 4465 30415 4485
rect 30435 4465 30450 4485
rect 30400 4435 30450 4465
rect 30400 4415 30415 4435
rect 30435 4415 30450 4435
rect 30400 4400 30450 4415
rect 30550 4735 30600 4750
rect 30550 4715 30565 4735
rect 30585 4715 30600 4735
rect 30550 4685 30600 4715
rect 30550 4665 30565 4685
rect 30585 4665 30600 4685
rect 30550 4635 30600 4665
rect 30550 4615 30565 4635
rect 30585 4615 30600 4635
rect 30550 4585 30600 4615
rect 30550 4565 30565 4585
rect 30585 4565 30600 4585
rect 30550 4535 30600 4565
rect 30550 4515 30565 4535
rect 30585 4515 30600 4535
rect 30550 4485 30600 4515
rect 30550 4465 30565 4485
rect 30585 4465 30600 4485
rect 30550 4435 30600 4465
rect 30700 4735 30750 4765
rect 31000 4785 31050 4800
rect 31000 4765 31015 4785
rect 31035 4765 31050 4785
rect 30700 4715 30715 4735
rect 30735 4715 30750 4735
rect 30700 4685 30750 4715
rect 30700 4665 30715 4685
rect 30735 4665 30750 4685
rect 30700 4635 30750 4665
rect 30700 4615 30715 4635
rect 30735 4615 30750 4635
rect 30700 4585 30750 4615
rect 30700 4565 30715 4585
rect 30735 4565 30750 4585
rect 30700 4535 30750 4565
rect 30700 4515 30715 4535
rect 30735 4515 30750 4535
rect 30700 4485 30750 4515
rect 30700 4465 30715 4485
rect 30735 4465 30750 4485
rect 30700 4450 30750 4465
rect 30850 4735 30900 4750
rect 30850 4715 30865 4735
rect 30885 4715 30900 4735
rect 30850 4685 30900 4715
rect 30850 4665 30865 4685
rect 30885 4665 30900 4685
rect 30850 4635 30900 4665
rect 30850 4615 30865 4635
rect 30885 4615 30900 4635
rect 30850 4585 30900 4615
rect 30850 4565 30865 4585
rect 30885 4565 30900 4585
rect 30850 4535 30900 4565
rect 30850 4515 30865 4535
rect 30885 4515 30900 4535
rect 30850 4485 30900 4515
rect 30850 4465 30865 4485
rect 30885 4465 30900 4485
rect 30550 4415 30565 4435
rect 30585 4415 30600 4435
rect 30550 4400 30600 4415
rect 30850 4435 30900 4465
rect 30850 4415 30865 4435
rect 30885 4415 30900 4435
rect 30850 4400 30900 4415
rect 29950 4385 30900 4400
rect 29950 4365 29965 4385
rect 29985 4365 30265 4385
rect 30285 4365 30415 4385
rect 30435 4365 30565 4385
rect 30585 4365 30865 4385
rect 30885 4365 30900 4385
rect 29950 4350 30900 4365
rect 31000 4735 31050 4765
rect 31300 4785 31350 4800
rect 31300 4765 31315 4785
rect 31335 4765 31350 4785
rect 31000 4715 31015 4735
rect 31035 4715 31050 4735
rect 31000 4685 31050 4715
rect 31000 4665 31015 4685
rect 31035 4665 31050 4685
rect 31000 4635 31050 4665
rect 31000 4615 31015 4635
rect 31035 4615 31050 4635
rect 31000 4585 31050 4615
rect 31000 4565 31015 4585
rect 31035 4565 31050 4585
rect 31000 4535 31050 4565
rect 31000 4515 31015 4535
rect 31035 4515 31050 4535
rect 31000 4485 31050 4515
rect 31000 4465 31015 4485
rect 31035 4465 31050 4485
rect 31000 4435 31050 4465
rect 31000 4415 31015 4435
rect 31035 4415 31050 4435
rect 31000 4385 31050 4415
rect 31000 4365 31015 4385
rect 31035 4365 31050 4385
rect 29350 4200 29400 4350
rect 29350 4185 29700 4200
rect 29350 4165 29365 4185
rect 29385 4165 29665 4185
rect 29685 4165 29700 4185
rect 29350 4150 29700 4165
rect 29350 4135 29400 4150
rect 29350 4115 29365 4135
rect 29385 4115 29400 4135
rect 29350 4085 29400 4115
rect 29650 4135 29700 4150
rect 29650 4115 29665 4135
rect 29685 4115 29700 4135
rect 29350 4065 29365 4085
rect 29385 4065 29400 4085
rect 29350 4035 29400 4065
rect 29350 4015 29365 4035
rect 29385 4015 29400 4035
rect 29350 3985 29400 4015
rect 29350 3965 29365 3985
rect 29385 3965 29400 3985
rect 29350 3935 29400 3965
rect 29350 3915 29365 3935
rect 29385 3915 29400 3935
rect 29350 3885 29400 3915
rect 29350 3865 29365 3885
rect 29385 3865 29400 3885
rect 29350 3835 29400 3865
rect 29350 3815 29365 3835
rect 29385 3815 29400 3835
rect 29350 3785 29400 3815
rect 29350 3765 29365 3785
rect 29385 3765 29400 3785
rect 29350 3735 29400 3765
rect 29350 3715 29365 3735
rect 29385 3715 29400 3735
rect 28750 3610 28760 3640
rect 28790 3610 28800 3640
rect 28150 3510 28160 3540
rect 28190 3510 28200 3540
rect 28150 3485 28200 3510
rect 28150 3465 28165 3485
rect 28185 3465 28200 3485
rect 28150 3440 28200 3465
rect 28150 3410 28160 3440
rect 28190 3410 28200 3440
rect 28150 3385 28200 3410
rect 28150 3365 28165 3385
rect 28185 3365 28200 3385
rect 28150 3340 28200 3365
rect 28150 3310 28160 3340
rect 28190 3310 28200 3340
rect 28150 3285 28200 3310
rect 28150 3265 28165 3285
rect 28185 3265 28200 3285
rect 28150 3240 28200 3265
rect 28150 3210 28160 3240
rect 28190 3210 28200 3240
rect 28150 3185 28200 3210
rect 28150 3165 28165 3185
rect 28185 3165 28200 3185
rect 28150 3140 28200 3165
rect 28150 3110 28160 3140
rect 28190 3110 28200 3140
rect 28150 3085 28200 3110
rect 28150 3065 28165 3085
rect 28185 3065 28200 3085
rect 24550 2960 24560 2990
rect 24590 2960 24600 2990
rect 24550 2950 24600 2960
rect 28150 2990 28200 3065
rect 28150 2960 28160 2990
rect 28190 2960 28200 2990
rect 28150 2950 28200 2960
rect 28750 3540 28800 3610
rect 28900 3640 28950 3650
rect 28900 3610 28910 3640
rect 28940 3610 28950 3640
rect 28900 3600 28950 3610
rect 29200 3640 29250 3650
rect 29200 3610 29210 3640
rect 29240 3610 29250 3640
rect 29200 3600 29250 3610
rect 29350 3640 29400 3715
rect 29500 4085 29550 4100
rect 29500 4065 29515 4085
rect 29535 4065 29550 4085
rect 29500 4035 29550 4065
rect 29500 4015 29515 4035
rect 29535 4015 29550 4035
rect 29500 3985 29550 4015
rect 29500 3965 29515 3985
rect 29535 3965 29550 3985
rect 29500 3935 29550 3965
rect 29500 3915 29515 3935
rect 29535 3915 29550 3935
rect 29500 3885 29550 3915
rect 29500 3865 29515 3885
rect 29535 3865 29550 3885
rect 29500 3835 29550 3865
rect 29500 3815 29515 3835
rect 29535 3815 29550 3835
rect 29500 3785 29550 3815
rect 29650 4085 29700 4115
rect 29650 4065 29665 4085
rect 29685 4065 29700 4085
rect 29650 4035 29700 4065
rect 29650 4015 29665 4035
rect 29685 4015 29700 4035
rect 29650 3985 29700 4015
rect 29650 3965 29665 3985
rect 29685 3965 29700 3985
rect 29650 3935 29700 3965
rect 29650 3915 29665 3935
rect 29685 3915 29700 3935
rect 29650 3885 29700 3915
rect 29650 3865 29665 3885
rect 29685 3865 29700 3885
rect 29650 3835 29700 3865
rect 29650 3815 29665 3835
rect 29685 3815 29700 3835
rect 29650 3800 29700 3815
rect 29800 4185 29850 4200
rect 29800 4165 29815 4185
rect 29835 4165 29850 4185
rect 29800 4135 29850 4165
rect 29800 4115 29815 4135
rect 29835 4115 29850 4135
rect 29800 4085 29850 4115
rect 29800 4065 29815 4085
rect 29835 4065 29850 4085
rect 29800 4035 29850 4065
rect 29800 4015 29815 4035
rect 29835 4015 29850 4035
rect 29800 3985 29850 4015
rect 29800 3965 29815 3985
rect 29835 3965 29850 3985
rect 29800 3935 29850 3965
rect 29800 3915 29815 3935
rect 29835 3915 29850 3935
rect 29800 3885 29850 3915
rect 29800 3865 29815 3885
rect 29835 3865 29850 3885
rect 29800 3835 29850 3865
rect 29800 3815 29815 3835
rect 29835 3815 29850 3835
rect 29500 3765 29515 3785
rect 29535 3765 29550 3785
rect 29500 3750 29550 3765
rect 29800 3785 29850 3815
rect 29950 4185 30900 4200
rect 29950 4165 29965 4185
rect 29985 4165 30265 4185
rect 30285 4165 30415 4185
rect 30435 4165 30565 4185
rect 30585 4165 30865 4185
rect 30885 4165 30900 4185
rect 29950 4150 30900 4165
rect 29950 4135 30000 4150
rect 29950 4115 29965 4135
rect 29985 4115 30000 4135
rect 29950 4085 30000 4115
rect 30250 4135 30300 4150
rect 30250 4115 30265 4135
rect 30285 4115 30300 4135
rect 29950 4065 29965 4085
rect 29985 4065 30000 4085
rect 29950 4035 30000 4065
rect 29950 4015 29965 4035
rect 29985 4015 30000 4035
rect 29950 3985 30000 4015
rect 29950 3965 29965 3985
rect 29985 3965 30000 3985
rect 29950 3935 30000 3965
rect 29950 3915 29965 3935
rect 29985 3915 30000 3935
rect 29950 3885 30000 3915
rect 29950 3865 29965 3885
rect 29985 3865 30000 3885
rect 29950 3835 30000 3865
rect 29950 3815 29965 3835
rect 29985 3815 30000 3835
rect 29950 3800 30000 3815
rect 30100 4085 30150 4100
rect 30100 4065 30115 4085
rect 30135 4065 30150 4085
rect 30100 4035 30150 4065
rect 30100 4015 30115 4035
rect 30135 4015 30150 4035
rect 30100 3985 30150 4015
rect 30100 3965 30115 3985
rect 30135 3965 30150 3985
rect 30100 3935 30150 3965
rect 30100 3915 30115 3935
rect 30135 3915 30150 3935
rect 30100 3885 30150 3915
rect 30100 3865 30115 3885
rect 30135 3865 30150 3885
rect 30100 3835 30150 3865
rect 30100 3815 30115 3835
rect 30135 3815 30150 3835
rect 29800 3765 29815 3785
rect 29835 3765 29850 3785
rect 29800 3750 29850 3765
rect 30100 3785 30150 3815
rect 30250 4085 30300 4115
rect 30250 4065 30265 4085
rect 30285 4065 30300 4085
rect 30250 4035 30300 4065
rect 30250 4015 30265 4035
rect 30285 4015 30300 4035
rect 30250 3985 30300 4015
rect 30250 3965 30265 3985
rect 30285 3965 30300 3985
rect 30250 3935 30300 3965
rect 30250 3915 30265 3935
rect 30285 3915 30300 3935
rect 30250 3885 30300 3915
rect 30250 3865 30265 3885
rect 30285 3865 30300 3885
rect 30250 3835 30300 3865
rect 30250 3815 30265 3835
rect 30285 3815 30300 3835
rect 30250 3800 30300 3815
rect 30400 4135 30450 4150
rect 30400 4115 30415 4135
rect 30435 4115 30450 4135
rect 30400 4085 30450 4115
rect 30400 4065 30415 4085
rect 30435 4065 30450 4085
rect 30400 4035 30450 4065
rect 30400 4015 30415 4035
rect 30435 4015 30450 4035
rect 30400 3985 30450 4015
rect 30400 3965 30415 3985
rect 30435 3965 30450 3985
rect 30400 3935 30450 3965
rect 30400 3915 30415 3935
rect 30435 3915 30450 3935
rect 30400 3885 30450 3915
rect 30400 3865 30415 3885
rect 30435 3865 30450 3885
rect 30400 3835 30450 3865
rect 30400 3815 30415 3835
rect 30435 3815 30450 3835
rect 30100 3765 30115 3785
rect 30135 3765 30150 3785
rect 30100 3750 30150 3765
rect 30400 3785 30450 3815
rect 30550 4135 30600 4150
rect 30550 4115 30565 4135
rect 30585 4115 30600 4135
rect 30550 4085 30600 4115
rect 30850 4135 30900 4150
rect 30850 4115 30865 4135
rect 30885 4115 30900 4135
rect 30550 4065 30565 4085
rect 30585 4065 30600 4085
rect 30550 4035 30600 4065
rect 30550 4015 30565 4035
rect 30585 4015 30600 4035
rect 30550 3985 30600 4015
rect 30550 3965 30565 3985
rect 30585 3965 30600 3985
rect 30550 3935 30600 3965
rect 30550 3915 30565 3935
rect 30585 3915 30600 3935
rect 30550 3885 30600 3915
rect 30550 3865 30565 3885
rect 30585 3865 30600 3885
rect 30550 3835 30600 3865
rect 30550 3815 30565 3835
rect 30585 3815 30600 3835
rect 30550 3800 30600 3815
rect 30700 4085 30750 4100
rect 30700 4065 30715 4085
rect 30735 4065 30750 4085
rect 30700 4035 30750 4065
rect 30700 4015 30715 4035
rect 30735 4015 30750 4035
rect 30700 3985 30750 4015
rect 30700 3965 30715 3985
rect 30735 3965 30750 3985
rect 30700 3935 30750 3965
rect 30700 3915 30715 3935
rect 30735 3915 30750 3935
rect 30700 3885 30750 3915
rect 30700 3865 30715 3885
rect 30735 3865 30750 3885
rect 30700 3835 30750 3865
rect 30700 3815 30715 3835
rect 30735 3815 30750 3835
rect 30400 3765 30415 3785
rect 30435 3765 30450 3785
rect 30400 3750 30450 3765
rect 30700 3785 30750 3815
rect 30850 4085 30900 4115
rect 30850 4065 30865 4085
rect 30885 4065 30900 4085
rect 30850 4035 30900 4065
rect 30850 4015 30865 4035
rect 30885 4015 30900 4035
rect 30850 3985 30900 4015
rect 30850 3965 30865 3985
rect 30885 3965 30900 3985
rect 30850 3935 30900 3965
rect 30850 3915 30865 3935
rect 30885 3915 30900 3935
rect 30850 3885 30900 3915
rect 30850 3865 30865 3885
rect 30885 3865 30900 3885
rect 30850 3835 30900 3865
rect 30850 3815 30865 3835
rect 30885 3815 30900 3835
rect 30850 3800 30900 3815
rect 31000 4185 31050 4365
rect 31150 4735 31200 4750
rect 31150 4715 31165 4735
rect 31185 4715 31200 4735
rect 31150 4685 31200 4715
rect 31150 4665 31165 4685
rect 31185 4665 31200 4685
rect 31150 4635 31200 4665
rect 31150 4615 31165 4635
rect 31185 4615 31200 4635
rect 31150 4585 31200 4615
rect 31150 4565 31165 4585
rect 31185 4565 31200 4585
rect 31150 4535 31200 4565
rect 31150 4515 31165 4535
rect 31185 4515 31200 4535
rect 31150 4485 31200 4515
rect 31150 4465 31165 4485
rect 31185 4465 31200 4485
rect 31150 4435 31200 4465
rect 31300 4735 31350 4765
rect 31300 4715 31315 4735
rect 31335 4715 31350 4735
rect 31300 4685 31350 4715
rect 31300 4665 31315 4685
rect 31335 4665 31350 4685
rect 31300 4635 31350 4665
rect 31300 4615 31315 4635
rect 31335 4615 31350 4635
rect 31300 4585 31350 4615
rect 31300 4565 31315 4585
rect 31335 4565 31350 4585
rect 31300 4535 31350 4565
rect 31300 4515 31315 4535
rect 31335 4515 31350 4535
rect 31300 4485 31350 4515
rect 31300 4465 31315 4485
rect 31335 4465 31350 4485
rect 31300 4450 31350 4465
rect 31450 4835 31500 4910
rect 31600 4940 31650 4950
rect 31600 4910 31610 4940
rect 31640 4910 31650 4940
rect 31600 4900 31650 4910
rect 31900 4940 31950 4950
rect 31900 4910 31910 4940
rect 31940 4910 31950 4940
rect 31900 4900 31950 4910
rect 32050 4940 32100 5010
rect 32050 4910 32060 4940
rect 32090 4910 32100 4940
rect 31450 4815 31465 4835
rect 31485 4815 31500 4835
rect 31450 4785 31500 4815
rect 31450 4765 31465 4785
rect 31485 4765 31500 4785
rect 31450 4735 31500 4765
rect 31450 4715 31465 4735
rect 31485 4715 31500 4735
rect 31450 4685 31500 4715
rect 31450 4665 31465 4685
rect 31485 4665 31500 4685
rect 31450 4635 31500 4665
rect 31450 4615 31465 4635
rect 31485 4615 31500 4635
rect 31450 4585 31500 4615
rect 31450 4565 31465 4585
rect 31485 4565 31500 4585
rect 31450 4535 31500 4565
rect 31450 4515 31465 4535
rect 31485 4515 31500 4535
rect 31450 4485 31500 4515
rect 31450 4465 31465 4485
rect 31485 4465 31500 4485
rect 31150 4415 31165 4435
rect 31185 4415 31200 4435
rect 31150 4400 31200 4415
rect 31450 4435 31500 4465
rect 31450 4415 31465 4435
rect 31485 4415 31500 4435
rect 31450 4400 31500 4415
rect 31150 4385 31500 4400
rect 31150 4365 31165 4385
rect 31185 4365 31465 4385
rect 31485 4365 31500 4385
rect 31150 4350 31500 4365
rect 31450 4200 31500 4350
rect 31000 4165 31015 4185
rect 31035 4165 31050 4185
rect 31000 4135 31050 4165
rect 31000 4115 31015 4135
rect 31035 4115 31050 4135
rect 31000 4085 31050 4115
rect 31000 4065 31015 4085
rect 31035 4065 31050 4085
rect 31000 4035 31050 4065
rect 31000 4015 31015 4035
rect 31035 4015 31050 4035
rect 31000 3985 31050 4015
rect 31000 3965 31015 3985
rect 31035 3965 31050 3985
rect 31000 3935 31050 3965
rect 31000 3915 31015 3935
rect 31035 3915 31050 3935
rect 31000 3885 31050 3915
rect 31000 3865 31015 3885
rect 31035 3865 31050 3885
rect 31000 3835 31050 3865
rect 31000 3815 31015 3835
rect 31035 3815 31050 3835
rect 30700 3765 30715 3785
rect 30735 3765 30750 3785
rect 30700 3750 30750 3765
rect 31000 3785 31050 3815
rect 31150 4185 31500 4200
rect 31150 4165 31165 4185
rect 31185 4165 31465 4185
rect 31485 4165 31500 4185
rect 31150 4150 31500 4165
rect 31150 4135 31200 4150
rect 31150 4115 31165 4135
rect 31185 4115 31200 4135
rect 31150 4085 31200 4115
rect 31450 4135 31500 4150
rect 31450 4115 31465 4135
rect 31485 4115 31500 4135
rect 31150 4065 31165 4085
rect 31185 4065 31200 4085
rect 31150 4035 31200 4065
rect 31150 4015 31165 4035
rect 31185 4015 31200 4035
rect 31150 3985 31200 4015
rect 31150 3965 31165 3985
rect 31185 3965 31200 3985
rect 31150 3935 31200 3965
rect 31150 3915 31165 3935
rect 31185 3915 31200 3935
rect 31150 3885 31200 3915
rect 31150 3865 31165 3885
rect 31185 3865 31200 3885
rect 31150 3835 31200 3865
rect 31150 3815 31165 3835
rect 31185 3815 31200 3835
rect 31150 3800 31200 3815
rect 31300 4085 31350 4100
rect 31300 4065 31315 4085
rect 31335 4065 31350 4085
rect 31300 4035 31350 4065
rect 31300 4015 31315 4035
rect 31335 4015 31350 4035
rect 31300 3985 31350 4015
rect 31300 3965 31315 3985
rect 31335 3965 31350 3985
rect 31300 3935 31350 3965
rect 31300 3915 31315 3935
rect 31335 3915 31350 3935
rect 31300 3885 31350 3915
rect 31300 3865 31315 3885
rect 31335 3865 31350 3885
rect 31300 3835 31350 3865
rect 31300 3815 31315 3835
rect 31335 3815 31350 3835
rect 31000 3765 31015 3785
rect 31035 3765 31050 3785
rect 31000 3750 31050 3765
rect 31300 3785 31350 3815
rect 31300 3765 31315 3785
rect 31335 3765 31350 3785
rect 31300 3750 31350 3765
rect 29500 3735 31350 3750
rect 29500 3715 29515 3735
rect 29535 3715 29815 3735
rect 29835 3715 30115 3735
rect 30135 3715 30415 3735
rect 30435 3715 30715 3735
rect 30735 3715 31015 3735
rect 31035 3715 31315 3735
rect 31335 3715 31350 3735
rect 29500 3700 31350 3715
rect 31450 4085 31500 4115
rect 31450 4065 31465 4085
rect 31485 4065 31500 4085
rect 31450 4035 31500 4065
rect 31450 4015 31465 4035
rect 31485 4015 31500 4035
rect 31450 3985 31500 4015
rect 31450 3965 31465 3985
rect 31485 3965 31500 3985
rect 31450 3935 31500 3965
rect 31450 3915 31465 3935
rect 31485 3915 31500 3935
rect 31450 3885 31500 3915
rect 31450 3865 31465 3885
rect 31485 3865 31500 3885
rect 31450 3835 31500 3865
rect 31450 3815 31465 3835
rect 31485 3815 31500 3835
rect 31450 3785 31500 3815
rect 31450 3765 31465 3785
rect 31485 3765 31500 3785
rect 31450 3735 31500 3765
rect 31450 3715 31465 3735
rect 31485 3715 31500 3735
rect 29350 3610 29360 3640
rect 29390 3610 29400 3640
rect 28750 3510 28760 3540
rect 28790 3510 28800 3540
rect 28750 3485 28800 3510
rect 28750 3465 28765 3485
rect 28785 3465 28800 3485
rect 28750 3440 28800 3465
rect 28750 3410 28760 3440
rect 28790 3410 28800 3440
rect 28750 3385 28800 3410
rect 28750 3365 28765 3385
rect 28785 3365 28800 3385
rect 28750 3340 28800 3365
rect 28750 3310 28760 3340
rect 28790 3310 28800 3340
rect 28750 3285 28800 3310
rect 28750 3265 28765 3285
rect 28785 3265 28800 3285
rect 28750 3240 28800 3265
rect 28750 3210 28760 3240
rect 28790 3210 28800 3240
rect 28750 3185 28800 3210
rect 28750 3165 28765 3185
rect 28785 3165 28800 3185
rect 28750 3140 28800 3165
rect 28750 3110 28760 3140
rect 28790 3110 28800 3140
rect 28750 3085 28800 3110
rect 28750 3065 28765 3085
rect 28785 3065 28800 3085
rect 28750 2990 28800 3065
rect 29350 3535 29400 3610
rect 29650 3640 29700 3650
rect 29650 3610 29660 3640
rect 29690 3610 29700 3640
rect 29650 3600 29700 3610
rect 29950 3640 30000 3650
rect 29950 3610 29960 3640
rect 29990 3610 30000 3640
rect 29950 3600 30000 3610
rect 30250 3640 30300 3650
rect 30250 3610 30260 3640
rect 30290 3610 30300 3640
rect 30250 3600 30300 3610
rect 30550 3640 30600 3650
rect 30550 3610 30560 3640
rect 30590 3610 30600 3640
rect 30550 3600 30600 3610
rect 30850 3640 30900 3650
rect 30850 3610 30860 3640
rect 30890 3610 30900 3640
rect 30850 3600 30900 3610
rect 31150 3640 31200 3650
rect 31150 3610 31160 3640
rect 31190 3610 31200 3640
rect 31150 3600 31200 3610
rect 31450 3640 31500 3715
rect 32050 4840 32100 4910
rect 32050 4810 32060 4840
rect 32090 4810 32100 4840
rect 32050 4785 32100 4810
rect 32050 4765 32065 4785
rect 32085 4765 32100 4785
rect 32050 4740 32100 4765
rect 32050 4710 32060 4740
rect 32090 4710 32100 4740
rect 32050 4685 32100 4710
rect 32050 4665 32065 4685
rect 32085 4665 32100 4685
rect 32050 4640 32100 4665
rect 32050 4610 32060 4640
rect 32090 4610 32100 4640
rect 32050 4585 32100 4610
rect 32050 4565 32065 4585
rect 32085 4565 32100 4585
rect 32050 4540 32100 4565
rect 32050 4510 32060 4540
rect 32090 4510 32100 4540
rect 32050 4485 32100 4510
rect 32050 4465 32065 4485
rect 32085 4465 32100 4485
rect 32050 4440 32100 4465
rect 32050 4410 32060 4440
rect 32090 4410 32100 4440
rect 32050 4385 32100 4410
rect 32050 4365 32065 4385
rect 32085 4365 32100 4385
rect 32050 4290 32100 4365
rect 32050 4260 32060 4290
rect 32090 4260 32100 4290
rect 32050 4185 32100 4260
rect 32050 4165 32065 4185
rect 32085 4165 32100 4185
rect 32050 4140 32100 4165
rect 32050 4110 32060 4140
rect 32090 4110 32100 4140
rect 32050 4085 32100 4110
rect 32050 4065 32065 4085
rect 32085 4065 32100 4085
rect 32050 4040 32100 4065
rect 32050 4010 32060 4040
rect 32090 4010 32100 4040
rect 32050 3985 32100 4010
rect 32050 3965 32065 3985
rect 32085 3965 32100 3985
rect 32050 3940 32100 3965
rect 32050 3910 32060 3940
rect 32090 3910 32100 3940
rect 32050 3885 32100 3910
rect 32050 3865 32065 3885
rect 32085 3865 32100 3885
rect 32050 3840 32100 3865
rect 32050 3810 32060 3840
rect 32090 3810 32100 3840
rect 32050 3785 32100 3810
rect 32050 3765 32065 3785
rect 32085 3765 32100 3785
rect 32050 3740 32100 3765
rect 32050 3710 32060 3740
rect 32090 3710 32100 3740
rect 31450 3610 31460 3640
rect 31490 3610 31500 3640
rect 29350 3515 29365 3535
rect 29385 3515 29400 3535
rect 29350 3485 29400 3515
rect 29350 3465 29365 3485
rect 29385 3465 29400 3485
rect 29350 3435 29400 3465
rect 29350 3415 29365 3435
rect 29385 3415 29400 3435
rect 29350 3385 29400 3415
rect 29350 3365 29365 3385
rect 29385 3365 29400 3385
rect 29350 3335 29400 3365
rect 29350 3315 29365 3335
rect 29385 3315 29400 3335
rect 29350 3285 29400 3315
rect 29350 3265 29365 3285
rect 29385 3265 29400 3285
rect 29350 3235 29400 3265
rect 29350 3215 29365 3235
rect 29385 3215 29400 3235
rect 29350 3185 29400 3215
rect 29350 3165 29365 3185
rect 29385 3165 29400 3185
rect 29350 3135 29400 3165
rect 29500 3535 31350 3550
rect 29500 3515 29515 3535
rect 29535 3515 29815 3535
rect 29835 3515 30115 3535
rect 30135 3515 30415 3535
rect 30435 3515 30715 3535
rect 30735 3515 31015 3535
rect 31035 3515 31315 3535
rect 31335 3515 31350 3535
rect 29500 3500 31350 3515
rect 29500 3485 29550 3500
rect 29500 3465 29515 3485
rect 29535 3465 29550 3485
rect 29500 3435 29550 3465
rect 29800 3485 29850 3500
rect 29800 3465 29815 3485
rect 29835 3465 29850 3485
rect 29500 3415 29515 3435
rect 29535 3415 29550 3435
rect 29500 3385 29550 3415
rect 29500 3365 29515 3385
rect 29535 3365 29550 3385
rect 29500 3335 29550 3365
rect 29500 3315 29515 3335
rect 29535 3315 29550 3335
rect 29500 3285 29550 3315
rect 29500 3265 29515 3285
rect 29535 3265 29550 3285
rect 29500 3235 29550 3265
rect 29500 3215 29515 3235
rect 29535 3215 29550 3235
rect 29500 3185 29550 3215
rect 29500 3165 29515 3185
rect 29535 3165 29550 3185
rect 29500 3150 29550 3165
rect 29650 3435 29700 3450
rect 29650 3415 29665 3435
rect 29685 3415 29700 3435
rect 29650 3385 29700 3415
rect 29650 3365 29665 3385
rect 29685 3365 29700 3385
rect 29650 3335 29700 3365
rect 29650 3315 29665 3335
rect 29685 3315 29700 3335
rect 29650 3285 29700 3315
rect 29650 3265 29665 3285
rect 29685 3265 29700 3285
rect 29650 3235 29700 3265
rect 29650 3215 29665 3235
rect 29685 3215 29700 3235
rect 29650 3185 29700 3215
rect 29650 3165 29665 3185
rect 29685 3165 29700 3185
rect 29350 3115 29365 3135
rect 29385 3115 29400 3135
rect 29350 3100 29400 3115
rect 29650 3135 29700 3165
rect 29650 3115 29665 3135
rect 29685 3115 29700 3135
rect 29650 3100 29700 3115
rect 29350 3085 29700 3100
rect 29350 3065 29365 3085
rect 29385 3065 29665 3085
rect 29685 3065 29700 3085
rect 29350 3050 29700 3065
rect 29800 3435 29850 3465
rect 30100 3485 30150 3500
rect 30100 3465 30115 3485
rect 30135 3465 30150 3485
rect 29800 3415 29815 3435
rect 29835 3415 29850 3435
rect 29800 3385 29850 3415
rect 29800 3365 29815 3385
rect 29835 3365 29850 3385
rect 29800 3335 29850 3365
rect 29800 3315 29815 3335
rect 29835 3315 29850 3335
rect 29800 3285 29850 3315
rect 29800 3265 29815 3285
rect 29835 3265 29850 3285
rect 29800 3235 29850 3265
rect 29800 3215 29815 3235
rect 29835 3215 29850 3235
rect 29800 3185 29850 3215
rect 29800 3165 29815 3185
rect 29835 3165 29850 3185
rect 29800 3135 29850 3165
rect 29800 3115 29815 3135
rect 29835 3115 29850 3135
rect 29800 3085 29850 3115
rect 29800 3065 29815 3085
rect 29835 3065 29850 3085
rect 29800 3050 29850 3065
rect 29950 3435 30000 3450
rect 29950 3415 29965 3435
rect 29985 3415 30000 3435
rect 29950 3385 30000 3415
rect 29950 3365 29965 3385
rect 29985 3365 30000 3385
rect 29950 3335 30000 3365
rect 29950 3315 29965 3335
rect 29985 3315 30000 3335
rect 29950 3285 30000 3315
rect 29950 3265 29965 3285
rect 29985 3265 30000 3285
rect 29950 3235 30000 3265
rect 29950 3215 29965 3235
rect 29985 3215 30000 3235
rect 29950 3185 30000 3215
rect 29950 3165 29965 3185
rect 29985 3165 30000 3185
rect 29950 3135 30000 3165
rect 30100 3435 30150 3465
rect 30400 3485 30450 3500
rect 30400 3465 30415 3485
rect 30435 3465 30450 3485
rect 30100 3415 30115 3435
rect 30135 3415 30150 3435
rect 30100 3385 30150 3415
rect 30100 3365 30115 3385
rect 30135 3365 30150 3385
rect 30100 3335 30150 3365
rect 30100 3315 30115 3335
rect 30135 3315 30150 3335
rect 30100 3285 30150 3315
rect 30100 3265 30115 3285
rect 30135 3265 30150 3285
rect 30100 3235 30150 3265
rect 30100 3215 30115 3235
rect 30135 3215 30150 3235
rect 30100 3185 30150 3215
rect 30100 3165 30115 3185
rect 30135 3165 30150 3185
rect 30100 3150 30150 3165
rect 30250 3435 30300 3450
rect 30250 3415 30265 3435
rect 30285 3415 30300 3435
rect 30250 3385 30300 3415
rect 30250 3365 30265 3385
rect 30285 3365 30300 3385
rect 30250 3335 30300 3365
rect 30250 3315 30265 3335
rect 30285 3315 30300 3335
rect 30250 3285 30300 3315
rect 30250 3265 30265 3285
rect 30285 3265 30300 3285
rect 30250 3235 30300 3265
rect 30250 3215 30265 3235
rect 30285 3215 30300 3235
rect 30250 3185 30300 3215
rect 30250 3165 30265 3185
rect 30285 3165 30300 3185
rect 29950 3115 29965 3135
rect 29985 3115 30000 3135
rect 29950 3100 30000 3115
rect 30250 3135 30300 3165
rect 30400 3435 30450 3465
rect 30700 3485 30750 3500
rect 30700 3465 30715 3485
rect 30735 3465 30750 3485
rect 30400 3415 30415 3435
rect 30435 3415 30450 3435
rect 30400 3385 30450 3415
rect 30400 3365 30415 3385
rect 30435 3365 30450 3385
rect 30400 3335 30450 3365
rect 30400 3315 30415 3335
rect 30435 3315 30450 3335
rect 30400 3285 30450 3315
rect 30400 3265 30415 3285
rect 30435 3265 30450 3285
rect 30400 3235 30450 3265
rect 30400 3215 30415 3235
rect 30435 3215 30450 3235
rect 30400 3185 30450 3215
rect 30400 3165 30415 3185
rect 30435 3165 30450 3185
rect 30400 3150 30450 3165
rect 30550 3435 30600 3450
rect 30550 3415 30565 3435
rect 30585 3415 30600 3435
rect 30550 3385 30600 3415
rect 30550 3365 30565 3385
rect 30585 3365 30600 3385
rect 30550 3335 30600 3365
rect 30550 3315 30565 3335
rect 30585 3315 30600 3335
rect 30550 3285 30600 3315
rect 30550 3265 30565 3285
rect 30585 3265 30600 3285
rect 30550 3235 30600 3265
rect 30550 3215 30565 3235
rect 30585 3215 30600 3235
rect 30550 3185 30600 3215
rect 30550 3165 30565 3185
rect 30585 3165 30600 3185
rect 30250 3115 30265 3135
rect 30285 3115 30300 3135
rect 30250 3100 30300 3115
rect 30550 3135 30600 3165
rect 30700 3435 30750 3465
rect 31000 3485 31050 3500
rect 31000 3465 31015 3485
rect 31035 3465 31050 3485
rect 30700 3415 30715 3435
rect 30735 3415 30750 3435
rect 30700 3385 30750 3415
rect 30700 3365 30715 3385
rect 30735 3365 30750 3385
rect 30700 3335 30750 3365
rect 30700 3315 30715 3335
rect 30735 3315 30750 3335
rect 30700 3285 30750 3315
rect 30700 3265 30715 3285
rect 30735 3265 30750 3285
rect 30700 3235 30750 3265
rect 30700 3215 30715 3235
rect 30735 3215 30750 3235
rect 30700 3185 30750 3215
rect 30700 3165 30715 3185
rect 30735 3165 30750 3185
rect 30700 3150 30750 3165
rect 30850 3435 30900 3450
rect 30850 3415 30865 3435
rect 30885 3415 30900 3435
rect 30850 3385 30900 3415
rect 30850 3365 30865 3385
rect 30885 3365 30900 3385
rect 30850 3335 30900 3365
rect 30850 3315 30865 3335
rect 30885 3315 30900 3335
rect 30850 3285 30900 3315
rect 30850 3265 30865 3285
rect 30885 3265 30900 3285
rect 30850 3235 30900 3265
rect 30850 3215 30865 3235
rect 30885 3215 30900 3235
rect 30850 3185 30900 3215
rect 30850 3165 30865 3185
rect 30885 3165 30900 3185
rect 30550 3115 30565 3135
rect 30585 3115 30600 3135
rect 30550 3100 30600 3115
rect 30850 3135 30900 3165
rect 30850 3115 30865 3135
rect 30885 3115 30900 3135
rect 30850 3100 30900 3115
rect 29950 3085 30900 3100
rect 29950 3065 29965 3085
rect 29985 3065 30265 3085
rect 30285 3065 30565 3085
rect 30585 3065 30865 3085
rect 30885 3065 30900 3085
rect 29950 3050 30900 3065
rect 31000 3435 31050 3465
rect 31300 3485 31350 3500
rect 31300 3465 31315 3485
rect 31335 3465 31350 3485
rect 31000 3415 31015 3435
rect 31035 3415 31050 3435
rect 31000 3385 31050 3415
rect 31000 3365 31015 3385
rect 31035 3365 31050 3385
rect 31000 3335 31050 3365
rect 31000 3315 31015 3335
rect 31035 3315 31050 3335
rect 31000 3285 31050 3315
rect 31000 3265 31015 3285
rect 31035 3265 31050 3285
rect 31000 3235 31050 3265
rect 31000 3215 31015 3235
rect 31035 3215 31050 3235
rect 31000 3185 31050 3215
rect 31000 3165 31015 3185
rect 31035 3165 31050 3185
rect 31000 3135 31050 3165
rect 31000 3115 31015 3135
rect 31035 3115 31050 3135
rect 31000 3085 31050 3115
rect 31000 3065 31015 3085
rect 31035 3065 31050 3085
rect 31000 3050 31050 3065
rect 31150 3435 31200 3450
rect 31150 3415 31165 3435
rect 31185 3415 31200 3435
rect 31150 3385 31200 3415
rect 31150 3365 31165 3385
rect 31185 3365 31200 3385
rect 31150 3335 31200 3365
rect 31150 3315 31165 3335
rect 31185 3315 31200 3335
rect 31150 3285 31200 3315
rect 31150 3265 31165 3285
rect 31185 3265 31200 3285
rect 31150 3235 31200 3265
rect 31150 3215 31165 3235
rect 31185 3215 31200 3235
rect 31150 3185 31200 3215
rect 31150 3165 31165 3185
rect 31185 3165 31200 3185
rect 31150 3135 31200 3165
rect 31300 3435 31350 3465
rect 31300 3415 31315 3435
rect 31335 3415 31350 3435
rect 31300 3385 31350 3415
rect 31300 3365 31315 3385
rect 31335 3365 31350 3385
rect 31300 3335 31350 3365
rect 31300 3315 31315 3335
rect 31335 3315 31350 3335
rect 31300 3285 31350 3315
rect 31300 3265 31315 3285
rect 31335 3265 31350 3285
rect 31300 3235 31350 3265
rect 31300 3215 31315 3235
rect 31335 3215 31350 3235
rect 31300 3185 31350 3215
rect 31300 3165 31315 3185
rect 31335 3165 31350 3185
rect 31300 3150 31350 3165
rect 31450 3535 31500 3610
rect 31600 3640 31650 3650
rect 31600 3610 31610 3640
rect 31640 3610 31650 3640
rect 31600 3600 31650 3610
rect 31900 3640 31950 3650
rect 31900 3610 31910 3640
rect 31940 3610 31950 3640
rect 31900 3600 31950 3610
rect 32050 3640 32100 3710
rect 32050 3610 32060 3640
rect 32090 3610 32100 3640
rect 31450 3515 31465 3535
rect 31485 3515 31500 3535
rect 31450 3485 31500 3515
rect 31450 3465 31465 3485
rect 31485 3465 31500 3485
rect 31450 3435 31500 3465
rect 31450 3415 31465 3435
rect 31485 3415 31500 3435
rect 31450 3385 31500 3415
rect 31450 3365 31465 3385
rect 31485 3365 31500 3385
rect 31450 3335 31500 3365
rect 31450 3315 31465 3335
rect 31485 3315 31500 3335
rect 31450 3285 31500 3315
rect 31450 3265 31465 3285
rect 31485 3265 31500 3285
rect 31450 3235 31500 3265
rect 31450 3215 31465 3235
rect 31485 3215 31500 3235
rect 31450 3185 31500 3215
rect 31450 3165 31465 3185
rect 31485 3165 31500 3185
rect 31150 3115 31165 3135
rect 31185 3115 31200 3135
rect 31150 3100 31200 3115
rect 31450 3135 31500 3165
rect 31450 3115 31465 3135
rect 31485 3115 31500 3135
rect 31450 3100 31500 3115
rect 31150 3085 31500 3100
rect 31150 3065 31165 3085
rect 31185 3065 31465 3085
rect 31485 3065 31500 3085
rect 31150 3050 31500 3065
rect 32050 3540 32100 3610
rect 32050 3510 32060 3540
rect 32090 3510 32100 3540
rect 32050 3485 32100 3510
rect 32050 3465 32065 3485
rect 32085 3465 32100 3485
rect 32050 3440 32100 3465
rect 32050 3410 32060 3440
rect 32090 3410 32100 3440
rect 32050 3385 32100 3410
rect 32050 3365 32065 3385
rect 32085 3365 32100 3385
rect 32050 3340 32100 3365
rect 32050 3310 32060 3340
rect 32090 3310 32100 3340
rect 32050 3285 32100 3310
rect 32050 3265 32065 3285
rect 32085 3265 32100 3285
rect 32050 3240 32100 3265
rect 32050 3210 32060 3240
rect 32090 3210 32100 3240
rect 32050 3185 32100 3210
rect 32050 3165 32065 3185
rect 32085 3165 32100 3185
rect 32050 3140 32100 3165
rect 32050 3110 32060 3140
rect 32090 3110 32100 3140
rect 32050 3085 32100 3110
rect 32050 3065 32065 3085
rect 32085 3065 32100 3085
rect 28750 2960 28760 2990
rect 28790 2960 28800 2990
rect 28750 2950 28800 2960
rect 32050 2990 32100 3065
rect 32050 2960 32060 2990
rect 32090 2960 32100 2990
rect 32050 2950 32100 2960
rect -650 1690 -600 1700
rect -650 1660 -640 1690
rect -610 1660 -600 1690
rect -650 1585 -600 1660
rect -50 1690 0 1700
rect -50 1660 -40 1690
rect -10 1660 0 1690
rect -650 1565 -635 1585
rect -615 1565 -600 1585
rect -650 1540 -600 1565
rect -650 1510 -640 1540
rect -610 1510 -600 1540
rect -650 1485 -600 1510
rect -650 1465 -635 1485
rect -615 1465 -600 1485
rect -650 1440 -600 1465
rect -650 1410 -640 1440
rect -610 1410 -600 1440
rect -650 1385 -600 1410
rect -650 1365 -635 1385
rect -615 1365 -600 1385
rect -650 1340 -600 1365
rect -650 1310 -640 1340
rect -610 1310 -600 1340
rect -650 1285 -600 1310
rect -650 1265 -635 1285
rect -615 1265 -600 1285
rect -650 1240 -600 1265
rect -650 1210 -640 1240
rect -610 1210 -600 1240
rect -650 1185 -600 1210
rect -650 1165 -635 1185
rect -615 1165 -600 1185
rect -650 1140 -600 1165
rect -650 1110 -640 1140
rect -610 1110 -600 1140
rect -650 1085 -600 1110
rect -650 1065 -635 1085
rect -615 1065 -600 1085
rect -650 1040 -600 1065
rect -650 1010 -640 1040
rect -610 1010 -600 1040
rect -650 985 -600 1010
rect -650 965 -635 985
rect -615 965 -600 985
rect -650 940 -600 965
rect -650 910 -640 940
rect -610 910 -600 940
rect -650 740 -600 910
rect -500 1585 -450 1600
rect -500 1565 -485 1585
rect -465 1565 -450 1585
rect -500 1535 -450 1565
rect -500 1515 -485 1535
rect -465 1515 -450 1535
rect -500 1485 -450 1515
rect -500 1465 -485 1485
rect -465 1465 -450 1485
rect -500 1435 -450 1465
rect -500 1415 -485 1435
rect -465 1415 -450 1435
rect -500 1385 -450 1415
rect -500 1365 -485 1385
rect -465 1365 -450 1385
rect -500 1335 -450 1365
rect -500 1315 -485 1335
rect -465 1315 -450 1335
rect -500 1285 -450 1315
rect -500 1265 -485 1285
rect -465 1265 -450 1285
rect -500 1235 -450 1265
rect -500 1215 -485 1235
rect -465 1215 -450 1235
rect -500 1185 -450 1215
rect -500 1165 -485 1185
rect -465 1165 -450 1185
rect -500 1135 -450 1165
rect -500 1115 -485 1135
rect -465 1115 -450 1135
rect -500 1085 -450 1115
rect -500 1065 -485 1085
rect -465 1065 -450 1085
rect -500 1035 -450 1065
rect -500 1015 -485 1035
rect -465 1015 -450 1035
rect -500 985 -450 1015
rect -500 965 -485 985
rect -465 965 -450 985
rect -500 935 -450 965
rect -500 915 -485 935
rect -465 915 -450 935
rect -500 900 -450 915
rect -350 1585 -300 1600
rect -350 1565 -335 1585
rect -315 1565 -300 1585
rect -350 1535 -300 1565
rect -350 1515 -335 1535
rect -315 1515 -300 1535
rect -350 1485 -300 1515
rect -350 1465 -335 1485
rect -315 1465 -300 1485
rect -350 1435 -300 1465
rect -350 1415 -335 1435
rect -315 1415 -300 1435
rect -350 1385 -300 1415
rect -350 1365 -335 1385
rect -315 1365 -300 1385
rect -350 1335 -300 1365
rect -350 1315 -335 1335
rect -315 1315 -300 1335
rect -350 1285 -300 1315
rect -350 1265 -335 1285
rect -315 1265 -300 1285
rect -350 1235 -300 1265
rect -350 1215 -335 1235
rect -315 1215 -300 1235
rect -350 1185 -300 1215
rect -350 1165 -335 1185
rect -315 1165 -300 1185
rect -350 1135 -300 1165
rect -350 1115 -335 1135
rect -315 1115 -300 1135
rect -350 1085 -300 1115
rect -350 1065 -335 1085
rect -315 1065 -300 1085
rect -350 1035 -300 1065
rect -350 1015 -335 1035
rect -315 1015 -300 1035
rect -350 985 -300 1015
rect -350 965 -335 985
rect -315 965 -300 985
rect -350 935 -300 965
rect -350 915 -335 935
rect -315 915 -300 935
rect -500 840 -450 850
rect -500 810 -490 840
rect -460 810 -450 840
rect -500 800 -450 810
rect -350 840 -300 915
rect -200 1585 -150 1600
rect -200 1565 -185 1585
rect -165 1565 -150 1585
rect -200 1535 -150 1565
rect -200 1515 -185 1535
rect -165 1515 -150 1535
rect -200 1485 -150 1515
rect -200 1465 -185 1485
rect -165 1465 -150 1485
rect -200 1435 -150 1465
rect -200 1415 -185 1435
rect -165 1415 -150 1435
rect -200 1385 -150 1415
rect -200 1365 -185 1385
rect -165 1365 -150 1385
rect -200 1335 -150 1365
rect -200 1315 -185 1335
rect -165 1315 -150 1335
rect -200 1285 -150 1315
rect -200 1265 -185 1285
rect -165 1265 -150 1285
rect -200 1235 -150 1265
rect -200 1215 -185 1235
rect -165 1215 -150 1235
rect -200 1185 -150 1215
rect -200 1165 -185 1185
rect -165 1165 -150 1185
rect -200 1135 -150 1165
rect -200 1115 -185 1135
rect -165 1115 -150 1135
rect -200 1085 -150 1115
rect -200 1065 -185 1085
rect -165 1065 -150 1085
rect -200 1035 -150 1065
rect -200 1015 -185 1035
rect -165 1015 -150 1035
rect -200 985 -150 1015
rect -200 965 -185 985
rect -165 965 -150 985
rect -200 935 -150 965
rect -200 915 -185 935
rect -165 915 -150 935
rect -200 900 -150 915
rect -50 1585 0 1660
rect 8350 1690 8400 1700
rect 8350 1660 8360 1690
rect 8390 1660 8400 1690
rect -50 1565 -35 1585
rect -15 1565 0 1585
rect -50 1540 0 1565
rect -50 1510 -40 1540
rect -10 1510 0 1540
rect -50 1485 0 1510
rect -50 1465 -35 1485
rect -15 1465 0 1485
rect -50 1440 0 1465
rect -50 1410 -40 1440
rect -10 1410 0 1440
rect -50 1385 0 1410
rect -50 1365 -35 1385
rect -15 1365 0 1385
rect -50 1340 0 1365
rect -50 1310 -40 1340
rect -10 1310 0 1340
rect -50 1285 0 1310
rect -50 1265 -35 1285
rect -15 1265 0 1285
rect -50 1240 0 1265
rect -50 1210 -40 1240
rect -10 1210 0 1240
rect -50 1185 0 1210
rect -50 1165 -35 1185
rect -15 1165 0 1185
rect -50 1140 0 1165
rect -50 1110 -40 1140
rect -10 1110 0 1140
rect -50 1085 0 1110
rect -50 1065 -35 1085
rect -15 1065 0 1085
rect -50 1040 0 1065
rect -50 1010 -40 1040
rect -10 1010 0 1040
rect -50 985 0 1010
rect -50 965 -35 985
rect -15 965 0 985
rect -50 940 0 965
rect -50 910 -40 940
rect -10 910 0 940
rect -350 810 -340 840
rect -310 810 -300 840
rect -650 710 -640 740
rect -610 710 -600 740
rect -650 685 -600 710
rect -650 665 -635 685
rect -615 665 -600 685
rect -650 640 -600 665
rect -650 610 -640 640
rect -610 610 -600 640
rect -650 585 -600 610
rect -650 565 -635 585
rect -615 565 -600 585
rect -650 540 -600 565
rect -650 510 -640 540
rect -610 510 -600 540
rect -650 485 -600 510
rect -650 465 -635 485
rect -615 465 -600 485
rect -650 440 -600 465
rect -650 410 -640 440
rect -610 410 -600 440
rect -650 385 -600 410
rect -650 365 -635 385
rect -615 365 -600 385
rect -650 340 -600 365
rect -650 310 -640 340
rect -610 310 -600 340
rect -650 285 -600 310
rect -650 265 -635 285
rect -615 265 -600 285
rect -650 240 -600 265
rect -650 210 -640 240
rect -610 210 -600 240
rect -650 185 -600 210
rect -650 165 -635 185
rect -615 165 -600 185
rect -650 140 -600 165
rect -650 110 -640 140
rect -610 110 -600 140
rect -650 85 -600 110
rect -650 65 -635 85
rect -615 65 -600 85
rect -650 -10 -600 65
rect -500 735 -450 750
rect -500 715 -485 735
rect -465 715 -450 735
rect -500 685 -450 715
rect -500 665 -485 685
rect -465 665 -450 685
rect -500 635 -450 665
rect -500 615 -485 635
rect -465 615 -450 635
rect -500 585 -450 615
rect -500 565 -485 585
rect -465 565 -450 585
rect -500 535 -450 565
rect -500 515 -485 535
rect -465 515 -450 535
rect -500 485 -450 515
rect -500 465 -485 485
rect -465 465 -450 485
rect -500 435 -450 465
rect -500 415 -485 435
rect -465 415 -450 435
rect -500 385 -450 415
rect -500 365 -485 385
rect -465 365 -450 385
rect -500 335 -450 365
rect -500 315 -485 335
rect -465 315 -450 335
rect -500 285 -450 315
rect -500 265 -485 285
rect -465 265 -450 285
rect -500 235 -450 265
rect -500 215 -485 235
rect -465 215 -450 235
rect -500 185 -450 215
rect -500 165 -485 185
rect -465 165 -450 185
rect -500 135 -450 165
rect -500 115 -485 135
rect -465 115 -450 135
rect -500 85 -450 115
rect -500 65 -485 85
rect -465 65 -450 85
rect -500 50 -450 65
rect -350 735 -300 810
rect -200 840 -150 850
rect -200 810 -190 840
rect -160 810 -150 840
rect -200 800 -150 810
rect -350 715 -335 735
rect -315 715 -300 735
rect -350 685 -300 715
rect -350 665 -335 685
rect -315 665 -300 685
rect -350 635 -300 665
rect -350 615 -335 635
rect -315 615 -300 635
rect -350 585 -300 615
rect -350 565 -335 585
rect -315 565 -300 585
rect -350 535 -300 565
rect -350 515 -335 535
rect -315 515 -300 535
rect -350 485 -300 515
rect -350 465 -335 485
rect -315 465 -300 485
rect -350 435 -300 465
rect -350 415 -335 435
rect -315 415 -300 435
rect -350 385 -300 415
rect -350 365 -335 385
rect -315 365 -300 385
rect -350 335 -300 365
rect -350 315 -335 335
rect -315 315 -300 335
rect -350 285 -300 315
rect -350 265 -335 285
rect -315 265 -300 285
rect -350 235 -300 265
rect -350 215 -335 235
rect -315 215 -300 235
rect -350 185 -300 215
rect -350 165 -335 185
rect -315 165 -300 185
rect -350 135 -300 165
rect -350 115 -335 135
rect -315 115 -300 135
rect -350 85 -300 115
rect -350 65 -335 85
rect -315 65 -300 85
rect -350 50 -300 65
rect -200 735 -150 750
rect -200 715 -185 735
rect -165 715 -150 735
rect -200 685 -150 715
rect -200 665 -185 685
rect -165 665 -150 685
rect -200 635 -150 665
rect -200 615 -185 635
rect -165 615 -150 635
rect -200 585 -150 615
rect -200 565 -185 585
rect -165 565 -150 585
rect -200 535 -150 565
rect -200 515 -185 535
rect -165 515 -150 535
rect -200 485 -150 515
rect -200 465 -185 485
rect -165 465 -150 485
rect -200 435 -150 465
rect -200 415 -185 435
rect -165 415 -150 435
rect -200 385 -150 415
rect -200 365 -185 385
rect -165 365 -150 385
rect -200 335 -150 365
rect -200 315 -185 335
rect -165 315 -150 335
rect -200 285 -150 315
rect -200 265 -185 285
rect -165 265 -150 285
rect -200 235 -150 265
rect -200 215 -185 235
rect -165 215 -150 235
rect -200 185 -150 215
rect -200 165 -185 185
rect -165 165 -150 185
rect -200 135 -150 165
rect -200 115 -185 135
rect -165 115 -150 135
rect -200 85 -150 115
rect -200 65 -185 85
rect -165 65 -150 85
rect -200 50 -150 65
rect -50 740 0 910
rect 1150 1585 7200 1600
rect 1150 1565 1165 1585
rect 1185 1565 1765 1585
rect 1785 1565 2365 1585
rect 2385 1565 2965 1585
rect 2985 1565 3565 1585
rect 3585 1565 3865 1585
rect 3885 1565 4165 1585
rect 4185 1565 4465 1585
rect 4485 1565 4765 1585
rect 4785 1565 5365 1585
rect 5385 1565 5965 1585
rect 5985 1565 6565 1585
rect 6585 1565 7165 1585
rect 7185 1565 7200 1585
rect 1150 1550 7200 1565
rect 1150 1535 1200 1550
rect 1150 1515 1165 1535
rect 1185 1515 1200 1535
rect 1150 1485 1200 1515
rect 1750 1535 1800 1550
rect 1750 1515 1765 1535
rect 1785 1515 1800 1535
rect 1150 1465 1165 1485
rect 1185 1465 1200 1485
rect 1150 1435 1200 1465
rect 1150 1415 1165 1435
rect 1185 1415 1200 1435
rect 1150 1385 1200 1415
rect 1150 1365 1165 1385
rect 1185 1365 1200 1385
rect 1150 1335 1200 1365
rect 1150 1315 1165 1335
rect 1185 1315 1200 1335
rect 1150 1285 1200 1315
rect 1150 1265 1165 1285
rect 1185 1265 1200 1285
rect 1150 1235 1200 1265
rect 1150 1215 1165 1235
rect 1185 1215 1200 1235
rect 1150 1185 1200 1215
rect 1150 1165 1165 1185
rect 1185 1165 1200 1185
rect 1150 1135 1200 1165
rect 1150 1115 1165 1135
rect 1185 1115 1200 1135
rect 1150 1085 1200 1115
rect 1150 1065 1165 1085
rect 1185 1065 1200 1085
rect 1150 1035 1200 1065
rect 1150 1015 1165 1035
rect 1185 1015 1200 1035
rect 1150 985 1200 1015
rect 1150 965 1165 985
rect 1185 965 1200 985
rect 1150 935 1200 965
rect 1150 915 1165 935
rect 1185 915 1200 935
rect 1150 900 1200 915
rect 1450 1485 1500 1500
rect 1450 1465 1465 1485
rect 1485 1465 1500 1485
rect 1450 1435 1500 1465
rect 1450 1415 1465 1435
rect 1485 1415 1500 1435
rect 1450 1385 1500 1415
rect 1450 1365 1465 1385
rect 1485 1365 1500 1385
rect 1450 1335 1500 1365
rect 1450 1315 1465 1335
rect 1485 1315 1500 1335
rect 1450 1285 1500 1315
rect 1450 1265 1465 1285
rect 1485 1265 1500 1285
rect 1450 1235 1500 1265
rect 1450 1215 1465 1235
rect 1485 1215 1500 1235
rect 1450 1185 1500 1215
rect 1450 1165 1465 1185
rect 1485 1165 1500 1185
rect 1450 1135 1500 1165
rect 1450 1115 1465 1135
rect 1485 1115 1500 1135
rect 1450 1085 1500 1115
rect 1450 1065 1465 1085
rect 1485 1065 1500 1085
rect 1450 1035 1500 1065
rect 1450 1015 1465 1035
rect 1485 1015 1500 1035
rect 1450 985 1500 1015
rect 1750 1485 1800 1515
rect 2350 1535 2400 1550
rect 2350 1515 2365 1535
rect 2385 1515 2400 1535
rect 1750 1465 1765 1485
rect 1785 1465 1800 1485
rect 1750 1435 1800 1465
rect 1750 1415 1765 1435
rect 1785 1415 1800 1435
rect 1750 1385 1800 1415
rect 1750 1365 1765 1385
rect 1785 1365 1800 1385
rect 1750 1335 1800 1365
rect 1750 1315 1765 1335
rect 1785 1315 1800 1335
rect 1750 1285 1800 1315
rect 1750 1265 1765 1285
rect 1785 1265 1800 1285
rect 1750 1235 1800 1265
rect 1750 1215 1765 1235
rect 1785 1215 1800 1235
rect 1750 1185 1800 1215
rect 1750 1165 1765 1185
rect 1785 1165 1800 1185
rect 1750 1135 1800 1165
rect 1750 1115 1765 1135
rect 1785 1115 1800 1135
rect 1750 1085 1800 1115
rect 1750 1065 1765 1085
rect 1785 1065 1800 1085
rect 1750 1035 1800 1065
rect 1750 1015 1765 1035
rect 1785 1015 1800 1035
rect 1750 1000 1800 1015
rect 2050 1485 2100 1500
rect 2050 1465 2065 1485
rect 2085 1465 2100 1485
rect 2050 1435 2100 1465
rect 2050 1415 2065 1435
rect 2085 1415 2100 1435
rect 2050 1385 2100 1415
rect 2050 1365 2065 1385
rect 2085 1365 2100 1385
rect 2050 1335 2100 1365
rect 2050 1315 2065 1335
rect 2085 1315 2100 1335
rect 2050 1285 2100 1315
rect 2050 1265 2065 1285
rect 2085 1265 2100 1285
rect 2050 1235 2100 1265
rect 2050 1215 2065 1235
rect 2085 1215 2100 1235
rect 2050 1185 2100 1215
rect 2050 1165 2065 1185
rect 2085 1165 2100 1185
rect 2050 1135 2100 1165
rect 2050 1115 2065 1135
rect 2085 1115 2100 1135
rect 2050 1085 2100 1115
rect 2050 1065 2065 1085
rect 2085 1065 2100 1085
rect 2050 1035 2100 1065
rect 2050 1015 2065 1035
rect 2085 1015 2100 1035
rect 1450 965 1465 985
rect 1485 965 1500 985
rect 1450 950 1500 965
rect 2050 985 2100 1015
rect 2350 1485 2400 1515
rect 2950 1535 3000 1550
rect 2950 1515 2965 1535
rect 2985 1515 3000 1535
rect 2350 1465 2365 1485
rect 2385 1465 2400 1485
rect 2350 1435 2400 1465
rect 2350 1415 2365 1435
rect 2385 1415 2400 1435
rect 2350 1385 2400 1415
rect 2350 1365 2365 1385
rect 2385 1365 2400 1385
rect 2350 1335 2400 1365
rect 2350 1315 2365 1335
rect 2385 1315 2400 1335
rect 2350 1285 2400 1315
rect 2350 1265 2365 1285
rect 2385 1265 2400 1285
rect 2350 1235 2400 1265
rect 2350 1215 2365 1235
rect 2385 1215 2400 1235
rect 2350 1185 2400 1215
rect 2350 1165 2365 1185
rect 2385 1165 2400 1185
rect 2350 1135 2400 1165
rect 2350 1115 2365 1135
rect 2385 1115 2400 1135
rect 2350 1085 2400 1115
rect 2350 1065 2365 1085
rect 2385 1065 2400 1085
rect 2350 1035 2400 1065
rect 2350 1015 2365 1035
rect 2385 1015 2400 1035
rect 2350 1000 2400 1015
rect 2650 1485 2700 1500
rect 2650 1465 2665 1485
rect 2685 1465 2700 1485
rect 2650 1435 2700 1465
rect 2650 1415 2665 1435
rect 2685 1415 2700 1435
rect 2650 1385 2700 1415
rect 2650 1365 2665 1385
rect 2685 1365 2700 1385
rect 2650 1335 2700 1365
rect 2650 1315 2665 1335
rect 2685 1315 2700 1335
rect 2650 1285 2700 1315
rect 2650 1265 2665 1285
rect 2685 1265 2700 1285
rect 2650 1235 2700 1265
rect 2650 1215 2665 1235
rect 2685 1215 2700 1235
rect 2650 1185 2700 1215
rect 2650 1165 2665 1185
rect 2685 1165 2700 1185
rect 2650 1135 2700 1165
rect 2650 1115 2665 1135
rect 2685 1115 2700 1135
rect 2650 1085 2700 1115
rect 2650 1065 2665 1085
rect 2685 1065 2700 1085
rect 2650 1035 2700 1065
rect 2650 1015 2665 1035
rect 2685 1015 2700 1035
rect 2050 965 2065 985
rect 2085 965 2100 985
rect 2050 950 2100 965
rect 2650 985 2700 1015
rect 2950 1485 3000 1515
rect 3550 1535 3600 1550
rect 3550 1515 3565 1535
rect 3585 1515 3600 1535
rect 2950 1465 2965 1485
rect 2985 1465 3000 1485
rect 2950 1435 3000 1465
rect 2950 1415 2965 1435
rect 2985 1415 3000 1435
rect 2950 1385 3000 1415
rect 2950 1365 2965 1385
rect 2985 1365 3000 1385
rect 2950 1335 3000 1365
rect 2950 1315 2965 1335
rect 2985 1315 3000 1335
rect 2950 1285 3000 1315
rect 2950 1265 2965 1285
rect 2985 1265 3000 1285
rect 2950 1235 3000 1265
rect 2950 1215 2965 1235
rect 2985 1215 3000 1235
rect 2950 1185 3000 1215
rect 2950 1165 2965 1185
rect 2985 1165 3000 1185
rect 2950 1135 3000 1165
rect 2950 1115 2965 1135
rect 2985 1115 3000 1135
rect 2950 1085 3000 1115
rect 2950 1065 2965 1085
rect 2985 1065 3000 1085
rect 2950 1035 3000 1065
rect 2950 1015 2965 1035
rect 2985 1015 3000 1035
rect 2950 1000 3000 1015
rect 3250 1485 3300 1500
rect 3250 1465 3265 1485
rect 3285 1465 3300 1485
rect 3250 1435 3300 1465
rect 3250 1415 3265 1435
rect 3285 1415 3300 1435
rect 3250 1385 3300 1415
rect 3250 1365 3265 1385
rect 3285 1365 3300 1385
rect 3250 1335 3300 1365
rect 3250 1315 3265 1335
rect 3285 1315 3300 1335
rect 3250 1285 3300 1315
rect 3250 1265 3265 1285
rect 3285 1265 3300 1285
rect 3250 1235 3300 1265
rect 3250 1215 3265 1235
rect 3285 1215 3300 1235
rect 3250 1185 3300 1215
rect 3250 1165 3265 1185
rect 3285 1165 3300 1185
rect 3250 1135 3300 1165
rect 3250 1115 3265 1135
rect 3285 1115 3300 1135
rect 3250 1085 3300 1115
rect 3250 1065 3265 1085
rect 3285 1065 3300 1085
rect 3250 1035 3300 1065
rect 3250 1015 3265 1035
rect 3285 1015 3300 1035
rect 2650 965 2665 985
rect 2685 965 2700 985
rect 2650 950 2700 965
rect 3250 985 3300 1015
rect 3250 965 3265 985
rect 3285 965 3300 985
rect 3250 950 3300 965
rect 1450 935 3300 950
rect 1450 915 1465 935
rect 1485 915 2065 935
rect 2085 915 2665 935
rect 2685 915 3265 935
rect 3285 915 3300 935
rect 1450 900 3300 915
rect 3550 1485 3600 1515
rect 3850 1535 3900 1550
rect 3850 1515 3865 1535
rect 3885 1515 3900 1535
rect 3550 1465 3565 1485
rect 3585 1465 3600 1485
rect 3550 1435 3600 1465
rect 3550 1415 3565 1435
rect 3585 1415 3600 1435
rect 3550 1385 3600 1415
rect 3550 1365 3565 1385
rect 3585 1365 3600 1385
rect 3550 1335 3600 1365
rect 3550 1315 3565 1335
rect 3585 1315 3600 1335
rect 3550 1285 3600 1315
rect 3550 1265 3565 1285
rect 3585 1265 3600 1285
rect 3550 1235 3600 1265
rect 3550 1215 3565 1235
rect 3585 1215 3600 1235
rect 3550 1185 3600 1215
rect 3550 1165 3565 1185
rect 3585 1165 3600 1185
rect 3550 1135 3600 1165
rect 3550 1115 3565 1135
rect 3585 1115 3600 1135
rect 3550 1085 3600 1115
rect 3550 1065 3565 1085
rect 3585 1065 3600 1085
rect 3550 1035 3600 1065
rect 3550 1015 3565 1035
rect 3585 1015 3600 1035
rect 3550 985 3600 1015
rect 3550 965 3565 985
rect 3585 965 3600 985
rect 3550 935 3600 965
rect 3550 915 3565 935
rect 3585 915 3600 935
rect 3550 900 3600 915
rect 3700 1485 3750 1500
rect 3700 1465 3715 1485
rect 3735 1465 3750 1485
rect 3700 1435 3750 1465
rect 3700 1415 3715 1435
rect 3735 1415 3750 1435
rect 3700 1385 3750 1415
rect 3700 1365 3715 1385
rect 3735 1365 3750 1385
rect 3700 1335 3750 1365
rect 3700 1315 3715 1335
rect 3735 1315 3750 1335
rect 3700 1285 3750 1315
rect 3700 1265 3715 1285
rect 3735 1265 3750 1285
rect 3700 1235 3750 1265
rect 3700 1215 3715 1235
rect 3735 1215 3750 1235
rect 3700 1185 3750 1215
rect 3700 1165 3715 1185
rect 3735 1165 3750 1185
rect 3700 1135 3750 1165
rect 3700 1115 3715 1135
rect 3735 1115 3750 1135
rect 3700 1085 3750 1115
rect 3700 1065 3715 1085
rect 3735 1065 3750 1085
rect 3700 1035 3750 1065
rect 3700 1015 3715 1035
rect 3735 1015 3750 1035
rect 3700 985 3750 1015
rect 3850 1485 3900 1515
rect 4150 1535 4200 1550
rect 4150 1515 4165 1535
rect 4185 1515 4200 1535
rect 3850 1465 3865 1485
rect 3885 1465 3900 1485
rect 3850 1435 3900 1465
rect 3850 1415 3865 1435
rect 3885 1415 3900 1435
rect 3850 1385 3900 1415
rect 3850 1365 3865 1385
rect 3885 1365 3900 1385
rect 3850 1335 3900 1365
rect 3850 1315 3865 1335
rect 3885 1315 3900 1335
rect 3850 1285 3900 1315
rect 3850 1265 3865 1285
rect 3885 1265 3900 1285
rect 3850 1235 3900 1265
rect 3850 1215 3865 1235
rect 3885 1215 3900 1235
rect 3850 1185 3900 1215
rect 3850 1165 3865 1185
rect 3885 1165 3900 1185
rect 3850 1135 3900 1165
rect 3850 1115 3865 1135
rect 3885 1115 3900 1135
rect 3850 1085 3900 1115
rect 3850 1065 3865 1085
rect 3885 1065 3900 1085
rect 3850 1035 3900 1065
rect 3850 1015 3865 1035
rect 3885 1015 3900 1035
rect 3850 1000 3900 1015
rect 4000 1485 4050 1500
rect 4000 1465 4015 1485
rect 4035 1465 4050 1485
rect 4000 1435 4050 1465
rect 4000 1415 4015 1435
rect 4035 1415 4050 1435
rect 4000 1385 4050 1415
rect 4000 1365 4015 1385
rect 4035 1365 4050 1385
rect 4000 1335 4050 1365
rect 4000 1315 4015 1335
rect 4035 1315 4050 1335
rect 4000 1285 4050 1315
rect 4000 1265 4015 1285
rect 4035 1265 4050 1285
rect 4000 1235 4050 1265
rect 4000 1215 4015 1235
rect 4035 1215 4050 1235
rect 4000 1185 4050 1215
rect 4000 1165 4015 1185
rect 4035 1165 4050 1185
rect 4000 1135 4050 1165
rect 4000 1115 4015 1135
rect 4035 1115 4050 1135
rect 4000 1085 4050 1115
rect 4000 1065 4015 1085
rect 4035 1065 4050 1085
rect 4000 1035 4050 1065
rect 4000 1015 4015 1035
rect 4035 1015 4050 1035
rect 3700 965 3715 985
rect 3735 965 3750 985
rect 3700 950 3750 965
rect 4000 985 4050 1015
rect 4000 965 4015 985
rect 4035 965 4050 985
rect 4000 950 4050 965
rect 3700 935 4050 950
rect 3700 915 3715 935
rect 3735 915 4015 935
rect 4035 915 4050 935
rect 3700 900 4050 915
rect 4150 1485 4200 1515
rect 4450 1535 4500 1550
rect 4450 1515 4465 1535
rect 4485 1515 4500 1535
rect 4150 1465 4165 1485
rect 4185 1465 4200 1485
rect 4150 1435 4200 1465
rect 4150 1415 4165 1435
rect 4185 1415 4200 1435
rect 4150 1385 4200 1415
rect 4150 1365 4165 1385
rect 4185 1365 4200 1385
rect 4150 1335 4200 1365
rect 4150 1315 4165 1335
rect 4185 1315 4200 1335
rect 4150 1285 4200 1315
rect 4150 1265 4165 1285
rect 4185 1265 4200 1285
rect 4150 1235 4200 1265
rect 4150 1215 4165 1235
rect 4185 1215 4200 1235
rect 4150 1185 4200 1215
rect 4150 1165 4165 1185
rect 4185 1165 4200 1185
rect 4150 1135 4200 1165
rect 4150 1115 4165 1135
rect 4185 1115 4200 1135
rect 4150 1085 4200 1115
rect 4150 1065 4165 1085
rect 4185 1065 4200 1085
rect 4150 1035 4200 1065
rect 4150 1015 4165 1035
rect 4185 1015 4200 1035
rect 4150 985 4200 1015
rect 4150 965 4165 985
rect 4185 965 4200 985
rect 4150 935 4200 965
rect 4150 915 4165 935
rect 4185 915 4200 935
rect 4150 900 4200 915
rect 4300 1485 4350 1500
rect 4300 1465 4315 1485
rect 4335 1465 4350 1485
rect 4300 1435 4350 1465
rect 4300 1415 4315 1435
rect 4335 1415 4350 1435
rect 4300 1385 4350 1415
rect 4300 1365 4315 1385
rect 4335 1365 4350 1385
rect 4300 1335 4350 1365
rect 4300 1315 4315 1335
rect 4335 1315 4350 1335
rect 4300 1285 4350 1315
rect 4300 1265 4315 1285
rect 4335 1265 4350 1285
rect 4300 1235 4350 1265
rect 4300 1215 4315 1235
rect 4335 1215 4350 1235
rect 4300 1185 4350 1215
rect 4300 1165 4315 1185
rect 4335 1165 4350 1185
rect 4300 1135 4350 1165
rect 4300 1115 4315 1135
rect 4335 1115 4350 1135
rect 4300 1085 4350 1115
rect 4300 1065 4315 1085
rect 4335 1065 4350 1085
rect 4300 1035 4350 1065
rect 4300 1015 4315 1035
rect 4335 1015 4350 1035
rect 4300 985 4350 1015
rect 4450 1485 4500 1515
rect 4750 1535 4800 1550
rect 4750 1515 4765 1535
rect 4785 1515 4800 1535
rect 4450 1465 4465 1485
rect 4485 1465 4500 1485
rect 4450 1435 4500 1465
rect 4450 1415 4465 1435
rect 4485 1415 4500 1435
rect 4450 1385 4500 1415
rect 4450 1365 4465 1385
rect 4485 1365 4500 1385
rect 4450 1335 4500 1365
rect 4450 1315 4465 1335
rect 4485 1315 4500 1335
rect 4450 1285 4500 1315
rect 4450 1265 4465 1285
rect 4485 1265 4500 1285
rect 4450 1235 4500 1265
rect 4450 1215 4465 1235
rect 4485 1215 4500 1235
rect 4450 1185 4500 1215
rect 4450 1165 4465 1185
rect 4485 1165 4500 1185
rect 4450 1135 4500 1165
rect 4450 1115 4465 1135
rect 4485 1115 4500 1135
rect 4450 1085 4500 1115
rect 4450 1065 4465 1085
rect 4485 1065 4500 1085
rect 4450 1035 4500 1065
rect 4450 1015 4465 1035
rect 4485 1015 4500 1035
rect 4450 1000 4500 1015
rect 4600 1485 4650 1500
rect 4600 1465 4615 1485
rect 4635 1465 4650 1485
rect 4600 1435 4650 1465
rect 4600 1415 4615 1435
rect 4635 1415 4650 1435
rect 4600 1385 4650 1415
rect 4600 1365 4615 1385
rect 4635 1365 4650 1385
rect 4600 1335 4650 1365
rect 4600 1315 4615 1335
rect 4635 1315 4650 1335
rect 4600 1285 4650 1315
rect 4600 1265 4615 1285
rect 4635 1265 4650 1285
rect 4600 1235 4650 1265
rect 4600 1215 4615 1235
rect 4635 1215 4650 1235
rect 4600 1185 4650 1215
rect 4600 1165 4615 1185
rect 4635 1165 4650 1185
rect 4600 1135 4650 1165
rect 4600 1115 4615 1135
rect 4635 1115 4650 1135
rect 4600 1085 4650 1115
rect 4600 1065 4615 1085
rect 4635 1065 4650 1085
rect 4600 1035 4650 1065
rect 4600 1015 4615 1035
rect 4635 1015 4650 1035
rect 4300 965 4315 985
rect 4335 965 4350 985
rect 4300 950 4350 965
rect 4600 985 4650 1015
rect 4600 965 4615 985
rect 4635 965 4650 985
rect 4600 950 4650 965
rect 4300 935 4650 950
rect 4300 915 4315 935
rect 4335 915 4615 935
rect 4635 915 4650 935
rect 4300 900 4650 915
rect 4750 1485 4800 1515
rect 5350 1535 5400 1550
rect 5350 1515 5365 1535
rect 5385 1515 5400 1535
rect 4750 1465 4765 1485
rect 4785 1465 4800 1485
rect 4750 1435 4800 1465
rect 4750 1415 4765 1435
rect 4785 1415 4800 1435
rect 4750 1385 4800 1415
rect 4750 1365 4765 1385
rect 4785 1365 4800 1385
rect 4750 1335 4800 1365
rect 4750 1315 4765 1335
rect 4785 1315 4800 1335
rect 4750 1285 4800 1315
rect 4750 1265 4765 1285
rect 4785 1265 4800 1285
rect 4750 1235 4800 1265
rect 4750 1215 4765 1235
rect 4785 1215 4800 1235
rect 4750 1185 4800 1215
rect 4750 1165 4765 1185
rect 4785 1165 4800 1185
rect 4750 1135 4800 1165
rect 4750 1115 4765 1135
rect 4785 1115 4800 1135
rect 4750 1085 4800 1115
rect 4750 1065 4765 1085
rect 4785 1065 4800 1085
rect 4750 1035 4800 1065
rect 4750 1015 4765 1035
rect 4785 1015 4800 1035
rect 4750 985 4800 1015
rect 4750 965 4765 985
rect 4785 965 4800 985
rect 4750 935 4800 965
rect 4750 915 4765 935
rect 4785 915 4800 935
rect 4750 900 4800 915
rect 5050 1485 5100 1500
rect 5050 1465 5065 1485
rect 5085 1465 5100 1485
rect 5050 1435 5100 1465
rect 5050 1415 5065 1435
rect 5085 1415 5100 1435
rect 5050 1385 5100 1415
rect 5050 1365 5065 1385
rect 5085 1365 5100 1385
rect 5050 1335 5100 1365
rect 5050 1315 5065 1335
rect 5085 1315 5100 1335
rect 5050 1285 5100 1315
rect 5050 1265 5065 1285
rect 5085 1265 5100 1285
rect 5050 1235 5100 1265
rect 5050 1215 5065 1235
rect 5085 1215 5100 1235
rect 5050 1185 5100 1215
rect 5050 1165 5065 1185
rect 5085 1165 5100 1185
rect 5050 1135 5100 1165
rect 5050 1115 5065 1135
rect 5085 1115 5100 1135
rect 5050 1085 5100 1115
rect 5050 1065 5065 1085
rect 5085 1065 5100 1085
rect 5050 1035 5100 1065
rect 5050 1015 5065 1035
rect 5085 1015 5100 1035
rect 5050 985 5100 1015
rect 5350 1485 5400 1515
rect 5950 1535 6000 1550
rect 5950 1515 5965 1535
rect 5985 1515 6000 1535
rect 5350 1465 5365 1485
rect 5385 1465 5400 1485
rect 5350 1435 5400 1465
rect 5350 1415 5365 1435
rect 5385 1415 5400 1435
rect 5350 1385 5400 1415
rect 5350 1365 5365 1385
rect 5385 1365 5400 1385
rect 5350 1335 5400 1365
rect 5350 1315 5365 1335
rect 5385 1315 5400 1335
rect 5350 1285 5400 1315
rect 5350 1265 5365 1285
rect 5385 1265 5400 1285
rect 5350 1235 5400 1265
rect 5350 1215 5365 1235
rect 5385 1215 5400 1235
rect 5350 1185 5400 1215
rect 5350 1165 5365 1185
rect 5385 1165 5400 1185
rect 5350 1135 5400 1165
rect 5350 1115 5365 1135
rect 5385 1115 5400 1135
rect 5350 1085 5400 1115
rect 5350 1065 5365 1085
rect 5385 1065 5400 1085
rect 5350 1035 5400 1065
rect 5350 1015 5365 1035
rect 5385 1015 5400 1035
rect 5350 1000 5400 1015
rect 5650 1485 5700 1500
rect 5650 1465 5665 1485
rect 5685 1465 5700 1485
rect 5650 1435 5700 1465
rect 5650 1415 5665 1435
rect 5685 1415 5700 1435
rect 5650 1385 5700 1415
rect 5650 1365 5665 1385
rect 5685 1365 5700 1385
rect 5650 1335 5700 1365
rect 5650 1315 5665 1335
rect 5685 1315 5700 1335
rect 5650 1285 5700 1315
rect 5650 1265 5665 1285
rect 5685 1265 5700 1285
rect 5650 1235 5700 1265
rect 5650 1215 5665 1235
rect 5685 1215 5700 1235
rect 5650 1185 5700 1215
rect 5650 1165 5665 1185
rect 5685 1165 5700 1185
rect 5650 1135 5700 1165
rect 5650 1115 5665 1135
rect 5685 1115 5700 1135
rect 5650 1085 5700 1115
rect 5650 1065 5665 1085
rect 5685 1065 5700 1085
rect 5650 1035 5700 1065
rect 5650 1015 5665 1035
rect 5685 1015 5700 1035
rect 5050 965 5065 985
rect 5085 965 5100 985
rect 5050 950 5100 965
rect 5650 985 5700 1015
rect 5950 1485 6000 1515
rect 6550 1535 6600 1550
rect 6550 1515 6565 1535
rect 6585 1515 6600 1535
rect 5950 1465 5965 1485
rect 5985 1465 6000 1485
rect 5950 1435 6000 1465
rect 5950 1415 5965 1435
rect 5985 1415 6000 1435
rect 5950 1385 6000 1415
rect 5950 1365 5965 1385
rect 5985 1365 6000 1385
rect 5950 1335 6000 1365
rect 5950 1315 5965 1335
rect 5985 1315 6000 1335
rect 5950 1285 6000 1315
rect 5950 1265 5965 1285
rect 5985 1265 6000 1285
rect 5950 1235 6000 1265
rect 5950 1215 5965 1235
rect 5985 1215 6000 1235
rect 5950 1185 6000 1215
rect 5950 1165 5965 1185
rect 5985 1165 6000 1185
rect 5950 1135 6000 1165
rect 5950 1115 5965 1135
rect 5985 1115 6000 1135
rect 5950 1085 6000 1115
rect 5950 1065 5965 1085
rect 5985 1065 6000 1085
rect 5950 1035 6000 1065
rect 5950 1015 5965 1035
rect 5985 1015 6000 1035
rect 5950 1000 6000 1015
rect 6250 1485 6300 1500
rect 6250 1465 6265 1485
rect 6285 1465 6300 1485
rect 6250 1435 6300 1465
rect 6250 1415 6265 1435
rect 6285 1415 6300 1435
rect 6250 1385 6300 1415
rect 6250 1365 6265 1385
rect 6285 1365 6300 1385
rect 6250 1335 6300 1365
rect 6250 1315 6265 1335
rect 6285 1315 6300 1335
rect 6250 1285 6300 1315
rect 6250 1265 6265 1285
rect 6285 1265 6300 1285
rect 6250 1235 6300 1265
rect 6250 1215 6265 1235
rect 6285 1215 6300 1235
rect 6250 1185 6300 1215
rect 6250 1165 6265 1185
rect 6285 1165 6300 1185
rect 6250 1135 6300 1165
rect 6250 1115 6265 1135
rect 6285 1115 6300 1135
rect 6250 1085 6300 1115
rect 6250 1065 6265 1085
rect 6285 1065 6300 1085
rect 6250 1035 6300 1065
rect 6250 1015 6265 1035
rect 6285 1015 6300 1035
rect 5650 965 5665 985
rect 5685 965 5700 985
rect 5650 950 5700 965
rect 6250 985 6300 1015
rect 6550 1485 6600 1515
rect 7150 1535 7200 1550
rect 7150 1515 7165 1535
rect 7185 1515 7200 1535
rect 6550 1465 6565 1485
rect 6585 1465 6600 1485
rect 6550 1435 6600 1465
rect 6550 1415 6565 1435
rect 6585 1415 6600 1435
rect 6550 1385 6600 1415
rect 6550 1365 6565 1385
rect 6585 1365 6600 1385
rect 6550 1335 6600 1365
rect 6550 1315 6565 1335
rect 6585 1315 6600 1335
rect 6550 1285 6600 1315
rect 6550 1265 6565 1285
rect 6585 1265 6600 1285
rect 6550 1235 6600 1265
rect 6550 1215 6565 1235
rect 6585 1215 6600 1235
rect 6550 1185 6600 1215
rect 6550 1165 6565 1185
rect 6585 1165 6600 1185
rect 6550 1135 6600 1165
rect 6550 1115 6565 1135
rect 6585 1115 6600 1135
rect 6550 1085 6600 1115
rect 6550 1065 6565 1085
rect 6585 1065 6600 1085
rect 6550 1035 6600 1065
rect 6550 1015 6565 1035
rect 6585 1015 6600 1035
rect 6550 1000 6600 1015
rect 6850 1485 6900 1500
rect 6850 1465 6865 1485
rect 6885 1465 6900 1485
rect 6850 1435 6900 1465
rect 6850 1415 6865 1435
rect 6885 1415 6900 1435
rect 6850 1385 6900 1415
rect 6850 1365 6865 1385
rect 6885 1365 6900 1385
rect 6850 1335 6900 1365
rect 6850 1315 6865 1335
rect 6885 1315 6900 1335
rect 6850 1285 6900 1315
rect 6850 1265 6865 1285
rect 6885 1265 6900 1285
rect 6850 1235 6900 1265
rect 6850 1215 6865 1235
rect 6885 1215 6900 1235
rect 6850 1185 6900 1215
rect 6850 1165 6865 1185
rect 6885 1165 6900 1185
rect 6850 1135 6900 1165
rect 6850 1115 6865 1135
rect 6885 1115 6900 1135
rect 6850 1085 6900 1115
rect 6850 1065 6865 1085
rect 6885 1065 6900 1085
rect 6850 1035 6900 1065
rect 6850 1015 6865 1035
rect 6885 1015 6900 1035
rect 6250 965 6265 985
rect 6285 965 6300 985
rect 6250 950 6300 965
rect 6850 985 6900 1015
rect 6850 965 6865 985
rect 6885 965 6900 985
rect 6850 950 6900 965
rect 5050 935 6900 950
rect 5050 915 5065 935
rect 5085 915 5665 935
rect 5685 915 6265 935
rect 6285 915 6865 935
rect 6885 915 6900 935
rect 5050 900 6900 915
rect 7150 1485 7200 1515
rect 7150 1465 7165 1485
rect 7185 1465 7200 1485
rect 7150 1435 7200 1465
rect 7150 1415 7165 1435
rect 7185 1415 7200 1435
rect 7150 1385 7200 1415
rect 7150 1365 7165 1385
rect 7185 1365 7200 1385
rect 7150 1335 7200 1365
rect 7150 1315 7165 1335
rect 7185 1315 7200 1335
rect 7150 1285 7200 1315
rect 7150 1265 7165 1285
rect 7185 1265 7200 1285
rect 7150 1235 7200 1265
rect 7150 1215 7165 1235
rect 7185 1215 7200 1235
rect 7150 1185 7200 1215
rect 7150 1165 7165 1185
rect 7185 1165 7200 1185
rect 7150 1135 7200 1165
rect 7150 1115 7165 1135
rect 7185 1115 7200 1135
rect 7150 1085 7200 1115
rect 7150 1065 7165 1085
rect 7185 1065 7200 1085
rect 7150 1035 7200 1065
rect 7150 1015 7165 1035
rect 7185 1015 7200 1035
rect 7150 985 7200 1015
rect 7150 965 7165 985
rect 7185 965 7200 985
rect 7150 935 7200 965
rect 7150 915 7165 935
rect 7185 915 7200 935
rect 7150 900 7200 915
rect 8350 1585 8400 1660
rect 10750 1690 10800 1700
rect 10750 1660 10760 1690
rect 10790 1660 10800 1690
rect 8350 1565 8365 1585
rect 8385 1565 8400 1585
rect 8350 1540 8400 1565
rect 8350 1510 8360 1540
rect 8390 1510 8400 1540
rect 8350 1485 8400 1510
rect 8350 1465 8365 1485
rect 8385 1465 8400 1485
rect 8350 1440 8400 1465
rect 8350 1410 8360 1440
rect 8390 1410 8400 1440
rect 8350 1385 8400 1410
rect 8350 1365 8365 1385
rect 8385 1365 8400 1385
rect 8350 1340 8400 1365
rect 8350 1310 8360 1340
rect 8390 1310 8400 1340
rect 8350 1285 8400 1310
rect 8350 1265 8365 1285
rect 8385 1265 8400 1285
rect 8350 1240 8400 1265
rect 8350 1210 8360 1240
rect 8390 1210 8400 1240
rect 8350 1185 8400 1210
rect 8350 1165 8365 1185
rect 8385 1165 8400 1185
rect 8350 1140 8400 1165
rect 8350 1110 8360 1140
rect 8390 1110 8400 1140
rect 8350 1085 8400 1110
rect 8350 1065 8365 1085
rect 8385 1065 8400 1085
rect 8350 1040 8400 1065
rect 8350 1010 8360 1040
rect 8390 1010 8400 1040
rect 8350 985 8400 1010
rect 8350 965 8365 985
rect 8385 965 8400 985
rect 8350 940 8400 965
rect 8350 910 8360 940
rect 8390 910 8400 940
rect 100 840 150 850
rect 100 810 110 840
rect 140 810 150 840
rect 100 800 150 810
rect 400 840 450 850
rect 400 810 410 840
rect 440 810 450 840
rect 400 800 450 810
rect 700 840 750 850
rect 700 810 710 840
rect 740 810 750 840
rect 700 800 750 810
rect 1000 840 1050 850
rect 1000 810 1010 840
rect 1040 810 1050 840
rect 1000 800 1050 810
rect 1300 840 1350 850
rect 1300 810 1310 840
rect 1340 810 1350 840
rect 1300 800 1350 810
rect 1600 840 1650 850
rect 1600 810 1610 840
rect 1640 810 1650 840
rect 1600 800 1650 810
rect 1900 840 1950 850
rect 1900 810 1910 840
rect 1940 810 1950 840
rect 1900 800 1950 810
rect 2200 840 2250 850
rect 2200 810 2210 840
rect 2240 810 2250 840
rect 2200 800 2250 810
rect 2350 840 2400 900
rect 2350 810 2360 840
rect 2390 810 2400 840
rect 2350 750 2400 810
rect 2500 840 2550 850
rect 2500 810 2510 840
rect 2540 810 2550 840
rect 2500 800 2550 810
rect 2800 840 2850 850
rect 2800 810 2810 840
rect 2840 810 2850 840
rect 2800 800 2850 810
rect 3100 840 3150 850
rect 3100 810 3110 840
rect 3140 810 3150 840
rect 3100 800 3150 810
rect 3400 840 3450 850
rect 3400 810 3410 840
rect 3440 810 3450 840
rect 3400 800 3450 810
rect 3700 840 3750 850
rect 3700 810 3710 840
rect 3740 810 3750 840
rect 3700 800 3750 810
rect 3850 840 3900 900
rect 3850 810 3860 840
rect 3890 810 3900 840
rect 3850 750 3900 810
rect 4000 840 4050 850
rect 4000 810 4010 840
rect 4040 810 4050 840
rect 4000 800 4050 810
rect 4300 840 4350 850
rect 4300 810 4310 840
rect 4340 810 4350 840
rect 4300 800 4350 810
rect 4450 840 4500 900
rect 4450 810 4460 840
rect 4490 810 4500 840
rect 4450 750 4500 810
rect 4600 840 4650 850
rect 4600 810 4610 840
rect 4640 810 4650 840
rect 4600 800 4650 810
rect 4900 840 4950 850
rect 4900 810 4910 840
rect 4940 810 4950 840
rect 4900 800 4950 810
rect 5200 840 5250 850
rect 5200 810 5210 840
rect 5240 810 5250 840
rect 5200 800 5250 810
rect 5500 840 5550 850
rect 5500 810 5510 840
rect 5540 810 5550 840
rect 5500 800 5550 810
rect 5800 840 5850 850
rect 5800 810 5810 840
rect 5840 810 5850 840
rect 5800 800 5850 810
rect 5950 840 6000 900
rect 5950 810 5960 840
rect 5990 810 6000 840
rect 5950 750 6000 810
rect 6100 840 6150 850
rect 6100 810 6110 840
rect 6140 810 6150 840
rect 6100 800 6150 810
rect 6400 840 6450 850
rect 6400 810 6410 840
rect 6440 810 6450 840
rect 6400 800 6450 810
rect 6700 840 6750 850
rect 6700 810 6710 840
rect 6740 810 6750 840
rect 6700 800 6750 810
rect 7000 840 7050 850
rect 7000 810 7010 840
rect 7040 810 7050 840
rect 7000 800 7050 810
rect 7300 840 7350 850
rect 7300 810 7310 840
rect 7340 810 7350 840
rect 7300 800 7350 810
rect 7600 840 7650 850
rect 7600 810 7610 840
rect 7640 810 7650 840
rect 7600 800 7650 810
rect 7900 840 7950 850
rect 7900 810 7910 840
rect 7940 810 7950 840
rect 7900 800 7950 810
rect 8200 840 8250 850
rect 8200 810 8210 840
rect 8240 810 8250 840
rect 8200 800 8250 810
rect -50 710 -40 740
rect -10 710 0 740
rect -50 685 0 710
rect -50 665 -35 685
rect -15 665 0 685
rect -50 640 0 665
rect -50 610 -40 640
rect -10 610 0 640
rect -50 585 0 610
rect -50 565 -35 585
rect -15 565 0 585
rect -50 540 0 565
rect -50 510 -40 540
rect -10 510 0 540
rect -50 485 0 510
rect -50 465 -35 485
rect -15 465 0 485
rect -50 440 0 465
rect -50 410 -40 440
rect -10 410 0 440
rect -50 385 0 410
rect -50 365 -35 385
rect -15 365 0 385
rect -50 340 0 365
rect -50 310 -40 340
rect -10 310 0 340
rect -50 285 0 310
rect -50 265 -35 285
rect -15 265 0 285
rect -50 240 0 265
rect -50 210 -40 240
rect -10 210 0 240
rect -50 185 0 210
rect -50 165 -35 185
rect -15 165 0 185
rect -50 140 0 165
rect -50 110 -40 140
rect -10 110 0 140
rect -50 85 0 110
rect -50 65 -35 85
rect -15 65 0 85
rect -650 -40 -640 -10
rect -610 -40 -600 -10
rect -650 -115 -600 -40
rect -50 -10 0 65
rect 1150 735 1200 750
rect 1150 715 1165 735
rect 1185 715 1200 735
rect 1150 685 1200 715
rect 1150 665 1165 685
rect 1185 665 1200 685
rect 1150 635 1200 665
rect 1150 615 1165 635
rect 1185 615 1200 635
rect 1150 585 1200 615
rect 1150 565 1165 585
rect 1185 565 1200 585
rect 1150 535 1200 565
rect 1150 515 1165 535
rect 1185 515 1200 535
rect 1150 485 1200 515
rect 1150 465 1165 485
rect 1185 465 1200 485
rect 1150 435 1200 465
rect 1150 415 1165 435
rect 1185 415 1200 435
rect 1150 385 1200 415
rect 1150 365 1165 385
rect 1185 365 1200 385
rect 1150 335 1200 365
rect 1150 315 1165 335
rect 1185 315 1200 335
rect 1150 285 1200 315
rect 1150 265 1165 285
rect 1185 265 1200 285
rect 1150 235 1200 265
rect 1150 215 1165 235
rect 1185 215 1200 235
rect 1150 185 1200 215
rect 1150 165 1165 185
rect 1185 165 1200 185
rect 1150 135 1200 165
rect 1450 735 3300 750
rect 1450 715 1465 735
rect 1485 715 2065 735
rect 2085 715 2665 735
rect 2685 715 3265 735
rect 3285 715 3300 735
rect 1450 700 3300 715
rect 1450 685 1500 700
rect 1450 665 1465 685
rect 1485 665 1500 685
rect 1450 635 1500 665
rect 2050 685 2100 700
rect 2050 665 2065 685
rect 2085 665 2100 685
rect 1450 615 1465 635
rect 1485 615 1500 635
rect 1450 585 1500 615
rect 1450 565 1465 585
rect 1485 565 1500 585
rect 1450 535 1500 565
rect 1450 515 1465 535
rect 1485 515 1500 535
rect 1450 485 1500 515
rect 1450 465 1465 485
rect 1485 465 1500 485
rect 1450 435 1500 465
rect 1450 415 1465 435
rect 1485 415 1500 435
rect 1450 385 1500 415
rect 1450 365 1465 385
rect 1485 365 1500 385
rect 1450 335 1500 365
rect 1450 315 1465 335
rect 1485 315 1500 335
rect 1450 285 1500 315
rect 1450 265 1465 285
rect 1485 265 1500 285
rect 1450 235 1500 265
rect 1450 215 1465 235
rect 1485 215 1500 235
rect 1450 185 1500 215
rect 1450 165 1465 185
rect 1485 165 1500 185
rect 1450 150 1500 165
rect 1750 635 1800 650
rect 1750 615 1765 635
rect 1785 615 1800 635
rect 1750 585 1800 615
rect 1750 565 1765 585
rect 1785 565 1800 585
rect 1750 535 1800 565
rect 1750 515 1765 535
rect 1785 515 1800 535
rect 1750 485 1800 515
rect 1750 465 1765 485
rect 1785 465 1800 485
rect 1750 435 1800 465
rect 1750 415 1765 435
rect 1785 415 1800 435
rect 1750 385 1800 415
rect 1750 365 1765 385
rect 1785 365 1800 385
rect 1750 335 1800 365
rect 1750 315 1765 335
rect 1785 315 1800 335
rect 1750 285 1800 315
rect 1750 265 1765 285
rect 1785 265 1800 285
rect 1750 235 1800 265
rect 1750 215 1765 235
rect 1785 215 1800 235
rect 1750 185 1800 215
rect 1750 165 1765 185
rect 1785 165 1800 185
rect 1150 115 1165 135
rect 1185 115 1200 135
rect 1150 100 1200 115
rect 1750 135 1800 165
rect 2050 635 2100 665
rect 2650 685 2700 700
rect 2650 665 2665 685
rect 2685 665 2700 685
rect 2050 615 2065 635
rect 2085 615 2100 635
rect 2050 585 2100 615
rect 2050 565 2065 585
rect 2085 565 2100 585
rect 2050 535 2100 565
rect 2050 515 2065 535
rect 2085 515 2100 535
rect 2050 485 2100 515
rect 2050 465 2065 485
rect 2085 465 2100 485
rect 2050 435 2100 465
rect 2050 415 2065 435
rect 2085 415 2100 435
rect 2050 385 2100 415
rect 2050 365 2065 385
rect 2085 365 2100 385
rect 2050 335 2100 365
rect 2050 315 2065 335
rect 2085 315 2100 335
rect 2050 285 2100 315
rect 2050 265 2065 285
rect 2085 265 2100 285
rect 2050 235 2100 265
rect 2050 215 2065 235
rect 2085 215 2100 235
rect 2050 185 2100 215
rect 2050 165 2065 185
rect 2085 165 2100 185
rect 2050 150 2100 165
rect 2350 635 2400 650
rect 2350 615 2365 635
rect 2385 615 2400 635
rect 2350 585 2400 615
rect 2350 565 2365 585
rect 2385 565 2400 585
rect 2350 535 2400 565
rect 2350 515 2365 535
rect 2385 515 2400 535
rect 2350 485 2400 515
rect 2350 465 2365 485
rect 2385 465 2400 485
rect 2350 435 2400 465
rect 2350 415 2365 435
rect 2385 415 2400 435
rect 2350 385 2400 415
rect 2350 365 2365 385
rect 2385 365 2400 385
rect 2350 335 2400 365
rect 2350 315 2365 335
rect 2385 315 2400 335
rect 2350 285 2400 315
rect 2350 265 2365 285
rect 2385 265 2400 285
rect 2350 235 2400 265
rect 2350 215 2365 235
rect 2385 215 2400 235
rect 2350 185 2400 215
rect 2350 165 2365 185
rect 2385 165 2400 185
rect 1750 115 1765 135
rect 1785 115 1800 135
rect 1750 100 1800 115
rect 2350 135 2400 165
rect 2650 635 2700 665
rect 3250 685 3300 700
rect 3250 665 3265 685
rect 3285 665 3300 685
rect 2650 615 2665 635
rect 2685 615 2700 635
rect 2650 585 2700 615
rect 2650 565 2665 585
rect 2685 565 2700 585
rect 2650 535 2700 565
rect 2650 515 2665 535
rect 2685 515 2700 535
rect 2650 485 2700 515
rect 2650 465 2665 485
rect 2685 465 2700 485
rect 2650 435 2700 465
rect 2650 415 2665 435
rect 2685 415 2700 435
rect 2650 385 2700 415
rect 2650 365 2665 385
rect 2685 365 2700 385
rect 2650 335 2700 365
rect 2650 315 2665 335
rect 2685 315 2700 335
rect 2650 285 2700 315
rect 2650 265 2665 285
rect 2685 265 2700 285
rect 2650 235 2700 265
rect 2650 215 2665 235
rect 2685 215 2700 235
rect 2650 185 2700 215
rect 2650 165 2665 185
rect 2685 165 2700 185
rect 2650 150 2700 165
rect 2950 635 3000 650
rect 2950 615 2965 635
rect 2985 615 3000 635
rect 2950 585 3000 615
rect 2950 565 2965 585
rect 2985 565 3000 585
rect 2950 535 3000 565
rect 2950 515 2965 535
rect 2985 515 3000 535
rect 2950 485 3000 515
rect 2950 465 2965 485
rect 2985 465 3000 485
rect 2950 435 3000 465
rect 2950 415 2965 435
rect 2985 415 3000 435
rect 2950 385 3000 415
rect 2950 365 2965 385
rect 2985 365 3000 385
rect 2950 335 3000 365
rect 2950 315 2965 335
rect 2985 315 3000 335
rect 2950 285 3000 315
rect 2950 265 2965 285
rect 2985 265 3000 285
rect 2950 235 3000 265
rect 2950 215 2965 235
rect 2985 215 3000 235
rect 2950 185 3000 215
rect 2950 165 2965 185
rect 2985 165 3000 185
rect 2350 115 2365 135
rect 2385 115 2400 135
rect 2350 100 2400 115
rect 2950 135 3000 165
rect 3250 635 3300 665
rect 3250 615 3265 635
rect 3285 615 3300 635
rect 3250 585 3300 615
rect 3250 565 3265 585
rect 3285 565 3300 585
rect 3250 535 3300 565
rect 3250 515 3265 535
rect 3285 515 3300 535
rect 3250 485 3300 515
rect 3250 465 3265 485
rect 3285 465 3300 485
rect 3250 435 3300 465
rect 3250 415 3265 435
rect 3285 415 3300 435
rect 3250 385 3300 415
rect 3250 365 3265 385
rect 3285 365 3300 385
rect 3250 335 3300 365
rect 3250 315 3265 335
rect 3285 315 3300 335
rect 3250 285 3300 315
rect 3250 265 3265 285
rect 3285 265 3300 285
rect 3250 235 3300 265
rect 3250 215 3265 235
rect 3285 215 3300 235
rect 3250 185 3300 215
rect 3250 165 3265 185
rect 3285 165 3300 185
rect 3250 150 3300 165
rect 3550 735 3600 750
rect 3550 715 3565 735
rect 3585 715 3600 735
rect 3550 685 3600 715
rect 3550 665 3565 685
rect 3585 665 3600 685
rect 3550 635 3600 665
rect 3550 615 3565 635
rect 3585 615 3600 635
rect 3550 585 3600 615
rect 3550 565 3565 585
rect 3585 565 3600 585
rect 3550 535 3600 565
rect 3550 515 3565 535
rect 3585 515 3600 535
rect 3550 485 3600 515
rect 3550 465 3565 485
rect 3585 465 3600 485
rect 3550 435 3600 465
rect 3550 415 3565 435
rect 3585 415 3600 435
rect 3550 385 3600 415
rect 3550 365 3565 385
rect 3585 365 3600 385
rect 3550 335 3600 365
rect 3550 315 3565 335
rect 3585 315 3600 335
rect 3550 285 3600 315
rect 3550 265 3565 285
rect 3585 265 3600 285
rect 3550 235 3600 265
rect 3550 215 3565 235
rect 3585 215 3600 235
rect 3550 185 3600 215
rect 3550 165 3565 185
rect 3585 165 3600 185
rect 2950 115 2965 135
rect 2985 115 3000 135
rect 2950 100 3000 115
rect 3550 135 3600 165
rect 3700 735 4050 750
rect 3700 715 3715 735
rect 3735 715 4015 735
rect 4035 715 4050 735
rect 3700 700 4050 715
rect 3700 685 3750 700
rect 3700 665 3715 685
rect 3735 665 3750 685
rect 3700 635 3750 665
rect 4000 685 4050 700
rect 4000 665 4015 685
rect 4035 665 4050 685
rect 3700 615 3715 635
rect 3735 615 3750 635
rect 3700 585 3750 615
rect 3700 565 3715 585
rect 3735 565 3750 585
rect 3700 535 3750 565
rect 3700 515 3715 535
rect 3735 515 3750 535
rect 3700 485 3750 515
rect 3700 465 3715 485
rect 3735 465 3750 485
rect 3700 435 3750 465
rect 3700 415 3715 435
rect 3735 415 3750 435
rect 3700 385 3750 415
rect 3700 365 3715 385
rect 3735 365 3750 385
rect 3700 335 3750 365
rect 3700 315 3715 335
rect 3735 315 3750 335
rect 3700 285 3750 315
rect 3700 265 3715 285
rect 3735 265 3750 285
rect 3700 235 3750 265
rect 3700 215 3715 235
rect 3735 215 3750 235
rect 3700 185 3750 215
rect 3700 165 3715 185
rect 3735 165 3750 185
rect 3700 150 3750 165
rect 3850 635 3900 650
rect 3850 615 3865 635
rect 3885 615 3900 635
rect 3850 585 3900 615
rect 3850 565 3865 585
rect 3885 565 3900 585
rect 3850 535 3900 565
rect 3850 515 3865 535
rect 3885 515 3900 535
rect 3850 485 3900 515
rect 3850 465 3865 485
rect 3885 465 3900 485
rect 3850 435 3900 465
rect 3850 415 3865 435
rect 3885 415 3900 435
rect 3850 385 3900 415
rect 3850 365 3865 385
rect 3885 365 3900 385
rect 3850 335 3900 365
rect 3850 315 3865 335
rect 3885 315 3900 335
rect 3850 285 3900 315
rect 3850 265 3865 285
rect 3885 265 3900 285
rect 3850 235 3900 265
rect 3850 215 3865 235
rect 3885 215 3900 235
rect 3850 185 3900 215
rect 3850 165 3865 185
rect 3885 165 3900 185
rect 3550 115 3565 135
rect 3585 115 3600 135
rect 3550 100 3600 115
rect 3850 135 3900 165
rect 4000 635 4050 665
rect 4000 615 4015 635
rect 4035 615 4050 635
rect 4000 585 4050 615
rect 4000 565 4015 585
rect 4035 565 4050 585
rect 4000 535 4050 565
rect 4000 515 4015 535
rect 4035 515 4050 535
rect 4000 485 4050 515
rect 4000 465 4015 485
rect 4035 465 4050 485
rect 4000 435 4050 465
rect 4000 415 4015 435
rect 4035 415 4050 435
rect 4000 385 4050 415
rect 4000 365 4015 385
rect 4035 365 4050 385
rect 4000 335 4050 365
rect 4000 315 4015 335
rect 4035 315 4050 335
rect 4000 285 4050 315
rect 4000 265 4015 285
rect 4035 265 4050 285
rect 4000 235 4050 265
rect 4000 215 4015 235
rect 4035 215 4050 235
rect 4000 185 4050 215
rect 4000 165 4015 185
rect 4035 165 4050 185
rect 4000 150 4050 165
rect 4150 735 4200 750
rect 4150 715 4165 735
rect 4185 715 4200 735
rect 4150 685 4200 715
rect 4150 665 4165 685
rect 4185 665 4200 685
rect 4150 635 4200 665
rect 4150 615 4165 635
rect 4185 615 4200 635
rect 4150 585 4200 615
rect 4150 565 4165 585
rect 4185 565 4200 585
rect 4150 535 4200 565
rect 4150 515 4165 535
rect 4185 515 4200 535
rect 4150 485 4200 515
rect 4150 465 4165 485
rect 4185 465 4200 485
rect 4150 435 4200 465
rect 4150 415 4165 435
rect 4185 415 4200 435
rect 4150 385 4200 415
rect 4150 365 4165 385
rect 4185 365 4200 385
rect 4150 335 4200 365
rect 4150 315 4165 335
rect 4185 315 4200 335
rect 4150 285 4200 315
rect 4150 265 4165 285
rect 4185 265 4200 285
rect 4150 235 4200 265
rect 4150 215 4165 235
rect 4185 215 4200 235
rect 4150 185 4200 215
rect 4150 165 4165 185
rect 4185 165 4200 185
rect 3850 115 3865 135
rect 3885 115 3900 135
rect 3850 100 3900 115
rect 4150 135 4200 165
rect 4300 735 4650 750
rect 4300 715 4315 735
rect 4335 715 4615 735
rect 4635 715 4650 735
rect 4300 700 4650 715
rect 4300 685 4350 700
rect 4300 665 4315 685
rect 4335 665 4350 685
rect 4300 635 4350 665
rect 4600 685 4650 700
rect 4600 665 4615 685
rect 4635 665 4650 685
rect 4300 615 4315 635
rect 4335 615 4350 635
rect 4300 585 4350 615
rect 4300 565 4315 585
rect 4335 565 4350 585
rect 4300 535 4350 565
rect 4300 515 4315 535
rect 4335 515 4350 535
rect 4300 485 4350 515
rect 4300 465 4315 485
rect 4335 465 4350 485
rect 4300 435 4350 465
rect 4300 415 4315 435
rect 4335 415 4350 435
rect 4300 385 4350 415
rect 4300 365 4315 385
rect 4335 365 4350 385
rect 4300 335 4350 365
rect 4300 315 4315 335
rect 4335 315 4350 335
rect 4300 285 4350 315
rect 4300 265 4315 285
rect 4335 265 4350 285
rect 4300 235 4350 265
rect 4300 215 4315 235
rect 4335 215 4350 235
rect 4300 185 4350 215
rect 4300 165 4315 185
rect 4335 165 4350 185
rect 4300 150 4350 165
rect 4450 635 4500 650
rect 4450 615 4465 635
rect 4485 615 4500 635
rect 4450 585 4500 615
rect 4450 565 4465 585
rect 4485 565 4500 585
rect 4450 535 4500 565
rect 4450 515 4465 535
rect 4485 515 4500 535
rect 4450 485 4500 515
rect 4450 465 4465 485
rect 4485 465 4500 485
rect 4450 435 4500 465
rect 4450 415 4465 435
rect 4485 415 4500 435
rect 4450 385 4500 415
rect 4450 365 4465 385
rect 4485 365 4500 385
rect 4450 335 4500 365
rect 4450 315 4465 335
rect 4485 315 4500 335
rect 4450 285 4500 315
rect 4450 265 4465 285
rect 4485 265 4500 285
rect 4450 235 4500 265
rect 4450 215 4465 235
rect 4485 215 4500 235
rect 4450 185 4500 215
rect 4450 165 4465 185
rect 4485 165 4500 185
rect 4150 115 4165 135
rect 4185 115 4200 135
rect 4150 100 4200 115
rect 4450 135 4500 165
rect 4600 635 4650 665
rect 4600 615 4615 635
rect 4635 615 4650 635
rect 4600 585 4650 615
rect 4600 565 4615 585
rect 4635 565 4650 585
rect 4600 535 4650 565
rect 4600 515 4615 535
rect 4635 515 4650 535
rect 4600 485 4650 515
rect 4600 465 4615 485
rect 4635 465 4650 485
rect 4600 435 4650 465
rect 4600 415 4615 435
rect 4635 415 4650 435
rect 4600 385 4650 415
rect 4600 365 4615 385
rect 4635 365 4650 385
rect 4600 335 4650 365
rect 4600 315 4615 335
rect 4635 315 4650 335
rect 4600 285 4650 315
rect 4600 265 4615 285
rect 4635 265 4650 285
rect 4600 235 4650 265
rect 4600 215 4615 235
rect 4635 215 4650 235
rect 4600 185 4650 215
rect 4600 165 4615 185
rect 4635 165 4650 185
rect 4600 150 4650 165
rect 4750 735 4800 750
rect 4750 715 4765 735
rect 4785 715 4800 735
rect 4750 685 4800 715
rect 4750 665 4765 685
rect 4785 665 4800 685
rect 4750 635 4800 665
rect 4750 615 4765 635
rect 4785 615 4800 635
rect 4750 585 4800 615
rect 4750 565 4765 585
rect 4785 565 4800 585
rect 4750 535 4800 565
rect 4750 515 4765 535
rect 4785 515 4800 535
rect 4750 485 4800 515
rect 4750 465 4765 485
rect 4785 465 4800 485
rect 4750 435 4800 465
rect 4750 415 4765 435
rect 4785 415 4800 435
rect 4750 385 4800 415
rect 4750 365 4765 385
rect 4785 365 4800 385
rect 4750 335 4800 365
rect 4750 315 4765 335
rect 4785 315 4800 335
rect 4750 285 4800 315
rect 4750 265 4765 285
rect 4785 265 4800 285
rect 4750 235 4800 265
rect 4750 215 4765 235
rect 4785 215 4800 235
rect 4750 185 4800 215
rect 4750 165 4765 185
rect 4785 165 4800 185
rect 4450 115 4465 135
rect 4485 115 4500 135
rect 4450 100 4500 115
rect 4750 135 4800 165
rect 5050 735 6900 750
rect 5050 715 5065 735
rect 5085 715 5665 735
rect 5685 715 6265 735
rect 6285 715 6865 735
rect 6885 715 6900 735
rect 5050 700 6900 715
rect 5050 685 5100 700
rect 5050 665 5065 685
rect 5085 665 5100 685
rect 5050 635 5100 665
rect 5650 685 5700 700
rect 5650 665 5665 685
rect 5685 665 5700 685
rect 5050 615 5065 635
rect 5085 615 5100 635
rect 5050 585 5100 615
rect 5050 565 5065 585
rect 5085 565 5100 585
rect 5050 535 5100 565
rect 5050 515 5065 535
rect 5085 515 5100 535
rect 5050 485 5100 515
rect 5050 465 5065 485
rect 5085 465 5100 485
rect 5050 435 5100 465
rect 5050 415 5065 435
rect 5085 415 5100 435
rect 5050 385 5100 415
rect 5050 365 5065 385
rect 5085 365 5100 385
rect 5050 335 5100 365
rect 5050 315 5065 335
rect 5085 315 5100 335
rect 5050 285 5100 315
rect 5050 265 5065 285
rect 5085 265 5100 285
rect 5050 235 5100 265
rect 5050 215 5065 235
rect 5085 215 5100 235
rect 5050 185 5100 215
rect 5050 165 5065 185
rect 5085 165 5100 185
rect 5050 150 5100 165
rect 5350 635 5400 650
rect 5350 615 5365 635
rect 5385 615 5400 635
rect 5350 585 5400 615
rect 5350 565 5365 585
rect 5385 565 5400 585
rect 5350 535 5400 565
rect 5350 515 5365 535
rect 5385 515 5400 535
rect 5350 485 5400 515
rect 5350 465 5365 485
rect 5385 465 5400 485
rect 5350 435 5400 465
rect 5350 415 5365 435
rect 5385 415 5400 435
rect 5350 385 5400 415
rect 5350 365 5365 385
rect 5385 365 5400 385
rect 5350 335 5400 365
rect 5350 315 5365 335
rect 5385 315 5400 335
rect 5350 285 5400 315
rect 5350 265 5365 285
rect 5385 265 5400 285
rect 5350 235 5400 265
rect 5350 215 5365 235
rect 5385 215 5400 235
rect 5350 185 5400 215
rect 5350 165 5365 185
rect 5385 165 5400 185
rect 4750 115 4765 135
rect 4785 115 4800 135
rect 4750 100 4800 115
rect 5350 135 5400 165
rect 5650 635 5700 665
rect 6250 685 6300 700
rect 6250 665 6265 685
rect 6285 665 6300 685
rect 5650 615 5665 635
rect 5685 615 5700 635
rect 5650 585 5700 615
rect 5650 565 5665 585
rect 5685 565 5700 585
rect 5650 535 5700 565
rect 5650 515 5665 535
rect 5685 515 5700 535
rect 5650 485 5700 515
rect 5650 465 5665 485
rect 5685 465 5700 485
rect 5650 435 5700 465
rect 5650 415 5665 435
rect 5685 415 5700 435
rect 5650 385 5700 415
rect 5650 365 5665 385
rect 5685 365 5700 385
rect 5650 335 5700 365
rect 5650 315 5665 335
rect 5685 315 5700 335
rect 5650 285 5700 315
rect 5650 265 5665 285
rect 5685 265 5700 285
rect 5650 235 5700 265
rect 5650 215 5665 235
rect 5685 215 5700 235
rect 5650 185 5700 215
rect 5650 165 5665 185
rect 5685 165 5700 185
rect 5650 150 5700 165
rect 5950 635 6000 650
rect 5950 615 5965 635
rect 5985 615 6000 635
rect 5950 585 6000 615
rect 5950 565 5965 585
rect 5985 565 6000 585
rect 5950 535 6000 565
rect 5950 515 5965 535
rect 5985 515 6000 535
rect 5950 485 6000 515
rect 5950 465 5965 485
rect 5985 465 6000 485
rect 5950 435 6000 465
rect 5950 415 5965 435
rect 5985 415 6000 435
rect 5950 385 6000 415
rect 5950 365 5965 385
rect 5985 365 6000 385
rect 5950 335 6000 365
rect 5950 315 5965 335
rect 5985 315 6000 335
rect 5950 285 6000 315
rect 5950 265 5965 285
rect 5985 265 6000 285
rect 5950 235 6000 265
rect 5950 215 5965 235
rect 5985 215 6000 235
rect 5950 185 6000 215
rect 5950 165 5965 185
rect 5985 165 6000 185
rect 5350 115 5365 135
rect 5385 115 5400 135
rect 5350 100 5400 115
rect 5950 135 6000 165
rect 6250 635 6300 665
rect 6850 685 6900 700
rect 6850 665 6865 685
rect 6885 665 6900 685
rect 6250 615 6265 635
rect 6285 615 6300 635
rect 6250 585 6300 615
rect 6250 565 6265 585
rect 6285 565 6300 585
rect 6250 535 6300 565
rect 6250 515 6265 535
rect 6285 515 6300 535
rect 6250 485 6300 515
rect 6250 465 6265 485
rect 6285 465 6300 485
rect 6250 435 6300 465
rect 6250 415 6265 435
rect 6285 415 6300 435
rect 6250 385 6300 415
rect 6250 365 6265 385
rect 6285 365 6300 385
rect 6250 335 6300 365
rect 6250 315 6265 335
rect 6285 315 6300 335
rect 6250 285 6300 315
rect 6250 265 6265 285
rect 6285 265 6300 285
rect 6250 235 6300 265
rect 6250 215 6265 235
rect 6285 215 6300 235
rect 6250 185 6300 215
rect 6250 165 6265 185
rect 6285 165 6300 185
rect 6250 150 6300 165
rect 6550 635 6600 650
rect 6550 615 6565 635
rect 6585 615 6600 635
rect 6550 585 6600 615
rect 6550 565 6565 585
rect 6585 565 6600 585
rect 6550 535 6600 565
rect 6550 515 6565 535
rect 6585 515 6600 535
rect 6550 485 6600 515
rect 6550 465 6565 485
rect 6585 465 6600 485
rect 6550 435 6600 465
rect 6550 415 6565 435
rect 6585 415 6600 435
rect 6550 385 6600 415
rect 6550 365 6565 385
rect 6585 365 6600 385
rect 6550 335 6600 365
rect 6550 315 6565 335
rect 6585 315 6600 335
rect 6550 285 6600 315
rect 6550 265 6565 285
rect 6585 265 6600 285
rect 6550 235 6600 265
rect 6550 215 6565 235
rect 6585 215 6600 235
rect 6550 185 6600 215
rect 6550 165 6565 185
rect 6585 165 6600 185
rect 5950 115 5965 135
rect 5985 115 6000 135
rect 5950 100 6000 115
rect 6550 135 6600 165
rect 6850 635 6900 665
rect 6850 615 6865 635
rect 6885 615 6900 635
rect 6850 585 6900 615
rect 6850 565 6865 585
rect 6885 565 6900 585
rect 6850 535 6900 565
rect 6850 515 6865 535
rect 6885 515 6900 535
rect 6850 485 6900 515
rect 6850 465 6865 485
rect 6885 465 6900 485
rect 6850 435 6900 465
rect 6850 415 6865 435
rect 6885 415 6900 435
rect 6850 385 6900 415
rect 6850 365 6865 385
rect 6885 365 6900 385
rect 6850 335 6900 365
rect 6850 315 6865 335
rect 6885 315 6900 335
rect 6850 285 6900 315
rect 6850 265 6865 285
rect 6885 265 6900 285
rect 6850 235 6900 265
rect 6850 215 6865 235
rect 6885 215 6900 235
rect 6850 185 6900 215
rect 6850 165 6865 185
rect 6885 165 6900 185
rect 6850 150 6900 165
rect 7150 735 7200 750
rect 7150 715 7165 735
rect 7185 715 7200 735
rect 7150 685 7200 715
rect 7150 665 7165 685
rect 7185 665 7200 685
rect 7150 635 7200 665
rect 7150 615 7165 635
rect 7185 615 7200 635
rect 7150 585 7200 615
rect 7150 565 7165 585
rect 7185 565 7200 585
rect 7150 535 7200 565
rect 7150 515 7165 535
rect 7185 515 7200 535
rect 7150 485 7200 515
rect 7150 465 7165 485
rect 7185 465 7200 485
rect 7150 435 7200 465
rect 7150 415 7165 435
rect 7185 415 7200 435
rect 7150 385 7200 415
rect 7150 365 7165 385
rect 7185 365 7200 385
rect 7150 335 7200 365
rect 7150 315 7165 335
rect 7185 315 7200 335
rect 7150 285 7200 315
rect 7150 265 7165 285
rect 7185 265 7200 285
rect 7150 235 7200 265
rect 7150 215 7165 235
rect 7185 215 7200 235
rect 7150 185 7200 215
rect 7150 165 7165 185
rect 7185 165 7200 185
rect 6550 115 6565 135
rect 6585 115 6600 135
rect 6550 100 6600 115
rect 7150 135 7200 165
rect 7150 115 7165 135
rect 7185 115 7200 135
rect 7150 100 7200 115
rect 1150 85 7200 100
rect 1150 65 1165 85
rect 1185 65 1765 85
rect 1785 65 2365 85
rect 2385 65 2965 85
rect 2985 65 3565 85
rect 3585 65 3865 85
rect 3885 65 4165 85
rect 4185 65 4465 85
rect 4485 65 4765 85
rect 4785 65 5365 85
rect 5385 65 5965 85
rect 5985 65 6565 85
rect 6585 65 7165 85
rect 7185 65 7200 85
rect 1150 50 7200 65
rect 8350 740 8400 910
rect 9550 1585 9600 1600
rect 9550 1565 9565 1585
rect 9585 1565 9600 1585
rect 9550 1535 9600 1565
rect 9550 1515 9565 1535
rect 9585 1515 9600 1535
rect 9550 1485 9600 1515
rect 9550 1465 9565 1485
rect 9585 1465 9600 1485
rect 9550 1435 9600 1465
rect 9550 1415 9565 1435
rect 9585 1415 9600 1435
rect 9550 1385 9600 1415
rect 9550 1365 9565 1385
rect 9585 1365 9600 1385
rect 9550 1335 9600 1365
rect 9550 1315 9565 1335
rect 9585 1315 9600 1335
rect 9550 1285 9600 1315
rect 9550 1265 9565 1285
rect 9585 1265 9600 1285
rect 9550 1235 9600 1265
rect 9550 1215 9565 1235
rect 9585 1215 9600 1235
rect 9550 1185 9600 1215
rect 9550 1165 9565 1185
rect 9585 1165 9600 1185
rect 9550 1135 9600 1165
rect 9550 1115 9565 1135
rect 9585 1115 9600 1135
rect 9550 1085 9600 1115
rect 9550 1065 9565 1085
rect 9585 1065 9600 1085
rect 9550 1035 9600 1065
rect 9550 1015 9565 1035
rect 9585 1015 9600 1035
rect 9550 985 9600 1015
rect 9550 965 9565 985
rect 9585 965 9600 985
rect 9550 935 9600 965
rect 9550 915 9565 935
rect 9585 915 9600 935
rect 8500 840 8550 850
rect 8500 810 8510 840
rect 8540 810 8550 840
rect 8500 800 8550 810
rect 8800 840 8850 850
rect 8800 810 8810 840
rect 8840 810 8850 840
rect 8800 800 8850 810
rect 9100 840 9150 850
rect 9100 810 9110 840
rect 9140 810 9150 840
rect 9100 800 9150 810
rect 9400 840 9450 850
rect 9400 810 9410 840
rect 9440 810 9450 840
rect 9400 800 9450 810
rect 9550 840 9600 915
rect 10750 1585 10800 1660
rect 15550 1690 15600 1700
rect 15550 1660 15560 1690
rect 15590 1660 15600 1690
rect 10750 1565 10765 1585
rect 10785 1565 10800 1585
rect 10750 1540 10800 1565
rect 10750 1510 10760 1540
rect 10790 1510 10800 1540
rect 10750 1485 10800 1510
rect 10750 1465 10765 1485
rect 10785 1465 10800 1485
rect 10750 1440 10800 1465
rect 10750 1410 10760 1440
rect 10790 1410 10800 1440
rect 10750 1385 10800 1410
rect 10750 1365 10765 1385
rect 10785 1365 10800 1385
rect 10750 1340 10800 1365
rect 10750 1310 10760 1340
rect 10790 1310 10800 1340
rect 10750 1285 10800 1310
rect 10750 1265 10765 1285
rect 10785 1265 10800 1285
rect 10750 1240 10800 1265
rect 10750 1210 10760 1240
rect 10790 1210 10800 1240
rect 10750 1185 10800 1210
rect 10750 1165 10765 1185
rect 10785 1165 10800 1185
rect 10750 1140 10800 1165
rect 10750 1110 10760 1140
rect 10790 1110 10800 1140
rect 10750 1085 10800 1110
rect 10750 1065 10765 1085
rect 10785 1065 10800 1085
rect 10750 1040 10800 1065
rect 10750 1010 10760 1040
rect 10790 1010 10800 1040
rect 10750 985 10800 1010
rect 10750 965 10765 985
rect 10785 965 10800 985
rect 10750 940 10800 965
rect 10750 910 10760 940
rect 10790 910 10800 940
rect 9550 810 9560 840
rect 9590 810 9600 840
rect 8350 710 8360 740
rect 8390 710 8400 740
rect 8350 685 8400 710
rect 8350 665 8365 685
rect 8385 665 8400 685
rect 8350 640 8400 665
rect 8350 610 8360 640
rect 8390 610 8400 640
rect 8350 585 8400 610
rect 8350 565 8365 585
rect 8385 565 8400 585
rect 8350 540 8400 565
rect 8350 510 8360 540
rect 8390 510 8400 540
rect 8350 485 8400 510
rect 8350 465 8365 485
rect 8385 465 8400 485
rect 8350 440 8400 465
rect 8350 410 8360 440
rect 8390 410 8400 440
rect 8350 385 8400 410
rect 8350 365 8365 385
rect 8385 365 8400 385
rect 8350 340 8400 365
rect 8350 310 8360 340
rect 8390 310 8400 340
rect 8350 285 8400 310
rect 8350 265 8365 285
rect 8385 265 8400 285
rect 8350 240 8400 265
rect 8350 210 8360 240
rect 8390 210 8400 240
rect 8350 185 8400 210
rect 8350 165 8365 185
rect 8385 165 8400 185
rect 8350 140 8400 165
rect 8350 110 8360 140
rect 8390 110 8400 140
rect 8350 85 8400 110
rect 8350 65 8365 85
rect 8385 65 8400 85
rect -50 -40 -40 -10
rect -10 -40 0 -10
rect -650 -135 -635 -115
rect -615 -135 -600 -115
rect -650 -160 -600 -135
rect -650 -190 -640 -160
rect -610 -190 -600 -160
rect -650 -215 -600 -190
rect -650 -235 -635 -215
rect -615 -235 -600 -215
rect -650 -260 -600 -235
rect -650 -290 -640 -260
rect -610 -290 -600 -260
rect -650 -315 -600 -290
rect -650 -335 -635 -315
rect -615 -335 -600 -315
rect -650 -360 -600 -335
rect -650 -390 -640 -360
rect -610 -390 -600 -360
rect -650 -415 -600 -390
rect -650 -435 -635 -415
rect -615 -435 -600 -415
rect -650 -460 -600 -435
rect -650 -490 -640 -460
rect -610 -490 -600 -460
rect -650 -515 -600 -490
rect -650 -535 -635 -515
rect -615 -535 -600 -515
rect -650 -560 -600 -535
rect -650 -590 -640 -560
rect -610 -590 -600 -560
rect -650 -615 -600 -590
rect -650 -635 -635 -615
rect -615 -635 -600 -615
rect -650 -660 -600 -635
rect -650 -690 -640 -660
rect -610 -690 -600 -660
rect -650 -715 -600 -690
rect -650 -735 -635 -715
rect -615 -735 -600 -715
rect -650 -760 -600 -735
rect -650 -790 -640 -760
rect -610 -790 -600 -760
rect -650 -960 -600 -790
rect -500 -115 -450 -100
rect -500 -135 -485 -115
rect -465 -135 -450 -115
rect -500 -165 -450 -135
rect -500 -185 -485 -165
rect -465 -185 -450 -165
rect -500 -215 -450 -185
rect -500 -235 -485 -215
rect -465 -235 -450 -215
rect -500 -265 -450 -235
rect -500 -285 -485 -265
rect -465 -285 -450 -265
rect -500 -315 -450 -285
rect -500 -335 -485 -315
rect -465 -335 -450 -315
rect -500 -365 -450 -335
rect -500 -385 -485 -365
rect -465 -385 -450 -365
rect -500 -415 -450 -385
rect -500 -435 -485 -415
rect -465 -435 -450 -415
rect -500 -465 -450 -435
rect -500 -485 -485 -465
rect -465 -485 -450 -465
rect -500 -515 -450 -485
rect -500 -535 -485 -515
rect -465 -535 -450 -515
rect -500 -565 -450 -535
rect -500 -585 -485 -565
rect -465 -585 -450 -565
rect -500 -615 -450 -585
rect -500 -635 -485 -615
rect -465 -635 -450 -615
rect -500 -665 -450 -635
rect -500 -685 -485 -665
rect -465 -685 -450 -665
rect -500 -715 -450 -685
rect -500 -735 -485 -715
rect -465 -735 -450 -715
rect -500 -765 -450 -735
rect -500 -785 -485 -765
rect -465 -785 -450 -765
rect -500 -800 -450 -785
rect -350 -115 -300 -100
rect -350 -135 -335 -115
rect -315 -135 -300 -115
rect -350 -165 -300 -135
rect -350 -185 -335 -165
rect -315 -185 -300 -165
rect -350 -215 -300 -185
rect -350 -235 -335 -215
rect -315 -235 -300 -215
rect -350 -265 -300 -235
rect -350 -285 -335 -265
rect -315 -285 -300 -265
rect -350 -315 -300 -285
rect -350 -335 -335 -315
rect -315 -335 -300 -315
rect -350 -365 -300 -335
rect -350 -385 -335 -365
rect -315 -385 -300 -365
rect -350 -415 -300 -385
rect -350 -435 -335 -415
rect -315 -435 -300 -415
rect -350 -465 -300 -435
rect -350 -485 -335 -465
rect -315 -485 -300 -465
rect -350 -515 -300 -485
rect -350 -535 -335 -515
rect -315 -535 -300 -515
rect -350 -565 -300 -535
rect -350 -585 -335 -565
rect -315 -585 -300 -565
rect -350 -615 -300 -585
rect -350 -635 -335 -615
rect -315 -635 -300 -615
rect -350 -665 -300 -635
rect -350 -685 -335 -665
rect -315 -685 -300 -665
rect -350 -715 -300 -685
rect -350 -735 -335 -715
rect -315 -735 -300 -715
rect -350 -765 -300 -735
rect -350 -785 -335 -765
rect -315 -785 -300 -765
rect -500 -860 -450 -850
rect -500 -890 -490 -860
rect -460 -890 -450 -860
rect -500 -900 -450 -890
rect -350 -860 -300 -785
rect -200 -115 -150 -100
rect -200 -135 -185 -115
rect -165 -135 -150 -115
rect -200 -165 -150 -135
rect -200 -185 -185 -165
rect -165 -185 -150 -165
rect -200 -215 -150 -185
rect -200 -235 -185 -215
rect -165 -235 -150 -215
rect -200 -265 -150 -235
rect -200 -285 -185 -265
rect -165 -285 -150 -265
rect -200 -315 -150 -285
rect -200 -335 -185 -315
rect -165 -335 -150 -315
rect -200 -365 -150 -335
rect -200 -385 -185 -365
rect -165 -385 -150 -365
rect -200 -415 -150 -385
rect -200 -435 -185 -415
rect -165 -435 -150 -415
rect -200 -465 -150 -435
rect -200 -485 -185 -465
rect -165 -485 -150 -465
rect -200 -515 -150 -485
rect -200 -535 -185 -515
rect -165 -535 -150 -515
rect -200 -565 -150 -535
rect -200 -585 -185 -565
rect -165 -585 -150 -565
rect -200 -615 -150 -585
rect -200 -635 -185 -615
rect -165 -635 -150 -615
rect -200 -665 -150 -635
rect -200 -685 -185 -665
rect -165 -685 -150 -665
rect -200 -715 -150 -685
rect -200 -735 -185 -715
rect -165 -735 -150 -715
rect -200 -765 -150 -735
rect -200 -785 -185 -765
rect -165 -785 -150 -765
rect -200 -800 -150 -785
rect -50 -115 0 -40
rect 8350 -10 8400 65
rect 9550 735 9600 810
rect 9700 840 9750 850
rect 9700 810 9710 840
rect 9740 810 9750 840
rect 9700 800 9750 810
rect 10000 840 10050 850
rect 10000 810 10010 840
rect 10040 810 10050 840
rect 10000 800 10050 810
rect 10300 840 10350 850
rect 10300 810 10310 840
rect 10340 810 10350 840
rect 10300 800 10350 810
rect 10600 840 10650 850
rect 10600 810 10610 840
rect 10640 810 10650 840
rect 10600 800 10650 810
rect 9550 715 9565 735
rect 9585 715 9600 735
rect 9550 685 9600 715
rect 9550 665 9565 685
rect 9585 665 9600 685
rect 9550 635 9600 665
rect 9550 615 9565 635
rect 9585 615 9600 635
rect 9550 585 9600 615
rect 9550 565 9565 585
rect 9585 565 9600 585
rect 9550 535 9600 565
rect 9550 515 9565 535
rect 9585 515 9600 535
rect 9550 485 9600 515
rect 9550 465 9565 485
rect 9585 465 9600 485
rect 9550 435 9600 465
rect 9550 415 9565 435
rect 9585 415 9600 435
rect 9550 385 9600 415
rect 9550 365 9565 385
rect 9585 365 9600 385
rect 9550 335 9600 365
rect 9550 315 9565 335
rect 9585 315 9600 335
rect 9550 285 9600 315
rect 9550 265 9565 285
rect 9585 265 9600 285
rect 9550 235 9600 265
rect 9550 215 9565 235
rect 9585 215 9600 235
rect 9550 185 9600 215
rect 9550 165 9565 185
rect 9585 165 9600 185
rect 9550 135 9600 165
rect 9550 115 9565 135
rect 9585 115 9600 135
rect 9550 85 9600 115
rect 9550 65 9565 85
rect 9585 65 9600 85
rect 9550 50 9600 65
rect 10750 740 10800 910
rect 11950 1585 14400 1600
rect 11950 1565 11965 1585
rect 11985 1565 12565 1585
rect 12585 1565 13165 1585
rect 13185 1565 13765 1585
rect 13785 1565 14365 1585
rect 14385 1565 14400 1585
rect 11950 1550 14400 1565
rect 11950 1535 12000 1550
rect 11950 1515 11965 1535
rect 11985 1515 12000 1535
rect 11950 1485 12000 1515
rect 12550 1535 12600 1550
rect 12550 1515 12565 1535
rect 12585 1515 12600 1535
rect 11950 1465 11965 1485
rect 11985 1465 12000 1485
rect 11950 1435 12000 1465
rect 11950 1415 11965 1435
rect 11985 1415 12000 1435
rect 11950 1385 12000 1415
rect 11950 1365 11965 1385
rect 11985 1365 12000 1385
rect 11950 1335 12000 1365
rect 11950 1315 11965 1335
rect 11985 1315 12000 1335
rect 11950 1285 12000 1315
rect 11950 1265 11965 1285
rect 11985 1265 12000 1285
rect 11950 1235 12000 1265
rect 11950 1215 11965 1235
rect 11985 1215 12000 1235
rect 11950 1185 12000 1215
rect 11950 1165 11965 1185
rect 11985 1165 12000 1185
rect 11950 1135 12000 1165
rect 11950 1115 11965 1135
rect 11985 1115 12000 1135
rect 11950 1085 12000 1115
rect 11950 1065 11965 1085
rect 11985 1065 12000 1085
rect 11950 1035 12000 1065
rect 11950 1015 11965 1035
rect 11985 1015 12000 1035
rect 11950 985 12000 1015
rect 11950 965 11965 985
rect 11985 965 12000 985
rect 11950 935 12000 965
rect 11950 915 11965 935
rect 11985 915 12000 935
rect 10900 840 10950 850
rect 10900 810 10910 840
rect 10940 810 10950 840
rect 10900 800 10950 810
rect 11200 840 11250 850
rect 11200 810 11210 840
rect 11240 810 11250 840
rect 11200 800 11250 810
rect 11500 840 11550 850
rect 11500 810 11510 840
rect 11540 810 11550 840
rect 11500 800 11550 810
rect 11800 840 11850 850
rect 11800 810 11810 840
rect 11840 810 11850 840
rect 11800 800 11850 810
rect 10750 710 10760 740
rect 10790 710 10800 740
rect 10750 685 10800 710
rect 10750 665 10765 685
rect 10785 665 10800 685
rect 10750 640 10800 665
rect 10750 610 10760 640
rect 10790 610 10800 640
rect 10750 585 10800 610
rect 10750 565 10765 585
rect 10785 565 10800 585
rect 10750 540 10800 565
rect 10750 510 10760 540
rect 10790 510 10800 540
rect 10750 485 10800 510
rect 10750 465 10765 485
rect 10785 465 10800 485
rect 10750 440 10800 465
rect 10750 410 10760 440
rect 10790 410 10800 440
rect 10750 385 10800 410
rect 10750 365 10765 385
rect 10785 365 10800 385
rect 10750 340 10800 365
rect 10750 310 10760 340
rect 10790 310 10800 340
rect 10750 285 10800 310
rect 10750 265 10765 285
rect 10785 265 10800 285
rect 10750 240 10800 265
rect 10750 210 10760 240
rect 10790 210 10800 240
rect 10750 185 10800 210
rect 10750 165 10765 185
rect 10785 165 10800 185
rect 10750 140 10800 165
rect 10750 110 10760 140
rect 10790 110 10800 140
rect 10750 85 10800 110
rect 10750 65 10765 85
rect 10785 65 10800 85
rect 8350 -40 8360 -10
rect 8390 -40 8400 -10
rect -50 -135 -35 -115
rect -15 -135 0 -115
rect -50 -160 0 -135
rect -50 -190 -40 -160
rect -10 -190 0 -160
rect -50 -215 0 -190
rect -50 -235 -35 -215
rect -15 -235 0 -215
rect -50 -260 0 -235
rect -50 -290 -40 -260
rect -10 -290 0 -260
rect -50 -315 0 -290
rect -50 -335 -35 -315
rect -15 -335 0 -315
rect -50 -360 0 -335
rect -50 -390 -40 -360
rect -10 -390 0 -360
rect -50 -415 0 -390
rect -50 -435 -35 -415
rect -15 -435 0 -415
rect -50 -460 0 -435
rect -50 -490 -40 -460
rect -10 -490 0 -460
rect -50 -515 0 -490
rect -50 -535 -35 -515
rect -15 -535 0 -515
rect -50 -560 0 -535
rect -50 -590 -40 -560
rect -10 -590 0 -560
rect -50 -615 0 -590
rect -50 -635 -35 -615
rect -15 -635 0 -615
rect -50 -660 0 -635
rect -50 -690 -40 -660
rect -10 -690 0 -660
rect -50 -715 0 -690
rect -50 -735 -35 -715
rect -15 -735 0 -715
rect -50 -760 0 -735
rect -50 -790 -40 -760
rect -10 -790 0 -760
rect -350 -890 -340 -860
rect -310 -890 -300 -860
rect -650 -990 -640 -960
rect -610 -990 -600 -960
rect -650 -1015 -600 -990
rect -650 -1035 -635 -1015
rect -615 -1035 -600 -1015
rect -650 -1060 -600 -1035
rect -650 -1090 -640 -1060
rect -610 -1090 -600 -1060
rect -650 -1115 -600 -1090
rect -650 -1135 -635 -1115
rect -615 -1135 -600 -1115
rect -650 -1160 -600 -1135
rect -650 -1190 -640 -1160
rect -610 -1190 -600 -1160
rect -650 -1215 -600 -1190
rect -650 -1235 -635 -1215
rect -615 -1235 -600 -1215
rect -650 -1260 -600 -1235
rect -650 -1290 -640 -1260
rect -610 -1290 -600 -1260
rect -650 -1315 -600 -1290
rect -650 -1335 -635 -1315
rect -615 -1335 -600 -1315
rect -650 -1360 -600 -1335
rect -650 -1390 -640 -1360
rect -610 -1390 -600 -1360
rect -650 -1415 -600 -1390
rect -650 -1435 -635 -1415
rect -615 -1435 -600 -1415
rect -650 -1460 -600 -1435
rect -650 -1490 -640 -1460
rect -610 -1490 -600 -1460
rect -650 -1515 -600 -1490
rect -650 -1535 -635 -1515
rect -615 -1535 -600 -1515
rect -650 -1560 -600 -1535
rect -650 -1590 -640 -1560
rect -610 -1590 -600 -1560
rect -650 -1615 -600 -1590
rect -650 -1635 -635 -1615
rect -615 -1635 -600 -1615
rect -650 -1710 -600 -1635
rect -500 -965 -450 -950
rect -500 -985 -485 -965
rect -465 -985 -450 -965
rect -500 -1015 -450 -985
rect -500 -1035 -485 -1015
rect -465 -1035 -450 -1015
rect -500 -1065 -450 -1035
rect -500 -1085 -485 -1065
rect -465 -1085 -450 -1065
rect -500 -1115 -450 -1085
rect -500 -1135 -485 -1115
rect -465 -1135 -450 -1115
rect -500 -1165 -450 -1135
rect -500 -1185 -485 -1165
rect -465 -1185 -450 -1165
rect -500 -1215 -450 -1185
rect -500 -1235 -485 -1215
rect -465 -1235 -450 -1215
rect -500 -1265 -450 -1235
rect -500 -1285 -485 -1265
rect -465 -1285 -450 -1265
rect -500 -1315 -450 -1285
rect -500 -1335 -485 -1315
rect -465 -1335 -450 -1315
rect -500 -1365 -450 -1335
rect -500 -1385 -485 -1365
rect -465 -1385 -450 -1365
rect -500 -1415 -450 -1385
rect -500 -1435 -485 -1415
rect -465 -1435 -450 -1415
rect -500 -1465 -450 -1435
rect -500 -1485 -485 -1465
rect -465 -1485 -450 -1465
rect -500 -1515 -450 -1485
rect -500 -1535 -485 -1515
rect -465 -1535 -450 -1515
rect -500 -1565 -450 -1535
rect -500 -1585 -485 -1565
rect -465 -1585 -450 -1565
rect -500 -1615 -450 -1585
rect -500 -1635 -485 -1615
rect -465 -1635 -450 -1615
rect -500 -1650 -450 -1635
rect -350 -965 -300 -890
rect -200 -860 -150 -850
rect -200 -890 -190 -860
rect -160 -890 -150 -860
rect -200 -900 -150 -890
rect -350 -985 -335 -965
rect -315 -985 -300 -965
rect -350 -1015 -300 -985
rect -350 -1035 -335 -1015
rect -315 -1035 -300 -1015
rect -350 -1065 -300 -1035
rect -350 -1085 -335 -1065
rect -315 -1085 -300 -1065
rect -350 -1115 -300 -1085
rect -350 -1135 -335 -1115
rect -315 -1135 -300 -1115
rect -350 -1165 -300 -1135
rect -350 -1185 -335 -1165
rect -315 -1185 -300 -1165
rect -350 -1215 -300 -1185
rect -350 -1235 -335 -1215
rect -315 -1235 -300 -1215
rect -350 -1265 -300 -1235
rect -350 -1285 -335 -1265
rect -315 -1285 -300 -1265
rect -350 -1315 -300 -1285
rect -350 -1335 -335 -1315
rect -315 -1335 -300 -1315
rect -350 -1365 -300 -1335
rect -350 -1385 -335 -1365
rect -315 -1385 -300 -1365
rect -350 -1415 -300 -1385
rect -350 -1435 -335 -1415
rect -315 -1435 -300 -1415
rect -350 -1465 -300 -1435
rect -350 -1485 -335 -1465
rect -315 -1485 -300 -1465
rect -350 -1515 -300 -1485
rect -350 -1535 -335 -1515
rect -315 -1535 -300 -1515
rect -350 -1565 -300 -1535
rect -350 -1585 -335 -1565
rect -315 -1585 -300 -1565
rect -350 -1615 -300 -1585
rect -350 -1635 -335 -1615
rect -315 -1635 -300 -1615
rect -350 -1650 -300 -1635
rect -200 -965 -150 -950
rect -200 -985 -185 -965
rect -165 -985 -150 -965
rect -200 -1015 -150 -985
rect -200 -1035 -185 -1015
rect -165 -1035 -150 -1015
rect -200 -1065 -150 -1035
rect -200 -1085 -185 -1065
rect -165 -1085 -150 -1065
rect -200 -1115 -150 -1085
rect -200 -1135 -185 -1115
rect -165 -1135 -150 -1115
rect -200 -1165 -150 -1135
rect -200 -1185 -185 -1165
rect -165 -1185 -150 -1165
rect -200 -1215 -150 -1185
rect -200 -1235 -185 -1215
rect -165 -1235 -150 -1215
rect -200 -1265 -150 -1235
rect -200 -1285 -185 -1265
rect -165 -1285 -150 -1265
rect -200 -1315 -150 -1285
rect -200 -1335 -185 -1315
rect -165 -1335 -150 -1315
rect -200 -1365 -150 -1335
rect -200 -1385 -185 -1365
rect -165 -1385 -150 -1365
rect -200 -1415 -150 -1385
rect -200 -1435 -185 -1415
rect -165 -1435 -150 -1415
rect -200 -1465 -150 -1435
rect -200 -1485 -185 -1465
rect -165 -1485 -150 -1465
rect -200 -1515 -150 -1485
rect -200 -1535 -185 -1515
rect -165 -1535 -150 -1515
rect -200 -1565 -150 -1535
rect -200 -1585 -185 -1565
rect -165 -1585 -150 -1565
rect -200 -1615 -150 -1585
rect -200 -1635 -185 -1615
rect -165 -1635 -150 -1615
rect -200 -1650 -150 -1635
rect -50 -960 0 -790
rect 1150 -115 7200 -100
rect 1150 -135 1165 -115
rect 1185 -135 1765 -115
rect 1785 -135 2365 -115
rect 2385 -135 2965 -115
rect 2985 -135 3565 -115
rect 3585 -135 3865 -115
rect 3885 -135 4165 -115
rect 4185 -135 4465 -115
rect 4485 -135 4765 -115
rect 4785 -135 5365 -115
rect 5385 -135 5965 -115
rect 5985 -135 6565 -115
rect 6585 -135 7165 -115
rect 7185 -135 7200 -115
rect 1150 -150 7200 -135
rect 1150 -165 1200 -150
rect 1150 -185 1165 -165
rect 1185 -185 1200 -165
rect 1150 -215 1200 -185
rect 1750 -165 1800 -150
rect 1750 -185 1765 -165
rect 1785 -185 1800 -165
rect 1150 -235 1165 -215
rect 1185 -235 1200 -215
rect 1150 -265 1200 -235
rect 1150 -285 1165 -265
rect 1185 -285 1200 -265
rect 1150 -315 1200 -285
rect 1150 -335 1165 -315
rect 1185 -335 1200 -315
rect 1150 -365 1200 -335
rect 1150 -385 1165 -365
rect 1185 -385 1200 -365
rect 1150 -415 1200 -385
rect 1150 -435 1165 -415
rect 1185 -435 1200 -415
rect 1150 -465 1200 -435
rect 1150 -485 1165 -465
rect 1185 -485 1200 -465
rect 1150 -515 1200 -485
rect 1150 -535 1165 -515
rect 1185 -535 1200 -515
rect 1150 -565 1200 -535
rect 1150 -585 1165 -565
rect 1185 -585 1200 -565
rect 1150 -615 1200 -585
rect 1150 -635 1165 -615
rect 1185 -635 1200 -615
rect 1150 -665 1200 -635
rect 1150 -685 1165 -665
rect 1185 -685 1200 -665
rect 1150 -715 1200 -685
rect 1150 -735 1165 -715
rect 1185 -735 1200 -715
rect 1150 -765 1200 -735
rect 1150 -785 1165 -765
rect 1185 -785 1200 -765
rect 1150 -800 1200 -785
rect 1450 -215 1500 -200
rect 1450 -235 1465 -215
rect 1485 -235 1500 -215
rect 1450 -265 1500 -235
rect 1450 -285 1465 -265
rect 1485 -285 1500 -265
rect 1450 -315 1500 -285
rect 1450 -335 1465 -315
rect 1485 -335 1500 -315
rect 1450 -365 1500 -335
rect 1450 -385 1465 -365
rect 1485 -385 1500 -365
rect 1450 -415 1500 -385
rect 1450 -435 1465 -415
rect 1485 -435 1500 -415
rect 1450 -465 1500 -435
rect 1450 -485 1465 -465
rect 1485 -485 1500 -465
rect 1450 -515 1500 -485
rect 1450 -535 1465 -515
rect 1485 -535 1500 -515
rect 1450 -565 1500 -535
rect 1450 -585 1465 -565
rect 1485 -585 1500 -565
rect 1450 -615 1500 -585
rect 1450 -635 1465 -615
rect 1485 -635 1500 -615
rect 1450 -665 1500 -635
rect 1450 -685 1465 -665
rect 1485 -685 1500 -665
rect 1450 -715 1500 -685
rect 1750 -215 1800 -185
rect 2350 -165 2400 -150
rect 2350 -185 2365 -165
rect 2385 -185 2400 -165
rect 1750 -235 1765 -215
rect 1785 -235 1800 -215
rect 1750 -265 1800 -235
rect 1750 -285 1765 -265
rect 1785 -285 1800 -265
rect 1750 -315 1800 -285
rect 1750 -335 1765 -315
rect 1785 -335 1800 -315
rect 1750 -365 1800 -335
rect 1750 -385 1765 -365
rect 1785 -385 1800 -365
rect 1750 -415 1800 -385
rect 1750 -435 1765 -415
rect 1785 -435 1800 -415
rect 1750 -465 1800 -435
rect 1750 -485 1765 -465
rect 1785 -485 1800 -465
rect 1750 -515 1800 -485
rect 1750 -535 1765 -515
rect 1785 -535 1800 -515
rect 1750 -565 1800 -535
rect 1750 -585 1765 -565
rect 1785 -585 1800 -565
rect 1750 -615 1800 -585
rect 1750 -635 1765 -615
rect 1785 -635 1800 -615
rect 1750 -665 1800 -635
rect 1750 -685 1765 -665
rect 1785 -685 1800 -665
rect 1750 -700 1800 -685
rect 2050 -215 2100 -200
rect 2050 -235 2065 -215
rect 2085 -235 2100 -215
rect 2050 -265 2100 -235
rect 2050 -285 2065 -265
rect 2085 -285 2100 -265
rect 2050 -315 2100 -285
rect 2050 -335 2065 -315
rect 2085 -335 2100 -315
rect 2050 -365 2100 -335
rect 2050 -385 2065 -365
rect 2085 -385 2100 -365
rect 2050 -415 2100 -385
rect 2050 -435 2065 -415
rect 2085 -435 2100 -415
rect 2050 -465 2100 -435
rect 2050 -485 2065 -465
rect 2085 -485 2100 -465
rect 2050 -515 2100 -485
rect 2050 -535 2065 -515
rect 2085 -535 2100 -515
rect 2050 -565 2100 -535
rect 2050 -585 2065 -565
rect 2085 -585 2100 -565
rect 2050 -615 2100 -585
rect 2050 -635 2065 -615
rect 2085 -635 2100 -615
rect 2050 -665 2100 -635
rect 2050 -685 2065 -665
rect 2085 -685 2100 -665
rect 1450 -735 1465 -715
rect 1485 -735 1500 -715
rect 1450 -750 1500 -735
rect 2050 -715 2100 -685
rect 2350 -215 2400 -185
rect 2950 -165 3000 -150
rect 2950 -185 2965 -165
rect 2985 -185 3000 -165
rect 2350 -235 2365 -215
rect 2385 -235 2400 -215
rect 2350 -265 2400 -235
rect 2350 -285 2365 -265
rect 2385 -285 2400 -265
rect 2350 -315 2400 -285
rect 2350 -335 2365 -315
rect 2385 -335 2400 -315
rect 2350 -365 2400 -335
rect 2350 -385 2365 -365
rect 2385 -385 2400 -365
rect 2350 -415 2400 -385
rect 2350 -435 2365 -415
rect 2385 -435 2400 -415
rect 2350 -465 2400 -435
rect 2350 -485 2365 -465
rect 2385 -485 2400 -465
rect 2350 -515 2400 -485
rect 2350 -535 2365 -515
rect 2385 -535 2400 -515
rect 2350 -565 2400 -535
rect 2350 -585 2365 -565
rect 2385 -585 2400 -565
rect 2350 -615 2400 -585
rect 2350 -635 2365 -615
rect 2385 -635 2400 -615
rect 2350 -665 2400 -635
rect 2350 -685 2365 -665
rect 2385 -685 2400 -665
rect 2350 -700 2400 -685
rect 2650 -215 2700 -200
rect 2650 -235 2665 -215
rect 2685 -235 2700 -215
rect 2650 -265 2700 -235
rect 2650 -285 2665 -265
rect 2685 -285 2700 -265
rect 2650 -315 2700 -285
rect 2650 -335 2665 -315
rect 2685 -335 2700 -315
rect 2650 -365 2700 -335
rect 2650 -385 2665 -365
rect 2685 -385 2700 -365
rect 2650 -415 2700 -385
rect 2650 -435 2665 -415
rect 2685 -435 2700 -415
rect 2650 -465 2700 -435
rect 2650 -485 2665 -465
rect 2685 -485 2700 -465
rect 2650 -515 2700 -485
rect 2650 -535 2665 -515
rect 2685 -535 2700 -515
rect 2650 -565 2700 -535
rect 2650 -585 2665 -565
rect 2685 -585 2700 -565
rect 2650 -615 2700 -585
rect 2650 -635 2665 -615
rect 2685 -635 2700 -615
rect 2650 -665 2700 -635
rect 2650 -685 2665 -665
rect 2685 -685 2700 -665
rect 2050 -735 2065 -715
rect 2085 -735 2100 -715
rect 2050 -750 2100 -735
rect 2650 -715 2700 -685
rect 2950 -215 3000 -185
rect 3550 -165 3600 -150
rect 3550 -185 3565 -165
rect 3585 -185 3600 -165
rect 2950 -235 2965 -215
rect 2985 -235 3000 -215
rect 2950 -265 3000 -235
rect 2950 -285 2965 -265
rect 2985 -285 3000 -265
rect 2950 -315 3000 -285
rect 2950 -335 2965 -315
rect 2985 -335 3000 -315
rect 2950 -365 3000 -335
rect 2950 -385 2965 -365
rect 2985 -385 3000 -365
rect 2950 -415 3000 -385
rect 2950 -435 2965 -415
rect 2985 -435 3000 -415
rect 2950 -465 3000 -435
rect 2950 -485 2965 -465
rect 2985 -485 3000 -465
rect 2950 -515 3000 -485
rect 2950 -535 2965 -515
rect 2985 -535 3000 -515
rect 2950 -565 3000 -535
rect 2950 -585 2965 -565
rect 2985 -585 3000 -565
rect 2950 -615 3000 -585
rect 2950 -635 2965 -615
rect 2985 -635 3000 -615
rect 2950 -665 3000 -635
rect 2950 -685 2965 -665
rect 2985 -685 3000 -665
rect 2950 -700 3000 -685
rect 3250 -215 3300 -200
rect 3250 -235 3265 -215
rect 3285 -235 3300 -215
rect 3250 -265 3300 -235
rect 3250 -285 3265 -265
rect 3285 -285 3300 -265
rect 3250 -315 3300 -285
rect 3250 -335 3265 -315
rect 3285 -335 3300 -315
rect 3250 -365 3300 -335
rect 3250 -385 3265 -365
rect 3285 -385 3300 -365
rect 3250 -415 3300 -385
rect 3250 -435 3265 -415
rect 3285 -435 3300 -415
rect 3250 -465 3300 -435
rect 3250 -485 3265 -465
rect 3285 -485 3300 -465
rect 3250 -515 3300 -485
rect 3250 -535 3265 -515
rect 3285 -535 3300 -515
rect 3250 -565 3300 -535
rect 3250 -585 3265 -565
rect 3285 -585 3300 -565
rect 3250 -615 3300 -585
rect 3250 -635 3265 -615
rect 3285 -635 3300 -615
rect 3250 -665 3300 -635
rect 3250 -685 3265 -665
rect 3285 -685 3300 -665
rect 2650 -735 2665 -715
rect 2685 -735 2700 -715
rect 2650 -750 2700 -735
rect 3250 -715 3300 -685
rect 3250 -735 3265 -715
rect 3285 -735 3300 -715
rect 3250 -750 3300 -735
rect 1450 -765 3300 -750
rect 1450 -785 1465 -765
rect 1485 -785 2065 -765
rect 2085 -785 2665 -765
rect 2685 -785 3265 -765
rect 3285 -785 3300 -765
rect 1450 -800 3300 -785
rect 3550 -215 3600 -185
rect 3850 -165 3900 -150
rect 3850 -185 3865 -165
rect 3885 -185 3900 -165
rect 3550 -235 3565 -215
rect 3585 -235 3600 -215
rect 3550 -265 3600 -235
rect 3550 -285 3565 -265
rect 3585 -285 3600 -265
rect 3550 -315 3600 -285
rect 3550 -335 3565 -315
rect 3585 -335 3600 -315
rect 3550 -365 3600 -335
rect 3550 -385 3565 -365
rect 3585 -385 3600 -365
rect 3550 -415 3600 -385
rect 3550 -435 3565 -415
rect 3585 -435 3600 -415
rect 3550 -465 3600 -435
rect 3550 -485 3565 -465
rect 3585 -485 3600 -465
rect 3550 -515 3600 -485
rect 3550 -535 3565 -515
rect 3585 -535 3600 -515
rect 3550 -565 3600 -535
rect 3550 -585 3565 -565
rect 3585 -585 3600 -565
rect 3550 -615 3600 -585
rect 3550 -635 3565 -615
rect 3585 -635 3600 -615
rect 3550 -665 3600 -635
rect 3550 -685 3565 -665
rect 3585 -685 3600 -665
rect 3550 -715 3600 -685
rect 3550 -735 3565 -715
rect 3585 -735 3600 -715
rect 3550 -765 3600 -735
rect 3550 -785 3565 -765
rect 3585 -785 3600 -765
rect 3550 -800 3600 -785
rect 3700 -215 3750 -200
rect 3700 -235 3715 -215
rect 3735 -235 3750 -215
rect 3700 -265 3750 -235
rect 3700 -285 3715 -265
rect 3735 -285 3750 -265
rect 3700 -315 3750 -285
rect 3700 -335 3715 -315
rect 3735 -335 3750 -315
rect 3700 -365 3750 -335
rect 3700 -385 3715 -365
rect 3735 -385 3750 -365
rect 3700 -415 3750 -385
rect 3700 -435 3715 -415
rect 3735 -435 3750 -415
rect 3700 -465 3750 -435
rect 3700 -485 3715 -465
rect 3735 -485 3750 -465
rect 3700 -515 3750 -485
rect 3700 -535 3715 -515
rect 3735 -535 3750 -515
rect 3700 -565 3750 -535
rect 3700 -585 3715 -565
rect 3735 -585 3750 -565
rect 3700 -615 3750 -585
rect 3700 -635 3715 -615
rect 3735 -635 3750 -615
rect 3700 -665 3750 -635
rect 3700 -685 3715 -665
rect 3735 -685 3750 -665
rect 3700 -715 3750 -685
rect 3850 -215 3900 -185
rect 4150 -165 4200 -150
rect 4150 -185 4165 -165
rect 4185 -185 4200 -165
rect 3850 -235 3865 -215
rect 3885 -235 3900 -215
rect 3850 -265 3900 -235
rect 3850 -285 3865 -265
rect 3885 -285 3900 -265
rect 3850 -315 3900 -285
rect 3850 -335 3865 -315
rect 3885 -335 3900 -315
rect 3850 -365 3900 -335
rect 3850 -385 3865 -365
rect 3885 -385 3900 -365
rect 3850 -415 3900 -385
rect 3850 -435 3865 -415
rect 3885 -435 3900 -415
rect 3850 -465 3900 -435
rect 3850 -485 3865 -465
rect 3885 -485 3900 -465
rect 3850 -515 3900 -485
rect 3850 -535 3865 -515
rect 3885 -535 3900 -515
rect 3850 -565 3900 -535
rect 3850 -585 3865 -565
rect 3885 -585 3900 -565
rect 3850 -615 3900 -585
rect 3850 -635 3865 -615
rect 3885 -635 3900 -615
rect 3850 -665 3900 -635
rect 3850 -685 3865 -665
rect 3885 -685 3900 -665
rect 3850 -700 3900 -685
rect 4000 -215 4050 -200
rect 4000 -235 4015 -215
rect 4035 -235 4050 -215
rect 4000 -265 4050 -235
rect 4000 -285 4015 -265
rect 4035 -285 4050 -265
rect 4000 -315 4050 -285
rect 4000 -335 4015 -315
rect 4035 -335 4050 -315
rect 4000 -365 4050 -335
rect 4000 -385 4015 -365
rect 4035 -385 4050 -365
rect 4000 -415 4050 -385
rect 4000 -435 4015 -415
rect 4035 -435 4050 -415
rect 4000 -465 4050 -435
rect 4000 -485 4015 -465
rect 4035 -485 4050 -465
rect 4000 -515 4050 -485
rect 4000 -535 4015 -515
rect 4035 -535 4050 -515
rect 4000 -565 4050 -535
rect 4000 -585 4015 -565
rect 4035 -585 4050 -565
rect 4000 -615 4050 -585
rect 4000 -635 4015 -615
rect 4035 -635 4050 -615
rect 4000 -665 4050 -635
rect 4000 -685 4015 -665
rect 4035 -685 4050 -665
rect 3700 -735 3715 -715
rect 3735 -735 3750 -715
rect 3700 -750 3750 -735
rect 4000 -715 4050 -685
rect 4000 -735 4015 -715
rect 4035 -735 4050 -715
rect 4000 -750 4050 -735
rect 3700 -765 4050 -750
rect 3700 -785 3715 -765
rect 3735 -785 4015 -765
rect 4035 -785 4050 -765
rect 3700 -800 4050 -785
rect 4150 -215 4200 -185
rect 4450 -165 4500 -150
rect 4450 -185 4465 -165
rect 4485 -185 4500 -165
rect 4150 -235 4165 -215
rect 4185 -235 4200 -215
rect 4150 -265 4200 -235
rect 4150 -285 4165 -265
rect 4185 -285 4200 -265
rect 4150 -315 4200 -285
rect 4150 -335 4165 -315
rect 4185 -335 4200 -315
rect 4150 -365 4200 -335
rect 4150 -385 4165 -365
rect 4185 -385 4200 -365
rect 4150 -415 4200 -385
rect 4150 -435 4165 -415
rect 4185 -435 4200 -415
rect 4150 -465 4200 -435
rect 4150 -485 4165 -465
rect 4185 -485 4200 -465
rect 4150 -515 4200 -485
rect 4150 -535 4165 -515
rect 4185 -535 4200 -515
rect 4150 -565 4200 -535
rect 4150 -585 4165 -565
rect 4185 -585 4200 -565
rect 4150 -615 4200 -585
rect 4150 -635 4165 -615
rect 4185 -635 4200 -615
rect 4150 -665 4200 -635
rect 4150 -685 4165 -665
rect 4185 -685 4200 -665
rect 4150 -715 4200 -685
rect 4150 -735 4165 -715
rect 4185 -735 4200 -715
rect 4150 -765 4200 -735
rect 4150 -785 4165 -765
rect 4185 -785 4200 -765
rect 4150 -800 4200 -785
rect 4300 -215 4350 -200
rect 4300 -235 4315 -215
rect 4335 -235 4350 -215
rect 4300 -265 4350 -235
rect 4300 -285 4315 -265
rect 4335 -285 4350 -265
rect 4300 -315 4350 -285
rect 4300 -335 4315 -315
rect 4335 -335 4350 -315
rect 4300 -365 4350 -335
rect 4300 -385 4315 -365
rect 4335 -385 4350 -365
rect 4300 -415 4350 -385
rect 4300 -435 4315 -415
rect 4335 -435 4350 -415
rect 4300 -465 4350 -435
rect 4300 -485 4315 -465
rect 4335 -485 4350 -465
rect 4300 -515 4350 -485
rect 4300 -535 4315 -515
rect 4335 -535 4350 -515
rect 4300 -565 4350 -535
rect 4300 -585 4315 -565
rect 4335 -585 4350 -565
rect 4300 -615 4350 -585
rect 4300 -635 4315 -615
rect 4335 -635 4350 -615
rect 4300 -665 4350 -635
rect 4300 -685 4315 -665
rect 4335 -685 4350 -665
rect 4300 -715 4350 -685
rect 4450 -215 4500 -185
rect 4750 -165 4800 -150
rect 4750 -185 4765 -165
rect 4785 -185 4800 -165
rect 4450 -235 4465 -215
rect 4485 -235 4500 -215
rect 4450 -265 4500 -235
rect 4450 -285 4465 -265
rect 4485 -285 4500 -265
rect 4450 -315 4500 -285
rect 4450 -335 4465 -315
rect 4485 -335 4500 -315
rect 4450 -365 4500 -335
rect 4450 -385 4465 -365
rect 4485 -385 4500 -365
rect 4450 -415 4500 -385
rect 4450 -435 4465 -415
rect 4485 -435 4500 -415
rect 4450 -465 4500 -435
rect 4450 -485 4465 -465
rect 4485 -485 4500 -465
rect 4450 -515 4500 -485
rect 4450 -535 4465 -515
rect 4485 -535 4500 -515
rect 4450 -565 4500 -535
rect 4450 -585 4465 -565
rect 4485 -585 4500 -565
rect 4450 -615 4500 -585
rect 4450 -635 4465 -615
rect 4485 -635 4500 -615
rect 4450 -665 4500 -635
rect 4450 -685 4465 -665
rect 4485 -685 4500 -665
rect 4450 -700 4500 -685
rect 4600 -215 4650 -200
rect 4600 -235 4615 -215
rect 4635 -235 4650 -215
rect 4600 -265 4650 -235
rect 4600 -285 4615 -265
rect 4635 -285 4650 -265
rect 4600 -315 4650 -285
rect 4600 -335 4615 -315
rect 4635 -335 4650 -315
rect 4600 -365 4650 -335
rect 4600 -385 4615 -365
rect 4635 -385 4650 -365
rect 4600 -415 4650 -385
rect 4600 -435 4615 -415
rect 4635 -435 4650 -415
rect 4600 -465 4650 -435
rect 4600 -485 4615 -465
rect 4635 -485 4650 -465
rect 4600 -515 4650 -485
rect 4600 -535 4615 -515
rect 4635 -535 4650 -515
rect 4600 -565 4650 -535
rect 4600 -585 4615 -565
rect 4635 -585 4650 -565
rect 4600 -615 4650 -585
rect 4600 -635 4615 -615
rect 4635 -635 4650 -615
rect 4600 -665 4650 -635
rect 4600 -685 4615 -665
rect 4635 -685 4650 -665
rect 4300 -735 4315 -715
rect 4335 -735 4350 -715
rect 4300 -750 4350 -735
rect 4600 -715 4650 -685
rect 4600 -735 4615 -715
rect 4635 -735 4650 -715
rect 4600 -750 4650 -735
rect 4300 -765 4650 -750
rect 4300 -785 4315 -765
rect 4335 -785 4615 -765
rect 4635 -785 4650 -765
rect 4300 -800 4650 -785
rect 4750 -215 4800 -185
rect 5350 -165 5400 -150
rect 5350 -185 5365 -165
rect 5385 -185 5400 -165
rect 4750 -235 4765 -215
rect 4785 -235 4800 -215
rect 4750 -265 4800 -235
rect 4750 -285 4765 -265
rect 4785 -285 4800 -265
rect 4750 -315 4800 -285
rect 4750 -335 4765 -315
rect 4785 -335 4800 -315
rect 4750 -365 4800 -335
rect 4750 -385 4765 -365
rect 4785 -385 4800 -365
rect 4750 -415 4800 -385
rect 4750 -435 4765 -415
rect 4785 -435 4800 -415
rect 4750 -465 4800 -435
rect 4750 -485 4765 -465
rect 4785 -485 4800 -465
rect 4750 -515 4800 -485
rect 4750 -535 4765 -515
rect 4785 -535 4800 -515
rect 4750 -565 4800 -535
rect 4750 -585 4765 -565
rect 4785 -585 4800 -565
rect 4750 -615 4800 -585
rect 4750 -635 4765 -615
rect 4785 -635 4800 -615
rect 4750 -665 4800 -635
rect 4750 -685 4765 -665
rect 4785 -685 4800 -665
rect 4750 -715 4800 -685
rect 4750 -735 4765 -715
rect 4785 -735 4800 -715
rect 4750 -765 4800 -735
rect 4750 -785 4765 -765
rect 4785 -785 4800 -765
rect 4750 -800 4800 -785
rect 5050 -215 5100 -200
rect 5050 -235 5065 -215
rect 5085 -235 5100 -215
rect 5050 -265 5100 -235
rect 5050 -285 5065 -265
rect 5085 -285 5100 -265
rect 5050 -315 5100 -285
rect 5050 -335 5065 -315
rect 5085 -335 5100 -315
rect 5050 -365 5100 -335
rect 5050 -385 5065 -365
rect 5085 -385 5100 -365
rect 5050 -415 5100 -385
rect 5050 -435 5065 -415
rect 5085 -435 5100 -415
rect 5050 -465 5100 -435
rect 5050 -485 5065 -465
rect 5085 -485 5100 -465
rect 5050 -515 5100 -485
rect 5050 -535 5065 -515
rect 5085 -535 5100 -515
rect 5050 -565 5100 -535
rect 5050 -585 5065 -565
rect 5085 -585 5100 -565
rect 5050 -615 5100 -585
rect 5050 -635 5065 -615
rect 5085 -635 5100 -615
rect 5050 -665 5100 -635
rect 5050 -685 5065 -665
rect 5085 -685 5100 -665
rect 5050 -715 5100 -685
rect 5350 -215 5400 -185
rect 5950 -165 6000 -150
rect 5950 -185 5965 -165
rect 5985 -185 6000 -165
rect 5350 -235 5365 -215
rect 5385 -235 5400 -215
rect 5350 -265 5400 -235
rect 5350 -285 5365 -265
rect 5385 -285 5400 -265
rect 5350 -315 5400 -285
rect 5350 -335 5365 -315
rect 5385 -335 5400 -315
rect 5350 -365 5400 -335
rect 5350 -385 5365 -365
rect 5385 -385 5400 -365
rect 5350 -415 5400 -385
rect 5350 -435 5365 -415
rect 5385 -435 5400 -415
rect 5350 -465 5400 -435
rect 5350 -485 5365 -465
rect 5385 -485 5400 -465
rect 5350 -515 5400 -485
rect 5350 -535 5365 -515
rect 5385 -535 5400 -515
rect 5350 -565 5400 -535
rect 5350 -585 5365 -565
rect 5385 -585 5400 -565
rect 5350 -615 5400 -585
rect 5350 -635 5365 -615
rect 5385 -635 5400 -615
rect 5350 -665 5400 -635
rect 5350 -685 5365 -665
rect 5385 -685 5400 -665
rect 5350 -700 5400 -685
rect 5650 -215 5700 -200
rect 5650 -235 5665 -215
rect 5685 -235 5700 -215
rect 5650 -265 5700 -235
rect 5650 -285 5665 -265
rect 5685 -285 5700 -265
rect 5650 -315 5700 -285
rect 5650 -335 5665 -315
rect 5685 -335 5700 -315
rect 5650 -365 5700 -335
rect 5650 -385 5665 -365
rect 5685 -385 5700 -365
rect 5650 -415 5700 -385
rect 5650 -435 5665 -415
rect 5685 -435 5700 -415
rect 5650 -465 5700 -435
rect 5650 -485 5665 -465
rect 5685 -485 5700 -465
rect 5650 -515 5700 -485
rect 5650 -535 5665 -515
rect 5685 -535 5700 -515
rect 5650 -565 5700 -535
rect 5650 -585 5665 -565
rect 5685 -585 5700 -565
rect 5650 -615 5700 -585
rect 5650 -635 5665 -615
rect 5685 -635 5700 -615
rect 5650 -665 5700 -635
rect 5650 -685 5665 -665
rect 5685 -685 5700 -665
rect 5050 -735 5065 -715
rect 5085 -735 5100 -715
rect 5050 -750 5100 -735
rect 5650 -715 5700 -685
rect 5950 -215 6000 -185
rect 6550 -165 6600 -150
rect 6550 -185 6565 -165
rect 6585 -185 6600 -165
rect 5950 -235 5965 -215
rect 5985 -235 6000 -215
rect 5950 -265 6000 -235
rect 5950 -285 5965 -265
rect 5985 -285 6000 -265
rect 5950 -315 6000 -285
rect 5950 -335 5965 -315
rect 5985 -335 6000 -315
rect 5950 -365 6000 -335
rect 5950 -385 5965 -365
rect 5985 -385 6000 -365
rect 5950 -415 6000 -385
rect 5950 -435 5965 -415
rect 5985 -435 6000 -415
rect 5950 -465 6000 -435
rect 5950 -485 5965 -465
rect 5985 -485 6000 -465
rect 5950 -515 6000 -485
rect 5950 -535 5965 -515
rect 5985 -535 6000 -515
rect 5950 -565 6000 -535
rect 5950 -585 5965 -565
rect 5985 -585 6000 -565
rect 5950 -615 6000 -585
rect 5950 -635 5965 -615
rect 5985 -635 6000 -615
rect 5950 -665 6000 -635
rect 5950 -685 5965 -665
rect 5985 -685 6000 -665
rect 5950 -700 6000 -685
rect 6250 -215 6300 -200
rect 6250 -235 6265 -215
rect 6285 -235 6300 -215
rect 6250 -265 6300 -235
rect 6250 -285 6265 -265
rect 6285 -285 6300 -265
rect 6250 -315 6300 -285
rect 6250 -335 6265 -315
rect 6285 -335 6300 -315
rect 6250 -365 6300 -335
rect 6250 -385 6265 -365
rect 6285 -385 6300 -365
rect 6250 -415 6300 -385
rect 6250 -435 6265 -415
rect 6285 -435 6300 -415
rect 6250 -465 6300 -435
rect 6250 -485 6265 -465
rect 6285 -485 6300 -465
rect 6250 -515 6300 -485
rect 6250 -535 6265 -515
rect 6285 -535 6300 -515
rect 6250 -565 6300 -535
rect 6250 -585 6265 -565
rect 6285 -585 6300 -565
rect 6250 -615 6300 -585
rect 6250 -635 6265 -615
rect 6285 -635 6300 -615
rect 6250 -665 6300 -635
rect 6250 -685 6265 -665
rect 6285 -685 6300 -665
rect 5650 -735 5665 -715
rect 5685 -735 5700 -715
rect 5650 -750 5700 -735
rect 6250 -715 6300 -685
rect 6550 -215 6600 -185
rect 7150 -165 7200 -150
rect 7150 -185 7165 -165
rect 7185 -185 7200 -165
rect 6550 -235 6565 -215
rect 6585 -235 6600 -215
rect 6550 -265 6600 -235
rect 6550 -285 6565 -265
rect 6585 -285 6600 -265
rect 6550 -315 6600 -285
rect 6550 -335 6565 -315
rect 6585 -335 6600 -315
rect 6550 -365 6600 -335
rect 6550 -385 6565 -365
rect 6585 -385 6600 -365
rect 6550 -415 6600 -385
rect 6550 -435 6565 -415
rect 6585 -435 6600 -415
rect 6550 -465 6600 -435
rect 6550 -485 6565 -465
rect 6585 -485 6600 -465
rect 6550 -515 6600 -485
rect 6550 -535 6565 -515
rect 6585 -535 6600 -515
rect 6550 -565 6600 -535
rect 6550 -585 6565 -565
rect 6585 -585 6600 -565
rect 6550 -615 6600 -585
rect 6550 -635 6565 -615
rect 6585 -635 6600 -615
rect 6550 -665 6600 -635
rect 6550 -685 6565 -665
rect 6585 -685 6600 -665
rect 6550 -700 6600 -685
rect 6850 -215 6900 -200
rect 6850 -235 6865 -215
rect 6885 -235 6900 -215
rect 6850 -265 6900 -235
rect 6850 -285 6865 -265
rect 6885 -285 6900 -265
rect 6850 -315 6900 -285
rect 6850 -335 6865 -315
rect 6885 -335 6900 -315
rect 6850 -365 6900 -335
rect 6850 -385 6865 -365
rect 6885 -385 6900 -365
rect 6850 -415 6900 -385
rect 6850 -435 6865 -415
rect 6885 -435 6900 -415
rect 6850 -465 6900 -435
rect 6850 -485 6865 -465
rect 6885 -485 6900 -465
rect 6850 -515 6900 -485
rect 6850 -535 6865 -515
rect 6885 -535 6900 -515
rect 6850 -565 6900 -535
rect 6850 -585 6865 -565
rect 6885 -585 6900 -565
rect 6850 -615 6900 -585
rect 6850 -635 6865 -615
rect 6885 -635 6900 -615
rect 6850 -665 6900 -635
rect 6850 -685 6865 -665
rect 6885 -685 6900 -665
rect 6250 -735 6265 -715
rect 6285 -735 6300 -715
rect 6250 -750 6300 -735
rect 6850 -715 6900 -685
rect 6850 -735 6865 -715
rect 6885 -735 6900 -715
rect 6850 -750 6900 -735
rect 5050 -765 6900 -750
rect 5050 -785 5065 -765
rect 5085 -785 5665 -765
rect 5685 -785 6265 -765
rect 6285 -785 6865 -765
rect 6885 -785 6900 -765
rect 5050 -800 6900 -785
rect 7150 -215 7200 -185
rect 7150 -235 7165 -215
rect 7185 -235 7200 -215
rect 7150 -265 7200 -235
rect 7150 -285 7165 -265
rect 7185 -285 7200 -265
rect 7150 -315 7200 -285
rect 7150 -335 7165 -315
rect 7185 -335 7200 -315
rect 7150 -365 7200 -335
rect 7150 -385 7165 -365
rect 7185 -385 7200 -365
rect 7150 -415 7200 -385
rect 7150 -435 7165 -415
rect 7185 -435 7200 -415
rect 7150 -465 7200 -435
rect 7150 -485 7165 -465
rect 7185 -485 7200 -465
rect 7150 -515 7200 -485
rect 7150 -535 7165 -515
rect 7185 -535 7200 -515
rect 7150 -565 7200 -535
rect 7150 -585 7165 -565
rect 7185 -585 7200 -565
rect 7150 -615 7200 -585
rect 7150 -635 7165 -615
rect 7185 -635 7200 -615
rect 7150 -665 7200 -635
rect 7150 -685 7165 -665
rect 7185 -685 7200 -665
rect 7150 -715 7200 -685
rect 7150 -735 7165 -715
rect 7185 -735 7200 -715
rect 7150 -765 7200 -735
rect 7150 -785 7165 -765
rect 7185 -785 7200 -765
rect 7150 -800 7200 -785
rect 8350 -115 8400 -40
rect 10750 -10 10800 65
rect 10750 -40 10760 -10
rect 10790 -40 10800 -10
rect 8350 -135 8365 -115
rect 8385 -135 8400 -115
rect 8350 -160 8400 -135
rect 8350 -190 8360 -160
rect 8390 -190 8400 -160
rect 8350 -215 8400 -190
rect 8350 -235 8365 -215
rect 8385 -235 8400 -215
rect 8350 -260 8400 -235
rect 8350 -290 8360 -260
rect 8390 -290 8400 -260
rect 8350 -315 8400 -290
rect 8350 -335 8365 -315
rect 8385 -335 8400 -315
rect 8350 -360 8400 -335
rect 8350 -390 8360 -360
rect 8390 -390 8400 -360
rect 8350 -415 8400 -390
rect 8350 -435 8365 -415
rect 8385 -435 8400 -415
rect 8350 -460 8400 -435
rect 8350 -490 8360 -460
rect 8390 -490 8400 -460
rect 8350 -515 8400 -490
rect 8350 -535 8365 -515
rect 8385 -535 8400 -515
rect 8350 -560 8400 -535
rect 8350 -590 8360 -560
rect 8390 -590 8400 -560
rect 8350 -615 8400 -590
rect 8350 -635 8365 -615
rect 8385 -635 8400 -615
rect 8350 -660 8400 -635
rect 8350 -690 8360 -660
rect 8390 -690 8400 -660
rect 8350 -715 8400 -690
rect 8350 -735 8365 -715
rect 8385 -735 8400 -715
rect 8350 -760 8400 -735
rect 8350 -790 8360 -760
rect 8390 -790 8400 -760
rect 100 -860 150 -850
rect 100 -890 110 -860
rect 140 -890 150 -860
rect 100 -900 150 -890
rect 400 -860 450 -850
rect 400 -890 410 -860
rect 440 -890 450 -860
rect 400 -900 450 -890
rect 700 -860 750 -850
rect 700 -890 710 -860
rect 740 -890 750 -860
rect 700 -900 750 -890
rect 1000 -860 1050 -850
rect 1000 -890 1010 -860
rect 1040 -890 1050 -860
rect 1000 -900 1050 -890
rect 1300 -860 1350 -850
rect 1300 -890 1310 -860
rect 1340 -890 1350 -860
rect 1300 -900 1350 -890
rect 1600 -860 1650 -850
rect 1600 -890 1610 -860
rect 1640 -890 1650 -860
rect 1600 -900 1650 -890
rect 1900 -860 1950 -850
rect 1900 -890 1910 -860
rect 1940 -890 1950 -860
rect 1900 -900 1950 -890
rect 2200 -860 2250 -850
rect 2200 -890 2210 -860
rect 2240 -890 2250 -860
rect 2200 -900 2250 -890
rect 2350 -860 2400 -800
rect 2350 -890 2360 -860
rect 2390 -890 2400 -860
rect 2350 -950 2400 -890
rect 2500 -860 2550 -850
rect 2500 -890 2510 -860
rect 2540 -890 2550 -860
rect 2500 -900 2550 -890
rect 2800 -860 2850 -850
rect 2800 -890 2810 -860
rect 2840 -890 2850 -860
rect 2800 -900 2850 -890
rect 3100 -860 3150 -850
rect 3100 -890 3110 -860
rect 3140 -890 3150 -860
rect 3100 -900 3150 -890
rect 3400 -860 3450 -850
rect 3400 -890 3410 -860
rect 3440 -890 3450 -860
rect 3400 -900 3450 -890
rect 3700 -860 3750 -850
rect 3700 -890 3710 -860
rect 3740 -890 3750 -860
rect 3700 -900 3750 -890
rect 3850 -860 3900 -800
rect 3850 -890 3860 -860
rect 3890 -890 3900 -860
rect 3850 -950 3900 -890
rect 4000 -860 4050 -850
rect 4000 -890 4010 -860
rect 4040 -890 4050 -860
rect 4000 -900 4050 -890
rect 4300 -860 4350 -850
rect 4300 -890 4310 -860
rect 4340 -890 4350 -860
rect 4300 -900 4350 -890
rect 4450 -860 4500 -800
rect 4450 -890 4460 -860
rect 4490 -890 4500 -860
rect 4450 -950 4500 -890
rect 4600 -860 4650 -850
rect 4600 -890 4610 -860
rect 4640 -890 4650 -860
rect 4600 -900 4650 -890
rect 4900 -860 4950 -850
rect 4900 -890 4910 -860
rect 4940 -890 4950 -860
rect 4900 -900 4950 -890
rect 5200 -860 5250 -850
rect 5200 -890 5210 -860
rect 5240 -890 5250 -860
rect 5200 -900 5250 -890
rect 5500 -860 5550 -850
rect 5500 -890 5510 -860
rect 5540 -890 5550 -860
rect 5500 -900 5550 -890
rect 5800 -860 5850 -850
rect 5800 -890 5810 -860
rect 5840 -890 5850 -860
rect 5800 -900 5850 -890
rect 5950 -860 6000 -800
rect 5950 -890 5960 -860
rect 5990 -890 6000 -860
rect 5950 -950 6000 -890
rect 6100 -860 6150 -850
rect 6100 -890 6110 -860
rect 6140 -890 6150 -860
rect 6100 -900 6150 -890
rect 6400 -860 6450 -850
rect 6400 -890 6410 -860
rect 6440 -890 6450 -860
rect 6400 -900 6450 -890
rect 6700 -860 6750 -850
rect 6700 -890 6710 -860
rect 6740 -890 6750 -860
rect 6700 -900 6750 -890
rect 7000 -860 7050 -850
rect 7000 -890 7010 -860
rect 7040 -890 7050 -860
rect 7000 -900 7050 -890
rect 7300 -860 7350 -850
rect 7300 -890 7310 -860
rect 7340 -890 7350 -860
rect 7300 -900 7350 -890
rect 7600 -860 7650 -850
rect 7600 -890 7610 -860
rect 7640 -890 7650 -860
rect 7600 -900 7650 -890
rect 7900 -860 7950 -850
rect 7900 -890 7910 -860
rect 7940 -890 7950 -860
rect 7900 -900 7950 -890
rect 8200 -860 8250 -850
rect 8200 -890 8210 -860
rect 8240 -890 8250 -860
rect 8200 -900 8250 -890
rect -50 -990 -40 -960
rect -10 -990 0 -960
rect -50 -1015 0 -990
rect -50 -1035 -35 -1015
rect -15 -1035 0 -1015
rect -50 -1060 0 -1035
rect -50 -1090 -40 -1060
rect -10 -1090 0 -1060
rect -50 -1115 0 -1090
rect -50 -1135 -35 -1115
rect -15 -1135 0 -1115
rect -50 -1160 0 -1135
rect -50 -1190 -40 -1160
rect -10 -1190 0 -1160
rect -50 -1215 0 -1190
rect -50 -1235 -35 -1215
rect -15 -1235 0 -1215
rect -50 -1260 0 -1235
rect -50 -1290 -40 -1260
rect -10 -1290 0 -1260
rect -50 -1315 0 -1290
rect -50 -1335 -35 -1315
rect -15 -1335 0 -1315
rect -50 -1360 0 -1335
rect -50 -1390 -40 -1360
rect -10 -1390 0 -1360
rect -50 -1415 0 -1390
rect -50 -1435 -35 -1415
rect -15 -1435 0 -1415
rect -50 -1460 0 -1435
rect -50 -1490 -40 -1460
rect -10 -1490 0 -1460
rect -50 -1515 0 -1490
rect -50 -1535 -35 -1515
rect -15 -1535 0 -1515
rect -50 -1560 0 -1535
rect -50 -1590 -40 -1560
rect -10 -1590 0 -1560
rect -50 -1615 0 -1590
rect -50 -1635 -35 -1615
rect -15 -1635 0 -1615
rect -650 -1740 -640 -1710
rect -610 -1740 -600 -1710
rect -650 -1750 -600 -1740
rect -50 -1710 0 -1635
rect 1150 -965 1200 -950
rect 1150 -985 1165 -965
rect 1185 -985 1200 -965
rect 1150 -1015 1200 -985
rect 1150 -1035 1165 -1015
rect 1185 -1035 1200 -1015
rect 1150 -1065 1200 -1035
rect 1150 -1085 1165 -1065
rect 1185 -1085 1200 -1065
rect 1150 -1115 1200 -1085
rect 1150 -1135 1165 -1115
rect 1185 -1135 1200 -1115
rect 1150 -1165 1200 -1135
rect 1150 -1185 1165 -1165
rect 1185 -1185 1200 -1165
rect 1150 -1215 1200 -1185
rect 1150 -1235 1165 -1215
rect 1185 -1235 1200 -1215
rect 1150 -1265 1200 -1235
rect 1150 -1285 1165 -1265
rect 1185 -1285 1200 -1265
rect 1150 -1315 1200 -1285
rect 1150 -1335 1165 -1315
rect 1185 -1335 1200 -1315
rect 1150 -1365 1200 -1335
rect 1150 -1385 1165 -1365
rect 1185 -1385 1200 -1365
rect 1150 -1415 1200 -1385
rect 1150 -1435 1165 -1415
rect 1185 -1435 1200 -1415
rect 1150 -1465 1200 -1435
rect 1150 -1485 1165 -1465
rect 1185 -1485 1200 -1465
rect 1150 -1515 1200 -1485
rect 1150 -1535 1165 -1515
rect 1185 -1535 1200 -1515
rect 1150 -1565 1200 -1535
rect 1450 -965 3300 -950
rect 1450 -985 1465 -965
rect 1485 -985 2065 -965
rect 2085 -985 2665 -965
rect 2685 -985 3265 -965
rect 3285 -985 3300 -965
rect 1450 -1000 3300 -985
rect 1450 -1015 1500 -1000
rect 1450 -1035 1465 -1015
rect 1485 -1035 1500 -1015
rect 1450 -1065 1500 -1035
rect 2050 -1015 2100 -1000
rect 2050 -1035 2065 -1015
rect 2085 -1035 2100 -1015
rect 1450 -1085 1465 -1065
rect 1485 -1085 1500 -1065
rect 1450 -1115 1500 -1085
rect 1450 -1135 1465 -1115
rect 1485 -1135 1500 -1115
rect 1450 -1165 1500 -1135
rect 1450 -1185 1465 -1165
rect 1485 -1185 1500 -1165
rect 1450 -1215 1500 -1185
rect 1450 -1235 1465 -1215
rect 1485 -1235 1500 -1215
rect 1450 -1265 1500 -1235
rect 1450 -1285 1465 -1265
rect 1485 -1285 1500 -1265
rect 1450 -1315 1500 -1285
rect 1450 -1335 1465 -1315
rect 1485 -1335 1500 -1315
rect 1450 -1365 1500 -1335
rect 1450 -1385 1465 -1365
rect 1485 -1385 1500 -1365
rect 1450 -1415 1500 -1385
rect 1450 -1435 1465 -1415
rect 1485 -1435 1500 -1415
rect 1450 -1465 1500 -1435
rect 1450 -1485 1465 -1465
rect 1485 -1485 1500 -1465
rect 1450 -1515 1500 -1485
rect 1450 -1535 1465 -1515
rect 1485 -1535 1500 -1515
rect 1450 -1550 1500 -1535
rect 1750 -1065 1800 -1050
rect 1750 -1085 1765 -1065
rect 1785 -1085 1800 -1065
rect 1750 -1115 1800 -1085
rect 1750 -1135 1765 -1115
rect 1785 -1135 1800 -1115
rect 1750 -1165 1800 -1135
rect 1750 -1185 1765 -1165
rect 1785 -1185 1800 -1165
rect 1750 -1215 1800 -1185
rect 1750 -1235 1765 -1215
rect 1785 -1235 1800 -1215
rect 1750 -1265 1800 -1235
rect 1750 -1285 1765 -1265
rect 1785 -1285 1800 -1265
rect 1750 -1315 1800 -1285
rect 1750 -1335 1765 -1315
rect 1785 -1335 1800 -1315
rect 1750 -1365 1800 -1335
rect 1750 -1385 1765 -1365
rect 1785 -1385 1800 -1365
rect 1750 -1415 1800 -1385
rect 1750 -1435 1765 -1415
rect 1785 -1435 1800 -1415
rect 1750 -1465 1800 -1435
rect 1750 -1485 1765 -1465
rect 1785 -1485 1800 -1465
rect 1750 -1515 1800 -1485
rect 1750 -1535 1765 -1515
rect 1785 -1535 1800 -1515
rect 1150 -1585 1165 -1565
rect 1185 -1585 1200 -1565
rect 1150 -1600 1200 -1585
rect 1750 -1565 1800 -1535
rect 2050 -1065 2100 -1035
rect 2650 -1015 2700 -1000
rect 2650 -1035 2665 -1015
rect 2685 -1035 2700 -1015
rect 2050 -1085 2065 -1065
rect 2085 -1085 2100 -1065
rect 2050 -1115 2100 -1085
rect 2050 -1135 2065 -1115
rect 2085 -1135 2100 -1115
rect 2050 -1165 2100 -1135
rect 2050 -1185 2065 -1165
rect 2085 -1185 2100 -1165
rect 2050 -1215 2100 -1185
rect 2050 -1235 2065 -1215
rect 2085 -1235 2100 -1215
rect 2050 -1265 2100 -1235
rect 2050 -1285 2065 -1265
rect 2085 -1285 2100 -1265
rect 2050 -1315 2100 -1285
rect 2050 -1335 2065 -1315
rect 2085 -1335 2100 -1315
rect 2050 -1365 2100 -1335
rect 2050 -1385 2065 -1365
rect 2085 -1385 2100 -1365
rect 2050 -1415 2100 -1385
rect 2050 -1435 2065 -1415
rect 2085 -1435 2100 -1415
rect 2050 -1465 2100 -1435
rect 2050 -1485 2065 -1465
rect 2085 -1485 2100 -1465
rect 2050 -1515 2100 -1485
rect 2050 -1535 2065 -1515
rect 2085 -1535 2100 -1515
rect 2050 -1550 2100 -1535
rect 2350 -1065 2400 -1050
rect 2350 -1085 2365 -1065
rect 2385 -1085 2400 -1065
rect 2350 -1115 2400 -1085
rect 2350 -1135 2365 -1115
rect 2385 -1135 2400 -1115
rect 2350 -1165 2400 -1135
rect 2350 -1185 2365 -1165
rect 2385 -1185 2400 -1165
rect 2350 -1215 2400 -1185
rect 2350 -1235 2365 -1215
rect 2385 -1235 2400 -1215
rect 2350 -1265 2400 -1235
rect 2350 -1285 2365 -1265
rect 2385 -1285 2400 -1265
rect 2350 -1315 2400 -1285
rect 2350 -1335 2365 -1315
rect 2385 -1335 2400 -1315
rect 2350 -1365 2400 -1335
rect 2350 -1385 2365 -1365
rect 2385 -1385 2400 -1365
rect 2350 -1415 2400 -1385
rect 2350 -1435 2365 -1415
rect 2385 -1435 2400 -1415
rect 2350 -1465 2400 -1435
rect 2350 -1485 2365 -1465
rect 2385 -1485 2400 -1465
rect 2350 -1515 2400 -1485
rect 2350 -1535 2365 -1515
rect 2385 -1535 2400 -1515
rect 1750 -1585 1765 -1565
rect 1785 -1585 1800 -1565
rect 1750 -1600 1800 -1585
rect 2350 -1565 2400 -1535
rect 2650 -1065 2700 -1035
rect 3250 -1015 3300 -1000
rect 3250 -1035 3265 -1015
rect 3285 -1035 3300 -1015
rect 2650 -1085 2665 -1065
rect 2685 -1085 2700 -1065
rect 2650 -1115 2700 -1085
rect 2650 -1135 2665 -1115
rect 2685 -1135 2700 -1115
rect 2650 -1165 2700 -1135
rect 2650 -1185 2665 -1165
rect 2685 -1185 2700 -1165
rect 2650 -1215 2700 -1185
rect 2650 -1235 2665 -1215
rect 2685 -1235 2700 -1215
rect 2650 -1265 2700 -1235
rect 2650 -1285 2665 -1265
rect 2685 -1285 2700 -1265
rect 2650 -1315 2700 -1285
rect 2650 -1335 2665 -1315
rect 2685 -1335 2700 -1315
rect 2650 -1365 2700 -1335
rect 2650 -1385 2665 -1365
rect 2685 -1385 2700 -1365
rect 2650 -1415 2700 -1385
rect 2650 -1435 2665 -1415
rect 2685 -1435 2700 -1415
rect 2650 -1465 2700 -1435
rect 2650 -1485 2665 -1465
rect 2685 -1485 2700 -1465
rect 2650 -1515 2700 -1485
rect 2650 -1535 2665 -1515
rect 2685 -1535 2700 -1515
rect 2650 -1550 2700 -1535
rect 2950 -1065 3000 -1050
rect 2950 -1085 2965 -1065
rect 2985 -1085 3000 -1065
rect 2950 -1115 3000 -1085
rect 2950 -1135 2965 -1115
rect 2985 -1135 3000 -1115
rect 2950 -1165 3000 -1135
rect 2950 -1185 2965 -1165
rect 2985 -1185 3000 -1165
rect 2950 -1215 3000 -1185
rect 2950 -1235 2965 -1215
rect 2985 -1235 3000 -1215
rect 2950 -1265 3000 -1235
rect 2950 -1285 2965 -1265
rect 2985 -1285 3000 -1265
rect 2950 -1315 3000 -1285
rect 2950 -1335 2965 -1315
rect 2985 -1335 3000 -1315
rect 2950 -1365 3000 -1335
rect 2950 -1385 2965 -1365
rect 2985 -1385 3000 -1365
rect 2950 -1415 3000 -1385
rect 2950 -1435 2965 -1415
rect 2985 -1435 3000 -1415
rect 2950 -1465 3000 -1435
rect 2950 -1485 2965 -1465
rect 2985 -1485 3000 -1465
rect 2950 -1515 3000 -1485
rect 2950 -1535 2965 -1515
rect 2985 -1535 3000 -1515
rect 2350 -1585 2365 -1565
rect 2385 -1585 2400 -1565
rect 2350 -1600 2400 -1585
rect 2950 -1565 3000 -1535
rect 3250 -1065 3300 -1035
rect 3250 -1085 3265 -1065
rect 3285 -1085 3300 -1065
rect 3250 -1115 3300 -1085
rect 3250 -1135 3265 -1115
rect 3285 -1135 3300 -1115
rect 3250 -1165 3300 -1135
rect 3250 -1185 3265 -1165
rect 3285 -1185 3300 -1165
rect 3250 -1215 3300 -1185
rect 3250 -1235 3265 -1215
rect 3285 -1235 3300 -1215
rect 3250 -1265 3300 -1235
rect 3250 -1285 3265 -1265
rect 3285 -1285 3300 -1265
rect 3250 -1315 3300 -1285
rect 3250 -1335 3265 -1315
rect 3285 -1335 3300 -1315
rect 3250 -1365 3300 -1335
rect 3250 -1385 3265 -1365
rect 3285 -1385 3300 -1365
rect 3250 -1415 3300 -1385
rect 3250 -1435 3265 -1415
rect 3285 -1435 3300 -1415
rect 3250 -1465 3300 -1435
rect 3250 -1485 3265 -1465
rect 3285 -1485 3300 -1465
rect 3250 -1515 3300 -1485
rect 3250 -1535 3265 -1515
rect 3285 -1535 3300 -1515
rect 3250 -1550 3300 -1535
rect 3550 -965 3600 -950
rect 3550 -985 3565 -965
rect 3585 -985 3600 -965
rect 3550 -1015 3600 -985
rect 3550 -1035 3565 -1015
rect 3585 -1035 3600 -1015
rect 3550 -1065 3600 -1035
rect 3550 -1085 3565 -1065
rect 3585 -1085 3600 -1065
rect 3550 -1115 3600 -1085
rect 3550 -1135 3565 -1115
rect 3585 -1135 3600 -1115
rect 3550 -1165 3600 -1135
rect 3550 -1185 3565 -1165
rect 3585 -1185 3600 -1165
rect 3550 -1215 3600 -1185
rect 3550 -1235 3565 -1215
rect 3585 -1235 3600 -1215
rect 3550 -1265 3600 -1235
rect 3550 -1285 3565 -1265
rect 3585 -1285 3600 -1265
rect 3550 -1315 3600 -1285
rect 3550 -1335 3565 -1315
rect 3585 -1335 3600 -1315
rect 3550 -1365 3600 -1335
rect 3550 -1385 3565 -1365
rect 3585 -1385 3600 -1365
rect 3550 -1415 3600 -1385
rect 3550 -1435 3565 -1415
rect 3585 -1435 3600 -1415
rect 3550 -1465 3600 -1435
rect 3550 -1485 3565 -1465
rect 3585 -1485 3600 -1465
rect 3550 -1515 3600 -1485
rect 3550 -1535 3565 -1515
rect 3585 -1535 3600 -1515
rect 2950 -1585 2965 -1565
rect 2985 -1585 3000 -1565
rect 2950 -1600 3000 -1585
rect 3550 -1565 3600 -1535
rect 3700 -965 4050 -950
rect 3700 -985 3715 -965
rect 3735 -985 4015 -965
rect 4035 -985 4050 -965
rect 3700 -1000 4050 -985
rect 3700 -1015 3750 -1000
rect 3700 -1035 3715 -1015
rect 3735 -1035 3750 -1015
rect 3700 -1065 3750 -1035
rect 4000 -1015 4050 -1000
rect 4000 -1035 4015 -1015
rect 4035 -1035 4050 -1015
rect 3700 -1085 3715 -1065
rect 3735 -1085 3750 -1065
rect 3700 -1115 3750 -1085
rect 3700 -1135 3715 -1115
rect 3735 -1135 3750 -1115
rect 3700 -1165 3750 -1135
rect 3700 -1185 3715 -1165
rect 3735 -1185 3750 -1165
rect 3700 -1215 3750 -1185
rect 3700 -1235 3715 -1215
rect 3735 -1235 3750 -1215
rect 3700 -1265 3750 -1235
rect 3700 -1285 3715 -1265
rect 3735 -1285 3750 -1265
rect 3700 -1315 3750 -1285
rect 3700 -1335 3715 -1315
rect 3735 -1335 3750 -1315
rect 3700 -1365 3750 -1335
rect 3700 -1385 3715 -1365
rect 3735 -1385 3750 -1365
rect 3700 -1415 3750 -1385
rect 3700 -1435 3715 -1415
rect 3735 -1435 3750 -1415
rect 3700 -1465 3750 -1435
rect 3700 -1485 3715 -1465
rect 3735 -1485 3750 -1465
rect 3700 -1515 3750 -1485
rect 3700 -1535 3715 -1515
rect 3735 -1535 3750 -1515
rect 3700 -1550 3750 -1535
rect 3850 -1065 3900 -1050
rect 3850 -1085 3865 -1065
rect 3885 -1085 3900 -1065
rect 3850 -1115 3900 -1085
rect 3850 -1135 3865 -1115
rect 3885 -1135 3900 -1115
rect 3850 -1165 3900 -1135
rect 3850 -1185 3865 -1165
rect 3885 -1185 3900 -1165
rect 3850 -1215 3900 -1185
rect 3850 -1235 3865 -1215
rect 3885 -1235 3900 -1215
rect 3850 -1265 3900 -1235
rect 3850 -1285 3865 -1265
rect 3885 -1285 3900 -1265
rect 3850 -1315 3900 -1285
rect 3850 -1335 3865 -1315
rect 3885 -1335 3900 -1315
rect 3850 -1365 3900 -1335
rect 3850 -1385 3865 -1365
rect 3885 -1385 3900 -1365
rect 3850 -1415 3900 -1385
rect 3850 -1435 3865 -1415
rect 3885 -1435 3900 -1415
rect 3850 -1465 3900 -1435
rect 3850 -1485 3865 -1465
rect 3885 -1485 3900 -1465
rect 3850 -1515 3900 -1485
rect 3850 -1535 3865 -1515
rect 3885 -1535 3900 -1515
rect 3550 -1585 3565 -1565
rect 3585 -1585 3600 -1565
rect 3550 -1600 3600 -1585
rect 3850 -1565 3900 -1535
rect 4000 -1065 4050 -1035
rect 4000 -1085 4015 -1065
rect 4035 -1085 4050 -1065
rect 4000 -1115 4050 -1085
rect 4000 -1135 4015 -1115
rect 4035 -1135 4050 -1115
rect 4000 -1165 4050 -1135
rect 4000 -1185 4015 -1165
rect 4035 -1185 4050 -1165
rect 4000 -1215 4050 -1185
rect 4000 -1235 4015 -1215
rect 4035 -1235 4050 -1215
rect 4000 -1265 4050 -1235
rect 4000 -1285 4015 -1265
rect 4035 -1285 4050 -1265
rect 4000 -1315 4050 -1285
rect 4000 -1335 4015 -1315
rect 4035 -1335 4050 -1315
rect 4000 -1365 4050 -1335
rect 4000 -1385 4015 -1365
rect 4035 -1385 4050 -1365
rect 4000 -1415 4050 -1385
rect 4000 -1435 4015 -1415
rect 4035 -1435 4050 -1415
rect 4000 -1465 4050 -1435
rect 4000 -1485 4015 -1465
rect 4035 -1485 4050 -1465
rect 4000 -1515 4050 -1485
rect 4000 -1535 4015 -1515
rect 4035 -1535 4050 -1515
rect 4000 -1550 4050 -1535
rect 4150 -965 4200 -950
rect 4150 -985 4165 -965
rect 4185 -985 4200 -965
rect 4150 -1015 4200 -985
rect 4150 -1035 4165 -1015
rect 4185 -1035 4200 -1015
rect 4150 -1065 4200 -1035
rect 4150 -1085 4165 -1065
rect 4185 -1085 4200 -1065
rect 4150 -1115 4200 -1085
rect 4150 -1135 4165 -1115
rect 4185 -1135 4200 -1115
rect 4150 -1165 4200 -1135
rect 4150 -1185 4165 -1165
rect 4185 -1185 4200 -1165
rect 4150 -1215 4200 -1185
rect 4150 -1235 4165 -1215
rect 4185 -1235 4200 -1215
rect 4150 -1265 4200 -1235
rect 4150 -1285 4165 -1265
rect 4185 -1285 4200 -1265
rect 4150 -1315 4200 -1285
rect 4150 -1335 4165 -1315
rect 4185 -1335 4200 -1315
rect 4150 -1365 4200 -1335
rect 4150 -1385 4165 -1365
rect 4185 -1385 4200 -1365
rect 4150 -1415 4200 -1385
rect 4150 -1435 4165 -1415
rect 4185 -1435 4200 -1415
rect 4150 -1465 4200 -1435
rect 4150 -1485 4165 -1465
rect 4185 -1485 4200 -1465
rect 4150 -1515 4200 -1485
rect 4150 -1535 4165 -1515
rect 4185 -1535 4200 -1515
rect 3850 -1585 3865 -1565
rect 3885 -1585 3900 -1565
rect 3850 -1600 3900 -1585
rect 4150 -1565 4200 -1535
rect 4300 -965 4650 -950
rect 4300 -985 4315 -965
rect 4335 -985 4615 -965
rect 4635 -985 4650 -965
rect 4300 -1000 4650 -985
rect 4300 -1015 4350 -1000
rect 4300 -1035 4315 -1015
rect 4335 -1035 4350 -1015
rect 4300 -1065 4350 -1035
rect 4600 -1015 4650 -1000
rect 4600 -1035 4615 -1015
rect 4635 -1035 4650 -1015
rect 4300 -1085 4315 -1065
rect 4335 -1085 4350 -1065
rect 4300 -1115 4350 -1085
rect 4300 -1135 4315 -1115
rect 4335 -1135 4350 -1115
rect 4300 -1165 4350 -1135
rect 4300 -1185 4315 -1165
rect 4335 -1185 4350 -1165
rect 4300 -1215 4350 -1185
rect 4300 -1235 4315 -1215
rect 4335 -1235 4350 -1215
rect 4300 -1265 4350 -1235
rect 4300 -1285 4315 -1265
rect 4335 -1285 4350 -1265
rect 4300 -1315 4350 -1285
rect 4300 -1335 4315 -1315
rect 4335 -1335 4350 -1315
rect 4300 -1365 4350 -1335
rect 4300 -1385 4315 -1365
rect 4335 -1385 4350 -1365
rect 4300 -1415 4350 -1385
rect 4300 -1435 4315 -1415
rect 4335 -1435 4350 -1415
rect 4300 -1465 4350 -1435
rect 4300 -1485 4315 -1465
rect 4335 -1485 4350 -1465
rect 4300 -1515 4350 -1485
rect 4300 -1535 4315 -1515
rect 4335 -1535 4350 -1515
rect 4300 -1550 4350 -1535
rect 4450 -1065 4500 -1050
rect 4450 -1085 4465 -1065
rect 4485 -1085 4500 -1065
rect 4450 -1115 4500 -1085
rect 4450 -1135 4465 -1115
rect 4485 -1135 4500 -1115
rect 4450 -1165 4500 -1135
rect 4450 -1185 4465 -1165
rect 4485 -1185 4500 -1165
rect 4450 -1215 4500 -1185
rect 4450 -1235 4465 -1215
rect 4485 -1235 4500 -1215
rect 4450 -1265 4500 -1235
rect 4450 -1285 4465 -1265
rect 4485 -1285 4500 -1265
rect 4450 -1315 4500 -1285
rect 4450 -1335 4465 -1315
rect 4485 -1335 4500 -1315
rect 4450 -1365 4500 -1335
rect 4450 -1385 4465 -1365
rect 4485 -1385 4500 -1365
rect 4450 -1415 4500 -1385
rect 4450 -1435 4465 -1415
rect 4485 -1435 4500 -1415
rect 4450 -1465 4500 -1435
rect 4450 -1485 4465 -1465
rect 4485 -1485 4500 -1465
rect 4450 -1515 4500 -1485
rect 4450 -1535 4465 -1515
rect 4485 -1535 4500 -1515
rect 4150 -1585 4165 -1565
rect 4185 -1585 4200 -1565
rect 4150 -1600 4200 -1585
rect 4450 -1565 4500 -1535
rect 4600 -1065 4650 -1035
rect 4600 -1085 4615 -1065
rect 4635 -1085 4650 -1065
rect 4600 -1115 4650 -1085
rect 4600 -1135 4615 -1115
rect 4635 -1135 4650 -1115
rect 4600 -1165 4650 -1135
rect 4600 -1185 4615 -1165
rect 4635 -1185 4650 -1165
rect 4600 -1215 4650 -1185
rect 4600 -1235 4615 -1215
rect 4635 -1235 4650 -1215
rect 4600 -1265 4650 -1235
rect 4600 -1285 4615 -1265
rect 4635 -1285 4650 -1265
rect 4600 -1315 4650 -1285
rect 4600 -1335 4615 -1315
rect 4635 -1335 4650 -1315
rect 4600 -1365 4650 -1335
rect 4600 -1385 4615 -1365
rect 4635 -1385 4650 -1365
rect 4600 -1415 4650 -1385
rect 4600 -1435 4615 -1415
rect 4635 -1435 4650 -1415
rect 4600 -1465 4650 -1435
rect 4600 -1485 4615 -1465
rect 4635 -1485 4650 -1465
rect 4600 -1515 4650 -1485
rect 4600 -1535 4615 -1515
rect 4635 -1535 4650 -1515
rect 4600 -1550 4650 -1535
rect 4750 -965 4800 -950
rect 4750 -985 4765 -965
rect 4785 -985 4800 -965
rect 4750 -1015 4800 -985
rect 4750 -1035 4765 -1015
rect 4785 -1035 4800 -1015
rect 4750 -1065 4800 -1035
rect 4750 -1085 4765 -1065
rect 4785 -1085 4800 -1065
rect 4750 -1115 4800 -1085
rect 4750 -1135 4765 -1115
rect 4785 -1135 4800 -1115
rect 4750 -1165 4800 -1135
rect 4750 -1185 4765 -1165
rect 4785 -1185 4800 -1165
rect 4750 -1215 4800 -1185
rect 4750 -1235 4765 -1215
rect 4785 -1235 4800 -1215
rect 4750 -1265 4800 -1235
rect 4750 -1285 4765 -1265
rect 4785 -1285 4800 -1265
rect 4750 -1315 4800 -1285
rect 4750 -1335 4765 -1315
rect 4785 -1335 4800 -1315
rect 4750 -1365 4800 -1335
rect 4750 -1385 4765 -1365
rect 4785 -1385 4800 -1365
rect 4750 -1415 4800 -1385
rect 4750 -1435 4765 -1415
rect 4785 -1435 4800 -1415
rect 4750 -1465 4800 -1435
rect 4750 -1485 4765 -1465
rect 4785 -1485 4800 -1465
rect 4750 -1515 4800 -1485
rect 4750 -1535 4765 -1515
rect 4785 -1535 4800 -1515
rect 4450 -1585 4465 -1565
rect 4485 -1585 4500 -1565
rect 4450 -1600 4500 -1585
rect 4750 -1565 4800 -1535
rect 5050 -965 6900 -950
rect 5050 -985 5065 -965
rect 5085 -985 5665 -965
rect 5685 -985 6265 -965
rect 6285 -985 6865 -965
rect 6885 -985 6900 -965
rect 5050 -1000 6900 -985
rect 5050 -1015 5100 -1000
rect 5050 -1035 5065 -1015
rect 5085 -1035 5100 -1015
rect 5050 -1065 5100 -1035
rect 5650 -1015 5700 -1000
rect 5650 -1035 5665 -1015
rect 5685 -1035 5700 -1015
rect 5050 -1085 5065 -1065
rect 5085 -1085 5100 -1065
rect 5050 -1115 5100 -1085
rect 5050 -1135 5065 -1115
rect 5085 -1135 5100 -1115
rect 5050 -1165 5100 -1135
rect 5050 -1185 5065 -1165
rect 5085 -1185 5100 -1165
rect 5050 -1215 5100 -1185
rect 5050 -1235 5065 -1215
rect 5085 -1235 5100 -1215
rect 5050 -1265 5100 -1235
rect 5050 -1285 5065 -1265
rect 5085 -1285 5100 -1265
rect 5050 -1315 5100 -1285
rect 5050 -1335 5065 -1315
rect 5085 -1335 5100 -1315
rect 5050 -1365 5100 -1335
rect 5050 -1385 5065 -1365
rect 5085 -1385 5100 -1365
rect 5050 -1415 5100 -1385
rect 5050 -1435 5065 -1415
rect 5085 -1435 5100 -1415
rect 5050 -1465 5100 -1435
rect 5050 -1485 5065 -1465
rect 5085 -1485 5100 -1465
rect 5050 -1515 5100 -1485
rect 5050 -1535 5065 -1515
rect 5085 -1535 5100 -1515
rect 5050 -1550 5100 -1535
rect 5350 -1065 5400 -1050
rect 5350 -1085 5365 -1065
rect 5385 -1085 5400 -1065
rect 5350 -1115 5400 -1085
rect 5350 -1135 5365 -1115
rect 5385 -1135 5400 -1115
rect 5350 -1165 5400 -1135
rect 5350 -1185 5365 -1165
rect 5385 -1185 5400 -1165
rect 5350 -1215 5400 -1185
rect 5350 -1235 5365 -1215
rect 5385 -1235 5400 -1215
rect 5350 -1265 5400 -1235
rect 5350 -1285 5365 -1265
rect 5385 -1285 5400 -1265
rect 5350 -1315 5400 -1285
rect 5350 -1335 5365 -1315
rect 5385 -1335 5400 -1315
rect 5350 -1365 5400 -1335
rect 5350 -1385 5365 -1365
rect 5385 -1385 5400 -1365
rect 5350 -1415 5400 -1385
rect 5350 -1435 5365 -1415
rect 5385 -1435 5400 -1415
rect 5350 -1465 5400 -1435
rect 5350 -1485 5365 -1465
rect 5385 -1485 5400 -1465
rect 5350 -1515 5400 -1485
rect 5350 -1535 5365 -1515
rect 5385 -1535 5400 -1515
rect 4750 -1585 4765 -1565
rect 4785 -1585 4800 -1565
rect 4750 -1600 4800 -1585
rect 5350 -1565 5400 -1535
rect 5650 -1065 5700 -1035
rect 6250 -1015 6300 -1000
rect 6250 -1035 6265 -1015
rect 6285 -1035 6300 -1015
rect 5650 -1085 5665 -1065
rect 5685 -1085 5700 -1065
rect 5650 -1115 5700 -1085
rect 5650 -1135 5665 -1115
rect 5685 -1135 5700 -1115
rect 5650 -1165 5700 -1135
rect 5650 -1185 5665 -1165
rect 5685 -1185 5700 -1165
rect 5650 -1215 5700 -1185
rect 5650 -1235 5665 -1215
rect 5685 -1235 5700 -1215
rect 5650 -1265 5700 -1235
rect 5650 -1285 5665 -1265
rect 5685 -1285 5700 -1265
rect 5650 -1315 5700 -1285
rect 5650 -1335 5665 -1315
rect 5685 -1335 5700 -1315
rect 5650 -1365 5700 -1335
rect 5650 -1385 5665 -1365
rect 5685 -1385 5700 -1365
rect 5650 -1415 5700 -1385
rect 5650 -1435 5665 -1415
rect 5685 -1435 5700 -1415
rect 5650 -1465 5700 -1435
rect 5650 -1485 5665 -1465
rect 5685 -1485 5700 -1465
rect 5650 -1515 5700 -1485
rect 5650 -1535 5665 -1515
rect 5685 -1535 5700 -1515
rect 5650 -1550 5700 -1535
rect 5950 -1065 6000 -1050
rect 5950 -1085 5965 -1065
rect 5985 -1085 6000 -1065
rect 5950 -1115 6000 -1085
rect 5950 -1135 5965 -1115
rect 5985 -1135 6000 -1115
rect 5950 -1165 6000 -1135
rect 5950 -1185 5965 -1165
rect 5985 -1185 6000 -1165
rect 5950 -1215 6000 -1185
rect 5950 -1235 5965 -1215
rect 5985 -1235 6000 -1215
rect 5950 -1265 6000 -1235
rect 5950 -1285 5965 -1265
rect 5985 -1285 6000 -1265
rect 5950 -1315 6000 -1285
rect 5950 -1335 5965 -1315
rect 5985 -1335 6000 -1315
rect 5950 -1365 6000 -1335
rect 5950 -1385 5965 -1365
rect 5985 -1385 6000 -1365
rect 5950 -1415 6000 -1385
rect 5950 -1435 5965 -1415
rect 5985 -1435 6000 -1415
rect 5950 -1465 6000 -1435
rect 5950 -1485 5965 -1465
rect 5985 -1485 6000 -1465
rect 5950 -1515 6000 -1485
rect 5950 -1535 5965 -1515
rect 5985 -1535 6000 -1515
rect 5350 -1585 5365 -1565
rect 5385 -1585 5400 -1565
rect 5350 -1600 5400 -1585
rect 5950 -1565 6000 -1535
rect 6250 -1065 6300 -1035
rect 6850 -1015 6900 -1000
rect 6850 -1035 6865 -1015
rect 6885 -1035 6900 -1015
rect 6250 -1085 6265 -1065
rect 6285 -1085 6300 -1065
rect 6250 -1115 6300 -1085
rect 6250 -1135 6265 -1115
rect 6285 -1135 6300 -1115
rect 6250 -1165 6300 -1135
rect 6250 -1185 6265 -1165
rect 6285 -1185 6300 -1165
rect 6250 -1215 6300 -1185
rect 6250 -1235 6265 -1215
rect 6285 -1235 6300 -1215
rect 6250 -1265 6300 -1235
rect 6250 -1285 6265 -1265
rect 6285 -1285 6300 -1265
rect 6250 -1315 6300 -1285
rect 6250 -1335 6265 -1315
rect 6285 -1335 6300 -1315
rect 6250 -1365 6300 -1335
rect 6250 -1385 6265 -1365
rect 6285 -1385 6300 -1365
rect 6250 -1415 6300 -1385
rect 6250 -1435 6265 -1415
rect 6285 -1435 6300 -1415
rect 6250 -1465 6300 -1435
rect 6250 -1485 6265 -1465
rect 6285 -1485 6300 -1465
rect 6250 -1515 6300 -1485
rect 6250 -1535 6265 -1515
rect 6285 -1535 6300 -1515
rect 6250 -1550 6300 -1535
rect 6550 -1065 6600 -1050
rect 6550 -1085 6565 -1065
rect 6585 -1085 6600 -1065
rect 6550 -1115 6600 -1085
rect 6550 -1135 6565 -1115
rect 6585 -1135 6600 -1115
rect 6550 -1165 6600 -1135
rect 6550 -1185 6565 -1165
rect 6585 -1185 6600 -1165
rect 6550 -1215 6600 -1185
rect 6550 -1235 6565 -1215
rect 6585 -1235 6600 -1215
rect 6550 -1265 6600 -1235
rect 6550 -1285 6565 -1265
rect 6585 -1285 6600 -1265
rect 6550 -1315 6600 -1285
rect 6550 -1335 6565 -1315
rect 6585 -1335 6600 -1315
rect 6550 -1365 6600 -1335
rect 6550 -1385 6565 -1365
rect 6585 -1385 6600 -1365
rect 6550 -1415 6600 -1385
rect 6550 -1435 6565 -1415
rect 6585 -1435 6600 -1415
rect 6550 -1465 6600 -1435
rect 6550 -1485 6565 -1465
rect 6585 -1485 6600 -1465
rect 6550 -1515 6600 -1485
rect 6550 -1535 6565 -1515
rect 6585 -1535 6600 -1515
rect 5950 -1585 5965 -1565
rect 5985 -1585 6000 -1565
rect 5950 -1600 6000 -1585
rect 6550 -1565 6600 -1535
rect 6850 -1065 6900 -1035
rect 6850 -1085 6865 -1065
rect 6885 -1085 6900 -1065
rect 6850 -1115 6900 -1085
rect 6850 -1135 6865 -1115
rect 6885 -1135 6900 -1115
rect 6850 -1165 6900 -1135
rect 6850 -1185 6865 -1165
rect 6885 -1185 6900 -1165
rect 6850 -1215 6900 -1185
rect 6850 -1235 6865 -1215
rect 6885 -1235 6900 -1215
rect 6850 -1265 6900 -1235
rect 6850 -1285 6865 -1265
rect 6885 -1285 6900 -1265
rect 6850 -1315 6900 -1285
rect 6850 -1335 6865 -1315
rect 6885 -1335 6900 -1315
rect 6850 -1365 6900 -1335
rect 6850 -1385 6865 -1365
rect 6885 -1385 6900 -1365
rect 6850 -1415 6900 -1385
rect 6850 -1435 6865 -1415
rect 6885 -1435 6900 -1415
rect 6850 -1465 6900 -1435
rect 6850 -1485 6865 -1465
rect 6885 -1485 6900 -1465
rect 6850 -1515 6900 -1485
rect 6850 -1535 6865 -1515
rect 6885 -1535 6900 -1515
rect 6850 -1550 6900 -1535
rect 7150 -965 7200 -950
rect 7150 -985 7165 -965
rect 7185 -985 7200 -965
rect 7150 -1015 7200 -985
rect 7150 -1035 7165 -1015
rect 7185 -1035 7200 -1015
rect 7150 -1065 7200 -1035
rect 7150 -1085 7165 -1065
rect 7185 -1085 7200 -1065
rect 7150 -1115 7200 -1085
rect 7150 -1135 7165 -1115
rect 7185 -1135 7200 -1115
rect 7150 -1165 7200 -1135
rect 7150 -1185 7165 -1165
rect 7185 -1185 7200 -1165
rect 7150 -1215 7200 -1185
rect 7150 -1235 7165 -1215
rect 7185 -1235 7200 -1215
rect 7150 -1265 7200 -1235
rect 7150 -1285 7165 -1265
rect 7185 -1285 7200 -1265
rect 7150 -1315 7200 -1285
rect 7150 -1335 7165 -1315
rect 7185 -1335 7200 -1315
rect 7150 -1365 7200 -1335
rect 7150 -1385 7165 -1365
rect 7185 -1385 7200 -1365
rect 7150 -1415 7200 -1385
rect 7150 -1435 7165 -1415
rect 7185 -1435 7200 -1415
rect 7150 -1465 7200 -1435
rect 7150 -1485 7165 -1465
rect 7185 -1485 7200 -1465
rect 7150 -1515 7200 -1485
rect 7150 -1535 7165 -1515
rect 7185 -1535 7200 -1515
rect 6550 -1585 6565 -1565
rect 6585 -1585 6600 -1565
rect 6550 -1600 6600 -1585
rect 7150 -1565 7200 -1535
rect 7150 -1585 7165 -1565
rect 7185 -1585 7200 -1565
rect 7150 -1600 7200 -1585
rect 1150 -1615 7200 -1600
rect 1150 -1635 1165 -1615
rect 1185 -1635 1765 -1615
rect 1785 -1635 2365 -1615
rect 2385 -1635 2965 -1615
rect 2985 -1635 3565 -1615
rect 3585 -1635 3865 -1615
rect 3885 -1635 4165 -1615
rect 4185 -1635 4465 -1615
rect 4485 -1635 4765 -1615
rect 4785 -1635 5365 -1615
rect 5385 -1635 5965 -1615
rect 5985 -1635 6565 -1615
rect 6585 -1635 7165 -1615
rect 7185 -1635 7200 -1615
rect 1150 -1650 7200 -1635
rect 8350 -960 8400 -790
rect 9550 -115 9600 -100
rect 9550 -135 9565 -115
rect 9585 -135 9600 -115
rect 9550 -165 9600 -135
rect 9550 -185 9565 -165
rect 9585 -185 9600 -165
rect 9550 -215 9600 -185
rect 9550 -235 9565 -215
rect 9585 -235 9600 -215
rect 9550 -265 9600 -235
rect 9550 -285 9565 -265
rect 9585 -285 9600 -265
rect 9550 -315 9600 -285
rect 9550 -335 9565 -315
rect 9585 -335 9600 -315
rect 9550 -365 9600 -335
rect 9550 -385 9565 -365
rect 9585 -385 9600 -365
rect 9550 -415 9600 -385
rect 9550 -435 9565 -415
rect 9585 -435 9600 -415
rect 9550 -465 9600 -435
rect 9550 -485 9565 -465
rect 9585 -485 9600 -465
rect 9550 -515 9600 -485
rect 9550 -535 9565 -515
rect 9585 -535 9600 -515
rect 9550 -565 9600 -535
rect 9550 -585 9565 -565
rect 9585 -585 9600 -565
rect 9550 -615 9600 -585
rect 9550 -635 9565 -615
rect 9585 -635 9600 -615
rect 9550 -665 9600 -635
rect 9550 -685 9565 -665
rect 9585 -685 9600 -665
rect 9550 -715 9600 -685
rect 9550 -735 9565 -715
rect 9585 -735 9600 -715
rect 9550 -765 9600 -735
rect 9550 -785 9565 -765
rect 9585 -785 9600 -765
rect 8500 -860 8550 -850
rect 8500 -890 8510 -860
rect 8540 -890 8550 -860
rect 8500 -900 8550 -890
rect 8800 -860 8850 -850
rect 8800 -890 8810 -860
rect 8840 -890 8850 -860
rect 8800 -900 8850 -890
rect 9100 -860 9150 -850
rect 9100 -890 9110 -860
rect 9140 -890 9150 -860
rect 9100 -900 9150 -890
rect 9400 -860 9450 -850
rect 9400 -890 9410 -860
rect 9440 -890 9450 -860
rect 9400 -900 9450 -890
rect 9550 -860 9600 -785
rect 10750 -115 10800 -40
rect 10750 -135 10765 -115
rect 10785 -135 10800 -115
rect 10750 -160 10800 -135
rect 10750 -190 10760 -160
rect 10790 -190 10800 -160
rect 10750 -215 10800 -190
rect 10750 -235 10765 -215
rect 10785 -235 10800 -215
rect 10750 -260 10800 -235
rect 10750 -290 10760 -260
rect 10790 -290 10800 -260
rect 10750 -315 10800 -290
rect 10750 -335 10765 -315
rect 10785 -335 10800 -315
rect 10750 -360 10800 -335
rect 10750 -390 10760 -360
rect 10790 -390 10800 -360
rect 10750 -415 10800 -390
rect 10750 -435 10765 -415
rect 10785 -435 10800 -415
rect 10750 -460 10800 -435
rect 10750 -490 10760 -460
rect 10790 -490 10800 -460
rect 10750 -515 10800 -490
rect 10750 -535 10765 -515
rect 10785 -535 10800 -515
rect 10750 -560 10800 -535
rect 10750 -590 10760 -560
rect 10790 -590 10800 -560
rect 10750 -615 10800 -590
rect 10750 -635 10765 -615
rect 10785 -635 10800 -615
rect 10750 -660 10800 -635
rect 10750 -690 10760 -660
rect 10790 -690 10800 -660
rect 10750 -715 10800 -690
rect 10750 -735 10765 -715
rect 10785 -735 10800 -715
rect 10750 -760 10800 -735
rect 10750 -790 10760 -760
rect 10790 -790 10800 -760
rect 9550 -890 9560 -860
rect 9590 -890 9600 -860
rect 8350 -990 8360 -960
rect 8390 -990 8400 -960
rect 8350 -1015 8400 -990
rect 8350 -1035 8365 -1015
rect 8385 -1035 8400 -1015
rect 8350 -1060 8400 -1035
rect 8350 -1090 8360 -1060
rect 8390 -1090 8400 -1060
rect 8350 -1115 8400 -1090
rect 8350 -1135 8365 -1115
rect 8385 -1135 8400 -1115
rect 8350 -1160 8400 -1135
rect 8350 -1190 8360 -1160
rect 8390 -1190 8400 -1160
rect 8350 -1215 8400 -1190
rect 8350 -1235 8365 -1215
rect 8385 -1235 8400 -1215
rect 8350 -1260 8400 -1235
rect 8350 -1290 8360 -1260
rect 8390 -1290 8400 -1260
rect 8350 -1315 8400 -1290
rect 8350 -1335 8365 -1315
rect 8385 -1335 8400 -1315
rect 8350 -1360 8400 -1335
rect 8350 -1390 8360 -1360
rect 8390 -1390 8400 -1360
rect 8350 -1415 8400 -1390
rect 8350 -1435 8365 -1415
rect 8385 -1435 8400 -1415
rect 8350 -1460 8400 -1435
rect 8350 -1490 8360 -1460
rect 8390 -1490 8400 -1460
rect 8350 -1515 8400 -1490
rect 8350 -1535 8365 -1515
rect 8385 -1535 8400 -1515
rect 8350 -1560 8400 -1535
rect 8350 -1590 8360 -1560
rect 8390 -1590 8400 -1560
rect 8350 -1615 8400 -1590
rect 8350 -1635 8365 -1615
rect 8385 -1635 8400 -1615
rect -50 -1740 -40 -1710
rect -10 -1740 0 -1710
rect -50 -1750 0 -1740
rect 8350 -1710 8400 -1635
rect 9550 -965 9600 -890
rect 9700 -860 9750 -850
rect 9700 -890 9710 -860
rect 9740 -890 9750 -860
rect 9700 -900 9750 -890
rect 10000 -860 10050 -850
rect 10000 -890 10010 -860
rect 10040 -890 10050 -860
rect 10000 -900 10050 -890
rect 10300 -860 10350 -850
rect 10300 -890 10310 -860
rect 10340 -890 10350 -860
rect 10300 -900 10350 -890
rect 10600 -860 10650 -850
rect 10600 -890 10610 -860
rect 10640 -890 10650 -860
rect 10600 -900 10650 -890
rect 9550 -985 9565 -965
rect 9585 -985 9600 -965
rect 9550 -1015 9600 -985
rect 9550 -1035 9565 -1015
rect 9585 -1035 9600 -1015
rect 9550 -1065 9600 -1035
rect 9550 -1085 9565 -1065
rect 9585 -1085 9600 -1065
rect 9550 -1115 9600 -1085
rect 9550 -1135 9565 -1115
rect 9585 -1135 9600 -1115
rect 9550 -1165 9600 -1135
rect 9550 -1185 9565 -1165
rect 9585 -1185 9600 -1165
rect 9550 -1215 9600 -1185
rect 9550 -1235 9565 -1215
rect 9585 -1235 9600 -1215
rect 9550 -1265 9600 -1235
rect 9550 -1285 9565 -1265
rect 9585 -1285 9600 -1265
rect 9550 -1315 9600 -1285
rect 9550 -1335 9565 -1315
rect 9585 -1335 9600 -1315
rect 9550 -1365 9600 -1335
rect 9550 -1385 9565 -1365
rect 9585 -1385 9600 -1365
rect 9550 -1415 9600 -1385
rect 9550 -1435 9565 -1415
rect 9585 -1435 9600 -1415
rect 9550 -1465 9600 -1435
rect 9550 -1485 9565 -1465
rect 9585 -1485 9600 -1465
rect 9550 -1515 9600 -1485
rect 9550 -1535 9565 -1515
rect 9585 -1535 9600 -1515
rect 9550 -1565 9600 -1535
rect 9550 -1585 9565 -1565
rect 9585 -1585 9600 -1565
rect 9550 -1615 9600 -1585
rect 9550 -1635 9565 -1615
rect 9585 -1635 9600 -1615
rect 9550 -1650 9600 -1635
rect 10750 -960 10800 -790
rect 11950 735 12000 915
rect 12250 1485 12300 1500
rect 12250 1465 12265 1485
rect 12285 1465 12300 1485
rect 12250 1435 12300 1465
rect 12250 1415 12265 1435
rect 12285 1415 12300 1435
rect 12250 1385 12300 1415
rect 12250 1365 12265 1385
rect 12285 1365 12300 1385
rect 12250 1335 12300 1365
rect 12250 1315 12265 1335
rect 12285 1315 12300 1335
rect 12250 1285 12300 1315
rect 12250 1265 12265 1285
rect 12285 1265 12300 1285
rect 12250 1235 12300 1265
rect 12250 1215 12265 1235
rect 12285 1215 12300 1235
rect 12250 1185 12300 1215
rect 12250 1165 12265 1185
rect 12285 1165 12300 1185
rect 12250 1135 12300 1165
rect 12250 1115 12265 1135
rect 12285 1115 12300 1135
rect 12250 1085 12300 1115
rect 12250 1065 12265 1085
rect 12285 1065 12300 1085
rect 12250 1035 12300 1065
rect 12250 1015 12265 1035
rect 12285 1015 12300 1035
rect 12250 985 12300 1015
rect 12550 1485 12600 1515
rect 13150 1535 13200 1550
rect 13150 1515 13165 1535
rect 13185 1515 13200 1535
rect 12550 1465 12565 1485
rect 12585 1465 12600 1485
rect 12550 1435 12600 1465
rect 12550 1415 12565 1435
rect 12585 1415 12600 1435
rect 12550 1385 12600 1415
rect 12550 1365 12565 1385
rect 12585 1365 12600 1385
rect 12550 1335 12600 1365
rect 12550 1315 12565 1335
rect 12585 1315 12600 1335
rect 12550 1285 12600 1315
rect 12550 1265 12565 1285
rect 12585 1265 12600 1285
rect 12550 1235 12600 1265
rect 12550 1215 12565 1235
rect 12585 1215 12600 1235
rect 12550 1185 12600 1215
rect 12550 1165 12565 1185
rect 12585 1165 12600 1185
rect 12550 1135 12600 1165
rect 12550 1115 12565 1135
rect 12585 1115 12600 1135
rect 12550 1085 12600 1115
rect 12550 1065 12565 1085
rect 12585 1065 12600 1085
rect 12550 1035 12600 1065
rect 12550 1015 12565 1035
rect 12585 1015 12600 1035
rect 12550 1000 12600 1015
rect 12850 1485 12900 1500
rect 12850 1465 12865 1485
rect 12885 1465 12900 1485
rect 12850 1435 12900 1465
rect 12850 1415 12865 1435
rect 12885 1415 12900 1435
rect 12850 1385 12900 1415
rect 12850 1365 12865 1385
rect 12885 1365 12900 1385
rect 12850 1335 12900 1365
rect 12850 1315 12865 1335
rect 12885 1315 12900 1335
rect 12850 1285 12900 1315
rect 12850 1265 12865 1285
rect 12885 1265 12900 1285
rect 12850 1235 12900 1265
rect 12850 1215 12865 1235
rect 12885 1215 12900 1235
rect 12850 1185 12900 1215
rect 12850 1165 12865 1185
rect 12885 1165 12900 1185
rect 12850 1135 12900 1165
rect 12850 1115 12865 1135
rect 12885 1115 12900 1135
rect 12850 1085 12900 1115
rect 12850 1065 12865 1085
rect 12885 1065 12900 1085
rect 12850 1035 12900 1065
rect 12850 1015 12865 1035
rect 12885 1015 12900 1035
rect 12250 965 12265 985
rect 12285 965 12300 985
rect 12250 950 12300 965
rect 12850 985 12900 1015
rect 12850 965 12865 985
rect 12885 965 12900 985
rect 12850 950 12900 965
rect 12250 935 12900 950
rect 12250 915 12265 935
rect 12285 915 12865 935
rect 12885 915 12900 935
rect 12250 900 12900 915
rect 13150 1485 13200 1515
rect 13750 1535 13800 1550
rect 13750 1515 13765 1535
rect 13785 1515 13800 1535
rect 13150 1465 13165 1485
rect 13185 1465 13200 1485
rect 13150 1435 13200 1465
rect 13150 1415 13165 1435
rect 13185 1415 13200 1435
rect 13150 1385 13200 1415
rect 13150 1365 13165 1385
rect 13185 1365 13200 1385
rect 13150 1335 13200 1365
rect 13150 1315 13165 1335
rect 13185 1315 13200 1335
rect 13150 1285 13200 1315
rect 13150 1265 13165 1285
rect 13185 1265 13200 1285
rect 13150 1235 13200 1265
rect 13150 1215 13165 1235
rect 13185 1215 13200 1235
rect 13150 1185 13200 1215
rect 13150 1165 13165 1185
rect 13185 1165 13200 1185
rect 13150 1135 13200 1165
rect 13150 1115 13165 1135
rect 13185 1115 13200 1135
rect 13150 1085 13200 1115
rect 13150 1065 13165 1085
rect 13185 1065 13200 1085
rect 13150 1035 13200 1065
rect 13150 1015 13165 1035
rect 13185 1015 13200 1035
rect 12100 840 12150 850
rect 12100 810 12110 840
rect 12140 810 12150 840
rect 12100 800 12150 810
rect 12400 840 12450 850
rect 12400 810 12410 840
rect 12440 810 12450 840
rect 12400 800 12450 810
rect 12550 840 12600 900
rect 12550 810 12560 840
rect 12590 810 12600 840
rect 12550 750 12600 810
rect 12700 840 12750 850
rect 12700 810 12710 840
rect 12740 810 12750 840
rect 12700 800 12750 810
rect 13000 840 13050 850
rect 13000 810 13010 840
rect 13040 810 13050 840
rect 13000 800 13050 810
rect 13150 840 13200 1015
rect 13450 1485 13500 1500
rect 13450 1465 13465 1485
rect 13485 1465 13500 1485
rect 13450 1435 13500 1465
rect 13450 1415 13465 1435
rect 13485 1415 13500 1435
rect 13450 1385 13500 1415
rect 13450 1365 13465 1385
rect 13485 1365 13500 1385
rect 13450 1335 13500 1365
rect 13450 1315 13465 1335
rect 13485 1315 13500 1335
rect 13450 1285 13500 1315
rect 13450 1265 13465 1285
rect 13485 1265 13500 1285
rect 13450 1235 13500 1265
rect 13450 1215 13465 1235
rect 13485 1215 13500 1235
rect 13450 1185 13500 1215
rect 13450 1165 13465 1185
rect 13485 1165 13500 1185
rect 13450 1135 13500 1165
rect 13450 1115 13465 1135
rect 13485 1115 13500 1135
rect 13450 1085 13500 1115
rect 13450 1065 13465 1085
rect 13485 1065 13500 1085
rect 13450 1035 13500 1065
rect 13450 1015 13465 1035
rect 13485 1015 13500 1035
rect 13450 985 13500 1015
rect 13750 1485 13800 1515
rect 14350 1535 14400 1550
rect 14350 1515 14365 1535
rect 14385 1515 14400 1535
rect 13750 1465 13765 1485
rect 13785 1465 13800 1485
rect 13750 1435 13800 1465
rect 13750 1415 13765 1435
rect 13785 1415 13800 1435
rect 13750 1385 13800 1415
rect 13750 1365 13765 1385
rect 13785 1365 13800 1385
rect 13750 1335 13800 1365
rect 13750 1315 13765 1335
rect 13785 1315 13800 1335
rect 13750 1285 13800 1315
rect 13750 1265 13765 1285
rect 13785 1265 13800 1285
rect 13750 1235 13800 1265
rect 13750 1215 13765 1235
rect 13785 1215 13800 1235
rect 13750 1185 13800 1215
rect 13750 1165 13765 1185
rect 13785 1165 13800 1185
rect 13750 1135 13800 1165
rect 13750 1115 13765 1135
rect 13785 1115 13800 1135
rect 13750 1085 13800 1115
rect 13750 1065 13765 1085
rect 13785 1065 13800 1085
rect 13750 1035 13800 1065
rect 13750 1015 13765 1035
rect 13785 1015 13800 1035
rect 13750 1000 13800 1015
rect 14050 1485 14100 1500
rect 14050 1465 14065 1485
rect 14085 1465 14100 1485
rect 14050 1435 14100 1465
rect 14050 1415 14065 1435
rect 14085 1415 14100 1435
rect 14050 1385 14100 1415
rect 14050 1365 14065 1385
rect 14085 1365 14100 1385
rect 14050 1335 14100 1365
rect 14050 1315 14065 1335
rect 14085 1315 14100 1335
rect 14050 1285 14100 1315
rect 14050 1265 14065 1285
rect 14085 1265 14100 1285
rect 14050 1235 14100 1265
rect 14050 1215 14065 1235
rect 14085 1215 14100 1235
rect 14050 1185 14100 1215
rect 14050 1165 14065 1185
rect 14085 1165 14100 1185
rect 14050 1135 14100 1165
rect 14050 1115 14065 1135
rect 14085 1115 14100 1135
rect 14050 1085 14100 1115
rect 14050 1065 14065 1085
rect 14085 1065 14100 1085
rect 14050 1035 14100 1065
rect 14050 1015 14065 1035
rect 14085 1015 14100 1035
rect 13450 965 13465 985
rect 13485 965 13500 985
rect 13450 950 13500 965
rect 14050 985 14100 1015
rect 14050 965 14065 985
rect 14085 965 14100 985
rect 14050 950 14100 965
rect 13450 935 14100 950
rect 13450 915 13465 935
rect 13485 915 14065 935
rect 14085 915 14100 935
rect 13450 900 14100 915
rect 14350 1485 14400 1515
rect 14350 1465 14365 1485
rect 14385 1465 14400 1485
rect 14350 1435 14400 1465
rect 14350 1415 14365 1435
rect 14385 1415 14400 1435
rect 14350 1385 14400 1415
rect 14350 1365 14365 1385
rect 14385 1365 14400 1385
rect 14350 1335 14400 1365
rect 14350 1315 14365 1335
rect 14385 1315 14400 1335
rect 14350 1285 14400 1315
rect 14350 1265 14365 1285
rect 14385 1265 14400 1285
rect 14350 1235 14400 1265
rect 14350 1215 14365 1235
rect 14385 1215 14400 1235
rect 14350 1185 14400 1215
rect 14350 1165 14365 1185
rect 14385 1165 14400 1185
rect 14350 1135 14400 1165
rect 14350 1115 14365 1135
rect 14385 1115 14400 1135
rect 14350 1085 14400 1115
rect 14350 1065 14365 1085
rect 14385 1065 14400 1085
rect 14350 1035 14400 1065
rect 14350 1015 14365 1035
rect 14385 1015 14400 1035
rect 14350 985 14400 1015
rect 14350 965 14365 985
rect 14385 965 14400 985
rect 14350 935 14400 965
rect 14350 915 14365 935
rect 14385 915 14400 935
rect 13150 810 13160 840
rect 13190 810 13200 840
rect 11950 715 11965 735
rect 11985 715 12000 735
rect 11950 685 12000 715
rect 11950 665 11965 685
rect 11985 665 12000 685
rect 11950 635 12000 665
rect 11950 615 11965 635
rect 11985 615 12000 635
rect 11950 585 12000 615
rect 11950 565 11965 585
rect 11985 565 12000 585
rect 11950 535 12000 565
rect 11950 515 11965 535
rect 11985 515 12000 535
rect 11950 485 12000 515
rect 11950 465 11965 485
rect 11985 465 12000 485
rect 11950 435 12000 465
rect 11950 415 11965 435
rect 11985 415 12000 435
rect 11950 385 12000 415
rect 11950 365 11965 385
rect 11985 365 12000 385
rect 11950 335 12000 365
rect 11950 315 11965 335
rect 11985 315 12000 335
rect 11950 285 12000 315
rect 11950 265 11965 285
rect 11985 265 12000 285
rect 11950 235 12000 265
rect 11950 215 11965 235
rect 11985 215 12000 235
rect 11950 185 12000 215
rect 11950 165 11965 185
rect 11985 165 12000 185
rect 11950 135 12000 165
rect 12250 735 12900 750
rect 12250 715 12265 735
rect 12285 715 12865 735
rect 12885 715 12900 735
rect 12250 700 12900 715
rect 12250 685 12300 700
rect 12250 665 12265 685
rect 12285 665 12300 685
rect 12250 635 12300 665
rect 12850 685 12900 700
rect 12850 665 12865 685
rect 12885 665 12900 685
rect 12250 615 12265 635
rect 12285 615 12300 635
rect 12250 585 12300 615
rect 12250 565 12265 585
rect 12285 565 12300 585
rect 12250 535 12300 565
rect 12250 515 12265 535
rect 12285 515 12300 535
rect 12250 485 12300 515
rect 12250 465 12265 485
rect 12285 465 12300 485
rect 12250 435 12300 465
rect 12250 415 12265 435
rect 12285 415 12300 435
rect 12250 385 12300 415
rect 12250 365 12265 385
rect 12285 365 12300 385
rect 12250 335 12300 365
rect 12250 315 12265 335
rect 12285 315 12300 335
rect 12250 285 12300 315
rect 12250 265 12265 285
rect 12285 265 12300 285
rect 12250 235 12300 265
rect 12250 215 12265 235
rect 12285 215 12300 235
rect 12250 185 12300 215
rect 12250 165 12265 185
rect 12285 165 12300 185
rect 12250 150 12300 165
rect 12550 635 12600 650
rect 12550 615 12565 635
rect 12585 615 12600 635
rect 12550 585 12600 615
rect 12550 565 12565 585
rect 12585 565 12600 585
rect 12550 535 12600 565
rect 12550 515 12565 535
rect 12585 515 12600 535
rect 12550 485 12600 515
rect 12550 465 12565 485
rect 12585 465 12600 485
rect 12550 435 12600 465
rect 12550 415 12565 435
rect 12585 415 12600 435
rect 12550 385 12600 415
rect 12550 365 12565 385
rect 12585 365 12600 385
rect 12550 335 12600 365
rect 12550 315 12565 335
rect 12585 315 12600 335
rect 12550 285 12600 315
rect 12550 265 12565 285
rect 12585 265 12600 285
rect 12550 235 12600 265
rect 12550 215 12565 235
rect 12585 215 12600 235
rect 12550 185 12600 215
rect 12550 165 12565 185
rect 12585 165 12600 185
rect 11950 115 11965 135
rect 11985 115 12000 135
rect 11950 100 12000 115
rect 12550 135 12600 165
rect 12850 635 12900 665
rect 12850 615 12865 635
rect 12885 615 12900 635
rect 12850 585 12900 615
rect 12850 565 12865 585
rect 12885 565 12900 585
rect 12850 535 12900 565
rect 12850 515 12865 535
rect 12885 515 12900 535
rect 12850 485 12900 515
rect 12850 465 12865 485
rect 12885 465 12900 485
rect 12850 435 12900 465
rect 12850 415 12865 435
rect 12885 415 12900 435
rect 12850 385 12900 415
rect 12850 365 12865 385
rect 12885 365 12900 385
rect 12850 335 12900 365
rect 12850 315 12865 335
rect 12885 315 12900 335
rect 12850 285 12900 315
rect 12850 265 12865 285
rect 12885 265 12900 285
rect 12850 235 12900 265
rect 12850 215 12865 235
rect 12885 215 12900 235
rect 12850 185 12900 215
rect 12850 165 12865 185
rect 12885 165 12900 185
rect 12850 150 12900 165
rect 13150 635 13200 810
rect 13300 840 13350 850
rect 13300 810 13310 840
rect 13340 810 13350 840
rect 13300 800 13350 810
rect 13600 840 13650 850
rect 13600 810 13610 840
rect 13640 810 13650 840
rect 13600 800 13650 810
rect 13750 840 13800 900
rect 13750 810 13760 840
rect 13790 810 13800 840
rect 13750 750 13800 810
rect 13900 840 13950 850
rect 13900 810 13910 840
rect 13940 810 13950 840
rect 13900 800 13950 810
rect 14200 840 14250 850
rect 14200 810 14210 840
rect 14240 810 14250 840
rect 14200 800 14250 810
rect 13150 615 13165 635
rect 13185 615 13200 635
rect 13150 585 13200 615
rect 13150 565 13165 585
rect 13185 565 13200 585
rect 13150 535 13200 565
rect 13150 515 13165 535
rect 13185 515 13200 535
rect 13150 485 13200 515
rect 13150 465 13165 485
rect 13185 465 13200 485
rect 13150 435 13200 465
rect 13150 415 13165 435
rect 13185 415 13200 435
rect 13150 385 13200 415
rect 13150 365 13165 385
rect 13185 365 13200 385
rect 13150 335 13200 365
rect 13150 315 13165 335
rect 13185 315 13200 335
rect 13150 285 13200 315
rect 13150 265 13165 285
rect 13185 265 13200 285
rect 13150 235 13200 265
rect 13150 215 13165 235
rect 13185 215 13200 235
rect 13150 185 13200 215
rect 13150 165 13165 185
rect 13185 165 13200 185
rect 12550 115 12565 135
rect 12585 115 12600 135
rect 12550 100 12600 115
rect 13150 135 13200 165
rect 13450 735 14100 750
rect 13450 715 13465 735
rect 13485 715 14065 735
rect 14085 715 14100 735
rect 13450 700 14100 715
rect 13450 685 13500 700
rect 13450 665 13465 685
rect 13485 665 13500 685
rect 13450 635 13500 665
rect 14050 685 14100 700
rect 14050 665 14065 685
rect 14085 665 14100 685
rect 13450 615 13465 635
rect 13485 615 13500 635
rect 13450 585 13500 615
rect 13450 565 13465 585
rect 13485 565 13500 585
rect 13450 535 13500 565
rect 13450 515 13465 535
rect 13485 515 13500 535
rect 13450 485 13500 515
rect 13450 465 13465 485
rect 13485 465 13500 485
rect 13450 435 13500 465
rect 13450 415 13465 435
rect 13485 415 13500 435
rect 13450 385 13500 415
rect 13450 365 13465 385
rect 13485 365 13500 385
rect 13450 335 13500 365
rect 13450 315 13465 335
rect 13485 315 13500 335
rect 13450 285 13500 315
rect 13450 265 13465 285
rect 13485 265 13500 285
rect 13450 235 13500 265
rect 13450 215 13465 235
rect 13485 215 13500 235
rect 13450 185 13500 215
rect 13450 165 13465 185
rect 13485 165 13500 185
rect 13450 150 13500 165
rect 13750 635 13800 650
rect 13750 615 13765 635
rect 13785 615 13800 635
rect 13750 585 13800 615
rect 13750 565 13765 585
rect 13785 565 13800 585
rect 13750 535 13800 565
rect 13750 515 13765 535
rect 13785 515 13800 535
rect 13750 485 13800 515
rect 13750 465 13765 485
rect 13785 465 13800 485
rect 13750 435 13800 465
rect 13750 415 13765 435
rect 13785 415 13800 435
rect 13750 385 13800 415
rect 13750 365 13765 385
rect 13785 365 13800 385
rect 13750 335 13800 365
rect 13750 315 13765 335
rect 13785 315 13800 335
rect 13750 285 13800 315
rect 13750 265 13765 285
rect 13785 265 13800 285
rect 13750 235 13800 265
rect 13750 215 13765 235
rect 13785 215 13800 235
rect 13750 185 13800 215
rect 13750 165 13765 185
rect 13785 165 13800 185
rect 13150 115 13165 135
rect 13185 115 13200 135
rect 13150 100 13200 115
rect 13750 135 13800 165
rect 14050 635 14100 665
rect 14050 615 14065 635
rect 14085 615 14100 635
rect 14050 585 14100 615
rect 14050 565 14065 585
rect 14085 565 14100 585
rect 14050 535 14100 565
rect 14050 515 14065 535
rect 14085 515 14100 535
rect 14050 485 14100 515
rect 14050 465 14065 485
rect 14085 465 14100 485
rect 14050 435 14100 465
rect 14050 415 14065 435
rect 14085 415 14100 435
rect 14050 385 14100 415
rect 14050 365 14065 385
rect 14085 365 14100 385
rect 14050 335 14100 365
rect 14050 315 14065 335
rect 14085 315 14100 335
rect 14050 285 14100 315
rect 14050 265 14065 285
rect 14085 265 14100 285
rect 14050 235 14100 265
rect 14050 215 14065 235
rect 14085 215 14100 235
rect 14050 185 14100 215
rect 14050 165 14065 185
rect 14085 165 14100 185
rect 14050 150 14100 165
rect 14350 735 14400 915
rect 15550 1585 15600 1660
rect 17950 1690 18000 1700
rect 17950 1660 17960 1690
rect 17990 1660 18000 1690
rect 15550 1565 15565 1585
rect 15585 1565 15600 1585
rect 15550 1540 15600 1565
rect 15550 1510 15560 1540
rect 15590 1510 15600 1540
rect 15550 1485 15600 1510
rect 15550 1465 15565 1485
rect 15585 1465 15600 1485
rect 15550 1440 15600 1465
rect 15550 1410 15560 1440
rect 15590 1410 15600 1440
rect 15550 1385 15600 1410
rect 15550 1365 15565 1385
rect 15585 1365 15600 1385
rect 15550 1340 15600 1365
rect 15550 1310 15560 1340
rect 15590 1310 15600 1340
rect 15550 1285 15600 1310
rect 15550 1265 15565 1285
rect 15585 1265 15600 1285
rect 15550 1240 15600 1265
rect 15550 1210 15560 1240
rect 15590 1210 15600 1240
rect 15550 1185 15600 1210
rect 15550 1165 15565 1185
rect 15585 1165 15600 1185
rect 15550 1140 15600 1165
rect 15550 1110 15560 1140
rect 15590 1110 15600 1140
rect 15550 1085 15600 1110
rect 15550 1065 15565 1085
rect 15585 1065 15600 1085
rect 15550 1040 15600 1065
rect 15550 1010 15560 1040
rect 15590 1010 15600 1040
rect 15550 985 15600 1010
rect 15550 965 15565 985
rect 15585 965 15600 985
rect 15550 940 15600 965
rect 15550 910 15560 940
rect 15590 910 15600 940
rect 14500 840 14550 850
rect 14500 810 14510 840
rect 14540 810 14550 840
rect 14500 800 14550 810
rect 14800 840 14850 850
rect 14800 810 14810 840
rect 14840 810 14850 840
rect 14800 800 14850 810
rect 15100 840 15150 850
rect 15100 810 15110 840
rect 15140 810 15150 840
rect 15100 800 15150 810
rect 15400 840 15450 850
rect 15400 810 15410 840
rect 15440 810 15450 840
rect 15400 800 15450 810
rect 14350 715 14365 735
rect 14385 715 14400 735
rect 14350 685 14400 715
rect 14350 665 14365 685
rect 14385 665 14400 685
rect 14350 635 14400 665
rect 14350 615 14365 635
rect 14385 615 14400 635
rect 14350 585 14400 615
rect 14350 565 14365 585
rect 14385 565 14400 585
rect 14350 535 14400 565
rect 14350 515 14365 535
rect 14385 515 14400 535
rect 14350 485 14400 515
rect 14350 465 14365 485
rect 14385 465 14400 485
rect 14350 435 14400 465
rect 14350 415 14365 435
rect 14385 415 14400 435
rect 14350 385 14400 415
rect 14350 365 14365 385
rect 14385 365 14400 385
rect 14350 335 14400 365
rect 14350 315 14365 335
rect 14385 315 14400 335
rect 14350 285 14400 315
rect 14350 265 14365 285
rect 14385 265 14400 285
rect 14350 235 14400 265
rect 14350 215 14365 235
rect 14385 215 14400 235
rect 14350 185 14400 215
rect 14350 165 14365 185
rect 14385 165 14400 185
rect 13750 115 13765 135
rect 13785 115 13800 135
rect 13750 100 13800 115
rect 14350 135 14400 165
rect 14350 115 14365 135
rect 14385 115 14400 135
rect 14350 100 14400 115
rect 11950 85 14400 100
rect 11950 65 11965 85
rect 11985 65 12565 85
rect 12585 65 13165 85
rect 13185 65 13765 85
rect 13785 65 14365 85
rect 14385 65 14400 85
rect 11950 50 14400 65
rect 11950 -100 12000 50
rect 13150 -100 13200 50
rect 14350 -100 14400 50
rect 11950 -115 14400 -100
rect 11950 -135 11965 -115
rect 11985 -135 12565 -115
rect 12585 -135 13165 -115
rect 13185 -135 13765 -115
rect 13785 -135 14365 -115
rect 14385 -135 14400 -115
rect 11950 -150 14400 -135
rect 11950 -165 12000 -150
rect 11950 -185 11965 -165
rect 11985 -185 12000 -165
rect 11950 -215 12000 -185
rect 12550 -165 12600 -150
rect 12550 -185 12565 -165
rect 12585 -185 12600 -165
rect 11950 -235 11965 -215
rect 11985 -235 12000 -215
rect 11950 -265 12000 -235
rect 11950 -285 11965 -265
rect 11985 -285 12000 -265
rect 11950 -315 12000 -285
rect 11950 -335 11965 -315
rect 11985 -335 12000 -315
rect 11950 -365 12000 -335
rect 11950 -385 11965 -365
rect 11985 -385 12000 -365
rect 11950 -415 12000 -385
rect 11950 -435 11965 -415
rect 11985 -435 12000 -415
rect 11950 -465 12000 -435
rect 11950 -485 11965 -465
rect 11985 -485 12000 -465
rect 11950 -515 12000 -485
rect 11950 -535 11965 -515
rect 11985 -535 12000 -515
rect 11950 -565 12000 -535
rect 11950 -585 11965 -565
rect 11985 -585 12000 -565
rect 11950 -615 12000 -585
rect 11950 -635 11965 -615
rect 11985 -635 12000 -615
rect 11950 -665 12000 -635
rect 11950 -685 11965 -665
rect 11985 -685 12000 -665
rect 11950 -715 12000 -685
rect 11950 -735 11965 -715
rect 11985 -735 12000 -715
rect 11950 -765 12000 -735
rect 11950 -785 11965 -765
rect 11985 -785 12000 -765
rect 10900 -860 10950 -850
rect 10900 -890 10910 -860
rect 10940 -890 10950 -860
rect 10900 -900 10950 -890
rect 11200 -860 11250 -850
rect 11200 -890 11210 -860
rect 11240 -890 11250 -860
rect 11200 -900 11250 -890
rect 11500 -860 11550 -850
rect 11500 -890 11510 -860
rect 11540 -890 11550 -860
rect 11500 -900 11550 -890
rect 11800 -860 11850 -850
rect 11800 -890 11810 -860
rect 11840 -890 11850 -860
rect 11800 -900 11850 -890
rect 10750 -990 10760 -960
rect 10790 -990 10800 -960
rect 10750 -1015 10800 -990
rect 10750 -1035 10765 -1015
rect 10785 -1035 10800 -1015
rect 10750 -1060 10800 -1035
rect 10750 -1090 10760 -1060
rect 10790 -1090 10800 -1060
rect 10750 -1115 10800 -1090
rect 10750 -1135 10765 -1115
rect 10785 -1135 10800 -1115
rect 10750 -1160 10800 -1135
rect 10750 -1190 10760 -1160
rect 10790 -1190 10800 -1160
rect 10750 -1215 10800 -1190
rect 10750 -1235 10765 -1215
rect 10785 -1235 10800 -1215
rect 10750 -1260 10800 -1235
rect 10750 -1290 10760 -1260
rect 10790 -1290 10800 -1260
rect 10750 -1315 10800 -1290
rect 10750 -1335 10765 -1315
rect 10785 -1335 10800 -1315
rect 10750 -1360 10800 -1335
rect 10750 -1390 10760 -1360
rect 10790 -1390 10800 -1360
rect 10750 -1415 10800 -1390
rect 10750 -1435 10765 -1415
rect 10785 -1435 10800 -1415
rect 10750 -1460 10800 -1435
rect 10750 -1490 10760 -1460
rect 10790 -1490 10800 -1460
rect 10750 -1515 10800 -1490
rect 10750 -1535 10765 -1515
rect 10785 -1535 10800 -1515
rect 10750 -1560 10800 -1535
rect 10750 -1590 10760 -1560
rect 10790 -1590 10800 -1560
rect 10750 -1615 10800 -1590
rect 10750 -1635 10765 -1615
rect 10785 -1635 10800 -1615
rect 8350 -1740 8360 -1710
rect 8390 -1740 8400 -1710
rect 8350 -1750 8400 -1740
rect 10750 -1710 10800 -1635
rect 11950 -965 12000 -785
rect 12250 -215 12300 -200
rect 12250 -235 12265 -215
rect 12285 -235 12300 -215
rect 12250 -265 12300 -235
rect 12250 -285 12265 -265
rect 12285 -285 12300 -265
rect 12250 -315 12300 -285
rect 12250 -335 12265 -315
rect 12285 -335 12300 -315
rect 12250 -365 12300 -335
rect 12250 -385 12265 -365
rect 12285 -385 12300 -365
rect 12250 -415 12300 -385
rect 12250 -435 12265 -415
rect 12285 -435 12300 -415
rect 12250 -465 12300 -435
rect 12250 -485 12265 -465
rect 12285 -485 12300 -465
rect 12250 -515 12300 -485
rect 12250 -535 12265 -515
rect 12285 -535 12300 -515
rect 12250 -565 12300 -535
rect 12250 -585 12265 -565
rect 12285 -585 12300 -565
rect 12250 -615 12300 -585
rect 12250 -635 12265 -615
rect 12285 -635 12300 -615
rect 12250 -665 12300 -635
rect 12250 -685 12265 -665
rect 12285 -685 12300 -665
rect 12250 -715 12300 -685
rect 12550 -215 12600 -185
rect 13150 -165 13200 -150
rect 13150 -185 13165 -165
rect 13185 -185 13200 -165
rect 12550 -235 12565 -215
rect 12585 -235 12600 -215
rect 12550 -265 12600 -235
rect 12550 -285 12565 -265
rect 12585 -285 12600 -265
rect 12550 -315 12600 -285
rect 12550 -335 12565 -315
rect 12585 -335 12600 -315
rect 12550 -365 12600 -335
rect 12550 -385 12565 -365
rect 12585 -385 12600 -365
rect 12550 -415 12600 -385
rect 12550 -435 12565 -415
rect 12585 -435 12600 -415
rect 12550 -465 12600 -435
rect 12550 -485 12565 -465
rect 12585 -485 12600 -465
rect 12550 -515 12600 -485
rect 12550 -535 12565 -515
rect 12585 -535 12600 -515
rect 12550 -565 12600 -535
rect 12550 -585 12565 -565
rect 12585 -585 12600 -565
rect 12550 -615 12600 -585
rect 12550 -635 12565 -615
rect 12585 -635 12600 -615
rect 12550 -665 12600 -635
rect 12550 -685 12565 -665
rect 12585 -685 12600 -665
rect 12550 -700 12600 -685
rect 12850 -215 12900 -200
rect 12850 -235 12865 -215
rect 12885 -235 12900 -215
rect 12850 -265 12900 -235
rect 12850 -285 12865 -265
rect 12885 -285 12900 -265
rect 12850 -315 12900 -285
rect 12850 -335 12865 -315
rect 12885 -335 12900 -315
rect 12850 -365 12900 -335
rect 12850 -385 12865 -365
rect 12885 -385 12900 -365
rect 12850 -415 12900 -385
rect 12850 -435 12865 -415
rect 12885 -435 12900 -415
rect 12850 -465 12900 -435
rect 12850 -485 12865 -465
rect 12885 -485 12900 -465
rect 12850 -515 12900 -485
rect 12850 -535 12865 -515
rect 12885 -535 12900 -515
rect 12850 -565 12900 -535
rect 12850 -585 12865 -565
rect 12885 -585 12900 -565
rect 12850 -615 12900 -585
rect 12850 -635 12865 -615
rect 12885 -635 12900 -615
rect 12850 -665 12900 -635
rect 12850 -685 12865 -665
rect 12885 -685 12900 -665
rect 12250 -735 12265 -715
rect 12285 -735 12300 -715
rect 12250 -750 12300 -735
rect 12850 -715 12900 -685
rect 12850 -735 12865 -715
rect 12885 -735 12900 -715
rect 12850 -750 12900 -735
rect 12250 -765 12900 -750
rect 12250 -785 12265 -765
rect 12285 -785 12865 -765
rect 12885 -785 12900 -765
rect 12250 -800 12900 -785
rect 13150 -215 13200 -185
rect 13750 -165 13800 -150
rect 13750 -185 13765 -165
rect 13785 -185 13800 -165
rect 13150 -235 13165 -215
rect 13185 -235 13200 -215
rect 13150 -265 13200 -235
rect 13150 -285 13165 -265
rect 13185 -285 13200 -265
rect 13150 -315 13200 -285
rect 13150 -335 13165 -315
rect 13185 -335 13200 -315
rect 13150 -365 13200 -335
rect 13150 -385 13165 -365
rect 13185 -385 13200 -365
rect 13150 -415 13200 -385
rect 13150 -435 13165 -415
rect 13185 -435 13200 -415
rect 13150 -465 13200 -435
rect 13150 -485 13165 -465
rect 13185 -485 13200 -465
rect 13150 -515 13200 -485
rect 13150 -535 13165 -515
rect 13185 -535 13200 -515
rect 13150 -565 13200 -535
rect 13150 -585 13165 -565
rect 13185 -585 13200 -565
rect 13150 -615 13200 -585
rect 13150 -635 13165 -615
rect 13185 -635 13200 -615
rect 13150 -665 13200 -635
rect 13150 -685 13165 -665
rect 13185 -685 13200 -665
rect 12100 -860 12150 -850
rect 12100 -890 12110 -860
rect 12140 -890 12150 -860
rect 12100 -900 12150 -890
rect 12400 -860 12450 -850
rect 12400 -890 12410 -860
rect 12440 -890 12450 -860
rect 12400 -900 12450 -890
rect 12550 -860 12600 -800
rect 12550 -890 12560 -860
rect 12590 -890 12600 -860
rect 12550 -950 12600 -890
rect 12700 -860 12750 -850
rect 12700 -890 12710 -860
rect 12740 -890 12750 -860
rect 12700 -900 12750 -890
rect 13000 -860 13050 -850
rect 13000 -890 13010 -860
rect 13040 -890 13050 -860
rect 13000 -900 13050 -890
rect 13150 -860 13200 -685
rect 13450 -215 13500 -200
rect 13450 -235 13465 -215
rect 13485 -235 13500 -215
rect 13450 -265 13500 -235
rect 13450 -285 13465 -265
rect 13485 -285 13500 -265
rect 13450 -315 13500 -285
rect 13450 -335 13465 -315
rect 13485 -335 13500 -315
rect 13450 -365 13500 -335
rect 13450 -385 13465 -365
rect 13485 -385 13500 -365
rect 13450 -415 13500 -385
rect 13450 -435 13465 -415
rect 13485 -435 13500 -415
rect 13450 -465 13500 -435
rect 13450 -485 13465 -465
rect 13485 -485 13500 -465
rect 13450 -515 13500 -485
rect 13450 -535 13465 -515
rect 13485 -535 13500 -515
rect 13450 -565 13500 -535
rect 13450 -585 13465 -565
rect 13485 -585 13500 -565
rect 13450 -615 13500 -585
rect 13450 -635 13465 -615
rect 13485 -635 13500 -615
rect 13450 -665 13500 -635
rect 13450 -685 13465 -665
rect 13485 -685 13500 -665
rect 13450 -715 13500 -685
rect 13750 -215 13800 -185
rect 14350 -165 14400 -150
rect 14350 -185 14365 -165
rect 14385 -185 14400 -165
rect 13750 -235 13765 -215
rect 13785 -235 13800 -215
rect 13750 -265 13800 -235
rect 13750 -285 13765 -265
rect 13785 -285 13800 -265
rect 13750 -315 13800 -285
rect 13750 -335 13765 -315
rect 13785 -335 13800 -315
rect 13750 -365 13800 -335
rect 13750 -385 13765 -365
rect 13785 -385 13800 -365
rect 13750 -415 13800 -385
rect 13750 -435 13765 -415
rect 13785 -435 13800 -415
rect 13750 -465 13800 -435
rect 13750 -485 13765 -465
rect 13785 -485 13800 -465
rect 13750 -515 13800 -485
rect 13750 -535 13765 -515
rect 13785 -535 13800 -515
rect 13750 -565 13800 -535
rect 13750 -585 13765 -565
rect 13785 -585 13800 -565
rect 13750 -615 13800 -585
rect 13750 -635 13765 -615
rect 13785 -635 13800 -615
rect 13750 -665 13800 -635
rect 13750 -685 13765 -665
rect 13785 -685 13800 -665
rect 13750 -700 13800 -685
rect 14050 -215 14100 -200
rect 14050 -235 14065 -215
rect 14085 -235 14100 -215
rect 14050 -265 14100 -235
rect 14050 -285 14065 -265
rect 14085 -285 14100 -265
rect 14050 -315 14100 -285
rect 14050 -335 14065 -315
rect 14085 -335 14100 -315
rect 14050 -365 14100 -335
rect 14050 -385 14065 -365
rect 14085 -385 14100 -365
rect 14050 -415 14100 -385
rect 14050 -435 14065 -415
rect 14085 -435 14100 -415
rect 14050 -465 14100 -435
rect 14050 -485 14065 -465
rect 14085 -485 14100 -465
rect 14050 -515 14100 -485
rect 14050 -535 14065 -515
rect 14085 -535 14100 -515
rect 14050 -565 14100 -535
rect 14050 -585 14065 -565
rect 14085 -585 14100 -565
rect 14050 -615 14100 -585
rect 14050 -635 14065 -615
rect 14085 -635 14100 -615
rect 14050 -665 14100 -635
rect 14050 -685 14065 -665
rect 14085 -685 14100 -665
rect 13450 -735 13465 -715
rect 13485 -735 13500 -715
rect 13450 -750 13500 -735
rect 14050 -715 14100 -685
rect 14050 -735 14065 -715
rect 14085 -735 14100 -715
rect 14050 -750 14100 -735
rect 13450 -765 14100 -750
rect 13450 -785 13465 -765
rect 13485 -785 14065 -765
rect 14085 -785 14100 -765
rect 13450 -800 14100 -785
rect 14350 -215 14400 -185
rect 14350 -235 14365 -215
rect 14385 -235 14400 -215
rect 14350 -265 14400 -235
rect 14350 -285 14365 -265
rect 14385 -285 14400 -265
rect 14350 -315 14400 -285
rect 14350 -335 14365 -315
rect 14385 -335 14400 -315
rect 14350 -365 14400 -335
rect 14350 -385 14365 -365
rect 14385 -385 14400 -365
rect 14350 -415 14400 -385
rect 14350 -435 14365 -415
rect 14385 -435 14400 -415
rect 14350 -465 14400 -435
rect 14350 -485 14365 -465
rect 14385 -485 14400 -465
rect 14350 -515 14400 -485
rect 14350 -535 14365 -515
rect 14385 -535 14400 -515
rect 14350 -565 14400 -535
rect 14350 -585 14365 -565
rect 14385 -585 14400 -565
rect 14350 -615 14400 -585
rect 14350 -635 14365 -615
rect 14385 -635 14400 -615
rect 14350 -665 14400 -635
rect 14350 -685 14365 -665
rect 14385 -685 14400 -665
rect 14350 -715 14400 -685
rect 14350 -735 14365 -715
rect 14385 -735 14400 -715
rect 14350 -765 14400 -735
rect 14350 -785 14365 -765
rect 14385 -785 14400 -765
rect 13150 -890 13160 -860
rect 13190 -890 13200 -860
rect 11950 -985 11965 -965
rect 11985 -985 12000 -965
rect 11950 -1015 12000 -985
rect 11950 -1035 11965 -1015
rect 11985 -1035 12000 -1015
rect 11950 -1065 12000 -1035
rect 11950 -1085 11965 -1065
rect 11985 -1085 12000 -1065
rect 11950 -1115 12000 -1085
rect 11950 -1135 11965 -1115
rect 11985 -1135 12000 -1115
rect 11950 -1165 12000 -1135
rect 11950 -1185 11965 -1165
rect 11985 -1185 12000 -1165
rect 11950 -1215 12000 -1185
rect 11950 -1235 11965 -1215
rect 11985 -1235 12000 -1215
rect 11950 -1265 12000 -1235
rect 11950 -1285 11965 -1265
rect 11985 -1285 12000 -1265
rect 11950 -1315 12000 -1285
rect 11950 -1335 11965 -1315
rect 11985 -1335 12000 -1315
rect 11950 -1365 12000 -1335
rect 11950 -1385 11965 -1365
rect 11985 -1385 12000 -1365
rect 11950 -1415 12000 -1385
rect 11950 -1435 11965 -1415
rect 11985 -1435 12000 -1415
rect 11950 -1465 12000 -1435
rect 11950 -1485 11965 -1465
rect 11985 -1485 12000 -1465
rect 11950 -1515 12000 -1485
rect 11950 -1535 11965 -1515
rect 11985 -1535 12000 -1515
rect 11950 -1565 12000 -1535
rect 12250 -965 12900 -950
rect 12250 -985 12265 -965
rect 12285 -985 12865 -965
rect 12885 -985 12900 -965
rect 12250 -1000 12900 -985
rect 12250 -1015 12300 -1000
rect 12250 -1035 12265 -1015
rect 12285 -1035 12300 -1015
rect 12250 -1065 12300 -1035
rect 12850 -1015 12900 -1000
rect 12850 -1035 12865 -1015
rect 12885 -1035 12900 -1015
rect 12250 -1085 12265 -1065
rect 12285 -1085 12300 -1065
rect 12250 -1115 12300 -1085
rect 12250 -1135 12265 -1115
rect 12285 -1135 12300 -1115
rect 12250 -1165 12300 -1135
rect 12250 -1185 12265 -1165
rect 12285 -1185 12300 -1165
rect 12250 -1215 12300 -1185
rect 12250 -1235 12265 -1215
rect 12285 -1235 12300 -1215
rect 12250 -1265 12300 -1235
rect 12250 -1285 12265 -1265
rect 12285 -1285 12300 -1265
rect 12250 -1315 12300 -1285
rect 12250 -1335 12265 -1315
rect 12285 -1335 12300 -1315
rect 12250 -1365 12300 -1335
rect 12250 -1385 12265 -1365
rect 12285 -1385 12300 -1365
rect 12250 -1415 12300 -1385
rect 12250 -1435 12265 -1415
rect 12285 -1435 12300 -1415
rect 12250 -1465 12300 -1435
rect 12250 -1485 12265 -1465
rect 12285 -1485 12300 -1465
rect 12250 -1515 12300 -1485
rect 12250 -1535 12265 -1515
rect 12285 -1535 12300 -1515
rect 12250 -1550 12300 -1535
rect 12550 -1065 12600 -1050
rect 12550 -1085 12565 -1065
rect 12585 -1085 12600 -1065
rect 12550 -1115 12600 -1085
rect 12550 -1135 12565 -1115
rect 12585 -1135 12600 -1115
rect 12550 -1165 12600 -1135
rect 12550 -1185 12565 -1165
rect 12585 -1185 12600 -1165
rect 12550 -1215 12600 -1185
rect 12550 -1235 12565 -1215
rect 12585 -1235 12600 -1215
rect 12550 -1265 12600 -1235
rect 12550 -1285 12565 -1265
rect 12585 -1285 12600 -1265
rect 12550 -1315 12600 -1285
rect 12550 -1335 12565 -1315
rect 12585 -1335 12600 -1315
rect 12550 -1365 12600 -1335
rect 12550 -1385 12565 -1365
rect 12585 -1385 12600 -1365
rect 12550 -1415 12600 -1385
rect 12550 -1435 12565 -1415
rect 12585 -1435 12600 -1415
rect 12550 -1465 12600 -1435
rect 12550 -1485 12565 -1465
rect 12585 -1485 12600 -1465
rect 12550 -1515 12600 -1485
rect 12550 -1535 12565 -1515
rect 12585 -1535 12600 -1515
rect 11950 -1585 11965 -1565
rect 11985 -1585 12000 -1565
rect 11950 -1600 12000 -1585
rect 12550 -1565 12600 -1535
rect 12850 -1065 12900 -1035
rect 12850 -1085 12865 -1065
rect 12885 -1085 12900 -1065
rect 12850 -1115 12900 -1085
rect 12850 -1135 12865 -1115
rect 12885 -1135 12900 -1115
rect 12850 -1165 12900 -1135
rect 12850 -1185 12865 -1165
rect 12885 -1185 12900 -1165
rect 12850 -1215 12900 -1185
rect 12850 -1235 12865 -1215
rect 12885 -1235 12900 -1215
rect 12850 -1265 12900 -1235
rect 12850 -1285 12865 -1265
rect 12885 -1285 12900 -1265
rect 12850 -1315 12900 -1285
rect 12850 -1335 12865 -1315
rect 12885 -1335 12900 -1315
rect 12850 -1365 12900 -1335
rect 12850 -1385 12865 -1365
rect 12885 -1385 12900 -1365
rect 12850 -1415 12900 -1385
rect 12850 -1435 12865 -1415
rect 12885 -1435 12900 -1415
rect 12850 -1465 12900 -1435
rect 12850 -1485 12865 -1465
rect 12885 -1485 12900 -1465
rect 12850 -1515 12900 -1485
rect 12850 -1535 12865 -1515
rect 12885 -1535 12900 -1515
rect 12850 -1550 12900 -1535
rect 13150 -1065 13200 -890
rect 13300 -860 13350 -850
rect 13300 -890 13310 -860
rect 13340 -890 13350 -860
rect 13300 -900 13350 -890
rect 13600 -860 13650 -850
rect 13600 -890 13610 -860
rect 13640 -890 13650 -860
rect 13600 -900 13650 -890
rect 13750 -860 13800 -800
rect 13750 -890 13760 -860
rect 13790 -890 13800 -860
rect 13750 -950 13800 -890
rect 13900 -860 13950 -850
rect 13900 -890 13910 -860
rect 13940 -890 13950 -860
rect 13900 -900 13950 -890
rect 14200 -860 14250 -850
rect 14200 -890 14210 -860
rect 14240 -890 14250 -860
rect 14200 -900 14250 -890
rect 13150 -1085 13165 -1065
rect 13185 -1085 13200 -1065
rect 13150 -1115 13200 -1085
rect 13150 -1135 13165 -1115
rect 13185 -1135 13200 -1115
rect 13150 -1165 13200 -1135
rect 13150 -1185 13165 -1165
rect 13185 -1185 13200 -1165
rect 13150 -1215 13200 -1185
rect 13150 -1235 13165 -1215
rect 13185 -1235 13200 -1215
rect 13150 -1265 13200 -1235
rect 13150 -1285 13165 -1265
rect 13185 -1285 13200 -1265
rect 13150 -1315 13200 -1285
rect 13150 -1335 13165 -1315
rect 13185 -1335 13200 -1315
rect 13150 -1365 13200 -1335
rect 13150 -1385 13165 -1365
rect 13185 -1385 13200 -1365
rect 13150 -1415 13200 -1385
rect 13150 -1435 13165 -1415
rect 13185 -1435 13200 -1415
rect 13150 -1465 13200 -1435
rect 13150 -1485 13165 -1465
rect 13185 -1485 13200 -1465
rect 13150 -1515 13200 -1485
rect 13150 -1535 13165 -1515
rect 13185 -1535 13200 -1515
rect 12550 -1585 12565 -1565
rect 12585 -1585 12600 -1565
rect 12550 -1600 12600 -1585
rect 13150 -1565 13200 -1535
rect 13450 -965 14100 -950
rect 13450 -985 13465 -965
rect 13485 -985 14065 -965
rect 14085 -985 14100 -965
rect 13450 -1000 14100 -985
rect 13450 -1015 13500 -1000
rect 13450 -1035 13465 -1015
rect 13485 -1035 13500 -1015
rect 13450 -1065 13500 -1035
rect 14050 -1015 14100 -1000
rect 14050 -1035 14065 -1015
rect 14085 -1035 14100 -1015
rect 13450 -1085 13465 -1065
rect 13485 -1085 13500 -1065
rect 13450 -1115 13500 -1085
rect 13450 -1135 13465 -1115
rect 13485 -1135 13500 -1115
rect 13450 -1165 13500 -1135
rect 13450 -1185 13465 -1165
rect 13485 -1185 13500 -1165
rect 13450 -1215 13500 -1185
rect 13450 -1235 13465 -1215
rect 13485 -1235 13500 -1215
rect 13450 -1265 13500 -1235
rect 13450 -1285 13465 -1265
rect 13485 -1285 13500 -1265
rect 13450 -1315 13500 -1285
rect 13450 -1335 13465 -1315
rect 13485 -1335 13500 -1315
rect 13450 -1365 13500 -1335
rect 13450 -1385 13465 -1365
rect 13485 -1385 13500 -1365
rect 13450 -1415 13500 -1385
rect 13450 -1435 13465 -1415
rect 13485 -1435 13500 -1415
rect 13450 -1465 13500 -1435
rect 13450 -1485 13465 -1465
rect 13485 -1485 13500 -1465
rect 13450 -1515 13500 -1485
rect 13450 -1535 13465 -1515
rect 13485 -1535 13500 -1515
rect 13450 -1550 13500 -1535
rect 13750 -1065 13800 -1050
rect 13750 -1085 13765 -1065
rect 13785 -1085 13800 -1065
rect 13750 -1115 13800 -1085
rect 13750 -1135 13765 -1115
rect 13785 -1135 13800 -1115
rect 13750 -1165 13800 -1135
rect 13750 -1185 13765 -1165
rect 13785 -1185 13800 -1165
rect 13750 -1215 13800 -1185
rect 13750 -1235 13765 -1215
rect 13785 -1235 13800 -1215
rect 13750 -1265 13800 -1235
rect 13750 -1285 13765 -1265
rect 13785 -1285 13800 -1265
rect 13750 -1315 13800 -1285
rect 13750 -1335 13765 -1315
rect 13785 -1335 13800 -1315
rect 13750 -1365 13800 -1335
rect 13750 -1385 13765 -1365
rect 13785 -1385 13800 -1365
rect 13750 -1415 13800 -1385
rect 13750 -1435 13765 -1415
rect 13785 -1435 13800 -1415
rect 13750 -1465 13800 -1435
rect 13750 -1485 13765 -1465
rect 13785 -1485 13800 -1465
rect 13750 -1515 13800 -1485
rect 13750 -1535 13765 -1515
rect 13785 -1535 13800 -1515
rect 13150 -1585 13165 -1565
rect 13185 -1585 13200 -1565
rect 13150 -1600 13200 -1585
rect 13750 -1565 13800 -1535
rect 14050 -1065 14100 -1035
rect 14050 -1085 14065 -1065
rect 14085 -1085 14100 -1065
rect 14050 -1115 14100 -1085
rect 14050 -1135 14065 -1115
rect 14085 -1135 14100 -1115
rect 14050 -1165 14100 -1135
rect 14050 -1185 14065 -1165
rect 14085 -1185 14100 -1165
rect 14050 -1215 14100 -1185
rect 14050 -1235 14065 -1215
rect 14085 -1235 14100 -1215
rect 14050 -1265 14100 -1235
rect 14050 -1285 14065 -1265
rect 14085 -1285 14100 -1265
rect 14050 -1315 14100 -1285
rect 14050 -1335 14065 -1315
rect 14085 -1335 14100 -1315
rect 14050 -1365 14100 -1335
rect 14050 -1385 14065 -1365
rect 14085 -1385 14100 -1365
rect 14050 -1415 14100 -1385
rect 14050 -1435 14065 -1415
rect 14085 -1435 14100 -1415
rect 14050 -1465 14100 -1435
rect 14050 -1485 14065 -1465
rect 14085 -1485 14100 -1465
rect 14050 -1515 14100 -1485
rect 14050 -1535 14065 -1515
rect 14085 -1535 14100 -1515
rect 14050 -1550 14100 -1535
rect 14350 -965 14400 -785
rect 15550 740 15600 910
rect 16750 1585 16800 1600
rect 16750 1565 16765 1585
rect 16785 1565 16800 1585
rect 16750 1535 16800 1565
rect 16750 1515 16765 1535
rect 16785 1515 16800 1535
rect 16750 1485 16800 1515
rect 16750 1465 16765 1485
rect 16785 1465 16800 1485
rect 16750 1435 16800 1465
rect 16750 1415 16765 1435
rect 16785 1415 16800 1435
rect 16750 1385 16800 1415
rect 16750 1365 16765 1385
rect 16785 1365 16800 1385
rect 16750 1335 16800 1365
rect 16750 1315 16765 1335
rect 16785 1315 16800 1335
rect 16750 1285 16800 1315
rect 16750 1265 16765 1285
rect 16785 1265 16800 1285
rect 16750 1235 16800 1265
rect 16750 1215 16765 1235
rect 16785 1215 16800 1235
rect 16750 1185 16800 1215
rect 16750 1165 16765 1185
rect 16785 1165 16800 1185
rect 16750 1135 16800 1165
rect 16750 1115 16765 1135
rect 16785 1115 16800 1135
rect 16750 1085 16800 1115
rect 16750 1065 16765 1085
rect 16785 1065 16800 1085
rect 16750 1035 16800 1065
rect 16750 1015 16765 1035
rect 16785 1015 16800 1035
rect 16750 985 16800 1015
rect 16750 965 16765 985
rect 16785 965 16800 985
rect 16750 935 16800 965
rect 16750 915 16765 935
rect 16785 915 16800 935
rect 15700 840 15750 850
rect 15700 810 15710 840
rect 15740 810 15750 840
rect 15700 800 15750 810
rect 16000 840 16050 850
rect 16000 810 16010 840
rect 16040 810 16050 840
rect 16000 800 16050 810
rect 16300 840 16350 850
rect 16300 810 16310 840
rect 16340 810 16350 840
rect 16300 800 16350 810
rect 16600 840 16650 850
rect 16600 810 16610 840
rect 16640 810 16650 840
rect 16600 800 16650 810
rect 16750 840 16800 915
rect 17950 1585 18000 1660
rect 20350 1690 20400 1700
rect 20350 1660 20360 1690
rect 20390 1660 20400 1690
rect 17950 1565 17965 1585
rect 17985 1565 18000 1585
rect 17950 1540 18000 1565
rect 17950 1510 17960 1540
rect 17990 1510 18000 1540
rect 17950 1485 18000 1510
rect 17950 1465 17965 1485
rect 17985 1465 18000 1485
rect 17950 1440 18000 1465
rect 17950 1410 17960 1440
rect 17990 1410 18000 1440
rect 17950 1385 18000 1410
rect 17950 1365 17965 1385
rect 17985 1365 18000 1385
rect 17950 1340 18000 1365
rect 17950 1310 17960 1340
rect 17990 1310 18000 1340
rect 17950 1285 18000 1310
rect 17950 1265 17965 1285
rect 17985 1265 18000 1285
rect 17950 1240 18000 1265
rect 17950 1210 17960 1240
rect 17990 1210 18000 1240
rect 17950 1185 18000 1210
rect 17950 1165 17965 1185
rect 17985 1165 18000 1185
rect 17950 1140 18000 1165
rect 17950 1110 17960 1140
rect 17990 1110 18000 1140
rect 17950 1085 18000 1110
rect 17950 1065 17965 1085
rect 17985 1065 18000 1085
rect 17950 1040 18000 1065
rect 17950 1010 17960 1040
rect 17990 1010 18000 1040
rect 17950 985 18000 1010
rect 17950 965 17965 985
rect 17985 965 18000 985
rect 17950 940 18000 965
rect 17950 910 17960 940
rect 17990 910 18000 940
rect 16750 810 16760 840
rect 16790 810 16800 840
rect 15550 710 15560 740
rect 15590 710 15600 740
rect 15550 685 15600 710
rect 15550 665 15565 685
rect 15585 665 15600 685
rect 15550 640 15600 665
rect 15550 610 15560 640
rect 15590 610 15600 640
rect 15550 585 15600 610
rect 15550 565 15565 585
rect 15585 565 15600 585
rect 15550 540 15600 565
rect 15550 510 15560 540
rect 15590 510 15600 540
rect 15550 485 15600 510
rect 15550 465 15565 485
rect 15585 465 15600 485
rect 15550 440 15600 465
rect 15550 410 15560 440
rect 15590 410 15600 440
rect 15550 385 15600 410
rect 15550 365 15565 385
rect 15585 365 15600 385
rect 15550 340 15600 365
rect 15550 310 15560 340
rect 15590 310 15600 340
rect 15550 285 15600 310
rect 15550 265 15565 285
rect 15585 265 15600 285
rect 15550 240 15600 265
rect 15550 210 15560 240
rect 15590 210 15600 240
rect 15550 185 15600 210
rect 15550 165 15565 185
rect 15585 165 15600 185
rect 15550 140 15600 165
rect 15550 110 15560 140
rect 15590 110 15600 140
rect 15550 85 15600 110
rect 15550 65 15565 85
rect 15585 65 15600 85
rect 15550 -10 15600 65
rect 16750 735 16800 810
rect 16900 840 16950 850
rect 16900 810 16910 840
rect 16940 810 16950 840
rect 16900 800 16950 810
rect 17200 840 17250 850
rect 17200 810 17210 840
rect 17240 810 17250 840
rect 17200 800 17250 810
rect 17500 840 17550 850
rect 17500 810 17510 840
rect 17540 810 17550 840
rect 17500 800 17550 810
rect 17800 840 17850 850
rect 17800 810 17810 840
rect 17840 810 17850 840
rect 17800 800 17850 810
rect 16750 715 16765 735
rect 16785 715 16800 735
rect 16750 685 16800 715
rect 16750 665 16765 685
rect 16785 665 16800 685
rect 16750 635 16800 665
rect 16750 615 16765 635
rect 16785 615 16800 635
rect 16750 585 16800 615
rect 16750 565 16765 585
rect 16785 565 16800 585
rect 16750 535 16800 565
rect 16750 515 16765 535
rect 16785 515 16800 535
rect 16750 485 16800 515
rect 16750 465 16765 485
rect 16785 465 16800 485
rect 16750 435 16800 465
rect 16750 415 16765 435
rect 16785 415 16800 435
rect 16750 385 16800 415
rect 16750 365 16765 385
rect 16785 365 16800 385
rect 16750 335 16800 365
rect 16750 315 16765 335
rect 16785 315 16800 335
rect 16750 285 16800 315
rect 16750 265 16765 285
rect 16785 265 16800 285
rect 16750 235 16800 265
rect 16750 215 16765 235
rect 16785 215 16800 235
rect 16750 185 16800 215
rect 16750 165 16765 185
rect 16785 165 16800 185
rect 16750 135 16800 165
rect 16750 115 16765 135
rect 16785 115 16800 135
rect 16750 85 16800 115
rect 16750 65 16765 85
rect 16785 65 16800 85
rect 16750 50 16800 65
rect 17950 740 18000 910
rect 19150 1585 19200 1600
rect 19150 1565 19165 1585
rect 19185 1565 19200 1585
rect 19150 1535 19200 1565
rect 19150 1515 19165 1535
rect 19185 1515 19200 1535
rect 19150 1485 19200 1515
rect 19150 1465 19165 1485
rect 19185 1465 19200 1485
rect 19150 1435 19200 1465
rect 19150 1415 19165 1435
rect 19185 1415 19200 1435
rect 19150 1385 19200 1415
rect 19150 1365 19165 1385
rect 19185 1365 19200 1385
rect 19150 1335 19200 1365
rect 19150 1315 19165 1335
rect 19185 1315 19200 1335
rect 19150 1285 19200 1315
rect 19150 1265 19165 1285
rect 19185 1265 19200 1285
rect 19150 1235 19200 1265
rect 19150 1215 19165 1235
rect 19185 1215 19200 1235
rect 19150 1185 19200 1215
rect 19150 1165 19165 1185
rect 19185 1165 19200 1185
rect 19150 1135 19200 1165
rect 19150 1115 19165 1135
rect 19185 1115 19200 1135
rect 19150 1085 19200 1115
rect 19150 1065 19165 1085
rect 19185 1065 19200 1085
rect 19150 1035 19200 1065
rect 19150 1015 19165 1035
rect 19185 1015 19200 1035
rect 19150 985 19200 1015
rect 19150 965 19165 985
rect 19185 965 19200 985
rect 19150 935 19200 965
rect 19150 915 19165 935
rect 19185 915 19200 935
rect 18100 840 18150 850
rect 18100 810 18110 840
rect 18140 810 18150 840
rect 18100 800 18150 810
rect 18400 840 18450 850
rect 18400 810 18410 840
rect 18440 810 18450 840
rect 18400 800 18450 810
rect 18700 840 18750 850
rect 18700 810 18710 840
rect 18740 810 18750 840
rect 18700 800 18750 810
rect 19000 840 19050 850
rect 19000 810 19010 840
rect 19040 810 19050 840
rect 19000 800 19050 810
rect 19150 840 19200 915
rect 20350 1585 20400 1660
rect 24550 1690 24600 1700
rect 24550 1660 24560 1690
rect 24590 1660 24600 1690
rect 20350 1565 20365 1585
rect 20385 1565 20400 1585
rect 20350 1540 20400 1565
rect 20350 1510 20360 1540
rect 20390 1510 20400 1540
rect 20350 1485 20400 1510
rect 20350 1465 20365 1485
rect 20385 1465 20400 1485
rect 20350 1440 20400 1465
rect 20350 1410 20360 1440
rect 20390 1410 20400 1440
rect 20350 1385 20400 1410
rect 20350 1365 20365 1385
rect 20385 1365 20400 1385
rect 20350 1340 20400 1365
rect 20350 1310 20360 1340
rect 20390 1310 20400 1340
rect 20350 1285 20400 1310
rect 20350 1265 20365 1285
rect 20385 1265 20400 1285
rect 20350 1240 20400 1265
rect 20350 1210 20360 1240
rect 20390 1210 20400 1240
rect 20350 1185 20400 1210
rect 20350 1165 20365 1185
rect 20385 1165 20400 1185
rect 20350 1140 20400 1165
rect 20350 1110 20360 1140
rect 20390 1110 20400 1140
rect 20350 1085 20400 1110
rect 20350 1065 20365 1085
rect 20385 1065 20400 1085
rect 20350 1040 20400 1065
rect 20350 1010 20360 1040
rect 20390 1010 20400 1040
rect 20350 985 20400 1010
rect 20350 965 20365 985
rect 20385 965 20400 985
rect 20350 940 20400 965
rect 20350 910 20360 940
rect 20390 910 20400 940
rect 19150 810 19160 840
rect 19190 810 19200 840
rect 17950 710 17960 740
rect 17990 710 18000 740
rect 17950 685 18000 710
rect 17950 665 17965 685
rect 17985 665 18000 685
rect 17950 640 18000 665
rect 17950 610 17960 640
rect 17990 610 18000 640
rect 17950 585 18000 610
rect 17950 565 17965 585
rect 17985 565 18000 585
rect 17950 540 18000 565
rect 17950 510 17960 540
rect 17990 510 18000 540
rect 17950 485 18000 510
rect 17950 465 17965 485
rect 17985 465 18000 485
rect 17950 440 18000 465
rect 17950 410 17960 440
rect 17990 410 18000 440
rect 17950 385 18000 410
rect 17950 365 17965 385
rect 17985 365 18000 385
rect 17950 340 18000 365
rect 17950 310 17960 340
rect 17990 310 18000 340
rect 17950 285 18000 310
rect 17950 265 17965 285
rect 17985 265 18000 285
rect 17950 240 18000 265
rect 17950 210 17960 240
rect 17990 210 18000 240
rect 17950 185 18000 210
rect 17950 165 17965 185
rect 17985 165 18000 185
rect 17950 140 18000 165
rect 17950 110 17960 140
rect 17990 110 18000 140
rect 17950 85 18000 110
rect 17950 65 17965 85
rect 17985 65 18000 85
rect 15550 -40 15560 -10
rect 15590 -40 15600 -10
rect 15550 -115 15600 -40
rect 17950 -10 18000 65
rect 19150 735 19200 810
rect 19300 840 19350 850
rect 19300 810 19310 840
rect 19340 810 19350 840
rect 19300 800 19350 810
rect 19600 840 19650 850
rect 19600 810 19610 840
rect 19640 810 19650 840
rect 19600 800 19650 810
rect 19900 840 19950 850
rect 19900 810 19910 840
rect 19940 810 19950 840
rect 19900 800 19950 810
rect 20200 840 20250 850
rect 20200 810 20210 840
rect 20240 810 20250 840
rect 20200 800 20250 810
rect 19150 715 19165 735
rect 19185 715 19200 735
rect 19150 685 19200 715
rect 19150 665 19165 685
rect 19185 665 19200 685
rect 19150 635 19200 665
rect 19150 615 19165 635
rect 19185 615 19200 635
rect 19150 585 19200 615
rect 19150 565 19165 585
rect 19185 565 19200 585
rect 19150 535 19200 565
rect 19150 515 19165 535
rect 19185 515 19200 535
rect 19150 485 19200 515
rect 19150 465 19165 485
rect 19185 465 19200 485
rect 19150 435 19200 465
rect 19150 415 19165 435
rect 19185 415 19200 435
rect 19150 385 19200 415
rect 19150 365 19165 385
rect 19185 365 19200 385
rect 19150 335 19200 365
rect 19150 315 19165 335
rect 19185 315 19200 335
rect 19150 285 19200 315
rect 19150 265 19165 285
rect 19185 265 19200 285
rect 19150 235 19200 265
rect 19150 215 19165 235
rect 19185 215 19200 235
rect 19150 185 19200 215
rect 19150 165 19165 185
rect 19185 165 19200 185
rect 19150 135 19200 165
rect 19150 115 19165 135
rect 19185 115 19200 135
rect 19150 85 19200 115
rect 19150 65 19165 85
rect 19185 65 19200 85
rect 19150 50 19200 65
rect 20350 740 20400 910
rect 21550 1585 21600 1600
rect 21550 1565 21565 1585
rect 21585 1565 21600 1585
rect 21550 1535 21600 1565
rect 21550 1515 21565 1535
rect 21585 1515 21600 1535
rect 21550 1485 21600 1515
rect 21550 1465 21565 1485
rect 21585 1465 21600 1485
rect 21550 1435 21600 1465
rect 21550 1415 21565 1435
rect 21585 1415 21600 1435
rect 21550 1385 21600 1415
rect 21550 1365 21565 1385
rect 21585 1365 21600 1385
rect 21550 1335 21600 1365
rect 21550 1315 21565 1335
rect 21585 1315 21600 1335
rect 21550 1285 21600 1315
rect 21550 1265 21565 1285
rect 21585 1265 21600 1285
rect 21550 1235 21600 1265
rect 21550 1215 21565 1235
rect 21585 1215 21600 1235
rect 21550 1185 21600 1215
rect 21550 1165 21565 1185
rect 21585 1165 21600 1185
rect 21550 1135 21600 1165
rect 21550 1115 21565 1135
rect 21585 1115 21600 1135
rect 21550 1085 21600 1115
rect 21550 1065 21565 1085
rect 21585 1065 21600 1085
rect 21550 1035 21600 1065
rect 21550 1015 21565 1035
rect 21585 1015 21600 1035
rect 21550 985 21600 1015
rect 21550 965 21565 985
rect 21585 965 21600 985
rect 21550 935 21600 965
rect 21550 915 21565 935
rect 21585 915 21600 935
rect 20500 840 20550 850
rect 20500 810 20510 840
rect 20540 810 20550 840
rect 20500 800 20550 810
rect 20800 840 20850 850
rect 20800 810 20810 840
rect 20840 810 20850 840
rect 20800 800 20850 810
rect 21100 840 21150 850
rect 21100 810 21110 840
rect 21140 810 21150 840
rect 21100 800 21150 810
rect 21400 840 21450 850
rect 21400 810 21410 840
rect 21440 810 21450 840
rect 21400 800 21450 810
rect 20350 710 20360 740
rect 20390 710 20400 740
rect 20350 685 20400 710
rect 20350 665 20365 685
rect 20385 665 20400 685
rect 20350 640 20400 665
rect 20350 610 20360 640
rect 20390 610 20400 640
rect 20350 585 20400 610
rect 20350 565 20365 585
rect 20385 565 20400 585
rect 20350 540 20400 565
rect 20350 510 20360 540
rect 20390 510 20400 540
rect 20350 485 20400 510
rect 20350 465 20365 485
rect 20385 465 20400 485
rect 20350 440 20400 465
rect 20350 410 20360 440
rect 20390 410 20400 440
rect 20350 385 20400 410
rect 20350 365 20365 385
rect 20385 365 20400 385
rect 20350 340 20400 365
rect 20350 310 20360 340
rect 20390 310 20400 340
rect 20350 285 20400 310
rect 20350 265 20365 285
rect 20385 265 20400 285
rect 20350 240 20400 265
rect 20350 210 20360 240
rect 20390 210 20400 240
rect 20350 185 20400 210
rect 20350 165 20365 185
rect 20385 165 20400 185
rect 20350 140 20400 165
rect 20350 110 20360 140
rect 20390 110 20400 140
rect 20350 85 20400 110
rect 20350 65 20365 85
rect 20385 65 20400 85
rect 17950 -40 17960 -10
rect 17990 -40 18000 -10
rect 15550 -135 15565 -115
rect 15585 -135 15600 -115
rect 15550 -160 15600 -135
rect 15550 -190 15560 -160
rect 15590 -190 15600 -160
rect 15550 -215 15600 -190
rect 15550 -235 15565 -215
rect 15585 -235 15600 -215
rect 15550 -260 15600 -235
rect 15550 -290 15560 -260
rect 15590 -290 15600 -260
rect 15550 -315 15600 -290
rect 15550 -335 15565 -315
rect 15585 -335 15600 -315
rect 15550 -360 15600 -335
rect 15550 -390 15560 -360
rect 15590 -390 15600 -360
rect 15550 -415 15600 -390
rect 15550 -435 15565 -415
rect 15585 -435 15600 -415
rect 15550 -460 15600 -435
rect 15550 -490 15560 -460
rect 15590 -490 15600 -460
rect 15550 -515 15600 -490
rect 15550 -535 15565 -515
rect 15585 -535 15600 -515
rect 15550 -560 15600 -535
rect 15550 -590 15560 -560
rect 15590 -590 15600 -560
rect 15550 -615 15600 -590
rect 15550 -635 15565 -615
rect 15585 -635 15600 -615
rect 15550 -660 15600 -635
rect 15550 -690 15560 -660
rect 15590 -690 15600 -660
rect 15550 -715 15600 -690
rect 15550 -735 15565 -715
rect 15585 -735 15600 -715
rect 15550 -760 15600 -735
rect 15550 -790 15560 -760
rect 15590 -790 15600 -760
rect 14500 -860 14550 -850
rect 14500 -890 14510 -860
rect 14540 -890 14550 -860
rect 14500 -900 14550 -890
rect 14800 -860 14850 -850
rect 14800 -890 14810 -860
rect 14840 -890 14850 -860
rect 14800 -900 14850 -890
rect 15100 -860 15150 -850
rect 15100 -890 15110 -860
rect 15140 -890 15150 -860
rect 15100 -900 15150 -890
rect 15400 -860 15450 -850
rect 15400 -890 15410 -860
rect 15440 -890 15450 -860
rect 15400 -900 15450 -890
rect 14350 -985 14365 -965
rect 14385 -985 14400 -965
rect 14350 -1015 14400 -985
rect 14350 -1035 14365 -1015
rect 14385 -1035 14400 -1015
rect 14350 -1065 14400 -1035
rect 14350 -1085 14365 -1065
rect 14385 -1085 14400 -1065
rect 14350 -1115 14400 -1085
rect 14350 -1135 14365 -1115
rect 14385 -1135 14400 -1115
rect 14350 -1165 14400 -1135
rect 14350 -1185 14365 -1165
rect 14385 -1185 14400 -1165
rect 14350 -1215 14400 -1185
rect 14350 -1235 14365 -1215
rect 14385 -1235 14400 -1215
rect 14350 -1265 14400 -1235
rect 14350 -1285 14365 -1265
rect 14385 -1285 14400 -1265
rect 14350 -1315 14400 -1285
rect 14350 -1335 14365 -1315
rect 14385 -1335 14400 -1315
rect 14350 -1365 14400 -1335
rect 14350 -1385 14365 -1365
rect 14385 -1385 14400 -1365
rect 14350 -1415 14400 -1385
rect 14350 -1435 14365 -1415
rect 14385 -1435 14400 -1415
rect 14350 -1465 14400 -1435
rect 14350 -1485 14365 -1465
rect 14385 -1485 14400 -1465
rect 14350 -1515 14400 -1485
rect 14350 -1535 14365 -1515
rect 14385 -1535 14400 -1515
rect 13750 -1585 13765 -1565
rect 13785 -1585 13800 -1565
rect 13750 -1600 13800 -1585
rect 14350 -1565 14400 -1535
rect 14350 -1585 14365 -1565
rect 14385 -1585 14400 -1565
rect 14350 -1600 14400 -1585
rect 11950 -1615 14400 -1600
rect 11950 -1635 11965 -1615
rect 11985 -1635 12565 -1615
rect 12585 -1635 13165 -1615
rect 13185 -1635 13765 -1615
rect 13785 -1635 14365 -1615
rect 14385 -1635 14400 -1615
rect 11950 -1650 14400 -1635
rect 15550 -960 15600 -790
rect 16750 -115 16800 -100
rect 16750 -135 16765 -115
rect 16785 -135 16800 -115
rect 16750 -165 16800 -135
rect 16750 -185 16765 -165
rect 16785 -185 16800 -165
rect 16750 -215 16800 -185
rect 16750 -235 16765 -215
rect 16785 -235 16800 -215
rect 16750 -265 16800 -235
rect 16750 -285 16765 -265
rect 16785 -285 16800 -265
rect 16750 -315 16800 -285
rect 16750 -335 16765 -315
rect 16785 -335 16800 -315
rect 16750 -365 16800 -335
rect 16750 -385 16765 -365
rect 16785 -385 16800 -365
rect 16750 -415 16800 -385
rect 16750 -435 16765 -415
rect 16785 -435 16800 -415
rect 16750 -465 16800 -435
rect 16750 -485 16765 -465
rect 16785 -485 16800 -465
rect 16750 -515 16800 -485
rect 16750 -535 16765 -515
rect 16785 -535 16800 -515
rect 16750 -565 16800 -535
rect 16750 -585 16765 -565
rect 16785 -585 16800 -565
rect 16750 -615 16800 -585
rect 16750 -635 16765 -615
rect 16785 -635 16800 -615
rect 16750 -665 16800 -635
rect 16750 -685 16765 -665
rect 16785 -685 16800 -665
rect 16750 -715 16800 -685
rect 16750 -735 16765 -715
rect 16785 -735 16800 -715
rect 16750 -765 16800 -735
rect 16750 -785 16765 -765
rect 16785 -785 16800 -765
rect 15700 -860 15750 -850
rect 15700 -890 15710 -860
rect 15740 -890 15750 -860
rect 15700 -900 15750 -890
rect 16000 -860 16050 -850
rect 16000 -890 16010 -860
rect 16040 -890 16050 -860
rect 16000 -900 16050 -890
rect 16300 -860 16350 -850
rect 16300 -890 16310 -860
rect 16340 -890 16350 -860
rect 16300 -900 16350 -890
rect 16600 -860 16650 -850
rect 16600 -890 16610 -860
rect 16640 -890 16650 -860
rect 16600 -900 16650 -890
rect 16750 -860 16800 -785
rect 17950 -115 18000 -40
rect 20350 -10 20400 65
rect 20350 -40 20360 -10
rect 20390 -40 20400 -10
rect 17950 -135 17965 -115
rect 17985 -135 18000 -115
rect 17950 -160 18000 -135
rect 17950 -190 17960 -160
rect 17990 -190 18000 -160
rect 17950 -215 18000 -190
rect 17950 -235 17965 -215
rect 17985 -235 18000 -215
rect 17950 -260 18000 -235
rect 17950 -290 17960 -260
rect 17990 -290 18000 -260
rect 17950 -315 18000 -290
rect 17950 -335 17965 -315
rect 17985 -335 18000 -315
rect 17950 -360 18000 -335
rect 17950 -390 17960 -360
rect 17990 -390 18000 -360
rect 17950 -415 18000 -390
rect 17950 -435 17965 -415
rect 17985 -435 18000 -415
rect 17950 -460 18000 -435
rect 17950 -490 17960 -460
rect 17990 -490 18000 -460
rect 17950 -515 18000 -490
rect 17950 -535 17965 -515
rect 17985 -535 18000 -515
rect 17950 -560 18000 -535
rect 17950 -590 17960 -560
rect 17990 -590 18000 -560
rect 17950 -615 18000 -590
rect 17950 -635 17965 -615
rect 17985 -635 18000 -615
rect 17950 -660 18000 -635
rect 17950 -690 17960 -660
rect 17990 -690 18000 -660
rect 17950 -715 18000 -690
rect 17950 -735 17965 -715
rect 17985 -735 18000 -715
rect 17950 -760 18000 -735
rect 17950 -790 17960 -760
rect 17990 -790 18000 -760
rect 16750 -890 16760 -860
rect 16790 -890 16800 -860
rect 15550 -990 15560 -960
rect 15590 -990 15600 -960
rect 15550 -1015 15600 -990
rect 15550 -1035 15565 -1015
rect 15585 -1035 15600 -1015
rect 15550 -1060 15600 -1035
rect 15550 -1090 15560 -1060
rect 15590 -1090 15600 -1060
rect 15550 -1115 15600 -1090
rect 15550 -1135 15565 -1115
rect 15585 -1135 15600 -1115
rect 15550 -1160 15600 -1135
rect 15550 -1190 15560 -1160
rect 15590 -1190 15600 -1160
rect 15550 -1215 15600 -1190
rect 15550 -1235 15565 -1215
rect 15585 -1235 15600 -1215
rect 15550 -1260 15600 -1235
rect 15550 -1290 15560 -1260
rect 15590 -1290 15600 -1260
rect 15550 -1315 15600 -1290
rect 15550 -1335 15565 -1315
rect 15585 -1335 15600 -1315
rect 15550 -1360 15600 -1335
rect 15550 -1390 15560 -1360
rect 15590 -1390 15600 -1360
rect 15550 -1415 15600 -1390
rect 15550 -1435 15565 -1415
rect 15585 -1435 15600 -1415
rect 15550 -1460 15600 -1435
rect 15550 -1490 15560 -1460
rect 15590 -1490 15600 -1460
rect 15550 -1515 15600 -1490
rect 15550 -1535 15565 -1515
rect 15585 -1535 15600 -1515
rect 15550 -1560 15600 -1535
rect 15550 -1590 15560 -1560
rect 15590 -1590 15600 -1560
rect 15550 -1615 15600 -1590
rect 15550 -1635 15565 -1615
rect 15585 -1635 15600 -1615
rect 10750 -1740 10760 -1710
rect 10790 -1740 10800 -1710
rect 10750 -1750 10800 -1740
rect 15550 -1710 15600 -1635
rect 16750 -965 16800 -890
rect 16900 -860 16950 -850
rect 16900 -890 16910 -860
rect 16940 -890 16950 -860
rect 16900 -900 16950 -890
rect 17200 -860 17250 -850
rect 17200 -890 17210 -860
rect 17240 -890 17250 -860
rect 17200 -900 17250 -890
rect 17500 -860 17550 -850
rect 17500 -890 17510 -860
rect 17540 -890 17550 -860
rect 17500 -900 17550 -890
rect 17800 -860 17850 -850
rect 17800 -890 17810 -860
rect 17840 -890 17850 -860
rect 17800 -900 17850 -890
rect 16750 -985 16765 -965
rect 16785 -985 16800 -965
rect 16750 -1015 16800 -985
rect 16750 -1035 16765 -1015
rect 16785 -1035 16800 -1015
rect 16750 -1065 16800 -1035
rect 16750 -1085 16765 -1065
rect 16785 -1085 16800 -1065
rect 16750 -1115 16800 -1085
rect 16750 -1135 16765 -1115
rect 16785 -1135 16800 -1115
rect 16750 -1165 16800 -1135
rect 16750 -1185 16765 -1165
rect 16785 -1185 16800 -1165
rect 16750 -1215 16800 -1185
rect 16750 -1235 16765 -1215
rect 16785 -1235 16800 -1215
rect 16750 -1265 16800 -1235
rect 16750 -1285 16765 -1265
rect 16785 -1285 16800 -1265
rect 16750 -1315 16800 -1285
rect 16750 -1335 16765 -1315
rect 16785 -1335 16800 -1315
rect 16750 -1365 16800 -1335
rect 16750 -1385 16765 -1365
rect 16785 -1385 16800 -1365
rect 16750 -1415 16800 -1385
rect 16750 -1435 16765 -1415
rect 16785 -1435 16800 -1415
rect 16750 -1465 16800 -1435
rect 16750 -1485 16765 -1465
rect 16785 -1485 16800 -1465
rect 16750 -1515 16800 -1485
rect 16750 -1535 16765 -1515
rect 16785 -1535 16800 -1515
rect 16750 -1565 16800 -1535
rect 16750 -1585 16765 -1565
rect 16785 -1585 16800 -1565
rect 16750 -1615 16800 -1585
rect 16750 -1635 16765 -1615
rect 16785 -1635 16800 -1615
rect 16750 -1650 16800 -1635
rect 17950 -960 18000 -790
rect 19150 -115 19200 -100
rect 19150 -135 19165 -115
rect 19185 -135 19200 -115
rect 19150 -165 19200 -135
rect 19150 -185 19165 -165
rect 19185 -185 19200 -165
rect 19150 -215 19200 -185
rect 19150 -235 19165 -215
rect 19185 -235 19200 -215
rect 19150 -265 19200 -235
rect 19150 -285 19165 -265
rect 19185 -285 19200 -265
rect 19150 -315 19200 -285
rect 19150 -335 19165 -315
rect 19185 -335 19200 -315
rect 19150 -365 19200 -335
rect 19150 -385 19165 -365
rect 19185 -385 19200 -365
rect 19150 -415 19200 -385
rect 19150 -435 19165 -415
rect 19185 -435 19200 -415
rect 19150 -465 19200 -435
rect 19150 -485 19165 -465
rect 19185 -485 19200 -465
rect 19150 -515 19200 -485
rect 19150 -535 19165 -515
rect 19185 -535 19200 -515
rect 19150 -565 19200 -535
rect 19150 -585 19165 -565
rect 19185 -585 19200 -565
rect 19150 -615 19200 -585
rect 19150 -635 19165 -615
rect 19185 -635 19200 -615
rect 19150 -665 19200 -635
rect 19150 -685 19165 -665
rect 19185 -685 19200 -665
rect 19150 -715 19200 -685
rect 19150 -735 19165 -715
rect 19185 -735 19200 -715
rect 19150 -765 19200 -735
rect 19150 -785 19165 -765
rect 19185 -785 19200 -765
rect 18100 -860 18150 -850
rect 18100 -890 18110 -860
rect 18140 -890 18150 -860
rect 18100 -900 18150 -890
rect 18400 -860 18450 -850
rect 18400 -890 18410 -860
rect 18440 -890 18450 -860
rect 18400 -900 18450 -890
rect 18700 -860 18750 -850
rect 18700 -890 18710 -860
rect 18740 -890 18750 -860
rect 18700 -900 18750 -890
rect 19000 -860 19050 -850
rect 19000 -890 19010 -860
rect 19040 -890 19050 -860
rect 19000 -900 19050 -890
rect 19150 -860 19200 -785
rect 20350 -115 20400 -40
rect 20350 -135 20365 -115
rect 20385 -135 20400 -115
rect 20350 -160 20400 -135
rect 20350 -190 20360 -160
rect 20390 -190 20400 -160
rect 20350 -215 20400 -190
rect 20350 -235 20365 -215
rect 20385 -235 20400 -215
rect 20350 -260 20400 -235
rect 20350 -290 20360 -260
rect 20390 -290 20400 -260
rect 20350 -315 20400 -290
rect 20350 -335 20365 -315
rect 20385 -335 20400 -315
rect 20350 -360 20400 -335
rect 20350 -390 20360 -360
rect 20390 -390 20400 -360
rect 20350 -415 20400 -390
rect 20350 -435 20365 -415
rect 20385 -435 20400 -415
rect 20350 -460 20400 -435
rect 20350 -490 20360 -460
rect 20390 -490 20400 -460
rect 20350 -515 20400 -490
rect 20350 -535 20365 -515
rect 20385 -535 20400 -515
rect 20350 -560 20400 -535
rect 20350 -590 20360 -560
rect 20390 -590 20400 -560
rect 20350 -615 20400 -590
rect 20350 -635 20365 -615
rect 20385 -635 20400 -615
rect 20350 -660 20400 -635
rect 20350 -690 20360 -660
rect 20390 -690 20400 -660
rect 20350 -715 20400 -690
rect 20350 -735 20365 -715
rect 20385 -735 20400 -715
rect 20350 -760 20400 -735
rect 20350 -790 20360 -760
rect 20390 -790 20400 -760
rect 19150 -890 19160 -860
rect 19190 -890 19200 -860
rect 17950 -990 17960 -960
rect 17990 -990 18000 -960
rect 17950 -1015 18000 -990
rect 17950 -1035 17965 -1015
rect 17985 -1035 18000 -1015
rect 17950 -1060 18000 -1035
rect 17950 -1090 17960 -1060
rect 17990 -1090 18000 -1060
rect 17950 -1115 18000 -1090
rect 17950 -1135 17965 -1115
rect 17985 -1135 18000 -1115
rect 17950 -1160 18000 -1135
rect 17950 -1190 17960 -1160
rect 17990 -1190 18000 -1160
rect 17950 -1215 18000 -1190
rect 17950 -1235 17965 -1215
rect 17985 -1235 18000 -1215
rect 17950 -1260 18000 -1235
rect 17950 -1290 17960 -1260
rect 17990 -1290 18000 -1260
rect 17950 -1315 18000 -1290
rect 17950 -1335 17965 -1315
rect 17985 -1335 18000 -1315
rect 17950 -1360 18000 -1335
rect 17950 -1390 17960 -1360
rect 17990 -1390 18000 -1360
rect 17950 -1415 18000 -1390
rect 17950 -1435 17965 -1415
rect 17985 -1435 18000 -1415
rect 17950 -1460 18000 -1435
rect 17950 -1490 17960 -1460
rect 17990 -1490 18000 -1460
rect 17950 -1515 18000 -1490
rect 17950 -1535 17965 -1515
rect 17985 -1535 18000 -1515
rect 17950 -1560 18000 -1535
rect 17950 -1590 17960 -1560
rect 17990 -1590 18000 -1560
rect 17950 -1615 18000 -1590
rect 17950 -1635 17965 -1615
rect 17985 -1635 18000 -1615
rect 15550 -1740 15560 -1710
rect 15590 -1740 15600 -1710
rect 15550 -1750 15600 -1740
rect 17950 -1710 18000 -1635
rect 19150 -965 19200 -890
rect 19300 -860 19350 -850
rect 19300 -890 19310 -860
rect 19340 -890 19350 -860
rect 19300 -900 19350 -890
rect 19600 -860 19650 -850
rect 19600 -890 19610 -860
rect 19640 -890 19650 -860
rect 19600 -900 19650 -890
rect 19900 -860 19950 -850
rect 19900 -890 19910 -860
rect 19940 -890 19950 -860
rect 19900 -900 19950 -890
rect 20200 -860 20250 -850
rect 20200 -890 20210 -860
rect 20240 -890 20250 -860
rect 20200 -900 20250 -890
rect 19150 -985 19165 -965
rect 19185 -985 19200 -965
rect 19150 -1015 19200 -985
rect 19150 -1035 19165 -1015
rect 19185 -1035 19200 -1015
rect 19150 -1065 19200 -1035
rect 19150 -1085 19165 -1065
rect 19185 -1085 19200 -1065
rect 19150 -1115 19200 -1085
rect 19150 -1135 19165 -1115
rect 19185 -1135 19200 -1115
rect 19150 -1165 19200 -1135
rect 19150 -1185 19165 -1165
rect 19185 -1185 19200 -1165
rect 19150 -1215 19200 -1185
rect 19150 -1235 19165 -1215
rect 19185 -1235 19200 -1215
rect 19150 -1265 19200 -1235
rect 19150 -1285 19165 -1265
rect 19185 -1285 19200 -1265
rect 19150 -1315 19200 -1285
rect 19150 -1335 19165 -1315
rect 19185 -1335 19200 -1315
rect 19150 -1365 19200 -1335
rect 19150 -1385 19165 -1365
rect 19185 -1385 19200 -1365
rect 19150 -1415 19200 -1385
rect 19150 -1435 19165 -1415
rect 19185 -1435 19200 -1415
rect 19150 -1465 19200 -1435
rect 19150 -1485 19165 -1465
rect 19185 -1485 19200 -1465
rect 19150 -1515 19200 -1485
rect 19150 -1535 19165 -1515
rect 19185 -1535 19200 -1515
rect 19150 -1565 19200 -1535
rect 19150 -1585 19165 -1565
rect 19185 -1585 19200 -1565
rect 19150 -1615 19200 -1585
rect 19150 -1635 19165 -1615
rect 19185 -1635 19200 -1615
rect 19150 -1650 19200 -1635
rect 20350 -960 20400 -790
rect 21550 735 21600 915
rect 22450 1585 22500 1600
rect 22450 1565 22465 1585
rect 22485 1565 22500 1585
rect 22450 1535 22500 1565
rect 22450 1515 22465 1535
rect 22485 1515 22500 1535
rect 22450 1485 22500 1515
rect 22450 1465 22465 1485
rect 22485 1465 22500 1485
rect 22450 1435 22500 1465
rect 22450 1415 22465 1435
rect 22485 1415 22500 1435
rect 22450 1385 22500 1415
rect 22450 1365 22465 1385
rect 22485 1365 22500 1385
rect 22450 1335 22500 1365
rect 22450 1315 22465 1335
rect 22485 1315 22500 1335
rect 22450 1285 22500 1315
rect 22450 1265 22465 1285
rect 22485 1265 22500 1285
rect 22450 1235 22500 1265
rect 22450 1215 22465 1235
rect 22485 1215 22500 1235
rect 22450 1185 22500 1215
rect 22450 1165 22465 1185
rect 22485 1165 22500 1185
rect 22450 1135 22500 1165
rect 22450 1115 22465 1135
rect 22485 1115 22500 1135
rect 22450 1085 22500 1115
rect 22450 1065 22465 1085
rect 22485 1065 22500 1085
rect 22450 1035 22500 1065
rect 22450 1015 22465 1035
rect 22485 1015 22500 1035
rect 22450 985 22500 1015
rect 22450 965 22465 985
rect 22485 965 22500 985
rect 22450 935 22500 965
rect 22450 915 22465 935
rect 22485 915 22500 935
rect 21700 840 21750 850
rect 21700 810 21710 840
rect 21740 810 21750 840
rect 21700 800 21750 810
rect 22000 840 22050 850
rect 22000 810 22010 840
rect 22040 810 22050 840
rect 22000 800 22050 810
rect 22300 840 22350 850
rect 22300 810 22310 840
rect 22340 810 22350 840
rect 22300 800 22350 810
rect 22450 840 22500 915
rect 23350 1585 23400 1600
rect 23350 1565 23365 1585
rect 23385 1565 23400 1585
rect 23350 1535 23400 1565
rect 23350 1515 23365 1535
rect 23385 1515 23400 1535
rect 23350 1485 23400 1515
rect 23350 1465 23365 1485
rect 23385 1465 23400 1485
rect 23350 1435 23400 1465
rect 23350 1415 23365 1435
rect 23385 1415 23400 1435
rect 23350 1385 23400 1415
rect 23350 1365 23365 1385
rect 23385 1365 23400 1385
rect 23350 1335 23400 1365
rect 23350 1315 23365 1335
rect 23385 1315 23400 1335
rect 23350 1285 23400 1315
rect 23350 1265 23365 1285
rect 23385 1265 23400 1285
rect 23350 1235 23400 1265
rect 23350 1215 23365 1235
rect 23385 1215 23400 1235
rect 23350 1185 23400 1215
rect 23350 1165 23365 1185
rect 23385 1165 23400 1185
rect 23350 1135 23400 1165
rect 23350 1115 23365 1135
rect 23385 1115 23400 1135
rect 23350 1085 23400 1115
rect 23350 1065 23365 1085
rect 23385 1065 23400 1085
rect 23350 1035 23400 1065
rect 23350 1015 23365 1035
rect 23385 1015 23400 1035
rect 23350 985 23400 1015
rect 23350 965 23365 985
rect 23385 965 23400 985
rect 23350 935 23400 965
rect 23350 915 23365 935
rect 23385 915 23400 935
rect 22450 810 22460 840
rect 22490 810 22500 840
rect 21550 715 21565 735
rect 21585 715 21600 735
rect 21550 685 21600 715
rect 21550 665 21565 685
rect 21585 665 21600 685
rect 21550 635 21600 665
rect 21550 615 21565 635
rect 21585 615 21600 635
rect 21550 585 21600 615
rect 21550 565 21565 585
rect 21585 565 21600 585
rect 21550 535 21600 565
rect 21550 515 21565 535
rect 21585 515 21600 535
rect 21550 485 21600 515
rect 21550 465 21565 485
rect 21585 465 21600 485
rect 21550 435 21600 465
rect 21550 415 21565 435
rect 21585 415 21600 435
rect 21550 385 21600 415
rect 21550 365 21565 385
rect 21585 365 21600 385
rect 21550 335 21600 365
rect 21550 315 21565 335
rect 21585 315 21600 335
rect 21550 285 21600 315
rect 21550 265 21565 285
rect 21585 265 21600 285
rect 21550 235 21600 265
rect 21550 215 21565 235
rect 21585 215 21600 235
rect 21550 185 21600 215
rect 21550 165 21565 185
rect 21585 165 21600 185
rect 21550 135 21600 165
rect 21550 115 21565 135
rect 21585 115 21600 135
rect 21550 85 21600 115
rect 21550 65 21565 85
rect 21585 65 21600 85
rect 21550 -115 21600 65
rect 22450 735 22500 810
rect 22600 840 22650 850
rect 22600 810 22610 840
rect 22640 810 22650 840
rect 22600 800 22650 810
rect 22900 840 22950 850
rect 22900 810 22910 840
rect 22940 810 22950 840
rect 22900 800 22950 810
rect 23200 840 23250 850
rect 23200 810 23210 840
rect 23240 810 23250 840
rect 23200 800 23250 810
rect 22450 715 22465 735
rect 22485 715 22500 735
rect 22450 685 22500 715
rect 22450 665 22465 685
rect 22485 665 22500 685
rect 22450 635 22500 665
rect 22450 615 22465 635
rect 22485 615 22500 635
rect 22450 585 22500 615
rect 22450 565 22465 585
rect 22485 565 22500 585
rect 22450 535 22500 565
rect 22450 515 22465 535
rect 22485 515 22500 535
rect 22450 485 22500 515
rect 22450 465 22465 485
rect 22485 465 22500 485
rect 22450 435 22500 465
rect 22450 415 22465 435
rect 22485 415 22500 435
rect 22450 385 22500 415
rect 22450 365 22465 385
rect 22485 365 22500 385
rect 22450 335 22500 365
rect 22450 315 22465 335
rect 22485 315 22500 335
rect 22450 285 22500 315
rect 22450 265 22465 285
rect 22485 265 22500 285
rect 22450 235 22500 265
rect 22450 215 22465 235
rect 22485 215 22500 235
rect 22450 185 22500 215
rect 22450 165 22465 185
rect 22485 165 22500 185
rect 22450 135 22500 165
rect 22450 115 22465 135
rect 22485 115 22500 135
rect 22450 85 22500 115
rect 22450 65 22465 85
rect 22485 65 22500 85
rect 22450 50 22500 65
rect 23350 735 23400 915
rect 24550 1585 24600 1660
rect 28750 1690 28800 1700
rect 28750 1660 28760 1690
rect 28790 1660 28800 1690
rect 24550 1565 24565 1585
rect 24585 1565 24600 1585
rect 24550 1540 24600 1565
rect 24550 1510 24560 1540
rect 24590 1510 24600 1540
rect 24550 1485 24600 1510
rect 24550 1465 24565 1485
rect 24585 1465 24600 1485
rect 24550 1440 24600 1465
rect 24550 1410 24560 1440
rect 24590 1410 24600 1440
rect 24550 1385 24600 1410
rect 24550 1365 24565 1385
rect 24585 1365 24600 1385
rect 24550 1340 24600 1365
rect 24550 1310 24560 1340
rect 24590 1310 24600 1340
rect 24550 1285 24600 1310
rect 24550 1265 24565 1285
rect 24585 1265 24600 1285
rect 24550 1240 24600 1265
rect 24550 1210 24560 1240
rect 24590 1210 24600 1240
rect 24550 1185 24600 1210
rect 24550 1165 24565 1185
rect 24585 1165 24600 1185
rect 24550 1140 24600 1165
rect 24550 1110 24560 1140
rect 24590 1110 24600 1140
rect 24550 1085 24600 1110
rect 24550 1065 24565 1085
rect 24585 1065 24600 1085
rect 24550 1040 24600 1065
rect 24550 1010 24560 1040
rect 24590 1010 24600 1040
rect 24550 985 24600 1010
rect 24550 965 24565 985
rect 24585 965 24600 985
rect 24550 940 24600 965
rect 24550 910 24560 940
rect 24590 910 24600 940
rect 23500 840 23550 850
rect 23500 810 23510 840
rect 23540 810 23550 840
rect 23500 800 23550 810
rect 23800 840 23850 850
rect 23800 810 23810 840
rect 23840 810 23850 840
rect 23800 800 23850 810
rect 24100 840 24150 850
rect 24100 810 24110 840
rect 24140 810 24150 840
rect 24100 800 24150 810
rect 24400 840 24450 850
rect 24400 810 24410 840
rect 24440 810 24450 840
rect 24400 800 24450 810
rect 23350 715 23365 735
rect 23385 715 23400 735
rect 23350 685 23400 715
rect 23350 665 23365 685
rect 23385 665 23400 685
rect 23350 635 23400 665
rect 23350 615 23365 635
rect 23385 615 23400 635
rect 23350 585 23400 615
rect 23350 565 23365 585
rect 23385 565 23400 585
rect 23350 535 23400 565
rect 23350 515 23365 535
rect 23385 515 23400 535
rect 23350 485 23400 515
rect 23350 465 23365 485
rect 23385 465 23400 485
rect 23350 435 23400 465
rect 23350 415 23365 435
rect 23385 415 23400 435
rect 23350 385 23400 415
rect 23350 365 23365 385
rect 23385 365 23400 385
rect 23350 335 23400 365
rect 23350 315 23365 335
rect 23385 315 23400 335
rect 23350 285 23400 315
rect 23350 265 23365 285
rect 23385 265 23400 285
rect 23350 235 23400 265
rect 23350 215 23365 235
rect 23385 215 23400 235
rect 23350 185 23400 215
rect 23350 165 23365 185
rect 23385 165 23400 185
rect 23350 135 23400 165
rect 23350 115 23365 135
rect 23385 115 23400 135
rect 23350 85 23400 115
rect 23350 65 23365 85
rect 23385 65 23400 85
rect 21550 -135 21565 -115
rect 21585 -135 21600 -115
rect 21550 -165 21600 -135
rect 21550 -185 21565 -165
rect 21585 -185 21600 -165
rect 21550 -215 21600 -185
rect 21550 -235 21565 -215
rect 21585 -235 21600 -215
rect 21550 -265 21600 -235
rect 21550 -285 21565 -265
rect 21585 -285 21600 -265
rect 21550 -315 21600 -285
rect 21550 -335 21565 -315
rect 21585 -335 21600 -315
rect 21550 -365 21600 -335
rect 21550 -385 21565 -365
rect 21585 -385 21600 -365
rect 21550 -415 21600 -385
rect 21550 -435 21565 -415
rect 21585 -435 21600 -415
rect 21550 -465 21600 -435
rect 21550 -485 21565 -465
rect 21585 -485 21600 -465
rect 21550 -515 21600 -485
rect 21550 -535 21565 -515
rect 21585 -535 21600 -515
rect 21550 -565 21600 -535
rect 21550 -585 21565 -565
rect 21585 -585 21600 -565
rect 21550 -615 21600 -585
rect 21550 -635 21565 -615
rect 21585 -635 21600 -615
rect 21550 -665 21600 -635
rect 21550 -685 21565 -665
rect 21585 -685 21600 -665
rect 21550 -715 21600 -685
rect 21550 -735 21565 -715
rect 21585 -735 21600 -715
rect 21550 -765 21600 -735
rect 21550 -785 21565 -765
rect 21585 -785 21600 -765
rect 20500 -860 20550 -850
rect 20500 -890 20510 -860
rect 20540 -890 20550 -860
rect 20500 -900 20550 -890
rect 20800 -860 20850 -850
rect 20800 -890 20810 -860
rect 20840 -890 20850 -860
rect 20800 -900 20850 -890
rect 21100 -860 21150 -850
rect 21100 -890 21110 -860
rect 21140 -890 21150 -860
rect 21100 -900 21150 -890
rect 21400 -860 21450 -850
rect 21400 -890 21410 -860
rect 21440 -890 21450 -860
rect 21400 -900 21450 -890
rect 20350 -990 20360 -960
rect 20390 -990 20400 -960
rect 20350 -1015 20400 -990
rect 20350 -1035 20365 -1015
rect 20385 -1035 20400 -1015
rect 20350 -1060 20400 -1035
rect 20350 -1090 20360 -1060
rect 20390 -1090 20400 -1060
rect 20350 -1115 20400 -1090
rect 20350 -1135 20365 -1115
rect 20385 -1135 20400 -1115
rect 20350 -1160 20400 -1135
rect 20350 -1190 20360 -1160
rect 20390 -1190 20400 -1160
rect 20350 -1215 20400 -1190
rect 20350 -1235 20365 -1215
rect 20385 -1235 20400 -1215
rect 20350 -1260 20400 -1235
rect 20350 -1290 20360 -1260
rect 20390 -1290 20400 -1260
rect 20350 -1315 20400 -1290
rect 20350 -1335 20365 -1315
rect 20385 -1335 20400 -1315
rect 20350 -1360 20400 -1335
rect 20350 -1390 20360 -1360
rect 20390 -1390 20400 -1360
rect 20350 -1415 20400 -1390
rect 20350 -1435 20365 -1415
rect 20385 -1435 20400 -1415
rect 20350 -1460 20400 -1435
rect 20350 -1490 20360 -1460
rect 20390 -1490 20400 -1460
rect 20350 -1515 20400 -1490
rect 20350 -1535 20365 -1515
rect 20385 -1535 20400 -1515
rect 20350 -1560 20400 -1535
rect 20350 -1590 20360 -1560
rect 20390 -1590 20400 -1560
rect 20350 -1615 20400 -1590
rect 20350 -1635 20365 -1615
rect 20385 -1635 20400 -1615
rect 17950 -1740 17960 -1710
rect 17990 -1740 18000 -1710
rect 17950 -1750 18000 -1740
rect 20350 -1710 20400 -1635
rect 21550 -965 21600 -785
rect 22450 -115 22500 -100
rect 22450 -135 22465 -115
rect 22485 -135 22500 -115
rect 22450 -165 22500 -135
rect 22450 -185 22465 -165
rect 22485 -185 22500 -165
rect 22450 -215 22500 -185
rect 22450 -235 22465 -215
rect 22485 -235 22500 -215
rect 22450 -265 22500 -235
rect 22450 -285 22465 -265
rect 22485 -285 22500 -265
rect 22450 -315 22500 -285
rect 22450 -335 22465 -315
rect 22485 -335 22500 -315
rect 22450 -365 22500 -335
rect 22450 -385 22465 -365
rect 22485 -385 22500 -365
rect 22450 -415 22500 -385
rect 22450 -435 22465 -415
rect 22485 -435 22500 -415
rect 22450 -465 22500 -435
rect 22450 -485 22465 -465
rect 22485 -485 22500 -465
rect 22450 -515 22500 -485
rect 22450 -535 22465 -515
rect 22485 -535 22500 -515
rect 22450 -565 22500 -535
rect 22450 -585 22465 -565
rect 22485 -585 22500 -565
rect 22450 -615 22500 -585
rect 22450 -635 22465 -615
rect 22485 -635 22500 -615
rect 22450 -665 22500 -635
rect 22450 -685 22465 -665
rect 22485 -685 22500 -665
rect 22450 -715 22500 -685
rect 22450 -735 22465 -715
rect 22485 -735 22500 -715
rect 22450 -765 22500 -735
rect 22450 -785 22465 -765
rect 22485 -785 22500 -765
rect 21700 -860 21750 -850
rect 21700 -890 21710 -860
rect 21740 -890 21750 -860
rect 21700 -900 21750 -890
rect 22000 -860 22050 -850
rect 22000 -890 22010 -860
rect 22040 -890 22050 -860
rect 22000 -900 22050 -890
rect 22300 -860 22350 -850
rect 22300 -890 22310 -860
rect 22340 -890 22350 -860
rect 22300 -900 22350 -890
rect 22450 -860 22500 -785
rect 23350 -115 23400 65
rect 23350 -135 23365 -115
rect 23385 -135 23400 -115
rect 23350 -165 23400 -135
rect 23350 -185 23365 -165
rect 23385 -185 23400 -165
rect 23350 -215 23400 -185
rect 23350 -235 23365 -215
rect 23385 -235 23400 -215
rect 23350 -265 23400 -235
rect 23350 -285 23365 -265
rect 23385 -285 23400 -265
rect 23350 -315 23400 -285
rect 23350 -335 23365 -315
rect 23385 -335 23400 -315
rect 23350 -365 23400 -335
rect 23350 -385 23365 -365
rect 23385 -385 23400 -365
rect 23350 -415 23400 -385
rect 23350 -435 23365 -415
rect 23385 -435 23400 -415
rect 23350 -465 23400 -435
rect 23350 -485 23365 -465
rect 23385 -485 23400 -465
rect 23350 -515 23400 -485
rect 23350 -535 23365 -515
rect 23385 -535 23400 -515
rect 23350 -565 23400 -535
rect 23350 -585 23365 -565
rect 23385 -585 23400 -565
rect 23350 -615 23400 -585
rect 23350 -635 23365 -615
rect 23385 -635 23400 -615
rect 23350 -665 23400 -635
rect 23350 -685 23365 -665
rect 23385 -685 23400 -665
rect 23350 -715 23400 -685
rect 23350 -735 23365 -715
rect 23385 -735 23400 -715
rect 23350 -765 23400 -735
rect 23350 -785 23365 -765
rect 23385 -785 23400 -765
rect 22450 -890 22460 -860
rect 22490 -890 22500 -860
rect 21550 -985 21565 -965
rect 21585 -985 21600 -965
rect 21550 -1015 21600 -985
rect 21550 -1035 21565 -1015
rect 21585 -1035 21600 -1015
rect 21550 -1065 21600 -1035
rect 21550 -1085 21565 -1065
rect 21585 -1085 21600 -1065
rect 21550 -1115 21600 -1085
rect 21550 -1135 21565 -1115
rect 21585 -1135 21600 -1115
rect 21550 -1165 21600 -1135
rect 21550 -1185 21565 -1165
rect 21585 -1185 21600 -1165
rect 21550 -1215 21600 -1185
rect 21550 -1235 21565 -1215
rect 21585 -1235 21600 -1215
rect 21550 -1265 21600 -1235
rect 21550 -1285 21565 -1265
rect 21585 -1285 21600 -1265
rect 21550 -1315 21600 -1285
rect 21550 -1335 21565 -1315
rect 21585 -1335 21600 -1315
rect 21550 -1365 21600 -1335
rect 21550 -1385 21565 -1365
rect 21585 -1385 21600 -1365
rect 21550 -1415 21600 -1385
rect 21550 -1435 21565 -1415
rect 21585 -1435 21600 -1415
rect 21550 -1465 21600 -1435
rect 21550 -1485 21565 -1465
rect 21585 -1485 21600 -1465
rect 21550 -1515 21600 -1485
rect 21550 -1535 21565 -1515
rect 21585 -1535 21600 -1515
rect 21550 -1565 21600 -1535
rect 21550 -1585 21565 -1565
rect 21585 -1585 21600 -1565
rect 21550 -1615 21600 -1585
rect 21550 -1635 21565 -1615
rect 21585 -1635 21600 -1615
rect 21550 -1650 21600 -1635
rect 22450 -965 22500 -890
rect 22600 -860 22650 -850
rect 22600 -890 22610 -860
rect 22640 -890 22650 -860
rect 22600 -900 22650 -890
rect 22900 -860 22950 -850
rect 22900 -890 22910 -860
rect 22940 -890 22950 -860
rect 22900 -900 22950 -890
rect 23200 -860 23250 -850
rect 23200 -890 23210 -860
rect 23240 -890 23250 -860
rect 23200 -900 23250 -890
rect 22450 -985 22465 -965
rect 22485 -985 22500 -965
rect 22450 -1015 22500 -985
rect 22450 -1035 22465 -1015
rect 22485 -1035 22500 -1015
rect 22450 -1065 22500 -1035
rect 22450 -1085 22465 -1065
rect 22485 -1085 22500 -1065
rect 22450 -1115 22500 -1085
rect 22450 -1135 22465 -1115
rect 22485 -1135 22500 -1115
rect 22450 -1165 22500 -1135
rect 22450 -1185 22465 -1165
rect 22485 -1185 22500 -1165
rect 22450 -1215 22500 -1185
rect 22450 -1235 22465 -1215
rect 22485 -1235 22500 -1215
rect 22450 -1265 22500 -1235
rect 22450 -1285 22465 -1265
rect 22485 -1285 22500 -1265
rect 22450 -1315 22500 -1285
rect 22450 -1335 22465 -1315
rect 22485 -1335 22500 -1315
rect 22450 -1365 22500 -1335
rect 22450 -1385 22465 -1365
rect 22485 -1385 22500 -1365
rect 22450 -1415 22500 -1385
rect 22450 -1435 22465 -1415
rect 22485 -1435 22500 -1415
rect 22450 -1465 22500 -1435
rect 22450 -1485 22465 -1465
rect 22485 -1485 22500 -1465
rect 22450 -1515 22500 -1485
rect 22450 -1535 22465 -1515
rect 22485 -1535 22500 -1515
rect 22450 -1565 22500 -1535
rect 22450 -1585 22465 -1565
rect 22485 -1585 22500 -1565
rect 22450 -1615 22500 -1585
rect 22450 -1635 22465 -1615
rect 22485 -1635 22500 -1615
rect 22450 -1650 22500 -1635
rect 23350 -965 23400 -785
rect 24550 740 24600 910
rect 25750 1585 25800 1600
rect 25750 1565 25765 1585
rect 25785 1565 25800 1585
rect 25750 1535 25800 1565
rect 25750 1515 25765 1535
rect 25785 1515 25800 1535
rect 25750 1485 25800 1515
rect 25750 1465 25765 1485
rect 25785 1465 25800 1485
rect 25750 1435 25800 1465
rect 25750 1415 25765 1435
rect 25785 1415 25800 1435
rect 25750 1385 25800 1415
rect 25750 1365 25765 1385
rect 25785 1365 25800 1385
rect 25750 1335 25800 1365
rect 25750 1315 25765 1335
rect 25785 1315 25800 1335
rect 25750 1285 25800 1315
rect 25750 1265 25765 1285
rect 25785 1265 25800 1285
rect 25750 1235 25800 1265
rect 25750 1215 25765 1235
rect 25785 1215 25800 1235
rect 25750 1185 25800 1215
rect 25750 1165 25765 1185
rect 25785 1165 25800 1185
rect 25750 1135 25800 1165
rect 25750 1115 25765 1135
rect 25785 1115 25800 1135
rect 25750 1085 25800 1115
rect 25750 1065 25765 1085
rect 25785 1065 25800 1085
rect 25750 1035 25800 1065
rect 25750 1015 25765 1035
rect 25785 1015 25800 1035
rect 25750 985 25800 1015
rect 25750 965 25765 985
rect 25785 965 25800 985
rect 25750 935 25800 965
rect 25750 915 25765 935
rect 25785 915 25800 935
rect 24700 840 24750 850
rect 24700 810 24710 840
rect 24740 810 24750 840
rect 24700 800 24750 810
rect 25000 840 25050 850
rect 25000 810 25010 840
rect 25040 810 25050 840
rect 25000 800 25050 810
rect 25300 840 25350 850
rect 25300 810 25310 840
rect 25340 810 25350 840
rect 25300 800 25350 810
rect 25600 840 25650 850
rect 25600 810 25610 840
rect 25640 810 25650 840
rect 25600 800 25650 810
rect 25750 840 25800 915
rect 26650 1585 26700 1600
rect 26650 1565 26665 1585
rect 26685 1565 26700 1585
rect 26650 1535 26700 1565
rect 26650 1515 26665 1535
rect 26685 1515 26700 1535
rect 26650 1485 26700 1515
rect 26650 1465 26665 1485
rect 26685 1465 26700 1485
rect 26650 1435 26700 1465
rect 26650 1415 26665 1435
rect 26685 1415 26700 1435
rect 26650 1385 26700 1415
rect 26650 1365 26665 1385
rect 26685 1365 26700 1385
rect 26650 1335 26700 1365
rect 26650 1315 26665 1335
rect 26685 1315 26700 1335
rect 26650 1285 26700 1315
rect 26650 1265 26665 1285
rect 26685 1265 26700 1285
rect 26650 1235 26700 1265
rect 26650 1215 26665 1235
rect 26685 1215 26700 1235
rect 26650 1185 26700 1215
rect 26650 1165 26665 1185
rect 26685 1165 26700 1185
rect 26650 1135 26700 1165
rect 26650 1115 26665 1135
rect 26685 1115 26700 1135
rect 26650 1085 26700 1115
rect 26650 1065 26665 1085
rect 26685 1065 26700 1085
rect 26650 1035 26700 1065
rect 26650 1015 26665 1035
rect 26685 1015 26700 1035
rect 26650 985 26700 1015
rect 26650 965 26665 985
rect 26685 965 26700 985
rect 26650 935 26700 965
rect 26650 915 26665 935
rect 26685 915 26700 935
rect 25750 810 25760 840
rect 25790 810 25800 840
rect 24550 710 24560 740
rect 24590 710 24600 740
rect 24550 685 24600 710
rect 24550 665 24565 685
rect 24585 665 24600 685
rect 24550 640 24600 665
rect 24550 610 24560 640
rect 24590 610 24600 640
rect 24550 585 24600 610
rect 24550 565 24565 585
rect 24585 565 24600 585
rect 24550 540 24600 565
rect 24550 510 24560 540
rect 24590 510 24600 540
rect 24550 485 24600 510
rect 24550 465 24565 485
rect 24585 465 24600 485
rect 24550 440 24600 465
rect 24550 410 24560 440
rect 24590 410 24600 440
rect 24550 385 24600 410
rect 24550 365 24565 385
rect 24585 365 24600 385
rect 24550 340 24600 365
rect 24550 310 24560 340
rect 24590 310 24600 340
rect 24550 285 24600 310
rect 24550 265 24565 285
rect 24585 265 24600 285
rect 24550 240 24600 265
rect 24550 210 24560 240
rect 24590 210 24600 240
rect 24550 185 24600 210
rect 24550 165 24565 185
rect 24585 165 24600 185
rect 24550 140 24600 165
rect 24550 110 24560 140
rect 24590 110 24600 140
rect 24550 85 24600 110
rect 24550 65 24565 85
rect 24585 65 24600 85
rect 24550 -10 24600 65
rect 25750 735 25800 810
rect 25900 840 25950 850
rect 25900 810 25910 840
rect 25940 810 25950 840
rect 25900 800 25950 810
rect 26200 840 26250 850
rect 26200 810 26210 840
rect 26240 810 26250 840
rect 26200 800 26250 810
rect 26500 840 26550 850
rect 26500 810 26510 840
rect 26540 810 26550 840
rect 26500 800 26550 810
rect 26650 840 26700 915
rect 27550 1585 27600 1600
rect 27550 1565 27565 1585
rect 27585 1565 27600 1585
rect 27550 1535 27600 1565
rect 27550 1515 27565 1535
rect 27585 1515 27600 1535
rect 27550 1485 27600 1515
rect 27550 1465 27565 1485
rect 27585 1465 27600 1485
rect 27550 1435 27600 1465
rect 27550 1415 27565 1435
rect 27585 1415 27600 1435
rect 27550 1385 27600 1415
rect 27550 1365 27565 1385
rect 27585 1365 27600 1385
rect 27550 1335 27600 1365
rect 27550 1315 27565 1335
rect 27585 1315 27600 1335
rect 27550 1285 27600 1315
rect 27550 1265 27565 1285
rect 27585 1265 27600 1285
rect 27550 1235 27600 1265
rect 27550 1215 27565 1235
rect 27585 1215 27600 1235
rect 27550 1185 27600 1215
rect 27550 1165 27565 1185
rect 27585 1165 27600 1185
rect 27550 1135 27600 1165
rect 27550 1115 27565 1135
rect 27585 1115 27600 1135
rect 27550 1085 27600 1115
rect 27550 1065 27565 1085
rect 27585 1065 27600 1085
rect 27550 1035 27600 1065
rect 27550 1015 27565 1035
rect 27585 1015 27600 1035
rect 27550 985 27600 1015
rect 27550 965 27565 985
rect 27585 965 27600 985
rect 27550 935 27600 965
rect 27550 915 27565 935
rect 27585 915 27600 935
rect 26650 810 26660 840
rect 26690 810 26700 840
rect 25750 715 25765 735
rect 25785 715 25800 735
rect 25750 685 25800 715
rect 25750 665 25765 685
rect 25785 665 25800 685
rect 25750 635 25800 665
rect 25750 615 25765 635
rect 25785 615 25800 635
rect 25750 585 25800 615
rect 25750 565 25765 585
rect 25785 565 25800 585
rect 25750 535 25800 565
rect 25750 515 25765 535
rect 25785 515 25800 535
rect 25750 485 25800 515
rect 25750 465 25765 485
rect 25785 465 25800 485
rect 25750 435 25800 465
rect 25750 415 25765 435
rect 25785 415 25800 435
rect 25750 385 25800 415
rect 25750 365 25765 385
rect 25785 365 25800 385
rect 25750 335 25800 365
rect 25750 315 25765 335
rect 25785 315 25800 335
rect 25750 285 25800 315
rect 25750 265 25765 285
rect 25785 265 25800 285
rect 25750 235 25800 265
rect 25750 215 25765 235
rect 25785 215 25800 235
rect 25750 185 25800 215
rect 25750 165 25765 185
rect 25785 165 25800 185
rect 25750 135 25800 165
rect 25750 115 25765 135
rect 25785 115 25800 135
rect 25750 85 25800 115
rect 25750 65 25765 85
rect 25785 65 25800 85
rect 25750 50 25800 65
rect 26650 735 26700 810
rect 26800 840 26850 850
rect 26800 810 26810 840
rect 26840 810 26850 840
rect 26800 800 26850 810
rect 27100 840 27150 850
rect 27100 810 27110 840
rect 27140 810 27150 840
rect 27100 800 27150 810
rect 27400 840 27450 850
rect 27400 810 27410 840
rect 27440 810 27450 840
rect 27400 800 27450 810
rect 27550 840 27600 915
rect 28750 1585 28800 1660
rect 28750 1565 28765 1585
rect 28785 1565 28800 1585
rect 28750 1540 28800 1565
rect 28750 1510 28760 1540
rect 28790 1510 28800 1540
rect 28750 1485 28800 1510
rect 28750 1465 28765 1485
rect 28785 1465 28800 1485
rect 28750 1440 28800 1465
rect 28750 1410 28760 1440
rect 28790 1410 28800 1440
rect 28750 1385 28800 1410
rect 28750 1365 28765 1385
rect 28785 1365 28800 1385
rect 28750 1340 28800 1365
rect 28750 1310 28760 1340
rect 28790 1310 28800 1340
rect 28750 1285 28800 1310
rect 28750 1265 28765 1285
rect 28785 1265 28800 1285
rect 28750 1240 28800 1265
rect 28750 1210 28760 1240
rect 28790 1210 28800 1240
rect 28750 1185 28800 1210
rect 28750 1165 28765 1185
rect 28785 1165 28800 1185
rect 28750 1140 28800 1165
rect 28750 1110 28760 1140
rect 28790 1110 28800 1140
rect 28750 1085 28800 1110
rect 28750 1065 28765 1085
rect 28785 1065 28800 1085
rect 28750 1040 28800 1065
rect 28750 1010 28760 1040
rect 28790 1010 28800 1040
rect 28750 985 28800 1010
rect 28750 965 28765 985
rect 28785 965 28800 985
rect 28750 940 28800 965
rect 28750 910 28760 940
rect 28790 910 28800 940
rect 27550 810 27560 840
rect 27590 810 27600 840
rect 26650 715 26665 735
rect 26685 715 26700 735
rect 26650 685 26700 715
rect 26650 665 26665 685
rect 26685 665 26700 685
rect 26650 635 26700 665
rect 26650 615 26665 635
rect 26685 615 26700 635
rect 26650 585 26700 615
rect 26650 565 26665 585
rect 26685 565 26700 585
rect 26650 535 26700 565
rect 26650 515 26665 535
rect 26685 515 26700 535
rect 26650 485 26700 515
rect 26650 465 26665 485
rect 26685 465 26700 485
rect 26650 435 26700 465
rect 26650 415 26665 435
rect 26685 415 26700 435
rect 26650 385 26700 415
rect 26650 365 26665 385
rect 26685 365 26700 385
rect 26650 335 26700 365
rect 26650 315 26665 335
rect 26685 315 26700 335
rect 26650 285 26700 315
rect 26650 265 26665 285
rect 26685 265 26700 285
rect 26650 235 26700 265
rect 26650 215 26665 235
rect 26685 215 26700 235
rect 26650 185 26700 215
rect 26650 165 26665 185
rect 26685 165 26700 185
rect 26650 135 26700 165
rect 26650 115 26665 135
rect 26685 115 26700 135
rect 26650 85 26700 115
rect 26650 65 26665 85
rect 26685 65 26700 85
rect 26650 50 26700 65
rect 27550 735 27600 810
rect 27700 840 27750 850
rect 27700 810 27710 840
rect 27740 810 27750 840
rect 27700 800 27750 810
rect 28000 840 28050 850
rect 28000 810 28010 840
rect 28040 810 28050 840
rect 28000 800 28050 810
rect 28300 840 28350 850
rect 28300 810 28310 840
rect 28340 810 28350 840
rect 28300 800 28350 810
rect 28600 840 28650 850
rect 28600 810 28610 840
rect 28640 810 28650 840
rect 28600 800 28650 810
rect 27550 715 27565 735
rect 27585 715 27600 735
rect 27550 685 27600 715
rect 27550 665 27565 685
rect 27585 665 27600 685
rect 27550 635 27600 665
rect 27550 615 27565 635
rect 27585 615 27600 635
rect 27550 585 27600 615
rect 27550 565 27565 585
rect 27585 565 27600 585
rect 27550 535 27600 565
rect 27550 515 27565 535
rect 27585 515 27600 535
rect 27550 485 27600 515
rect 27550 465 27565 485
rect 27585 465 27600 485
rect 27550 435 27600 465
rect 27550 415 27565 435
rect 27585 415 27600 435
rect 27550 385 27600 415
rect 27550 365 27565 385
rect 27585 365 27600 385
rect 27550 335 27600 365
rect 27550 315 27565 335
rect 27585 315 27600 335
rect 27550 285 27600 315
rect 27550 265 27565 285
rect 27585 265 27600 285
rect 27550 235 27600 265
rect 27550 215 27565 235
rect 27585 215 27600 235
rect 27550 185 27600 215
rect 27550 165 27565 185
rect 27585 165 27600 185
rect 27550 135 27600 165
rect 27550 115 27565 135
rect 27585 115 27600 135
rect 27550 85 27600 115
rect 27550 65 27565 85
rect 27585 65 27600 85
rect 27550 50 27600 65
rect 28750 740 28800 910
rect 28750 710 28760 740
rect 28790 710 28800 740
rect 28750 685 28800 710
rect 28750 665 28765 685
rect 28785 665 28800 685
rect 28750 640 28800 665
rect 28750 610 28760 640
rect 28790 610 28800 640
rect 28750 585 28800 610
rect 28750 565 28765 585
rect 28785 565 28800 585
rect 28750 540 28800 565
rect 28750 510 28760 540
rect 28790 510 28800 540
rect 28750 485 28800 510
rect 28750 465 28765 485
rect 28785 465 28800 485
rect 28750 440 28800 465
rect 28750 410 28760 440
rect 28790 410 28800 440
rect 28750 385 28800 410
rect 28750 365 28765 385
rect 28785 365 28800 385
rect 28750 340 28800 365
rect 28750 310 28760 340
rect 28790 310 28800 340
rect 28750 285 28800 310
rect 28750 265 28765 285
rect 28785 265 28800 285
rect 28750 240 28800 265
rect 28750 210 28760 240
rect 28790 210 28800 240
rect 28750 185 28800 210
rect 28750 165 28765 185
rect 28785 165 28800 185
rect 28750 140 28800 165
rect 28750 110 28760 140
rect 28790 110 28800 140
rect 28750 85 28800 110
rect 28750 65 28765 85
rect 28785 65 28800 85
rect 24550 -40 24560 -10
rect 24590 -40 24600 -10
rect 24550 -115 24600 -40
rect 28750 -10 28800 65
rect 28750 -40 28760 -10
rect 28790 -40 28800 -10
rect 24550 -135 24565 -115
rect 24585 -135 24600 -115
rect 24550 -160 24600 -135
rect 24550 -190 24560 -160
rect 24590 -190 24600 -160
rect 24550 -215 24600 -190
rect 24550 -235 24565 -215
rect 24585 -235 24600 -215
rect 24550 -260 24600 -235
rect 24550 -290 24560 -260
rect 24590 -290 24600 -260
rect 24550 -315 24600 -290
rect 24550 -335 24565 -315
rect 24585 -335 24600 -315
rect 24550 -360 24600 -335
rect 24550 -390 24560 -360
rect 24590 -390 24600 -360
rect 24550 -415 24600 -390
rect 24550 -435 24565 -415
rect 24585 -435 24600 -415
rect 24550 -460 24600 -435
rect 24550 -490 24560 -460
rect 24590 -490 24600 -460
rect 24550 -515 24600 -490
rect 24550 -535 24565 -515
rect 24585 -535 24600 -515
rect 24550 -560 24600 -535
rect 24550 -590 24560 -560
rect 24590 -590 24600 -560
rect 24550 -615 24600 -590
rect 24550 -635 24565 -615
rect 24585 -635 24600 -615
rect 24550 -660 24600 -635
rect 24550 -690 24560 -660
rect 24590 -690 24600 -660
rect 24550 -715 24600 -690
rect 24550 -735 24565 -715
rect 24585 -735 24600 -715
rect 24550 -760 24600 -735
rect 24550 -790 24560 -760
rect 24590 -790 24600 -760
rect 23500 -860 23550 -850
rect 23500 -890 23510 -860
rect 23540 -890 23550 -860
rect 23500 -900 23550 -890
rect 23800 -860 23850 -850
rect 23800 -890 23810 -860
rect 23840 -890 23850 -860
rect 23800 -900 23850 -890
rect 24100 -860 24150 -850
rect 24100 -890 24110 -860
rect 24140 -890 24150 -860
rect 24100 -900 24150 -890
rect 24400 -860 24450 -850
rect 24400 -890 24410 -860
rect 24440 -890 24450 -860
rect 24400 -900 24450 -890
rect 23350 -985 23365 -965
rect 23385 -985 23400 -965
rect 23350 -1015 23400 -985
rect 23350 -1035 23365 -1015
rect 23385 -1035 23400 -1015
rect 23350 -1065 23400 -1035
rect 23350 -1085 23365 -1065
rect 23385 -1085 23400 -1065
rect 23350 -1115 23400 -1085
rect 23350 -1135 23365 -1115
rect 23385 -1135 23400 -1115
rect 23350 -1165 23400 -1135
rect 23350 -1185 23365 -1165
rect 23385 -1185 23400 -1165
rect 23350 -1215 23400 -1185
rect 23350 -1235 23365 -1215
rect 23385 -1235 23400 -1215
rect 23350 -1265 23400 -1235
rect 23350 -1285 23365 -1265
rect 23385 -1285 23400 -1265
rect 23350 -1315 23400 -1285
rect 23350 -1335 23365 -1315
rect 23385 -1335 23400 -1315
rect 23350 -1365 23400 -1335
rect 23350 -1385 23365 -1365
rect 23385 -1385 23400 -1365
rect 23350 -1415 23400 -1385
rect 23350 -1435 23365 -1415
rect 23385 -1435 23400 -1415
rect 23350 -1465 23400 -1435
rect 23350 -1485 23365 -1465
rect 23385 -1485 23400 -1465
rect 23350 -1515 23400 -1485
rect 23350 -1535 23365 -1515
rect 23385 -1535 23400 -1515
rect 23350 -1565 23400 -1535
rect 23350 -1585 23365 -1565
rect 23385 -1585 23400 -1565
rect 23350 -1615 23400 -1585
rect 23350 -1635 23365 -1615
rect 23385 -1635 23400 -1615
rect 23350 -1650 23400 -1635
rect 24550 -960 24600 -790
rect 25750 -115 25800 -100
rect 25750 -135 25765 -115
rect 25785 -135 25800 -115
rect 25750 -165 25800 -135
rect 25750 -185 25765 -165
rect 25785 -185 25800 -165
rect 25750 -215 25800 -185
rect 25750 -235 25765 -215
rect 25785 -235 25800 -215
rect 25750 -265 25800 -235
rect 25750 -285 25765 -265
rect 25785 -285 25800 -265
rect 25750 -315 25800 -285
rect 25750 -335 25765 -315
rect 25785 -335 25800 -315
rect 25750 -365 25800 -335
rect 25750 -385 25765 -365
rect 25785 -385 25800 -365
rect 25750 -415 25800 -385
rect 25750 -435 25765 -415
rect 25785 -435 25800 -415
rect 25750 -465 25800 -435
rect 25750 -485 25765 -465
rect 25785 -485 25800 -465
rect 25750 -515 25800 -485
rect 25750 -535 25765 -515
rect 25785 -535 25800 -515
rect 25750 -565 25800 -535
rect 25750 -585 25765 -565
rect 25785 -585 25800 -565
rect 25750 -615 25800 -585
rect 25750 -635 25765 -615
rect 25785 -635 25800 -615
rect 25750 -665 25800 -635
rect 25750 -685 25765 -665
rect 25785 -685 25800 -665
rect 25750 -715 25800 -685
rect 25750 -735 25765 -715
rect 25785 -735 25800 -715
rect 25750 -765 25800 -735
rect 25750 -785 25765 -765
rect 25785 -785 25800 -765
rect 24700 -860 24750 -850
rect 24700 -890 24710 -860
rect 24740 -890 24750 -860
rect 24700 -900 24750 -890
rect 25000 -860 25050 -850
rect 25000 -890 25010 -860
rect 25040 -890 25050 -860
rect 25000 -900 25050 -890
rect 25300 -860 25350 -850
rect 25300 -890 25310 -860
rect 25340 -890 25350 -860
rect 25300 -900 25350 -890
rect 25600 -860 25650 -850
rect 25600 -890 25610 -860
rect 25640 -890 25650 -860
rect 25600 -900 25650 -890
rect 25750 -860 25800 -785
rect 26650 -115 26700 -100
rect 26650 -135 26665 -115
rect 26685 -135 26700 -115
rect 26650 -165 26700 -135
rect 26650 -185 26665 -165
rect 26685 -185 26700 -165
rect 26650 -215 26700 -185
rect 26650 -235 26665 -215
rect 26685 -235 26700 -215
rect 26650 -265 26700 -235
rect 26650 -285 26665 -265
rect 26685 -285 26700 -265
rect 26650 -315 26700 -285
rect 26650 -335 26665 -315
rect 26685 -335 26700 -315
rect 26650 -365 26700 -335
rect 26650 -385 26665 -365
rect 26685 -385 26700 -365
rect 26650 -415 26700 -385
rect 26650 -435 26665 -415
rect 26685 -435 26700 -415
rect 26650 -465 26700 -435
rect 26650 -485 26665 -465
rect 26685 -485 26700 -465
rect 26650 -515 26700 -485
rect 26650 -535 26665 -515
rect 26685 -535 26700 -515
rect 26650 -565 26700 -535
rect 26650 -585 26665 -565
rect 26685 -585 26700 -565
rect 26650 -615 26700 -585
rect 26650 -635 26665 -615
rect 26685 -635 26700 -615
rect 26650 -665 26700 -635
rect 26650 -685 26665 -665
rect 26685 -685 26700 -665
rect 26650 -715 26700 -685
rect 26650 -735 26665 -715
rect 26685 -735 26700 -715
rect 26650 -765 26700 -735
rect 26650 -785 26665 -765
rect 26685 -785 26700 -765
rect 25750 -890 25760 -860
rect 25790 -890 25800 -860
rect 24550 -990 24560 -960
rect 24590 -990 24600 -960
rect 24550 -1015 24600 -990
rect 24550 -1035 24565 -1015
rect 24585 -1035 24600 -1015
rect 24550 -1060 24600 -1035
rect 24550 -1090 24560 -1060
rect 24590 -1090 24600 -1060
rect 24550 -1115 24600 -1090
rect 24550 -1135 24565 -1115
rect 24585 -1135 24600 -1115
rect 24550 -1160 24600 -1135
rect 24550 -1190 24560 -1160
rect 24590 -1190 24600 -1160
rect 24550 -1215 24600 -1190
rect 24550 -1235 24565 -1215
rect 24585 -1235 24600 -1215
rect 24550 -1260 24600 -1235
rect 24550 -1290 24560 -1260
rect 24590 -1290 24600 -1260
rect 24550 -1315 24600 -1290
rect 24550 -1335 24565 -1315
rect 24585 -1335 24600 -1315
rect 24550 -1360 24600 -1335
rect 24550 -1390 24560 -1360
rect 24590 -1390 24600 -1360
rect 24550 -1415 24600 -1390
rect 24550 -1435 24565 -1415
rect 24585 -1435 24600 -1415
rect 24550 -1460 24600 -1435
rect 24550 -1490 24560 -1460
rect 24590 -1490 24600 -1460
rect 24550 -1515 24600 -1490
rect 24550 -1535 24565 -1515
rect 24585 -1535 24600 -1515
rect 24550 -1560 24600 -1535
rect 24550 -1590 24560 -1560
rect 24590 -1590 24600 -1560
rect 24550 -1615 24600 -1590
rect 24550 -1635 24565 -1615
rect 24585 -1635 24600 -1615
rect 20350 -1740 20360 -1710
rect 20390 -1740 20400 -1710
rect 20350 -1750 20400 -1740
rect 24550 -1710 24600 -1635
rect 25750 -965 25800 -890
rect 25900 -860 25950 -850
rect 25900 -890 25910 -860
rect 25940 -890 25950 -860
rect 25900 -900 25950 -890
rect 26200 -860 26250 -850
rect 26200 -890 26210 -860
rect 26240 -890 26250 -860
rect 26200 -900 26250 -890
rect 26500 -860 26550 -850
rect 26500 -890 26510 -860
rect 26540 -890 26550 -860
rect 26500 -900 26550 -890
rect 26650 -860 26700 -785
rect 27550 -115 27600 -100
rect 27550 -135 27565 -115
rect 27585 -135 27600 -115
rect 27550 -165 27600 -135
rect 27550 -185 27565 -165
rect 27585 -185 27600 -165
rect 27550 -215 27600 -185
rect 27550 -235 27565 -215
rect 27585 -235 27600 -215
rect 27550 -265 27600 -235
rect 27550 -285 27565 -265
rect 27585 -285 27600 -265
rect 27550 -315 27600 -285
rect 27550 -335 27565 -315
rect 27585 -335 27600 -315
rect 27550 -365 27600 -335
rect 27550 -385 27565 -365
rect 27585 -385 27600 -365
rect 27550 -415 27600 -385
rect 27550 -435 27565 -415
rect 27585 -435 27600 -415
rect 27550 -465 27600 -435
rect 27550 -485 27565 -465
rect 27585 -485 27600 -465
rect 27550 -515 27600 -485
rect 27550 -535 27565 -515
rect 27585 -535 27600 -515
rect 27550 -565 27600 -535
rect 27550 -585 27565 -565
rect 27585 -585 27600 -565
rect 27550 -615 27600 -585
rect 27550 -635 27565 -615
rect 27585 -635 27600 -615
rect 27550 -665 27600 -635
rect 27550 -685 27565 -665
rect 27585 -685 27600 -665
rect 27550 -715 27600 -685
rect 27550 -735 27565 -715
rect 27585 -735 27600 -715
rect 27550 -765 27600 -735
rect 27550 -785 27565 -765
rect 27585 -785 27600 -765
rect 26650 -890 26660 -860
rect 26690 -890 26700 -860
rect 25750 -985 25765 -965
rect 25785 -985 25800 -965
rect 25750 -1015 25800 -985
rect 25750 -1035 25765 -1015
rect 25785 -1035 25800 -1015
rect 25750 -1065 25800 -1035
rect 25750 -1085 25765 -1065
rect 25785 -1085 25800 -1065
rect 25750 -1115 25800 -1085
rect 25750 -1135 25765 -1115
rect 25785 -1135 25800 -1115
rect 25750 -1165 25800 -1135
rect 25750 -1185 25765 -1165
rect 25785 -1185 25800 -1165
rect 25750 -1215 25800 -1185
rect 25750 -1235 25765 -1215
rect 25785 -1235 25800 -1215
rect 25750 -1265 25800 -1235
rect 25750 -1285 25765 -1265
rect 25785 -1285 25800 -1265
rect 25750 -1315 25800 -1285
rect 25750 -1335 25765 -1315
rect 25785 -1335 25800 -1315
rect 25750 -1365 25800 -1335
rect 25750 -1385 25765 -1365
rect 25785 -1385 25800 -1365
rect 25750 -1415 25800 -1385
rect 25750 -1435 25765 -1415
rect 25785 -1435 25800 -1415
rect 25750 -1465 25800 -1435
rect 25750 -1485 25765 -1465
rect 25785 -1485 25800 -1465
rect 25750 -1515 25800 -1485
rect 25750 -1535 25765 -1515
rect 25785 -1535 25800 -1515
rect 25750 -1565 25800 -1535
rect 25750 -1585 25765 -1565
rect 25785 -1585 25800 -1565
rect 25750 -1615 25800 -1585
rect 25750 -1635 25765 -1615
rect 25785 -1635 25800 -1615
rect 25750 -1650 25800 -1635
rect 26650 -965 26700 -890
rect 26800 -860 26850 -850
rect 26800 -890 26810 -860
rect 26840 -890 26850 -860
rect 26800 -900 26850 -890
rect 27100 -860 27150 -850
rect 27100 -890 27110 -860
rect 27140 -890 27150 -860
rect 27100 -900 27150 -890
rect 27400 -860 27450 -850
rect 27400 -890 27410 -860
rect 27440 -890 27450 -860
rect 27400 -900 27450 -890
rect 27550 -860 27600 -785
rect 28750 -115 28800 -40
rect 28750 -135 28765 -115
rect 28785 -135 28800 -115
rect 28750 -160 28800 -135
rect 28750 -190 28760 -160
rect 28790 -190 28800 -160
rect 28750 -215 28800 -190
rect 28750 -235 28765 -215
rect 28785 -235 28800 -215
rect 28750 -260 28800 -235
rect 28750 -290 28760 -260
rect 28790 -290 28800 -260
rect 28750 -315 28800 -290
rect 28750 -335 28765 -315
rect 28785 -335 28800 -315
rect 28750 -360 28800 -335
rect 28750 -390 28760 -360
rect 28790 -390 28800 -360
rect 28750 -415 28800 -390
rect 28750 -435 28765 -415
rect 28785 -435 28800 -415
rect 28750 -460 28800 -435
rect 28750 -490 28760 -460
rect 28790 -490 28800 -460
rect 28750 -515 28800 -490
rect 28750 -535 28765 -515
rect 28785 -535 28800 -515
rect 28750 -560 28800 -535
rect 28750 -590 28760 -560
rect 28790 -590 28800 -560
rect 28750 -615 28800 -590
rect 28750 -635 28765 -615
rect 28785 -635 28800 -615
rect 28750 -660 28800 -635
rect 28750 -690 28760 -660
rect 28790 -690 28800 -660
rect 28750 -715 28800 -690
rect 28750 -735 28765 -715
rect 28785 -735 28800 -715
rect 28750 -760 28800 -735
rect 28750 -790 28760 -760
rect 28790 -790 28800 -760
rect 27550 -890 27560 -860
rect 27590 -890 27600 -860
rect 26650 -985 26665 -965
rect 26685 -985 26700 -965
rect 26650 -1015 26700 -985
rect 26650 -1035 26665 -1015
rect 26685 -1035 26700 -1015
rect 26650 -1065 26700 -1035
rect 26650 -1085 26665 -1065
rect 26685 -1085 26700 -1065
rect 26650 -1115 26700 -1085
rect 26650 -1135 26665 -1115
rect 26685 -1135 26700 -1115
rect 26650 -1165 26700 -1135
rect 26650 -1185 26665 -1165
rect 26685 -1185 26700 -1165
rect 26650 -1215 26700 -1185
rect 26650 -1235 26665 -1215
rect 26685 -1235 26700 -1215
rect 26650 -1265 26700 -1235
rect 26650 -1285 26665 -1265
rect 26685 -1285 26700 -1265
rect 26650 -1315 26700 -1285
rect 26650 -1335 26665 -1315
rect 26685 -1335 26700 -1315
rect 26650 -1365 26700 -1335
rect 26650 -1385 26665 -1365
rect 26685 -1385 26700 -1365
rect 26650 -1415 26700 -1385
rect 26650 -1435 26665 -1415
rect 26685 -1435 26700 -1415
rect 26650 -1465 26700 -1435
rect 26650 -1485 26665 -1465
rect 26685 -1485 26700 -1465
rect 26650 -1515 26700 -1485
rect 26650 -1535 26665 -1515
rect 26685 -1535 26700 -1515
rect 26650 -1565 26700 -1535
rect 26650 -1585 26665 -1565
rect 26685 -1585 26700 -1565
rect 26650 -1615 26700 -1585
rect 26650 -1635 26665 -1615
rect 26685 -1635 26700 -1615
rect 26650 -1650 26700 -1635
rect 27550 -965 27600 -890
rect 27700 -860 27750 -850
rect 27700 -890 27710 -860
rect 27740 -890 27750 -860
rect 27700 -900 27750 -890
rect 28000 -860 28050 -850
rect 28000 -890 28010 -860
rect 28040 -890 28050 -860
rect 28000 -900 28050 -890
rect 28300 -860 28350 -850
rect 28300 -890 28310 -860
rect 28340 -890 28350 -860
rect 28300 -900 28350 -890
rect 28600 -860 28650 -850
rect 28600 -890 28610 -860
rect 28640 -890 28650 -860
rect 28600 -900 28650 -890
rect 27550 -985 27565 -965
rect 27585 -985 27600 -965
rect 27550 -1015 27600 -985
rect 27550 -1035 27565 -1015
rect 27585 -1035 27600 -1015
rect 27550 -1065 27600 -1035
rect 27550 -1085 27565 -1065
rect 27585 -1085 27600 -1065
rect 27550 -1115 27600 -1085
rect 27550 -1135 27565 -1115
rect 27585 -1135 27600 -1115
rect 27550 -1165 27600 -1135
rect 27550 -1185 27565 -1165
rect 27585 -1185 27600 -1165
rect 27550 -1215 27600 -1185
rect 27550 -1235 27565 -1215
rect 27585 -1235 27600 -1215
rect 27550 -1265 27600 -1235
rect 27550 -1285 27565 -1265
rect 27585 -1285 27600 -1265
rect 27550 -1315 27600 -1285
rect 27550 -1335 27565 -1315
rect 27585 -1335 27600 -1315
rect 27550 -1365 27600 -1335
rect 27550 -1385 27565 -1365
rect 27585 -1385 27600 -1365
rect 27550 -1415 27600 -1385
rect 27550 -1435 27565 -1415
rect 27585 -1435 27600 -1415
rect 27550 -1465 27600 -1435
rect 27550 -1485 27565 -1465
rect 27585 -1485 27600 -1465
rect 27550 -1515 27600 -1485
rect 27550 -1535 27565 -1515
rect 27585 -1535 27600 -1515
rect 27550 -1565 27600 -1535
rect 27550 -1585 27565 -1565
rect 27585 -1585 27600 -1565
rect 27550 -1615 27600 -1585
rect 27550 -1635 27565 -1615
rect 27585 -1635 27600 -1615
rect 27550 -1650 27600 -1635
rect 28750 -960 28800 -790
rect 28750 -990 28760 -960
rect 28790 -990 28800 -960
rect 28750 -1015 28800 -990
rect 28750 -1035 28765 -1015
rect 28785 -1035 28800 -1015
rect 28750 -1060 28800 -1035
rect 28750 -1090 28760 -1060
rect 28790 -1090 28800 -1060
rect 28750 -1115 28800 -1090
rect 28750 -1135 28765 -1115
rect 28785 -1135 28800 -1115
rect 28750 -1160 28800 -1135
rect 28750 -1190 28760 -1160
rect 28790 -1190 28800 -1160
rect 28750 -1215 28800 -1190
rect 28750 -1235 28765 -1215
rect 28785 -1235 28800 -1215
rect 28750 -1260 28800 -1235
rect 28750 -1290 28760 -1260
rect 28790 -1290 28800 -1260
rect 28750 -1315 28800 -1290
rect 28750 -1335 28765 -1315
rect 28785 -1335 28800 -1315
rect 28750 -1360 28800 -1335
rect 28750 -1390 28760 -1360
rect 28790 -1390 28800 -1360
rect 28750 -1415 28800 -1390
rect 28750 -1435 28765 -1415
rect 28785 -1435 28800 -1415
rect 28750 -1460 28800 -1435
rect 28750 -1490 28760 -1460
rect 28790 -1490 28800 -1460
rect 28750 -1515 28800 -1490
rect 28750 -1535 28765 -1515
rect 28785 -1535 28800 -1515
rect 28750 -1560 28800 -1535
rect 28750 -1590 28760 -1560
rect 28790 -1590 28800 -1560
rect 28750 -1615 28800 -1590
rect 28750 -1635 28765 -1615
rect 28785 -1635 28800 -1615
rect 24550 -1740 24560 -1710
rect 24590 -1740 24600 -1710
rect 24550 -1750 24600 -1740
rect 28750 -1710 28800 -1635
rect 28750 -1740 28760 -1710
rect 28790 -1740 28800 -1710
rect 28750 -1750 28800 -1740
<< via1 >>
rect -640 5585 -610 5590
rect -640 5565 -635 5585
rect -635 5565 -615 5585
rect -615 5565 -610 5585
rect -640 5560 -610 5565
rect -40 5560 -10 5590
rect -640 5435 -610 5440
rect -640 5415 -635 5435
rect -635 5415 -615 5435
rect -615 5415 -610 5435
rect -640 5410 -610 5415
rect -640 5335 -610 5340
rect -640 5315 -635 5335
rect -635 5315 -615 5335
rect -615 5315 -610 5335
rect -640 5310 -610 5315
rect -640 5235 -610 5240
rect -640 5215 -635 5235
rect -635 5215 -615 5235
rect -615 5215 -610 5235
rect -640 5210 -610 5215
rect -640 5135 -610 5140
rect -640 5115 -635 5135
rect -635 5115 -615 5135
rect -615 5115 -610 5135
rect -640 5110 -610 5115
rect -640 5035 -610 5040
rect -640 5015 -635 5035
rect -635 5015 -615 5035
rect -615 5015 -610 5035
rect -640 5010 -610 5015
rect 4160 5560 4190 5590
rect -490 4935 -460 4940
rect -490 4915 -485 4935
rect -485 4915 -465 4935
rect -465 4915 -460 4935
rect -490 4910 -460 4915
rect -340 4910 -310 4940
rect -190 4935 -160 4940
rect -190 4915 -185 4935
rect -185 4915 -165 4935
rect -165 4915 -160 4935
rect -190 4910 -160 4915
rect -640 4835 -610 4840
rect -640 4815 -635 4835
rect -635 4815 -615 4835
rect -615 4815 -610 4835
rect -640 4810 -610 4815
rect -640 4735 -610 4740
rect -640 4715 -635 4735
rect -635 4715 -615 4735
rect -615 4715 -610 4735
rect -640 4710 -610 4715
rect -640 4635 -610 4640
rect -640 4615 -635 4635
rect -635 4615 -615 4635
rect -615 4615 -610 4635
rect -640 4610 -610 4615
rect -640 4535 -610 4540
rect -640 4515 -635 4535
rect -635 4515 -615 4535
rect -615 4515 -610 4535
rect -640 4510 -610 4515
rect -640 4435 -610 4440
rect -640 4415 -635 4435
rect -635 4415 -615 4435
rect -615 4415 -610 4435
rect -640 4410 -610 4415
rect 110 4935 140 4940
rect 110 4915 115 4935
rect 115 4915 135 4935
rect 135 4915 140 4935
rect 110 4910 140 4915
rect 410 4935 440 4940
rect 410 4915 415 4935
rect 415 4915 435 4935
rect 435 4915 440 4935
rect 410 4910 440 4915
rect 710 4935 740 4940
rect 710 4915 715 4935
rect 715 4915 735 4935
rect 735 4915 740 4935
rect 710 4910 740 4915
rect 1010 4935 1040 4940
rect 1010 4915 1015 4935
rect 1015 4915 1035 4935
rect 1035 4915 1040 4935
rect 1010 4910 1040 4915
rect 1160 4910 1190 4940
rect 1310 4935 1340 4940
rect 1310 4915 1315 4935
rect 1315 4915 1335 4935
rect 1335 4915 1340 4935
rect 1310 4910 1340 4915
rect 1610 4935 1640 4940
rect 1610 4915 1615 4935
rect 1615 4915 1635 4935
rect 1635 4915 1640 4935
rect 1610 4910 1640 4915
rect -40 4810 -10 4840
rect -40 4735 -10 4740
rect -40 4715 -35 4735
rect -35 4715 -15 4735
rect -15 4715 -10 4735
rect -40 4710 -10 4715
rect -40 4635 -10 4640
rect -40 4615 -35 4635
rect -35 4615 -15 4635
rect -15 4615 -10 4635
rect -40 4610 -10 4615
rect -40 4535 -10 4540
rect -40 4515 -35 4535
rect -35 4515 -15 4535
rect -15 4515 -10 4535
rect -40 4510 -10 4515
rect -40 4435 -10 4440
rect -40 4415 -35 4435
rect -35 4415 -15 4435
rect -15 4415 -10 4435
rect -40 4410 -10 4415
rect -640 4285 -610 4290
rect -640 4265 -635 4285
rect -635 4265 -615 4285
rect -615 4265 -610 4285
rect -640 4260 -610 4265
rect 1910 4935 1940 4940
rect 1910 4915 1915 4935
rect 1915 4915 1935 4935
rect 1935 4915 1940 4935
rect 1910 4910 1940 4915
rect 2060 4910 2090 4940
rect 2210 4935 2240 4940
rect 2210 4915 2215 4935
rect 2215 4915 2235 4935
rect 2235 4915 2240 4935
rect 2210 4910 2240 4915
rect 8360 5585 8390 5590
rect 8360 5565 8365 5585
rect 8365 5565 8385 5585
rect 8385 5565 8390 5585
rect 8360 5560 8390 5565
rect 2510 4935 2540 4940
rect 2510 4915 2515 4935
rect 2515 4915 2535 4935
rect 2535 4915 2540 4935
rect 2510 4910 2540 4915
rect 2810 4935 2840 4940
rect 2810 4915 2815 4935
rect 2815 4915 2835 4935
rect 2835 4915 2840 4935
rect 2810 4910 2840 4915
rect 2960 4910 2990 4940
rect 3110 4935 3140 4940
rect 3110 4915 3115 4935
rect 3115 4915 3135 4935
rect 3135 4915 3140 4935
rect 3110 4910 3140 4915
rect 3410 4935 3440 4940
rect 3410 4915 3415 4935
rect 3415 4915 3435 4935
rect 3435 4915 3440 4935
rect 3410 4910 3440 4915
rect 3710 4935 3740 4940
rect 3710 4915 3715 4935
rect 3715 4915 3735 4935
rect 3735 4915 3740 4935
rect 3710 4910 3740 4915
rect 4010 4935 4040 4940
rect 4010 4915 4015 4935
rect 4015 4915 4035 4935
rect 4035 4915 4040 4935
rect 4010 4910 4040 4915
rect 4310 4935 4340 4940
rect 4310 4915 4315 4935
rect 4315 4915 4335 4935
rect 4335 4915 4340 4935
rect 4310 4910 4340 4915
rect 4610 4935 4640 4940
rect 4610 4915 4615 4935
rect 4615 4915 4635 4935
rect 4635 4915 4640 4935
rect 4610 4910 4640 4915
rect 4910 4935 4940 4940
rect 4910 4915 4915 4935
rect 4915 4915 4935 4935
rect 4935 4915 4940 4935
rect 4910 4910 4940 4915
rect 5210 4935 5240 4940
rect 5210 4915 5215 4935
rect 5215 4915 5235 4935
rect 5235 4915 5240 4935
rect 5210 4910 5240 4915
rect 5360 4910 5390 4940
rect 5510 4935 5540 4940
rect 5510 4915 5515 4935
rect 5515 4915 5535 4935
rect 5535 4915 5540 4935
rect 5510 4910 5540 4915
rect 5810 4935 5840 4940
rect 5810 4915 5815 4935
rect 5815 4915 5835 4935
rect 5835 4915 5840 4935
rect 5810 4910 5840 4915
rect 4160 4810 4190 4840
rect 4160 4735 4190 4740
rect 4160 4715 4165 4735
rect 4165 4715 4185 4735
rect 4185 4715 4190 4735
rect 4160 4710 4190 4715
rect 4160 4635 4190 4640
rect 4160 4615 4165 4635
rect 4165 4615 4185 4635
rect 4185 4615 4190 4635
rect 4160 4610 4190 4615
rect 4160 4535 4190 4540
rect 4160 4515 4165 4535
rect 4165 4515 4185 4535
rect 4185 4515 4190 4535
rect 4160 4510 4190 4515
rect 4160 4435 4190 4440
rect 4160 4415 4165 4435
rect 4165 4415 4185 4435
rect 4185 4415 4190 4435
rect 4160 4410 4190 4415
rect -40 4285 -10 4290
rect -40 4265 -35 4285
rect -35 4265 -15 4285
rect -15 4265 -10 4285
rect -40 4260 -10 4265
rect -640 4135 -610 4140
rect -640 4115 -635 4135
rect -635 4115 -615 4135
rect -615 4115 -610 4135
rect -640 4110 -610 4115
rect -640 4035 -610 4040
rect -640 4015 -635 4035
rect -635 4015 -615 4035
rect -615 4015 -610 4035
rect -640 4010 -610 4015
rect -640 3935 -610 3940
rect -640 3915 -635 3935
rect -635 3915 -615 3935
rect -615 3915 -610 3935
rect -640 3910 -610 3915
rect -640 3835 -610 3840
rect -640 3815 -635 3835
rect -635 3815 -615 3835
rect -615 3815 -610 3835
rect -640 3810 -610 3815
rect -640 3735 -610 3740
rect -640 3715 -635 3735
rect -635 3715 -615 3735
rect -615 3715 -610 3735
rect -640 3710 -610 3715
rect 6110 4935 6140 4940
rect 6110 4915 6115 4935
rect 6115 4915 6135 4935
rect 6135 4915 6140 4935
rect 6110 4910 6140 4915
rect 6260 4910 6290 4940
rect 6410 4935 6440 4940
rect 6410 4915 6415 4935
rect 6415 4915 6435 4935
rect 6435 4915 6440 4935
rect 6410 4910 6440 4915
rect 8660 5585 8690 5590
rect 8660 5565 8665 5585
rect 8665 5565 8685 5585
rect 8685 5565 8690 5585
rect 8660 5560 8690 5565
rect 8360 5435 8390 5440
rect 8360 5415 8365 5435
rect 8365 5415 8385 5435
rect 8385 5415 8390 5435
rect 8360 5410 8390 5415
rect 8360 5335 8390 5340
rect 8360 5315 8365 5335
rect 8365 5315 8385 5335
rect 8385 5315 8390 5335
rect 8360 5310 8390 5315
rect 8360 5235 8390 5240
rect 8360 5215 8365 5235
rect 8365 5215 8385 5235
rect 8385 5215 8390 5235
rect 8360 5210 8390 5215
rect 8360 5135 8390 5140
rect 8360 5115 8365 5135
rect 8365 5115 8385 5135
rect 8385 5115 8390 5135
rect 8360 5110 8390 5115
rect 8360 5035 8390 5040
rect 8360 5015 8365 5035
rect 8365 5015 8385 5035
rect 8385 5015 8390 5035
rect 8360 5010 8390 5015
rect 6710 4935 6740 4940
rect 6710 4915 6715 4935
rect 6715 4915 6735 4935
rect 6735 4915 6740 4935
rect 6710 4910 6740 4915
rect 7010 4935 7040 4940
rect 7010 4915 7015 4935
rect 7015 4915 7035 4935
rect 7035 4915 7040 4935
rect 7010 4910 7040 4915
rect 7160 4910 7190 4940
rect 7310 4935 7340 4940
rect 7310 4915 7315 4935
rect 7315 4915 7335 4935
rect 7335 4915 7340 4935
rect 7310 4910 7340 4915
rect 7610 4935 7640 4940
rect 7610 4915 7615 4935
rect 7615 4915 7635 4935
rect 7635 4915 7640 4935
rect 7610 4910 7640 4915
rect 7910 4935 7940 4940
rect 7910 4915 7915 4935
rect 7915 4915 7935 4935
rect 7935 4915 7940 4935
rect 7910 4910 7940 4915
rect 8210 4935 8240 4940
rect 8210 4915 8215 4935
rect 8215 4915 8235 4935
rect 8235 4915 8240 4935
rect 8210 4910 8240 4915
rect 8960 5585 8990 5590
rect 8960 5565 8965 5585
rect 8965 5565 8985 5585
rect 8985 5565 8990 5585
rect 8960 5560 8990 5565
rect 8660 5435 8690 5440
rect 8660 5415 8665 5435
rect 8665 5415 8685 5435
rect 8685 5415 8690 5435
rect 8660 5410 8690 5415
rect 8660 5335 8690 5340
rect 8660 5315 8665 5335
rect 8665 5315 8685 5335
rect 8685 5315 8690 5335
rect 8660 5310 8690 5315
rect 8660 5235 8690 5240
rect 8660 5215 8665 5235
rect 8665 5215 8685 5235
rect 8685 5215 8690 5235
rect 8660 5210 8690 5215
rect 8660 5135 8690 5140
rect 8660 5115 8665 5135
rect 8665 5115 8685 5135
rect 8685 5115 8690 5135
rect 8660 5110 8690 5115
rect 8660 5035 8690 5040
rect 8660 5015 8665 5035
rect 8665 5015 8685 5035
rect 8685 5015 8690 5035
rect 8660 5010 8690 5015
rect 8510 4935 8540 4940
rect 8510 4915 8515 4935
rect 8515 4915 8535 4935
rect 8535 4915 8540 4935
rect 8510 4910 8540 4915
rect 8360 4835 8390 4840
rect 8360 4815 8365 4835
rect 8365 4815 8385 4835
rect 8385 4815 8390 4835
rect 8360 4810 8390 4815
rect 8360 4735 8390 4740
rect 8360 4715 8365 4735
rect 8365 4715 8385 4735
rect 8385 4715 8390 4735
rect 8360 4710 8390 4715
rect 8360 4635 8390 4640
rect 8360 4615 8365 4635
rect 8365 4615 8385 4635
rect 8385 4615 8390 4635
rect 8360 4610 8390 4615
rect 8360 4535 8390 4540
rect 8360 4515 8365 4535
rect 8365 4515 8385 4535
rect 8385 4515 8390 4535
rect 8360 4510 8390 4515
rect 8360 4435 8390 4440
rect 8360 4415 8365 4435
rect 8365 4415 8385 4435
rect 8385 4415 8390 4435
rect 8360 4410 8390 4415
rect 4160 4285 4190 4290
rect 4160 4265 4165 4285
rect 4165 4265 4185 4285
rect 4185 4265 4190 4285
rect 4160 4260 4190 4265
rect -490 3635 -460 3640
rect -490 3615 -485 3635
rect -485 3615 -465 3635
rect -465 3615 -460 3635
rect -490 3610 -460 3615
rect -340 3610 -310 3640
rect -190 3635 -160 3640
rect -190 3615 -185 3635
rect -185 3615 -165 3635
rect -165 3615 -160 3635
rect -190 3610 -160 3615
rect -640 3535 -610 3540
rect -640 3515 -635 3535
rect -635 3515 -615 3535
rect -615 3515 -610 3535
rect -640 3510 -610 3515
rect -640 3435 -610 3440
rect -640 3415 -635 3435
rect -635 3415 -615 3435
rect -615 3415 -610 3435
rect -640 3410 -610 3415
rect -640 3335 -610 3340
rect -640 3315 -635 3335
rect -635 3315 -615 3335
rect -615 3315 -610 3335
rect -640 3310 -610 3315
rect -640 3235 -610 3240
rect -640 3215 -635 3235
rect -635 3215 -615 3235
rect -615 3215 -610 3235
rect -640 3210 -610 3215
rect -640 3135 -610 3140
rect -640 3115 -635 3135
rect -635 3115 -615 3135
rect -615 3115 -610 3135
rect -640 3110 -610 3115
rect 110 3635 140 3640
rect 110 3615 115 3635
rect 115 3615 135 3635
rect 135 3615 140 3635
rect 110 3610 140 3615
rect 410 3635 440 3640
rect 410 3615 415 3635
rect 415 3615 435 3635
rect 435 3615 440 3635
rect 410 3610 440 3615
rect -40 3510 -10 3540
rect -40 3435 -10 3440
rect -40 3415 -35 3435
rect -35 3415 -15 3435
rect -15 3415 -10 3435
rect -40 3410 -10 3415
rect -40 3335 -10 3340
rect -40 3315 -35 3335
rect -35 3315 -15 3335
rect -15 3315 -10 3335
rect -40 3310 -10 3315
rect -40 3235 -10 3240
rect -40 3215 -35 3235
rect -35 3215 -15 3235
rect -15 3215 -10 3235
rect -40 3210 -10 3215
rect -40 3135 -10 3140
rect -40 3115 -35 3135
rect -35 3115 -15 3135
rect -15 3115 -10 3135
rect -40 3110 -10 3115
rect -640 2985 -610 2990
rect -640 2965 -635 2985
rect -635 2965 -615 2985
rect -615 2965 -610 2985
rect -640 2960 -610 2965
rect 710 3635 740 3640
rect 710 3615 715 3635
rect 715 3615 735 3635
rect 735 3615 740 3635
rect 710 3610 740 3615
rect 1010 3635 1040 3640
rect 1010 3615 1015 3635
rect 1015 3615 1035 3635
rect 1035 3615 1040 3635
rect 1010 3610 1040 3615
rect 1160 3610 1190 3640
rect 1310 3635 1340 3640
rect 1310 3615 1315 3635
rect 1315 3615 1335 3635
rect 1335 3615 1340 3635
rect 1310 3610 1340 3615
rect 1610 3635 1640 3640
rect 1610 3615 1615 3635
rect 1615 3615 1635 3635
rect 1635 3615 1640 3635
rect 1610 3610 1640 3615
rect 1910 3635 1940 3640
rect 1910 3615 1915 3635
rect 1915 3615 1935 3635
rect 1935 3615 1940 3635
rect 1910 3610 1940 3615
rect 2060 3610 2090 3640
rect 2210 3635 2240 3640
rect 2210 3615 2215 3635
rect 2215 3615 2235 3635
rect 2235 3615 2240 3635
rect 2210 3610 2240 3615
rect 2510 3635 2540 3640
rect 2510 3615 2515 3635
rect 2515 3615 2535 3635
rect 2535 3615 2540 3635
rect 2510 3610 2540 3615
rect 2810 3635 2840 3640
rect 2810 3615 2815 3635
rect 2815 3615 2835 3635
rect 2835 3615 2840 3635
rect 2810 3610 2840 3615
rect 2960 3610 2990 3640
rect 3110 3635 3140 3640
rect 3110 3615 3115 3635
rect 3115 3615 3135 3635
rect 3135 3615 3140 3635
rect 3110 3610 3140 3615
rect 3410 3635 3440 3640
rect 3410 3615 3415 3635
rect 3415 3615 3435 3635
rect 3435 3615 3440 3635
rect 3410 3610 3440 3615
rect 9260 5585 9290 5590
rect 9260 5565 9265 5585
rect 9265 5565 9285 5585
rect 9285 5565 9290 5585
rect 9260 5560 9290 5565
rect 8960 5435 8990 5440
rect 8960 5415 8965 5435
rect 8965 5415 8985 5435
rect 8985 5415 8990 5435
rect 8960 5410 8990 5415
rect 8960 5335 8990 5340
rect 8960 5315 8965 5335
rect 8965 5315 8985 5335
rect 8985 5315 8990 5335
rect 8960 5310 8990 5315
rect 8960 5235 8990 5240
rect 8960 5215 8965 5235
rect 8965 5215 8985 5235
rect 8985 5215 8990 5235
rect 8960 5210 8990 5215
rect 8960 5135 8990 5140
rect 8960 5115 8965 5135
rect 8965 5115 8985 5135
rect 8985 5115 8990 5135
rect 8960 5110 8990 5115
rect 8960 5035 8990 5040
rect 8960 5015 8965 5035
rect 8965 5015 8985 5035
rect 8985 5015 8990 5035
rect 8960 5010 8990 5015
rect 8810 4935 8840 4940
rect 8810 4915 8815 4935
rect 8815 4915 8835 4935
rect 8835 4915 8840 4935
rect 8810 4910 8840 4915
rect 8660 4835 8690 4840
rect 8660 4815 8665 4835
rect 8665 4815 8685 4835
rect 8685 4815 8690 4835
rect 8660 4810 8690 4815
rect 8660 4735 8690 4740
rect 8660 4715 8665 4735
rect 8665 4715 8685 4735
rect 8685 4715 8690 4735
rect 8660 4710 8690 4715
rect 8660 4635 8690 4640
rect 8660 4615 8665 4635
rect 8665 4615 8685 4635
rect 8685 4615 8690 4635
rect 8660 4610 8690 4615
rect 8660 4535 8690 4540
rect 8660 4515 8665 4535
rect 8665 4515 8685 4535
rect 8685 4515 8690 4535
rect 8660 4510 8690 4515
rect 8660 4435 8690 4440
rect 8660 4415 8665 4435
rect 8665 4415 8685 4435
rect 8685 4415 8690 4435
rect 8660 4410 8690 4415
rect 8360 4285 8390 4290
rect 8360 4265 8365 4285
rect 8365 4265 8385 4285
rect 8385 4265 8390 4285
rect 8360 4260 8390 4265
rect 3710 3635 3740 3640
rect 3710 3615 3715 3635
rect 3715 3615 3735 3635
rect 3735 3615 3740 3635
rect 3710 3610 3740 3615
rect 4010 3635 4040 3640
rect 4010 3615 4015 3635
rect 4015 3615 4035 3635
rect 4035 3615 4040 3635
rect 4010 3610 4040 3615
rect 4310 3635 4340 3640
rect 4310 3615 4315 3635
rect 4315 3615 4335 3635
rect 4335 3615 4340 3635
rect 4310 3610 4340 3615
rect 4610 3635 4640 3640
rect 4610 3615 4615 3635
rect 4615 3615 4635 3635
rect 4635 3615 4640 3635
rect 4610 3610 4640 3615
rect 4160 3510 4190 3540
rect 4160 3435 4190 3440
rect 4160 3415 4165 3435
rect 4165 3415 4185 3435
rect 4185 3415 4190 3435
rect 4160 3410 4190 3415
rect 4160 3335 4190 3340
rect 4160 3315 4165 3335
rect 4165 3315 4185 3335
rect 4185 3315 4190 3335
rect 4160 3310 4190 3315
rect 4160 3235 4190 3240
rect 4160 3215 4165 3235
rect 4165 3215 4185 3235
rect 4185 3215 4190 3235
rect 4160 3210 4190 3215
rect 4160 3135 4190 3140
rect 4160 3115 4165 3135
rect 4165 3115 4185 3135
rect 4185 3115 4190 3135
rect 4160 3110 4190 3115
rect -40 2985 -10 2990
rect -40 2965 -35 2985
rect -35 2965 -15 2985
rect -15 2965 -10 2985
rect -40 2960 -10 2965
rect 4910 3635 4940 3640
rect 4910 3615 4915 3635
rect 4915 3615 4935 3635
rect 4935 3615 4940 3635
rect 4910 3610 4940 3615
rect 5210 3635 5240 3640
rect 5210 3615 5215 3635
rect 5215 3615 5235 3635
rect 5235 3615 5240 3635
rect 5210 3610 5240 3615
rect 5360 3610 5390 3640
rect 5510 3635 5540 3640
rect 5510 3615 5515 3635
rect 5515 3615 5535 3635
rect 5535 3615 5540 3635
rect 5510 3610 5540 3615
rect 5810 3635 5840 3640
rect 5810 3615 5815 3635
rect 5815 3615 5835 3635
rect 5835 3615 5840 3635
rect 5810 3610 5840 3615
rect 6110 3635 6140 3640
rect 6110 3615 6115 3635
rect 6115 3615 6135 3635
rect 6135 3615 6140 3635
rect 6110 3610 6140 3615
rect 6260 3610 6290 3640
rect 6410 3635 6440 3640
rect 6410 3615 6415 3635
rect 6415 3615 6435 3635
rect 6435 3615 6440 3635
rect 6410 3610 6440 3615
rect 6710 3635 6740 3640
rect 6710 3615 6715 3635
rect 6715 3615 6735 3635
rect 6735 3615 6740 3635
rect 6710 3610 6740 3615
rect 7010 3635 7040 3640
rect 7010 3615 7015 3635
rect 7015 3615 7035 3635
rect 7035 3615 7040 3635
rect 7010 3610 7040 3615
rect 7160 3610 7190 3640
rect 7310 3635 7340 3640
rect 7310 3615 7315 3635
rect 7315 3615 7335 3635
rect 7335 3615 7340 3635
rect 7310 3610 7340 3615
rect 7610 3635 7640 3640
rect 7610 3615 7615 3635
rect 7615 3615 7635 3635
rect 7635 3615 7640 3635
rect 7610 3610 7640 3615
rect 9560 5585 9590 5590
rect 9560 5565 9565 5585
rect 9565 5565 9585 5585
rect 9585 5565 9590 5585
rect 9560 5560 9590 5565
rect 9260 5435 9290 5440
rect 9260 5415 9265 5435
rect 9265 5415 9285 5435
rect 9285 5415 9290 5435
rect 9260 5410 9290 5415
rect 9260 5335 9290 5340
rect 9260 5315 9265 5335
rect 9265 5315 9285 5335
rect 9285 5315 9290 5335
rect 9260 5310 9290 5315
rect 9260 5235 9290 5240
rect 9260 5215 9265 5235
rect 9265 5215 9285 5235
rect 9285 5215 9290 5235
rect 9260 5210 9290 5215
rect 9260 5135 9290 5140
rect 9260 5115 9265 5135
rect 9265 5115 9285 5135
rect 9285 5115 9290 5135
rect 9260 5110 9290 5115
rect 9260 5035 9290 5040
rect 9260 5015 9265 5035
rect 9265 5015 9285 5035
rect 9285 5015 9290 5035
rect 9260 5010 9290 5015
rect 9110 4935 9140 4940
rect 9110 4915 9115 4935
rect 9115 4915 9135 4935
rect 9135 4915 9140 4935
rect 9110 4910 9140 4915
rect 8960 4835 8990 4840
rect 8960 4815 8965 4835
rect 8965 4815 8985 4835
rect 8985 4815 8990 4835
rect 8960 4810 8990 4815
rect 8960 4735 8990 4740
rect 8960 4715 8965 4735
rect 8965 4715 8985 4735
rect 8985 4715 8990 4735
rect 8960 4710 8990 4715
rect 8960 4635 8990 4640
rect 8960 4615 8965 4635
rect 8965 4615 8985 4635
rect 8985 4615 8990 4635
rect 8960 4610 8990 4615
rect 8960 4535 8990 4540
rect 8960 4515 8965 4535
rect 8965 4515 8985 4535
rect 8985 4515 8990 4535
rect 8960 4510 8990 4515
rect 8960 4435 8990 4440
rect 8960 4415 8965 4435
rect 8965 4415 8985 4435
rect 8985 4415 8990 4435
rect 8960 4410 8990 4415
rect 8660 4285 8690 4290
rect 8660 4265 8665 4285
rect 8665 4265 8685 4285
rect 8685 4265 8690 4285
rect 8660 4260 8690 4265
rect 8360 4135 8390 4140
rect 8360 4115 8365 4135
rect 8365 4115 8385 4135
rect 8385 4115 8390 4135
rect 8360 4110 8390 4115
rect 8360 4035 8390 4040
rect 8360 4015 8365 4035
rect 8365 4015 8385 4035
rect 8385 4015 8390 4035
rect 8360 4010 8390 4015
rect 8360 3935 8390 3940
rect 8360 3915 8365 3935
rect 8365 3915 8385 3935
rect 8385 3915 8390 3935
rect 8360 3910 8390 3915
rect 8360 3835 8390 3840
rect 8360 3815 8365 3835
rect 8365 3815 8385 3835
rect 8385 3815 8390 3835
rect 8360 3810 8390 3815
rect 8360 3735 8390 3740
rect 8360 3715 8365 3735
rect 8365 3715 8385 3735
rect 8385 3715 8390 3735
rect 8360 3710 8390 3715
rect 7910 3635 7940 3640
rect 7910 3615 7915 3635
rect 7915 3615 7935 3635
rect 7935 3615 7940 3635
rect 7910 3610 7940 3615
rect 8210 3635 8240 3640
rect 8210 3615 8215 3635
rect 8215 3615 8235 3635
rect 8235 3615 8240 3635
rect 8210 3610 8240 3615
rect 9860 5585 9890 5590
rect 9860 5565 9865 5585
rect 9865 5565 9885 5585
rect 9885 5565 9890 5585
rect 9860 5560 9890 5565
rect 9560 5435 9590 5440
rect 9560 5415 9565 5435
rect 9565 5415 9585 5435
rect 9585 5415 9590 5435
rect 9560 5410 9590 5415
rect 9560 5335 9590 5340
rect 9560 5315 9565 5335
rect 9565 5315 9585 5335
rect 9585 5315 9590 5335
rect 9560 5310 9590 5315
rect 9560 5235 9590 5240
rect 9560 5215 9565 5235
rect 9565 5215 9585 5235
rect 9585 5215 9590 5235
rect 9560 5210 9590 5215
rect 9560 5135 9590 5140
rect 9560 5115 9565 5135
rect 9565 5115 9585 5135
rect 9585 5115 9590 5135
rect 9560 5110 9590 5115
rect 9560 5035 9590 5040
rect 9560 5015 9565 5035
rect 9565 5015 9585 5035
rect 9585 5015 9590 5035
rect 9560 5010 9590 5015
rect 9410 4935 9440 4940
rect 9410 4915 9415 4935
rect 9415 4915 9435 4935
rect 9435 4915 9440 4935
rect 9410 4910 9440 4915
rect 9260 4835 9290 4840
rect 9260 4815 9265 4835
rect 9265 4815 9285 4835
rect 9285 4815 9290 4835
rect 9260 4810 9290 4815
rect 9260 4735 9290 4740
rect 9260 4715 9265 4735
rect 9265 4715 9285 4735
rect 9285 4715 9290 4735
rect 9260 4710 9290 4715
rect 9260 4635 9290 4640
rect 9260 4615 9265 4635
rect 9265 4615 9285 4635
rect 9285 4615 9290 4635
rect 9260 4610 9290 4615
rect 9260 4535 9290 4540
rect 9260 4515 9265 4535
rect 9265 4515 9285 4535
rect 9285 4515 9290 4535
rect 9260 4510 9290 4515
rect 9260 4435 9290 4440
rect 9260 4415 9265 4435
rect 9265 4415 9285 4435
rect 9285 4415 9290 4435
rect 9260 4410 9290 4415
rect 8960 4285 8990 4290
rect 8960 4265 8965 4285
rect 8965 4265 8985 4285
rect 8985 4265 8990 4285
rect 8960 4260 8990 4265
rect 8660 4135 8690 4140
rect 8660 4115 8665 4135
rect 8665 4115 8685 4135
rect 8685 4115 8690 4135
rect 8660 4110 8690 4115
rect 8660 4035 8690 4040
rect 8660 4015 8665 4035
rect 8665 4015 8685 4035
rect 8685 4015 8690 4035
rect 8660 4010 8690 4015
rect 8660 3935 8690 3940
rect 8660 3915 8665 3935
rect 8665 3915 8685 3935
rect 8685 3915 8690 3935
rect 8660 3910 8690 3915
rect 8660 3835 8690 3840
rect 8660 3815 8665 3835
rect 8665 3815 8685 3835
rect 8685 3815 8690 3835
rect 8660 3810 8690 3815
rect 8660 3735 8690 3740
rect 8660 3715 8665 3735
rect 8665 3715 8685 3735
rect 8685 3715 8690 3735
rect 8660 3710 8690 3715
rect 8510 3635 8540 3640
rect 8510 3615 8515 3635
rect 8515 3615 8535 3635
rect 8535 3615 8540 3635
rect 8510 3610 8540 3615
rect 8360 3535 8390 3540
rect 8360 3515 8365 3535
rect 8365 3515 8385 3535
rect 8385 3515 8390 3535
rect 8360 3510 8390 3515
rect 8360 3435 8390 3440
rect 8360 3415 8365 3435
rect 8365 3415 8385 3435
rect 8385 3415 8390 3435
rect 8360 3410 8390 3415
rect 8360 3335 8390 3340
rect 8360 3315 8365 3335
rect 8365 3315 8385 3335
rect 8385 3315 8390 3335
rect 8360 3310 8390 3315
rect 8360 3235 8390 3240
rect 8360 3215 8365 3235
rect 8365 3215 8385 3235
rect 8385 3215 8390 3235
rect 8360 3210 8390 3215
rect 8360 3135 8390 3140
rect 8360 3115 8365 3135
rect 8365 3115 8385 3135
rect 8385 3115 8390 3135
rect 8360 3110 8390 3115
rect 4160 2985 4190 2990
rect 4160 2965 4165 2985
rect 4165 2965 4185 2985
rect 4185 2965 4190 2985
rect 4160 2960 4190 2965
rect 10160 5585 10190 5590
rect 10160 5565 10165 5585
rect 10165 5565 10185 5585
rect 10185 5565 10190 5585
rect 10160 5560 10190 5565
rect 9860 5435 9890 5440
rect 9860 5415 9865 5435
rect 9865 5415 9885 5435
rect 9885 5415 9890 5435
rect 9860 5410 9890 5415
rect 9860 5335 9890 5340
rect 9860 5315 9865 5335
rect 9865 5315 9885 5335
rect 9885 5315 9890 5335
rect 9860 5310 9890 5315
rect 9860 5235 9890 5240
rect 9860 5215 9865 5235
rect 9865 5215 9885 5235
rect 9885 5215 9890 5235
rect 9860 5210 9890 5215
rect 9860 5135 9890 5140
rect 9860 5115 9865 5135
rect 9865 5115 9885 5135
rect 9885 5115 9890 5135
rect 9860 5110 9890 5115
rect 9860 5035 9890 5040
rect 9860 5015 9865 5035
rect 9865 5015 9885 5035
rect 9885 5015 9890 5035
rect 9860 5010 9890 5015
rect 9710 4935 9740 4940
rect 9710 4915 9715 4935
rect 9715 4915 9735 4935
rect 9735 4915 9740 4935
rect 9710 4910 9740 4915
rect 9560 4835 9590 4840
rect 9560 4815 9565 4835
rect 9565 4815 9585 4835
rect 9585 4815 9590 4835
rect 9560 4810 9590 4815
rect 9560 4735 9590 4740
rect 9560 4715 9565 4735
rect 9565 4715 9585 4735
rect 9585 4715 9590 4735
rect 9560 4710 9590 4715
rect 9560 4635 9590 4640
rect 9560 4615 9565 4635
rect 9565 4615 9585 4635
rect 9585 4615 9590 4635
rect 9560 4610 9590 4615
rect 9560 4535 9590 4540
rect 9560 4515 9565 4535
rect 9565 4515 9585 4535
rect 9585 4515 9590 4535
rect 9560 4510 9590 4515
rect 9560 4435 9590 4440
rect 9560 4415 9565 4435
rect 9565 4415 9585 4435
rect 9585 4415 9590 4435
rect 9560 4410 9590 4415
rect 9260 4285 9290 4290
rect 9260 4265 9265 4285
rect 9265 4265 9285 4285
rect 9285 4265 9290 4285
rect 9260 4260 9290 4265
rect 8960 4135 8990 4140
rect 8960 4115 8965 4135
rect 8965 4115 8985 4135
rect 8985 4115 8990 4135
rect 8960 4110 8990 4115
rect 8960 4035 8990 4040
rect 8960 4015 8965 4035
rect 8965 4015 8985 4035
rect 8985 4015 8990 4035
rect 8960 4010 8990 4015
rect 8960 3935 8990 3940
rect 8960 3915 8965 3935
rect 8965 3915 8985 3935
rect 8985 3915 8990 3935
rect 8960 3910 8990 3915
rect 8960 3835 8990 3840
rect 8960 3815 8965 3835
rect 8965 3815 8985 3835
rect 8985 3815 8990 3835
rect 8960 3810 8990 3815
rect 8960 3735 8990 3740
rect 8960 3715 8965 3735
rect 8965 3715 8985 3735
rect 8985 3715 8990 3735
rect 8960 3710 8990 3715
rect 8810 3635 8840 3640
rect 8810 3615 8815 3635
rect 8815 3615 8835 3635
rect 8835 3615 8840 3635
rect 8810 3610 8840 3615
rect 8660 3535 8690 3540
rect 8660 3515 8665 3535
rect 8665 3515 8685 3535
rect 8685 3515 8690 3535
rect 8660 3510 8690 3515
rect 8660 3435 8690 3440
rect 8660 3415 8665 3435
rect 8665 3415 8685 3435
rect 8685 3415 8690 3435
rect 8660 3410 8690 3415
rect 8660 3335 8690 3340
rect 8660 3315 8665 3335
rect 8665 3315 8685 3335
rect 8685 3315 8690 3335
rect 8660 3310 8690 3315
rect 8660 3235 8690 3240
rect 8660 3215 8665 3235
rect 8665 3215 8685 3235
rect 8685 3215 8690 3235
rect 8660 3210 8690 3215
rect 8660 3135 8690 3140
rect 8660 3115 8665 3135
rect 8665 3115 8685 3135
rect 8685 3115 8690 3135
rect 8660 3110 8690 3115
rect 8360 2985 8390 2990
rect 8360 2965 8365 2985
rect 8365 2965 8385 2985
rect 8385 2965 8390 2985
rect 8360 2960 8390 2965
rect 10460 5585 10490 5590
rect 10460 5565 10465 5585
rect 10465 5565 10485 5585
rect 10485 5565 10490 5585
rect 10460 5560 10490 5565
rect 10160 5435 10190 5440
rect 10160 5415 10165 5435
rect 10165 5415 10185 5435
rect 10185 5415 10190 5435
rect 10160 5410 10190 5415
rect 10160 5335 10190 5340
rect 10160 5315 10165 5335
rect 10165 5315 10185 5335
rect 10185 5315 10190 5335
rect 10160 5310 10190 5315
rect 10160 5235 10190 5240
rect 10160 5215 10165 5235
rect 10165 5215 10185 5235
rect 10185 5215 10190 5235
rect 10160 5210 10190 5215
rect 10160 5135 10190 5140
rect 10160 5115 10165 5135
rect 10165 5115 10185 5135
rect 10185 5115 10190 5135
rect 10160 5110 10190 5115
rect 10160 5035 10190 5040
rect 10160 5015 10165 5035
rect 10165 5015 10185 5035
rect 10185 5015 10190 5035
rect 10160 5010 10190 5015
rect 10010 4935 10040 4940
rect 10010 4915 10015 4935
rect 10015 4915 10035 4935
rect 10035 4915 10040 4935
rect 10010 4910 10040 4915
rect 9860 4835 9890 4840
rect 9860 4815 9865 4835
rect 9865 4815 9885 4835
rect 9885 4815 9890 4835
rect 9860 4810 9890 4815
rect 9860 4735 9890 4740
rect 9860 4715 9865 4735
rect 9865 4715 9885 4735
rect 9885 4715 9890 4735
rect 9860 4710 9890 4715
rect 9860 4635 9890 4640
rect 9860 4615 9865 4635
rect 9865 4615 9885 4635
rect 9885 4615 9890 4635
rect 9860 4610 9890 4615
rect 9860 4535 9890 4540
rect 9860 4515 9865 4535
rect 9865 4515 9885 4535
rect 9885 4515 9890 4535
rect 9860 4510 9890 4515
rect 9860 4435 9890 4440
rect 9860 4415 9865 4435
rect 9865 4415 9885 4435
rect 9885 4415 9890 4435
rect 9860 4410 9890 4415
rect 9560 4285 9590 4290
rect 9560 4265 9565 4285
rect 9565 4265 9585 4285
rect 9585 4265 9590 4285
rect 9560 4260 9590 4265
rect 9260 4135 9290 4140
rect 9260 4115 9265 4135
rect 9265 4115 9285 4135
rect 9285 4115 9290 4135
rect 9260 4110 9290 4115
rect 9260 4035 9290 4040
rect 9260 4015 9265 4035
rect 9265 4015 9285 4035
rect 9285 4015 9290 4035
rect 9260 4010 9290 4015
rect 9260 3935 9290 3940
rect 9260 3915 9265 3935
rect 9265 3915 9285 3935
rect 9285 3915 9290 3935
rect 9260 3910 9290 3915
rect 9260 3835 9290 3840
rect 9260 3815 9265 3835
rect 9265 3815 9285 3835
rect 9285 3815 9290 3835
rect 9260 3810 9290 3815
rect 9260 3735 9290 3740
rect 9260 3715 9265 3735
rect 9265 3715 9285 3735
rect 9285 3715 9290 3735
rect 9260 3710 9290 3715
rect 9110 3635 9140 3640
rect 9110 3615 9115 3635
rect 9115 3615 9135 3635
rect 9135 3615 9140 3635
rect 9110 3610 9140 3615
rect 8960 3535 8990 3540
rect 8960 3515 8965 3535
rect 8965 3515 8985 3535
rect 8985 3515 8990 3535
rect 8960 3510 8990 3515
rect 8960 3435 8990 3440
rect 8960 3415 8965 3435
rect 8965 3415 8985 3435
rect 8985 3415 8990 3435
rect 8960 3410 8990 3415
rect 8960 3335 8990 3340
rect 8960 3315 8965 3335
rect 8965 3315 8985 3335
rect 8985 3315 8990 3335
rect 8960 3310 8990 3315
rect 8960 3235 8990 3240
rect 8960 3215 8965 3235
rect 8965 3215 8985 3235
rect 8985 3215 8990 3235
rect 8960 3210 8990 3215
rect 8960 3135 8990 3140
rect 8960 3115 8965 3135
rect 8965 3115 8985 3135
rect 8985 3115 8990 3135
rect 8960 3110 8990 3115
rect 8660 2985 8690 2990
rect 8660 2965 8665 2985
rect 8665 2965 8685 2985
rect 8685 2965 8690 2985
rect 8660 2960 8690 2965
rect 10760 5585 10790 5590
rect 10760 5565 10765 5585
rect 10765 5565 10785 5585
rect 10785 5565 10790 5585
rect 10760 5560 10790 5565
rect 10460 5435 10490 5440
rect 10460 5415 10465 5435
rect 10465 5415 10485 5435
rect 10485 5415 10490 5435
rect 10460 5410 10490 5415
rect 10460 5335 10490 5340
rect 10460 5315 10465 5335
rect 10465 5315 10485 5335
rect 10485 5315 10490 5335
rect 10460 5310 10490 5315
rect 10460 5235 10490 5240
rect 10460 5215 10465 5235
rect 10465 5215 10485 5235
rect 10485 5215 10490 5235
rect 10460 5210 10490 5215
rect 10460 5135 10490 5140
rect 10460 5115 10465 5135
rect 10465 5115 10485 5135
rect 10485 5115 10490 5135
rect 10460 5110 10490 5115
rect 10460 5035 10490 5040
rect 10460 5015 10465 5035
rect 10465 5015 10485 5035
rect 10485 5015 10490 5035
rect 10460 5010 10490 5015
rect 10310 4935 10340 4940
rect 10310 4915 10315 4935
rect 10315 4915 10335 4935
rect 10335 4915 10340 4935
rect 10310 4910 10340 4915
rect 10160 4835 10190 4840
rect 10160 4815 10165 4835
rect 10165 4815 10185 4835
rect 10185 4815 10190 4835
rect 10160 4810 10190 4815
rect 10160 4735 10190 4740
rect 10160 4715 10165 4735
rect 10165 4715 10185 4735
rect 10185 4715 10190 4735
rect 10160 4710 10190 4715
rect 10160 4635 10190 4640
rect 10160 4615 10165 4635
rect 10165 4615 10185 4635
rect 10185 4615 10190 4635
rect 10160 4610 10190 4615
rect 10160 4535 10190 4540
rect 10160 4515 10165 4535
rect 10165 4515 10185 4535
rect 10185 4515 10190 4535
rect 10160 4510 10190 4515
rect 10160 4435 10190 4440
rect 10160 4415 10165 4435
rect 10165 4415 10185 4435
rect 10185 4415 10190 4435
rect 10160 4410 10190 4415
rect 9860 4285 9890 4290
rect 9860 4265 9865 4285
rect 9865 4265 9885 4285
rect 9885 4265 9890 4285
rect 9860 4260 9890 4265
rect 9560 4135 9590 4140
rect 9560 4115 9565 4135
rect 9565 4115 9585 4135
rect 9585 4115 9590 4135
rect 9560 4110 9590 4115
rect 9560 4035 9590 4040
rect 9560 4015 9565 4035
rect 9565 4015 9585 4035
rect 9585 4015 9590 4035
rect 9560 4010 9590 4015
rect 9560 3935 9590 3940
rect 9560 3915 9565 3935
rect 9565 3915 9585 3935
rect 9585 3915 9590 3935
rect 9560 3910 9590 3915
rect 9560 3835 9590 3840
rect 9560 3815 9565 3835
rect 9565 3815 9585 3835
rect 9585 3815 9590 3835
rect 9560 3810 9590 3815
rect 9560 3735 9590 3740
rect 9560 3715 9565 3735
rect 9565 3715 9585 3735
rect 9585 3715 9590 3735
rect 9560 3710 9590 3715
rect 9410 3635 9440 3640
rect 9410 3615 9415 3635
rect 9415 3615 9435 3635
rect 9435 3615 9440 3635
rect 9410 3610 9440 3615
rect 9260 3535 9290 3540
rect 9260 3515 9265 3535
rect 9265 3515 9285 3535
rect 9285 3515 9290 3535
rect 9260 3510 9290 3515
rect 9260 3435 9290 3440
rect 9260 3415 9265 3435
rect 9265 3415 9285 3435
rect 9285 3415 9290 3435
rect 9260 3410 9290 3415
rect 9260 3335 9290 3340
rect 9260 3315 9265 3335
rect 9265 3315 9285 3335
rect 9285 3315 9290 3335
rect 9260 3310 9290 3315
rect 9260 3235 9290 3240
rect 9260 3215 9265 3235
rect 9265 3215 9285 3235
rect 9285 3215 9290 3235
rect 9260 3210 9290 3215
rect 9260 3135 9290 3140
rect 9260 3115 9265 3135
rect 9265 3115 9285 3135
rect 9285 3115 9290 3135
rect 9260 3110 9290 3115
rect 8960 2985 8990 2990
rect 8960 2965 8965 2985
rect 8965 2965 8985 2985
rect 8985 2965 8990 2985
rect 8960 2960 8990 2965
rect 11960 5585 11990 5590
rect 11960 5565 11965 5585
rect 11965 5565 11985 5585
rect 11985 5565 11990 5585
rect 11960 5560 11990 5565
rect 10760 5435 10790 5440
rect 10760 5415 10765 5435
rect 10765 5415 10785 5435
rect 10785 5415 10790 5435
rect 10760 5410 10790 5415
rect 10760 5335 10790 5340
rect 10760 5315 10765 5335
rect 10765 5315 10785 5335
rect 10785 5315 10790 5335
rect 10760 5310 10790 5315
rect 10760 5235 10790 5240
rect 10760 5215 10765 5235
rect 10765 5215 10785 5235
rect 10785 5215 10790 5235
rect 10760 5210 10790 5215
rect 10760 5135 10790 5140
rect 10760 5115 10765 5135
rect 10765 5115 10785 5135
rect 10785 5115 10790 5135
rect 10760 5110 10790 5115
rect 10760 5035 10790 5040
rect 10760 5015 10765 5035
rect 10765 5015 10785 5035
rect 10785 5015 10790 5035
rect 10760 5010 10790 5015
rect 10610 4935 10640 4940
rect 10610 4915 10615 4935
rect 10615 4915 10635 4935
rect 10635 4915 10640 4935
rect 10610 4910 10640 4915
rect 10460 4835 10490 4840
rect 10460 4815 10465 4835
rect 10465 4815 10485 4835
rect 10485 4815 10490 4835
rect 10460 4810 10490 4815
rect 10460 4735 10490 4740
rect 10460 4715 10465 4735
rect 10465 4715 10485 4735
rect 10485 4715 10490 4735
rect 10460 4710 10490 4715
rect 10460 4635 10490 4640
rect 10460 4615 10465 4635
rect 10465 4615 10485 4635
rect 10485 4615 10490 4635
rect 10460 4610 10490 4615
rect 10460 4535 10490 4540
rect 10460 4515 10465 4535
rect 10465 4515 10485 4535
rect 10485 4515 10490 4535
rect 10460 4510 10490 4515
rect 10460 4435 10490 4440
rect 10460 4415 10465 4435
rect 10465 4415 10485 4435
rect 10485 4415 10490 4435
rect 10460 4410 10490 4415
rect 10160 4285 10190 4290
rect 10160 4265 10165 4285
rect 10165 4265 10185 4285
rect 10185 4265 10190 4285
rect 10160 4260 10190 4265
rect 9860 4135 9890 4140
rect 9860 4115 9865 4135
rect 9865 4115 9885 4135
rect 9885 4115 9890 4135
rect 9860 4110 9890 4115
rect 9860 4035 9890 4040
rect 9860 4015 9865 4035
rect 9865 4015 9885 4035
rect 9885 4015 9890 4035
rect 9860 4010 9890 4015
rect 9860 3935 9890 3940
rect 9860 3915 9865 3935
rect 9865 3915 9885 3935
rect 9885 3915 9890 3935
rect 9860 3910 9890 3915
rect 9860 3835 9890 3840
rect 9860 3815 9865 3835
rect 9865 3815 9885 3835
rect 9885 3815 9890 3835
rect 9860 3810 9890 3815
rect 9860 3735 9890 3740
rect 9860 3715 9865 3735
rect 9865 3715 9885 3735
rect 9885 3715 9890 3735
rect 9860 3710 9890 3715
rect 9710 3635 9740 3640
rect 9710 3615 9715 3635
rect 9715 3615 9735 3635
rect 9735 3615 9740 3635
rect 9710 3610 9740 3615
rect 9560 3535 9590 3540
rect 9560 3515 9565 3535
rect 9565 3515 9585 3535
rect 9585 3515 9590 3535
rect 9560 3510 9590 3515
rect 9560 3435 9590 3440
rect 9560 3415 9565 3435
rect 9565 3415 9585 3435
rect 9585 3415 9590 3435
rect 9560 3410 9590 3415
rect 9560 3335 9590 3340
rect 9560 3315 9565 3335
rect 9565 3315 9585 3335
rect 9585 3315 9590 3335
rect 9560 3310 9590 3315
rect 9560 3235 9590 3240
rect 9560 3215 9565 3235
rect 9565 3215 9585 3235
rect 9585 3215 9590 3235
rect 9560 3210 9590 3215
rect 9560 3135 9590 3140
rect 9560 3115 9565 3135
rect 9565 3115 9585 3135
rect 9585 3115 9590 3135
rect 9560 3110 9590 3115
rect 9260 2985 9290 2990
rect 9260 2965 9265 2985
rect 9265 2965 9285 2985
rect 9285 2965 9290 2985
rect 9260 2960 9290 2965
rect 10910 4935 10940 4940
rect 10910 4915 10915 4935
rect 10915 4915 10935 4935
rect 10935 4915 10940 4935
rect 10910 4910 10940 4915
rect 11210 4935 11240 4940
rect 11210 4915 11215 4935
rect 11215 4915 11235 4935
rect 11235 4915 11240 4935
rect 11210 4910 11240 4915
rect 13160 5585 13190 5590
rect 13160 5565 13165 5585
rect 13165 5565 13185 5585
rect 13185 5565 13190 5585
rect 13160 5560 13190 5565
rect 11960 5435 11990 5440
rect 11960 5415 11965 5435
rect 11965 5415 11985 5435
rect 11985 5415 11990 5435
rect 11960 5410 11990 5415
rect 11960 5335 11990 5340
rect 11960 5315 11965 5335
rect 11965 5315 11985 5335
rect 11985 5315 11990 5335
rect 11960 5310 11990 5315
rect 11960 5235 11990 5240
rect 11960 5215 11965 5235
rect 11965 5215 11985 5235
rect 11985 5215 11990 5235
rect 11960 5210 11990 5215
rect 11960 5135 11990 5140
rect 11960 5115 11965 5135
rect 11965 5115 11985 5135
rect 11985 5115 11990 5135
rect 11960 5110 11990 5115
rect 11960 5035 11990 5040
rect 11960 5015 11965 5035
rect 11965 5015 11985 5035
rect 11985 5015 11990 5035
rect 11960 5010 11990 5015
rect 11360 4910 11390 4940
rect 10760 4835 10790 4840
rect 10760 4815 10765 4835
rect 10765 4815 10785 4835
rect 10785 4815 10790 4835
rect 10760 4810 10790 4815
rect 10760 4735 10790 4740
rect 10760 4715 10765 4735
rect 10765 4715 10785 4735
rect 10785 4715 10790 4735
rect 10760 4710 10790 4715
rect 10760 4635 10790 4640
rect 10760 4615 10765 4635
rect 10765 4615 10785 4635
rect 10785 4615 10790 4635
rect 10760 4610 10790 4615
rect 10760 4535 10790 4540
rect 10760 4515 10765 4535
rect 10765 4515 10785 4535
rect 10785 4515 10790 4535
rect 10760 4510 10790 4515
rect 10760 4435 10790 4440
rect 10760 4415 10765 4435
rect 10765 4415 10785 4435
rect 10785 4415 10790 4435
rect 10760 4410 10790 4415
rect 10460 4285 10490 4290
rect 10460 4265 10465 4285
rect 10465 4265 10485 4285
rect 10485 4265 10490 4285
rect 10460 4260 10490 4265
rect 10160 4135 10190 4140
rect 10160 4115 10165 4135
rect 10165 4115 10185 4135
rect 10185 4115 10190 4135
rect 10160 4110 10190 4115
rect 10160 4035 10190 4040
rect 10160 4015 10165 4035
rect 10165 4015 10185 4035
rect 10185 4015 10190 4035
rect 10160 4010 10190 4015
rect 10160 3935 10190 3940
rect 10160 3915 10165 3935
rect 10165 3915 10185 3935
rect 10185 3915 10190 3935
rect 10160 3910 10190 3915
rect 10160 3835 10190 3840
rect 10160 3815 10165 3835
rect 10165 3815 10185 3835
rect 10185 3815 10190 3835
rect 10160 3810 10190 3815
rect 10160 3735 10190 3740
rect 10160 3715 10165 3735
rect 10165 3715 10185 3735
rect 10185 3715 10190 3735
rect 10160 3710 10190 3715
rect 10010 3635 10040 3640
rect 10010 3615 10015 3635
rect 10015 3615 10035 3635
rect 10035 3615 10040 3635
rect 10010 3610 10040 3615
rect 9860 3535 9890 3540
rect 9860 3515 9865 3535
rect 9865 3515 9885 3535
rect 9885 3515 9890 3535
rect 9860 3510 9890 3515
rect 9860 3435 9890 3440
rect 9860 3415 9865 3435
rect 9865 3415 9885 3435
rect 9885 3415 9890 3435
rect 9860 3410 9890 3415
rect 9860 3335 9890 3340
rect 9860 3315 9865 3335
rect 9865 3315 9885 3335
rect 9885 3315 9890 3335
rect 9860 3310 9890 3315
rect 9860 3235 9890 3240
rect 9860 3215 9865 3235
rect 9865 3215 9885 3235
rect 9885 3215 9890 3235
rect 9860 3210 9890 3215
rect 9860 3135 9890 3140
rect 9860 3115 9865 3135
rect 9865 3115 9885 3135
rect 9885 3115 9890 3135
rect 9860 3110 9890 3115
rect 9560 2985 9590 2990
rect 9560 2965 9565 2985
rect 9565 2965 9585 2985
rect 9585 2965 9590 2985
rect 9560 2960 9590 2965
rect 10760 4285 10790 4290
rect 10760 4265 10765 4285
rect 10765 4265 10785 4285
rect 10785 4265 10790 4285
rect 10760 4260 10790 4265
rect 10460 4135 10490 4140
rect 10460 4115 10465 4135
rect 10465 4115 10485 4135
rect 10485 4115 10490 4135
rect 10460 4110 10490 4115
rect 10460 4035 10490 4040
rect 10460 4015 10465 4035
rect 10465 4015 10485 4035
rect 10485 4015 10490 4035
rect 10460 4010 10490 4015
rect 10460 3935 10490 3940
rect 10460 3915 10465 3935
rect 10465 3915 10485 3935
rect 10485 3915 10490 3935
rect 10460 3910 10490 3915
rect 10460 3835 10490 3840
rect 10460 3815 10465 3835
rect 10465 3815 10485 3835
rect 10485 3815 10490 3835
rect 10460 3810 10490 3815
rect 10460 3735 10490 3740
rect 10460 3715 10465 3735
rect 10465 3715 10485 3735
rect 10485 3715 10490 3735
rect 10460 3710 10490 3715
rect 10310 3635 10340 3640
rect 10310 3615 10315 3635
rect 10315 3615 10335 3635
rect 10335 3615 10340 3635
rect 10310 3610 10340 3615
rect 10160 3535 10190 3540
rect 10160 3515 10165 3535
rect 10165 3515 10185 3535
rect 10185 3515 10190 3535
rect 10160 3510 10190 3515
rect 10160 3435 10190 3440
rect 10160 3415 10165 3435
rect 10165 3415 10185 3435
rect 10185 3415 10190 3435
rect 10160 3410 10190 3415
rect 10160 3335 10190 3340
rect 10160 3315 10165 3335
rect 10165 3315 10185 3335
rect 10185 3315 10190 3335
rect 10160 3310 10190 3315
rect 10160 3235 10190 3240
rect 10160 3215 10165 3235
rect 10165 3215 10185 3235
rect 10185 3215 10190 3235
rect 10160 3210 10190 3215
rect 10160 3135 10190 3140
rect 10160 3115 10165 3135
rect 10165 3115 10185 3135
rect 10185 3115 10190 3135
rect 10160 3110 10190 3115
rect 9860 2985 9890 2990
rect 9860 2965 9865 2985
rect 9865 2965 9885 2985
rect 9885 2965 9890 2985
rect 9860 2960 9890 2965
rect 10760 4135 10790 4140
rect 10760 4115 10765 4135
rect 10765 4115 10785 4135
rect 10785 4115 10790 4135
rect 10760 4110 10790 4115
rect 10760 4035 10790 4040
rect 10760 4015 10765 4035
rect 10765 4015 10785 4035
rect 10785 4015 10790 4035
rect 10760 4010 10790 4015
rect 10760 3935 10790 3940
rect 10760 3915 10765 3935
rect 10765 3915 10785 3935
rect 10785 3915 10790 3935
rect 10760 3910 10790 3915
rect 10760 3835 10790 3840
rect 10760 3815 10765 3835
rect 10765 3815 10785 3835
rect 10785 3815 10790 3835
rect 10760 3810 10790 3815
rect 10760 3735 10790 3740
rect 10760 3715 10765 3735
rect 10765 3715 10785 3735
rect 10785 3715 10790 3735
rect 10760 3710 10790 3715
rect 10610 3635 10640 3640
rect 10610 3615 10615 3635
rect 10615 3615 10635 3635
rect 10635 3615 10640 3635
rect 10610 3610 10640 3615
rect 10460 3535 10490 3540
rect 10460 3515 10465 3535
rect 10465 3515 10485 3535
rect 10485 3515 10490 3535
rect 10460 3510 10490 3515
rect 10460 3435 10490 3440
rect 10460 3415 10465 3435
rect 10465 3415 10485 3435
rect 10485 3415 10490 3435
rect 10460 3410 10490 3415
rect 10460 3335 10490 3340
rect 10460 3315 10465 3335
rect 10465 3315 10485 3335
rect 10485 3315 10490 3335
rect 10460 3310 10490 3315
rect 10460 3235 10490 3240
rect 10460 3215 10465 3235
rect 10465 3215 10485 3235
rect 10485 3215 10490 3235
rect 10460 3210 10490 3215
rect 10460 3135 10490 3140
rect 10460 3115 10465 3135
rect 10465 3115 10485 3135
rect 10485 3115 10490 3135
rect 10460 3110 10490 3115
rect 10160 2985 10190 2990
rect 10160 2965 10165 2985
rect 10165 2965 10185 2985
rect 10185 2965 10190 2985
rect 10160 2960 10190 2965
rect 11510 4935 11540 4940
rect 11510 4915 11515 4935
rect 11515 4915 11535 4935
rect 11535 4915 11540 4935
rect 11510 4910 11540 4915
rect 11810 4935 11840 4940
rect 11810 4915 11815 4935
rect 11815 4915 11835 4935
rect 11835 4915 11840 4935
rect 11810 4910 11840 4915
rect 10910 3635 10940 3640
rect 10910 3615 10915 3635
rect 10915 3615 10935 3635
rect 10935 3615 10940 3635
rect 10910 3610 10940 3615
rect 11210 3635 11240 3640
rect 11210 3615 11215 3635
rect 11215 3615 11235 3635
rect 11235 3615 11240 3635
rect 11210 3610 11240 3615
rect 12110 4935 12140 4940
rect 12110 4915 12115 4935
rect 12115 4915 12135 4935
rect 12135 4915 12140 4935
rect 12110 4910 12140 4915
rect 12410 4935 12440 4940
rect 12410 4915 12415 4935
rect 12415 4915 12435 4935
rect 12435 4915 12440 4935
rect 12410 4910 12440 4915
rect 14360 5585 14390 5590
rect 14360 5565 14365 5585
rect 14365 5565 14385 5585
rect 14385 5565 14390 5585
rect 14360 5560 14390 5565
rect 13160 5435 13190 5440
rect 13160 5415 13165 5435
rect 13165 5415 13185 5435
rect 13185 5415 13190 5435
rect 13160 5410 13190 5415
rect 13160 5335 13190 5340
rect 13160 5315 13165 5335
rect 13165 5315 13185 5335
rect 13185 5315 13190 5335
rect 13160 5310 13190 5315
rect 13160 5235 13190 5240
rect 13160 5215 13165 5235
rect 13165 5215 13185 5235
rect 13185 5215 13190 5235
rect 13160 5210 13190 5215
rect 13160 5135 13190 5140
rect 13160 5115 13165 5135
rect 13165 5115 13185 5135
rect 13185 5115 13190 5135
rect 13160 5110 13190 5115
rect 13160 5035 13190 5040
rect 13160 5015 13165 5035
rect 13165 5015 13185 5035
rect 13185 5015 13190 5035
rect 13160 5010 13190 5015
rect 12560 4910 12590 4940
rect 11960 4835 11990 4840
rect 11960 4815 11965 4835
rect 11965 4815 11985 4835
rect 11985 4815 11990 4835
rect 11960 4810 11990 4815
rect 11960 4735 11990 4740
rect 11960 4715 11965 4735
rect 11965 4715 11985 4735
rect 11985 4715 11990 4735
rect 11960 4710 11990 4715
rect 11960 4635 11990 4640
rect 11960 4615 11965 4635
rect 11965 4615 11985 4635
rect 11985 4615 11990 4635
rect 11960 4610 11990 4615
rect 11960 4535 11990 4540
rect 11960 4515 11965 4535
rect 11965 4515 11985 4535
rect 11985 4515 11990 4535
rect 11960 4510 11990 4515
rect 11960 4435 11990 4440
rect 11960 4415 11965 4435
rect 11965 4415 11985 4435
rect 11985 4415 11990 4435
rect 11960 4410 11990 4415
rect 11960 4285 11990 4290
rect 11960 4265 11965 4285
rect 11965 4265 11985 4285
rect 11985 4265 11990 4285
rect 11960 4260 11990 4265
rect 11960 4135 11990 4140
rect 11960 4115 11965 4135
rect 11965 4115 11985 4135
rect 11985 4115 11990 4135
rect 11960 4110 11990 4115
rect 11960 4035 11990 4040
rect 11960 4015 11965 4035
rect 11965 4015 11985 4035
rect 11985 4015 11990 4035
rect 11960 4010 11990 4015
rect 11960 3935 11990 3940
rect 11960 3915 11965 3935
rect 11965 3915 11985 3935
rect 11985 3915 11990 3935
rect 11960 3910 11990 3915
rect 11960 3835 11990 3840
rect 11960 3815 11965 3835
rect 11965 3815 11985 3835
rect 11985 3815 11990 3835
rect 11960 3810 11990 3815
rect 11960 3735 11990 3740
rect 11960 3715 11965 3735
rect 11965 3715 11985 3735
rect 11985 3715 11990 3735
rect 11960 3710 11990 3715
rect 11360 3610 11390 3640
rect 10760 3535 10790 3540
rect 10760 3515 10765 3535
rect 10765 3515 10785 3535
rect 10785 3515 10790 3535
rect 10760 3510 10790 3515
rect 10760 3435 10790 3440
rect 10760 3415 10765 3435
rect 10765 3415 10785 3435
rect 10785 3415 10790 3435
rect 10760 3410 10790 3415
rect 10760 3335 10790 3340
rect 10760 3315 10765 3335
rect 10765 3315 10785 3335
rect 10785 3315 10790 3335
rect 10760 3310 10790 3315
rect 10760 3235 10790 3240
rect 10760 3215 10765 3235
rect 10765 3215 10785 3235
rect 10785 3215 10790 3235
rect 10760 3210 10790 3215
rect 10760 3135 10790 3140
rect 10760 3115 10765 3135
rect 10765 3115 10785 3135
rect 10785 3115 10790 3135
rect 10760 3110 10790 3115
rect 10460 2985 10490 2990
rect 10460 2965 10465 2985
rect 10465 2965 10485 2985
rect 10485 2965 10490 2985
rect 10460 2960 10490 2965
rect 11510 3635 11540 3640
rect 11510 3615 11515 3635
rect 11515 3615 11535 3635
rect 11535 3615 11540 3635
rect 11510 3610 11540 3615
rect 11810 3635 11840 3640
rect 11810 3615 11815 3635
rect 11815 3615 11835 3635
rect 11835 3615 11840 3635
rect 11810 3610 11840 3615
rect 12710 4935 12740 4940
rect 12710 4915 12715 4935
rect 12715 4915 12735 4935
rect 12735 4915 12740 4935
rect 12710 4910 12740 4915
rect 13010 4935 13040 4940
rect 13010 4915 13015 4935
rect 13015 4915 13035 4935
rect 13035 4915 13040 4935
rect 13010 4910 13040 4915
rect 12110 3635 12140 3640
rect 12110 3615 12115 3635
rect 12115 3615 12135 3635
rect 12135 3615 12140 3635
rect 12110 3610 12140 3615
rect 12410 3635 12440 3640
rect 12410 3615 12415 3635
rect 12415 3615 12435 3635
rect 12435 3615 12440 3635
rect 12410 3610 12440 3615
rect 13310 4935 13340 4940
rect 13310 4915 13315 4935
rect 13315 4915 13335 4935
rect 13335 4915 13340 4935
rect 13310 4910 13340 4915
rect 13610 4935 13640 4940
rect 13610 4915 13615 4935
rect 13615 4915 13635 4935
rect 13635 4915 13640 4935
rect 13610 4910 13640 4915
rect 15560 5585 15590 5590
rect 15560 5565 15565 5585
rect 15565 5565 15585 5585
rect 15585 5565 15590 5585
rect 15560 5560 15590 5565
rect 14360 5435 14390 5440
rect 14360 5415 14365 5435
rect 14365 5415 14385 5435
rect 14385 5415 14390 5435
rect 14360 5410 14390 5415
rect 14360 5335 14390 5340
rect 14360 5315 14365 5335
rect 14365 5315 14385 5335
rect 14385 5315 14390 5335
rect 14360 5310 14390 5315
rect 14360 5235 14390 5240
rect 14360 5215 14365 5235
rect 14365 5215 14385 5235
rect 14385 5215 14390 5235
rect 14360 5210 14390 5215
rect 14360 5135 14390 5140
rect 14360 5115 14365 5135
rect 14365 5115 14385 5135
rect 14385 5115 14390 5135
rect 14360 5110 14390 5115
rect 14360 5035 14390 5040
rect 14360 5015 14365 5035
rect 14365 5015 14385 5035
rect 14385 5015 14390 5035
rect 14360 5010 14390 5015
rect 13760 4910 13790 4940
rect 13160 4835 13190 4840
rect 13160 4815 13165 4835
rect 13165 4815 13185 4835
rect 13185 4815 13190 4835
rect 13160 4810 13190 4815
rect 13160 4735 13190 4740
rect 13160 4715 13165 4735
rect 13165 4715 13185 4735
rect 13185 4715 13190 4735
rect 13160 4710 13190 4715
rect 13160 4635 13190 4640
rect 13160 4615 13165 4635
rect 13165 4615 13185 4635
rect 13185 4615 13190 4635
rect 13160 4610 13190 4615
rect 13160 4535 13190 4540
rect 13160 4515 13165 4535
rect 13165 4515 13185 4535
rect 13185 4515 13190 4535
rect 13160 4510 13190 4515
rect 13160 4435 13190 4440
rect 13160 4415 13165 4435
rect 13165 4415 13185 4435
rect 13185 4415 13190 4435
rect 13160 4410 13190 4415
rect 13160 4285 13190 4290
rect 13160 4265 13165 4285
rect 13165 4265 13185 4285
rect 13185 4265 13190 4285
rect 13160 4260 13190 4265
rect 13160 4135 13190 4140
rect 13160 4115 13165 4135
rect 13165 4115 13185 4135
rect 13185 4115 13190 4135
rect 13160 4110 13190 4115
rect 13160 4035 13190 4040
rect 13160 4015 13165 4035
rect 13165 4015 13185 4035
rect 13185 4015 13190 4035
rect 13160 4010 13190 4015
rect 13160 3935 13190 3940
rect 13160 3915 13165 3935
rect 13165 3915 13185 3935
rect 13185 3915 13190 3935
rect 13160 3910 13190 3915
rect 13160 3835 13190 3840
rect 13160 3815 13165 3835
rect 13165 3815 13185 3835
rect 13185 3815 13190 3835
rect 13160 3810 13190 3815
rect 13160 3735 13190 3740
rect 13160 3715 13165 3735
rect 13165 3715 13185 3735
rect 13185 3715 13190 3735
rect 13160 3710 13190 3715
rect 12560 3610 12590 3640
rect 11960 3535 11990 3540
rect 11960 3515 11965 3535
rect 11965 3515 11985 3535
rect 11985 3515 11990 3535
rect 11960 3510 11990 3515
rect 11960 3435 11990 3440
rect 11960 3415 11965 3435
rect 11965 3415 11985 3435
rect 11985 3415 11990 3435
rect 11960 3410 11990 3415
rect 11960 3335 11990 3340
rect 11960 3315 11965 3335
rect 11965 3315 11985 3335
rect 11985 3315 11990 3335
rect 11960 3310 11990 3315
rect 11960 3235 11990 3240
rect 11960 3215 11965 3235
rect 11965 3215 11985 3235
rect 11985 3215 11990 3235
rect 11960 3210 11990 3215
rect 11960 3135 11990 3140
rect 11960 3115 11965 3135
rect 11965 3115 11985 3135
rect 11985 3115 11990 3135
rect 11960 3110 11990 3115
rect 10760 2985 10790 2990
rect 10760 2965 10765 2985
rect 10765 2965 10785 2985
rect 10785 2965 10790 2985
rect 10760 2960 10790 2965
rect 12710 3635 12740 3640
rect 12710 3615 12715 3635
rect 12715 3615 12735 3635
rect 12735 3615 12740 3635
rect 12710 3610 12740 3615
rect 13010 3635 13040 3640
rect 13010 3615 13015 3635
rect 13015 3615 13035 3635
rect 13035 3615 13040 3635
rect 13010 3610 13040 3615
rect 13910 4935 13940 4940
rect 13910 4915 13915 4935
rect 13915 4915 13935 4935
rect 13935 4915 13940 4935
rect 13910 4910 13940 4915
rect 14210 4935 14240 4940
rect 14210 4915 14215 4935
rect 14215 4915 14235 4935
rect 14235 4915 14240 4935
rect 14210 4910 14240 4915
rect 13310 3635 13340 3640
rect 13310 3615 13315 3635
rect 13315 3615 13335 3635
rect 13335 3615 13340 3635
rect 13310 3610 13340 3615
rect 13610 3635 13640 3640
rect 13610 3615 13615 3635
rect 13615 3615 13635 3635
rect 13635 3615 13640 3635
rect 13610 3610 13640 3615
rect 14510 4935 14540 4940
rect 14510 4915 14515 4935
rect 14515 4915 14535 4935
rect 14535 4915 14540 4935
rect 14510 4910 14540 4915
rect 14810 4935 14840 4940
rect 14810 4915 14815 4935
rect 14815 4915 14835 4935
rect 14835 4915 14840 4935
rect 14810 4910 14840 4915
rect 20360 5585 20390 5590
rect 20360 5565 20365 5585
rect 20365 5565 20385 5585
rect 20385 5565 20390 5585
rect 20360 5560 20390 5565
rect 15560 5435 15590 5440
rect 15560 5415 15565 5435
rect 15565 5415 15585 5435
rect 15585 5415 15590 5435
rect 15560 5410 15590 5415
rect 15560 5335 15590 5340
rect 15560 5315 15565 5335
rect 15565 5315 15585 5335
rect 15585 5315 15590 5335
rect 15560 5310 15590 5315
rect 15560 5235 15590 5240
rect 15560 5215 15565 5235
rect 15565 5215 15585 5235
rect 15585 5215 15590 5235
rect 15560 5210 15590 5215
rect 15560 5135 15590 5140
rect 15560 5115 15565 5135
rect 15565 5115 15585 5135
rect 15585 5115 15590 5135
rect 15560 5110 15590 5115
rect 15560 5035 15590 5040
rect 15560 5015 15565 5035
rect 15565 5015 15585 5035
rect 15585 5015 15590 5035
rect 15560 5010 15590 5015
rect 14960 4910 14990 4940
rect 14360 4835 14390 4840
rect 14360 4815 14365 4835
rect 14365 4815 14385 4835
rect 14385 4815 14390 4835
rect 14360 4810 14390 4815
rect 14360 4735 14390 4740
rect 14360 4715 14365 4735
rect 14365 4715 14385 4735
rect 14385 4715 14390 4735
rect 14360 4710 14390 4715
rect 14360 4635 14390 4640
rect 14360 4615 14365 4635
rect 14365 4615 14385 4635
rect 14385 4615 14390 4635
rect 14360 4610 14390 4615
rect 14360 4535 14390 4540
rect 14360 4515 14365 4535
rect 14365 4515 14385 4535
rect 14385 4515 14390 4535
rect 14360 4510 14390 4515
rect 14360 4435 14390 4440
rect 14360 4415 14365 4435
rect 14365 4415 14385 4435
rect 14385 4415 14390 4435
rect 14360 4410 14390 4415
rect 14360 4285 14390 4290
rect 14360 4265 14365 4285
rect 14365 4265 14385 4285
rect 14385 4265 14390 4285
rect 14360 4260 14390 4265
rect 14360 4135 14390 4140
rect 14360 4115 14365 4135
rect 14365 4115 14385 4135
rect 14385 4115 14390 4135
rect 14360 4110 14390 4115
rect 14360 4035 14390 4040
rect 14360 4015 14365 4035
rect 14365 4015 14385 4035
rect 14385 4015 14390 4035
rect 14360 4010 14390 4015
rect 14360 3935 14390 3940
rect 14360 3915 14365 3935
rect 14365 3915 14385 3935
rect 14385 3915 14390 3935
rect 14360 3910 14390 3915
rect 14360 3835 14390 3840
rect 14360 3815 14365 3835
rect 14365 3815 14385 3835
rect 14385 3815 14390 3835
rect 14360 3810 14390 3815
rect 14360 3735 14390 3740
rect 14360 3715 14365 3735
rect 14365 3715 14385 3735
rect 14385 3715 14390 3735
rect 14360 3710 14390 3715
rect 13760 3610 13790 3640
rect 13160 3535 13190 3540
rect 13160 3515 13165 3535
rect 13165 3515 13185 3535
rect 13185 3515 13190 3535
rect 13160 3510 13190 3515
rect 13160 3435 13190 3440
rect 13160 3415 13165 3435
rect 13165 3415 13185 3435
rect 13185 3415 13190 3435
rect 13160 3410 13190 3415
rect 13160 3335 13190 3340
rect 13160 3315 13165 3335
rect 13165 3315 13185 3335
rect 13185 3315 13190 3335
rect 13160 3310 13190 3315
rect 13160 3235 13190 3240
rect 13160 3215 13165 3235
rect 13165 3215 13185 3235
rect 13185 3215 13190 3235
rect 13160 3210 13190 3215
rect 13160 3135 13190 3140
rect 13160 3115 13165 3135
rect 13165 3115 13185 3135
rect 13185 3115 13190 3135
rect 13160 3110 13190 3115
rect 11960 2985 11990 2990
rect 11960 2965 11965 2985
rect 11965 2965 11985 2985
rect 11985 2965 11990 2985
rect 11960 2960 11990 2965
rect 13910 3635 13940 3640
rect 13910 3615 13915 3635
rect 13915 3615 13935 3635
rect 13935 3615 13940 3635
rect 13910 3610 13940 3615
rect 14210 3635 14240 3640
rect 14210 3615 14215 3635
rect 14215 3615 14235 3635
rect 14235 3615 14240 3635
rect 14210 3610 14240 3615
rect 15110 4935 15140 4940
rect 15110 4915 15115 4935
rect 15115 4915 15135 4935
rect 15135 4915 15140 4935
rect 15110 4910 15140 4915
rect 15410 4935 15440 4940
rect 15410 4915 15415 4935
rect 15415 4915 15435 4935
rect 15435 4915 15440 4935
rect 15410 4910 15440 4915
rect 14510 3635 14540 3640
rect 14510 3615 14515 3635
rect 14515 3615 14535 3635
rect 14535 3615 14540 3635
rect 14510 3610 14540 3615
rect 14810 3635 14840 3640
rect 14810 3615 14815 3635
rect 14815 3615 14835 3635
rect 14835 3615 14840 3635
rect 14810 3610 14840 3615
rect 15710 4935 15740 4940
rect 15710 4915 15715 4935
rect 15715 4915 15735 4935
rect 15735 4915 15740 4935
rect 15710 4910 15740 4915
rect 16010 4935 16040 4940
rect 16010 4915 16015 4935
rect 16015 4915 16035 4935
rect 16035 4915 16040 4935
rect 16010 4910 16040 4915
rect 15560 4835 15590 4840
rect 15560 4815 15565 4835
rect 15565 4815 15585 4835
rect 15585 4815 15590 4835
rect 15560 4810 15590 4815
rect 15560 4735 15590 4740
rect 15560 4715 15565 4735
rect 15565 4715 15585 4735
rect 15585 4715 15590 4735
rect 15560 4710 15590 4715
rect 15560 4635 15590 4640
rect 15560 4615 15565 4635
rect 15565 4615 15585 4635
rect 15585 4615 15590 4635
rect 15560 4610 15590 4615
rect 15560 4535 15590 4540
rect 15560 4515 15565 4535
rect 15565 4515 15585 4535
rect 15585 4515 15590 4535
rect 15560 4510 15590 4515
rect 15560 4435 15590 4440
rect 15560 4415 15565 4435
rect 15565 4415 15585 4435
rect 15585 4415 15590 4435
rect 15560 4410 15590 4415
rect 16310 4935 16340 4940
rect 16310 4915 16315 4935
rect 16315 4915 16335 4935
rect 16335 4915 16340 4935
rect 16310 4910 16340 4915
rect 16610 4935 16640 4940
rect 16610 4915 16615 4935
rect 16615 4915 16635 4935
rect 16635 4915 16640 4935
rect 16610 4910 16640 4915
rect 16760 4910 16790 4940
rect 16910 4935 16940 4940
rect 16910 4915 16915 4935
rect 16915 4915 16935 4935
rect 16935 4915 16940 4935
rect 16910 4910 16940 4915
rect 17210 4935 17240 4940
rect 17210 4915 17215 4935
rect 17215 4915 17235 4935
rect 17235 4915 17240 4935
rect 17210 4910 17240 4915
rect 17960 5335 17990 5340
rect 17960 5315 17965 5335
rect 17965 5315 17985 5335
rect 17985 5315 17990 5335
rect 17960 5310 17990 5315
rect 17960 5235 17990 5240
rect 17960 5215 17965 5235
rect 17965 5215 17985 5235
rect 17985 5215 17990 5235
rect 17960 5210 17990 5215
rect 17960 5135 17990 5140
rect 17960 5115 17965 5135
rect 17965 5115 17985 5135
rect 17985 5115 17990 5135
rect 17960 5110 17990 5115
rect 17960 5035 17990 5040
rect 17960 5015 17965 5035
rect 17965 5015 17985 5035
rect 17985 5015 17990 5035
rect 17960 5010 17990 5015
rect 17510 4935 17540 4940
rect 17510 4915 17515 4935
rect 17515 4915 17535 4935
rect 17535 4915 17540 4935
rect 17510 4910 17540 4915
rect 17810 4935 17840 4940
rect 17810 4915 17815 4935
rect 17815 4915 17835 4935
rect 17835 4915 17840 4935
rect 17810 4910 17840 4915
rect 18110 4935 18140 4940
rect 18110 4915 18115 4935
rect 18115 4915 18135 4935
rect 18135 4915 18140 4935
rect 18110 4910 18140 4915
rect 18410 4935 18440 4940
rect 18410 4915 18415 4935
rect 18415 4915 18435 4935
rect 18435 4915 18440 4935
rect 18410 4910 18440 4915
rect 17960 4835 17990 4840
rect 17960 4815 17965 4835
rect 17965 4815 17985 4835
rect 17985 4815 17990 4835
rect 17960 4810 17990 4815
rect 17960 4735 17990 4740
rect 17960 4715 17965 4735
rect 17965 4715 17985 4735
rect 17985 4715 17990 4735
rect 17960 4710 17990 4715
rect 17960 4635 17990 4640
rect 17960 4615 17965 4635
rect 17965 4615 17985 4635
rect 17985 4615 17990 4635
rect 17960 4610 17990 4615
rect 17960 4535 17990 4540
rect 17960 4515 17965 4535
rect 17965 4515 17985 4535
rect 17985 4515 17990 4535
rect 17960 4510 17990 4515
rect 18710 4935 18740 4940
rect 18710 4915 18715 4935
rect 18715 4915 18735 4935
rect 18735 4915 18740 4935
rect 18710 4910 18740 4915
rect 19010 4935 19040 4940
rect 19010 4915 19015 4935
rect 19015 4915 19035 4935
rect 19035 4915 19040 4935
rect 19010 4910 19040 4915
rect 19160 4910 19190 4940
rect 19310 4935 19340 4940
rect 19310 4915 19315 4935
rect 19315 4915 19335 4935
rect 19335 4915 19340 4935
rect 19310 4910 19340 4915
rect 19610 4935 19640 4940
rect 19610 4915 19615 4935
rect 19615 4915 19635 4935
rect 19635 4915 19640 4935
rect 19610 4910 19640 4915
rect 22460 5585 22490 5590
rect 22460 5565 22465 5585
rect 22465 5565 22485 5585
rect 22485 5565 22490 5585
rect 22460 5560 22490 5565
rect 20360 5435 20390 5440
rect 20360 5415 20365 5435
rect 20365 5415 20385 5435
rect 20385 5415 20390 5435
rect 20360 5410 20390 5415
rect 20360 5335 20390 5340
rect 20360 5315 20365 5335
rect 20365 5315 20385 5335
rect 20385 5315 20390 5335
rect 20360 5310 20390 5315
rect 20360 5235 20390 5240
rect 20360 5215 20365 5235
rect 20365 5215 20385 5235
rect 20385 5215 20390 5235
rect 20360 5210 20390 5215
rect 20360 5135 20390 5140
rect 20360 5115 20365 5135
rect 20365 5115 20385 5135
rect 20385 5115 20390 5135
rect 20360 5110 20390 5115
rect 20360 5035 20390 5040
rect 20360 5015 20365 5035
rect 20365 5015 20385 5035
rect 20385 5015 20390 5035
rect 20360 5010 20390 5015
rect 19910 4935 19940 4940
rect 19910 4915 19915 4935
rect 19915 4915 19935 4935
rect 19935 4915 19940 4935
rect 19910 4910 19940 4915
rect 20210 4935 20240 4940
rect 20210 4915 20215 4935
rect 20215 4915 20235 4935
rect 20235 4915 20240 4935
rect 20210 4910 20240 4915
rect 20510 4935 20540 4940
rect 20510 4915 20515 4935
rect 20515 4915 20535 4935
rect 20535 4915 20540 4935
rect 20510 4910 20540 4915
rect 20810 4935 20840 4940
rect 20810 4915 20815 4935
rect 20815 4915 20835 4935
rect 20835 4915 20840 4935
rect 20810 4910 20840 4915
rect 20960 4910 20990 4940
rect 20360 4835 20390 4840
rect 20360 4815 20365 4835
rect 20365 4815 20385 4835
rect 20385 4815 20390 4835
rect 20360 4810 20390 4815
rect 20360 4735 20390 4740
rect 20360 4715 20365 4735
rect 20365 4715 20385 4735
rect 20385 4715 20390 4735
rect 20360 4710 20390 4715
rect 20360 4635 20390 4640
rect 20360 4615 20365 4635
rect 20365 4615 20385 4635
rect 20385 4615 20390 4635
rect 20360 4610 20390 4615
rect 20360 4535 20390 4540
rect 20360 4515 20365 4535
rect 20365 4515 20385 4535
rect 20385 4515 20390 4535
rect 20360 4510 20390 4515
rect 20360 4435 20390 4440
rect 20360 4415 20365 4435
rect 20365 4415 20385 4435
rect 20385 4415 20390 4435
rect 20360 4410 20390 4415
rect 15560 4285 15590 4290
rect 15560 4265 15565 4285
rect 15565 4265 15585 4285
rect 15585 4265 15590 4285
rect 15560 4260 15590 4265
rect 20360 4285 20390 4290
rect 20360 4265 20365 4285
rect 20365 4265 20385 4285
rect 20385 4265 20390 4285
rect 20360 4260 20390 4265
rect 15560 4135 15590 4140
rect 15560 4115 15565 4135
rect 15565 4115 15585 4135
rect 15585 4115 15590 4135
rect 15560 4110 15590 4115
rect 15560 4035 15590 4040
rect 15560 4015 15565 4035
rect 15565 4015 15585 4035
rect 15585 4015 15590 4035
rect 15560 4010 15590 4015
rect 15560 3935 15590 3940
rect 15560 3915 15565 3935
rect 15565 3915 15585 3935
rect 15585 3915 15590 3935
rect 15560 3910 15590 3915
rect 15560 3835 15590 3840
rect 15560 3815 15565 3835
rect 15565 3815 15585 3835
rect 15585 3815 15590 3835
rect 15560 3810 15590 3815
rect 15560 3735 15590 3740
rect 15560 3715 15565 3735
rect 15565 3715 15585 3735
rect 15585 3715 15590 3735
rect 15560 3710 15590 3715
rect 14960 3610 14990 3640
rect 14360 3535 14390 3540
rect 14360 3515 14365 3535
rect 14365 3515 14385 3535
rect 14385 3515 14390 3535
rect 14360 3510 14390 3515
rect 14360 3435 14390 3440
rect 14360 3415 14365 3435
rect 14365 3415 14385 3435
rect 14385 3415 14390 3435
rect 14360 3410 14390 3415
rect 14360 3335 14390 3340
rect 14360 3315 14365 3335
rect 14365 3315 14385 3335
rect 14385 3315 14390 3335
rect 14360 3310 14390 3315
rect 14360 3235 14390 3240
rect 14360 3215 14365 3235
rect 14365 3215 14385 3235
rect 14385 3215 14390 3235
rect 14360 3210 14390 3215
rect 14360 3135 14390 3140
rect 14360 3115 14365 3135
rect 14365 3115 14385 3135
rect 14385 3115 14390 3135
rect 14360 3110 14390 3115
rect 13160 2985 13190 2990
rect 13160 2965 13165 2985
rect 13165 2965 13185 2985
rect 13185 2965 13190 2985
rect 13160 2960 13190 2965
rect 15110 3635 15140 3640
rect 15110 3615 15115 3635
rect 15115 3615 15135 3635
rect 15135 3615 15140 3635
rect 15110 3610 15140 3615
rect 15410 3635 15440 3640
rect 15410 3615 15415 3635
rect 15415 3615 15435 3635
rect 15435 3615 15440 3635
rect 15410 3610 15440 3615
rect 15710 3635 15740 3640
rect 15710 3615 15715 3635
rect 15715 3615 15735 3635
rect 15735 3615 15740 3635
rect 15710 3610 15740 3615
rect 16010 3635 16040 3640
rect 16010 3615 16015 3635
rect 16015 3615 16035 3635
rect 16035 3615 16040 3635
rect 16010 3610 16040 3615
rect 15560 3535 15590 3540
rect 15560 3515 15565 3535
rect 15565 3515 15585 3535
rect 15585 3515 15590 3535
rect 15560 3510 15590 3515
rect 15560 3435 15590 3440
rect 15560 3415 15565 3435
rect 15565 3415 15585 3435
rect 15585 3415 15590 3435
rect 15560 3410 15590 3415
rect 15560 3335 15590 3340
rect 15560 3315 15565 3335
rect 15565 3315 15585 3335
rect 15585 3315 15590 3335
rect 15560 3310 15590 3315
rect 15560 3235 15590 3240
rect 15560 3215 15565 3235
rect 15565 3215 15585 3235
rect 15585 3215 15590 3235
rect 15560 3210 15590 3215
rect 15560 3135 15590 3140
rect 15560 3115 15565 3135
rect 15565 3115 15585 3135
rect 15585 3115 15590 3135
rect 15560 3110 15590 3115
rect 14360 2985 14390 2990
rect 14360 2965 14365 2985
rect 14365 2965 14385 2985
rect 14385 2965 14390 2985
rect 14360 2960 14390 2965
rect 16310 3635 16340 3640
rect 16310 3615 16315 3635
rect 16315 3615 16335 3635
rect 16335 3615 16340 3635
rect 16310 3610 16340 3615
rect 16610 3635 16640 3640
rect 16610 3615 16615 3635
rect 16615 3615 16635 3635
rect 16635 3615 16640 3635
rect 16610 3610 16640 3615
rect 16760 3610 16790 3640
rect 16910 3635 16940 3640
rect 16910 3615 16915 3635
rect 16915 3615 16935 3635
rect 16935 3615 16940 3635
rect 16910 3610 16940 3615
rect 17210 3635 17240 3640
rect 17210 3615 17215 3635
rect 17215 3615 17235 3635
rect 17235 3615 17240 3635
rect 17210 3610 17240 3615
rect 17960 4035 17990 4040
rect 17960 4015 17965 4035
rect 17965 4015 17985 4035
rect 17985 4015 17990 4035
rect 17960 4010 17990 4015
rect 17960 3935 17990 3940
rect 17960 3915 17965 3935
rect 17965 3915 17985 3935
rect 17985 3915 17990 3935
rect 17960 3910 17990 3915
rect 17960 3835 17990 3840
rect 17960 3815 17965 3835
rect 17965 3815 17985 3835
rect 17985 3815 17990 3835
rect 17960 3810 17990 3815
rect 17960 3735 17990 3740
rect 17960 3715 17965 3735
rect 17965 3715 17985 3735
rect 17985 3715 17990 3735
rect 17960 3710 17990 3715
rect 17510 3635 17540 3640
rect 17510 3615 17515 3635
rect 17515 3615 17535 3635
rect 17535 3615 17540 3635
rect 17510 3610 17540 3615
rect 17810 3635 17840 3640
rect 17810 3615 17815 3635
rect 17815 3615 17835 3635
rect 17835 3615 17840 3635
rect 17810 3610 17840 3615
rect 18110 3635 18140 3640
rect 18110 3615 18115 3635
rect 18115 3615 18135 3635
rect 18135 3615 18140 3635
rect 18110 3610 18140 3615
rect 18410 3635 18440 3640
rect 18410 3615 18415 3635
rect 18415 3615 18435 3635
rect 18435 3615 18440 3635
rect 18410 3610 18440 3615
rect 17960 3535 17990 3540
rect 17960 3515 17965 3535
rect 17965 3515 17985 3535
rect 17985 3515 17990 3535
rect 17960 3510 17990 3515
rect 17960 3435 17990 3440
rect 17960 3415 17965 3435
rect 17965 3415 17985 3435
rect 17985 3415 17990 3435
rect 17960 3410 17990 3415
rect 17960 3335 17990 3340
rect 17960 3315 17965 3335
rect 17965 3315 17985 3335
rect 17985 3315 17990 3335
rect 17960 3310 17990 3315
rect 17960 3235 17990 3240
rect 17960 3215 17965 3235
rect 17965 3215 17985 3235
rect 17985 3215 17990 3235
rect 17960 3210 17990 3215
rect 18710 3635 18740 3640
rect 18710 3615 18715 3635
rect 18715 3615 18735 3635
rect 18735 3615 18740 3635
rect 18710 3610 18740 3615
rect 19010 3635 19040 3640
rect 19010 3615 19015 3635
rect 19015 3615 19035 3635
rect 19035 3615 19040 3635
rect 19010 3610 19040 3615
rect 19160 3610 19190 3640
rect 19310 3635 19340 3640
rect 19310 3615 19315 3635
rect 19315 3615 19335 3635
rect 19335 3615 19340 3635
rect 19310 3610 19340 3615
rect 19610 3635 19640 3640
rect 19610 3615 19615 3635
rect 19615 3615 19635 3635
rect 19635 3615 19640 3635
rect 19610 3610 19640 3615
rect 20360 4135 20390 4140
rect 20360 4115 20365 4135
rect 20365 4115 20385 4135
rect 20385 4115 20390 4135
rect 20360 4110 20390 4115
rect 20360 4035 20390 4040
rect 20360 4015 20365 4035
rect 20365 4015 20385 4035
rect 20385 4015 20390 4035
rect 20360 4010 20390 4015
rect 20360 3935 20390 3940
rect 20360 3915 20365 3935
rect 20365 3915 20385 3935
rect 20385 3915 20390 3935
rect 20360 3910 20390 3915
rect 20360 3835 20390 3840
rect 20360 3815 20365 3835
rect 20365 3815 20385 3835
rect 20385 3815 20390 3835
rect 20360 3810 20390 3815
rect 20360 3735 20390 3740
rect 20360 3715 20365 3735
rect 20365 3715 20385 3735
rect 20385 3715 20390 3735
rect 20360 3710 20390 3715
rect 19910 3635 19940 3640
rect 19910 3615 19915 3635
rect 19915 3615 19935 3635
rect 19935 3615 19940 3635
rect 19910 3610 19940 3615
rect 20210 3635 20240 3640
rect 20210 3615 20215 3635
rect 20215 3615 20235 3635
rect 20235 3615 20240 3635
rect 20210 3610 20240 3615
rect 21110 4935 21140 4940
rect 21110 4915 21115 4935
rect 21115 4915 21135 4935
rect 21135 4915 21140 4935
rect 21110 4910 21140 4915
rect 21410 4910 21440 4940
rect 20510 3635 20540 3640
rect 20510 3615 20515 3635
rect 20515 3615 20535 3635
rect 20535 3615 20540 3635
rect 20510 3610 20540 3615
rect 20810 3635 20840 3640
rect 20810 3615 20815 3635
rect 20815 3615 20835 3635
rect 20835 3615 20840 3635
rect 20810 3610 20840 3615
rect 21710 4935 21740 4940
rect 21710 4915 21715 4935
rect 21715 4915 21735 4935
rect 21735 4915 21740 4935
rect 21710 4910 21740 4915
rect 24560 5585 24590 5590
rect 24560 5565 24565 5585
rect 24565 5565 24585 5585
rect 24585 5565 24590 5585
rect 24560 5560 24590 5565
rect 22460 5435 22490 5440
rect 22460 5415 22465 5435
rect 22465 5415 22485 5435
rect 22485 5415 22490 5435
rect 22460 5410 22490 5415
rect 22460 5335 22490 5340
rect 22460 5315 22465 5335
rect 22465 5315 22485 5335
rect 22485 5315 22490 5335
rect 22460 5310 22490 5315
rect 22460 5235 22490 5240
rect 22460 5215 22465 5235
rect 22465 5215 22485 5235
rect 22485 5215 22490 5235
rect 22460 5210 22490 5215
rect 22460 5135 22490 5140
rect 22460 5115 22465 5135
rect 22465 5115 22485 5135
rect 22485 5115 22490 5135
rect 22460 5110 22490 5115
rect 22460 5035 22490 5040
rect 22460 5015 22465 5035
rect 22465 5015 22485 5035
rect 22485 5015 22490 5035
rect 22460 5010 22490 5015
rect 21860 4910 21890 4940
rect 20960 3610 20990 3640
rect 20360 3535 20390 3540
rect 20360 3515 20365 3535
rect 20365 3515 20385 3535
rect 20385 3515 20390 3535
rect 20360 3510 20390 3515
rect 20360 3435 20390 3440
rect 20360 3415 20365 3435
rect 20365 3415 20385 3435
rect 20385 3415 20390 3435
rect 20360 3410 20390 3415
rect 20360 3335 20390 3340
rect 20360 3315 20365 3335
rect 20365 3315 20385 3335
rect 20385 3315 20390 3335
rect 20360 3310 20390 3315
rect 20360 3235 20390 3240
rect 20360 3215 20365 3235
rect 20365 3215 20385 3235
rect 20385 3215 20390 3235
rect 20360 3210 20390 3215
rect 20360 3135 20390 3140
rect 20360 3115 20365 3135
rect 20365 3115 20385 3135
rect 20385 3115 20390 3135
rect 20360 3110 20390 3115
rect 15560 2985 15590 2990
rect 15560 2965 15565 2985
rect 15565 2965 15585 2985
rect 15585 2965 15590 2985
rect 15560 2960 15590 2965
rect 21110 3635 21140 3640
rect 21110 3615 21115 3635
rect 21115 3615 21135 3635
rect 21135 3615 21140 3635
rect 21110 3610 21140 3615
rect 22010 4935 22040 4940
rect 22010 4915 22015 4935
rect 22015 4915 22035 4935
rect 22035 4915 22040 4935
rect 22010 4910 22040 4915
rect 22310 4935 22340 4940
rect 22310 4915 22315 4935
rect 22315 4915 22335 4935
rect 22335 4915 22340 4935
rect 22310 4910 22340 4915
rect 21410 3610 21440 3640
rect 21710 3635 21740 3640
rect 21710 3615 21715 3635
rect 21715 3615 21735 3635
rect 21735 3615 21740 3635
rect 21710 3610 21740 3615
rect 22610 4935 22640 4940
rect 22610 4915 22615 4935
rect 22615 4915 22635 4935
rect 22635 4915 22640 4935
rect 22610 4910 22640 4915
rect 22910 4935 22940 4940
rect 22910 4915 22915 4935
rect 22915 4915 22935 4935
rect 22935 4915 22940 4935
rect 22910 4910 22940 4915
rect 23060 4910 23090 4940
rect 22460 4835 22490 4840
rect 22460 4815 22465 4835
rect 22465 4815 22485 4835
rect 22485 4815 22490 4835
rect 22460 4810 22490 4815
rect 22460 4735 22490 4740
rect 22460 4715 22465 4735
rect 22465 4715 22485 4735
rect 22485 4715 22490 4735
rect 22460 4710 22490 4715
rect 22460 4635 22490 4640
rect 22460 4615 22465 4635
rect 22465 4615 22485 4635
rect 22485 4615 22490 4635
rect 22460 4610 22490 4615
rect 22460 4535 22490 4540
rect 22460 4515 22465 4535
rect 22465 4515 22485 4535
rect 22485 4515 22490 4535
rect 22460 4510 22490 4515
rect 22460 4435 22490 4440
rect 22460 4415 22465 4435
rect 22465 4415 22485 4435
rect 22485 4415 22490 4435
rect 22460 4410 22490 4415
rect 22460 4285 22490 4290
rect 22460 4265 22465 4285
rect 22465 4265 22485 4285
rect 22485 4265 22490 4285
rect 22460 4260 22490 4265
rect 22460 4135 22490 4140
rect 22460 4115 22465 4135
rect 22465 4115 22485 4135
rect 22485 4115 22490 4135
rect 22460 4110 22490 4115
rect 22460 4035 22490 4040
rect 22460 4015 22465 4035
rect 22465 4015 22485 4035
rect 22485 4015 22490 4035
rect 22460 4010 22490 4015
rect 22460 3935 22490 3940
rect 22460 3915 22465 3935
rect 22465 3915 22485 3935
rect 22485 3915 22490 3935
rect 22460 3910 22490 3915
rect 22460 3835 22490 3840
rect 22460 3815 22465 3835
rect 22465 3815 22485 3835
rect 22485 3815 22490 3835
rect 22460 3810 22490 3815
rect 22460 3735 22490 3740
rect 22460 3715 22465 3735
rect 22465 3715 22485 3735
rect 22485 3715 22490 3735
rect 22460 3710 22490 3715
rect 21860 3610 21890 3640
rect 22010 3635 22040 3640
rect 22010 3615 22015 3635
rect 22015 3615 22035 3635
rect 22035 3615 22040 3635
rect 22010 3610 22040 3615
rect 22310 3635 22340 3640
rect 22310 3615 22315 3635
rect 22315 3615 22335 3635
rect 22335 3615 22340 3635
rect 22310 3610 22340 3615
rect 23210 4935 23240 4940
rect 23210 4915 23215 4935
rect 23215 4915 23235 4935
rect 23235 4915 23240 4935
rect 23210 4910 23240 4915
rect 23360 4935 23390 4940
rect 23360 4915 23365 4935
rect 23365 4915 23385 4935
rect 23385 4915 23390 4935
rect 23360 4910 23390 4915
rect 23510 4910 23540 4940
rect 22610 3635 22640 3640
rect 22610 3615 22615 3635
rect 22615 3615 22635 3635
rect 22635 3615 22640 3635
rect 22610 3610 22640 3615
rect 22910 3635 22940 3640
rect 22910 3615 22915 3635
rect 22915 3615 22935 3635
rect 22935 3615 22940 3635
rect 22910 3610 22940 3615
rect 23660 4935 23690 4940
rect 23660 4915 23665 4935
rect 23665 4915 23685 4935
rect 23685 4915 23690 4935
rect 23660 4910 23690 4915
rect 23810 4935 23840 4940
rect 23810 4915 23815 4935
rect 23815 4915 23835 4935
rect 23835 4915 23840 4935
rect 23810 4910 23840 4915
rect 26660 5585 26690 5590
rect 26660 5565 26665 5585
rect 26665 5565 26685 5585
rect 26685 5565 26690 5585
rect 26660 5560 26690 5565
rect 24560 5435 24590 5440
rect 24560 5415 24565 5435
rect 24565 5415 24585 5435
rect 24585 5415 24590 5435
rect 24560 5410 24590 5415
rect 24560 5335 24590 5340
rect 24560 5315 24565 5335
rect 24565 5315 24585 5335
rect 24585 5315 24590 5335
rect 24560 5310 24590 5315
rect 24560 5235 24590 5240
rect 24560 5215 24565 5235
rect 24565 5215 24585 5235
rect 24585 5215 24590 5235
rect 24560 5210 24590 5215
rect 24560 5135 24590 5140
rect 24560 5115 24565 5135
rect 24565 5115 24585 5135
rect 24585 5115 24590 5135
rect 24560 5110 24590 5115
rect 24560 5035 24590 5040
rect 24560 5015 24565 5035
rect 24565 5015 24585 5035
rect 24585 5015 24590 5035
rect 24560 5010 24590 5015
rect 23960 4910 23990 4940
rect 23060 3610 23090 3640
rect 22460 3535 22490 3540
rect 22460 3515 22465 3535
rect 22465 3515 22485 3535
rect 22485 3515 22490 3535
rect 22460 3510 22490 3515
rect 22460 3435 22490 3440
rect 22460 3415 22465 3435
rect 22465 3415 22485 3435
rect 22485 3415 22490 3435
rect 22460 3410 22490 3415
rect 22460 3335 22490 3340
rect 22460 3315 22465 3335
rect 22465 3315 22485 3335
rect 22485 3315 22490 3335
rect 22460 3310 22490 3315
rect 22460 3235 22490 3240
rect 22460 3215 22465 3235
rect 22465 3215 22485 3235
rect 22485 3215 22490 3235
rect 22460 3210 22490 3215
rect 22460 3135 22490 3140
rect 22460 3115 22465 3135
rect 22465 3115 22485 3135
rect 22485 3115 22490 3135
rect 22460 3110 22490 3115
rect 23210 3635 23240 3640
rect 23210 3615 23215 3635
rect 23215 3615 23235 3635
rect 23235 3615 23240 3635
rect 23210 3610 23240 3615
rect 23360 3635 23390 3640
rect 23360 3615 23365 3635
rect 23365 3615 23385 3635
rect 23385 3615 23390 3635
rect 23360 3610 23390 3615
rect 24110 4935 24140 4940
rect 24110 4915 24115 4935
rect 24115 4915 24135 4935
rect 24135 4915 24140 4935
rect 24110 4910 24140 4915
rect 24410 4935 24440 4940
rect 24410 4915 24415 4935
rect 24415 4915 24435 4935
rect 24435 4915 24440 4935
rect 24410 4910 24440 4915
rect 23510 3610 23540 3640
rect 23660 3635 23690 3640
rect 23660 3615 23665 3635
rect 23665 3615 23685 3635
rect 23685 3615 23690 3635
rect 23660 3610 23690 3615
rect 23810 3635 23840 3640
rect 23810 3615 23815 3635
rect 23815 3615 23835 3635
rect 23835 3615 23840 3635
rect 23810 3610 23840 3615
rect 24710 4935 24740 4940
rect 24710 4915 24715 4935
rect 24715 4915 24735 4935
rect 24735 4915 24740 4935
rect 24710 4910 24740 4915
rect 25010 4935 25040 4940
rect 25010 4915 25015 4935
rect 25015 4915 25035 4935
rect 25035 4915 25040 4935
rect 25010 4910 25040 4915
rect 24560 4835 24590 4840
rect 24560 4815 24565 4835
rect 24565 4815 24585 4835
rect 24585 4815 24590 4835
rect 24560 4810 24590 4815
rect 24560 4735 24590 4740
rect 24560 4715 24565 4735
rect 24565 4715 24585 4735
rect 24585 4715 24590 4735
rect 24560 4710 24590 4715
rect 24560 4635 24590 4640
rect 24560 4615 24565 4635
rect 24565 4615 24585 4635
rect 24585 4615 24590 4635
rect 24560 4610 24590 4615
rect 24560 4535 24590 4540
rect 24560 4515 24565 4535
rect 24565 4515 24585 4535
rect 24585 4515 24590 4535
rect 24560 4510 24590 4515
rect 24560 4435 24590 4440
rect 24560 4415 24565 4435
rect 24565 4415 24585 4435
rect 24585 4415 24590 4435
rect 24560 4410 24590 4415
rect 25460 4935 25490 4940
rect 25460 4915 25465 4935
rect 25465 4915 25485 4935
rect 25485 4915 25490 4935
rect 25460 4910 25490 4915
rect 25610 4910 25640 4940
rect 25760 4935 25790 4940
rect 25760 4915 25765 4935
rect 25765 4915 25785 4935
rect 25785 4915 25790 4935
rect 25760 4910 25790 4915
rect 24560 4285 24590 4290
rect 24560 4265 24565 4285
rect 24565 4265 24585 4285
rect 24585 4265 24590 4285
rect 24560 4260 24590 4265
rect 24560 4135 24590 4140
rect 24560 4115 24565 4135
rect 24565 4115 24585 4135
rect 24585 4115 24590 4135
rect 24560 4110 24590 4115
rect 24560 4035 24590 4040
rect 24560 4015 24565 4035
rect 24565 4015 24585 4035
rect 24585 4015 24590 4035
rect 24560 4010 24590 4015
rect 24560 3935 24590 3940
rect 24560 3915 24565 3935
rect 24565 3915 24585 3935
rect 24585 3915 24590 3935
rect 24560 3910 24590 3915
rect 24560 3835 24590 3840
rect 24560 3815 24565 3835
rect 24565 3815 24585 3835
rect 24585 3815 24590 3835
rect 24560 3810 24590 3815
rect 24560 3735 24590 3740
rect 24560 3715 24565 3735
rect 24565 3715 24585 3735
rect 24585 3715 24590 3735
rect 24560 3710 24590 3715
rect 23960 3610 23990 3640
rect 24110 3635 24140 3640
rect 24110 3615 24115 3635
rect 24115 3615 24135 3635
rect 24135 3615 24140 3635
rect 24110 3610 24140 3615
rect 24410 3635 24440 3640
rect 24410 3615 24415 3635
rect 24415 3615 24435 3635
rect 24435 3615 24440 3635
rect 24410 3610 24440 3615
rect 24710 3635 24740 3640
rect 24710 3615 24715 3635
rect 24715 3615 24735 3635
rect 24735 3615 24740 3635
rect 24710 3610 24740 3615
rect 25010 3635 25040 3640
rect 25010 3615 25015 3635
rect 25015 3615 25035 3635
rect 25035 3615 25040 3635
rect 25010 3610 25040 3615
rect 24560 3535 24590 3540
rect 24560 3515 24565 3535
rect 24565 3515 24585 3535
rect 24585 3515 24590 3535
rect 24560 3510 24590 3515
rect 24560 3435 24590 3440
rect 24560 3415 24565 3435
rect 24565 3415 24585 3435
rect 24585 3415 24590 3435
rect 24560 3410 24590 3415
rect 24560 3335 24590 3340
rect 24560 3315 24565 3335
rect 24565 3315 24585 3335
rect 24585 3315 24590 3335
rect 24560 3310 24590 3315
rect 24560 3235 24590 3240
rect 24560 3215 24565 3235
rect 24565 3215 24585 3235
rect 24585 3215 24590 3235
rect 24560 3210 24590 3215
rect 24560 3135 24590 3140
rect 24560 3115 24565 3135
rect 24565 3115 24585 3135
rect 24585 3115 24590 3135
rect 24560 3110 24590 3115
rect 20360 2985 20390 2990
rect 20360 2965 20365 2985
rect 20365 2965 20385 2985
rect 20385 2965 20390 2985
rect 20360 2960 20390 2965
rect 28160 5585 28190 5590
rect 28160 5565 28165 5585
rect 28165 5565 28185 5585
rect 28185 5565 28190 5585
rect 28160 5560 28190 5565
rect 26660 5435 26690 5440
rect 26660 5415 26665 5435
rect 26665 5415 26685 5435
rect 26685 5415 26690 5435
rect 26660 5410 26690 5415
rect 26660 5335 26690 5340
rect 26660 5315 26665 5335
rect 26665 5315 26685 5335
rect 26685 5315 26690 5335
rect 26660 5310 26690 5315
rect 26660 5235 26690 5240
rect 26660 5215 26665 5235
rect 26665 5215 26685 5235
rect 26685 5215 26690 5235
rect 26660 5210 26690 5215
rect 26660 5135 26690 5140
rect 26660 5115 26665 5135
rect 26665 5115 26685 5135
rect 26685 5115 26690 5135
rect 26660 5110 26690 5115
rect 26660 5035 26690 5040
rect 26660 5015 26665 5035
rect 26665 5015 26685 5035
rect 26685 5015 26690 5035
rect 26660 5010 26690 5015
rect 26210 4935 26240 4940
rect 26210 4915 26215 4935
rect 26215 4915 26235 4935
rect 26235 4915 26240 4935
rect 26210 4910 26240 4915
rect 26510 4935 26540 4940
rect 26510 4915 26515 4935
rect 26515 4915 26535 4935
rect 26535 4915 26540 4935
rect 26510 4910 26540 4915
rect 26810 4935 26840 4940
rect 26810 4915 26815 4935
rect 26815 4915 26835 4935
rect 26835 4915 26840 4935
rect 26810 4910 26840 4915
rect 27110 4935 27140 4940
rect 27110 4915 27115 4935
rect 27115 4915 27135 4935
rect 27135 4915 27140 4935
rect 27110 4910 27140 4915
rect 26660 4835 26690 4840
rect 26660 4815 26665 4835
rect 26665 4815 26685 4835
rect 26685 4815 26690 4835
rect 26660 4810 26690 4815
rect 26660 4735 26690 4740
rect 26660 4715 26665 4735
rect 26665 4715 26685 4735
rect 26685 4715 26690 4735
rect 26660 4710 26690 4715
rect 26660 4635 26690 4640
rect 26660 4615 26665 4635
rect 26665 4615 26685 4635
rect 26685 4615 26690 4635
rect 26660 4610 26690 4615
rect 26660 4535 26690 4540
rect 26660 4515 26665 4535
rect 26665 4515 26685 4535
rect 26685 4515 26690 4535
rect 26660 4510 26690 4515
rect 26660 4435 26690 4440
rect 26660 4415 26665 4435
rect 26665 4415 26685 4435
rect 26685 4415 26690 4435
rect 26660 4410 26690 4415
rect 27560 4935 27590 4940
rect 27560 4915 27565 4935
rect 27565 4915 27585 4935
rect 27585 4915 27590 4935
rect 27560 4910 27590 4915
rect 28160 5435 28190 5440
rect 28160 5415 28165 5435
rect 28165 5415 28185 5435
rect 28185 5415 28190 5435
rect 28160 5410 28190 5415
rect 28160 5335 28190 5340
rect 28160 5315 28165 5335
rect 28165 5315 28185 5335
rect 28185 5315 28190 5335
rect 28160 5310 28190 5315
rect 28160 5235 28190 5240
rect 28160 5215 28165 5235
rect 28165 5215 28185 5235
rect 28185 5215 28190 5235
rect 28160 5210 28190 5215
rect 28160 5135 28190 5140
rect 28160 5115 28165 5135
rect 28165 5115 28185 5135
rect 28185 5115 28190 5135
rect 28160 5110 28190 5115
rect 28160 5035 28190 5040
rect 28160 5015 28165 5035
rect 28165 5015 28185 5035
rect 28185 5015 28190 5035
rect 28160 5010 28190 5015
rect 27710 4910 27740 4940
rect 27860 4935 27890 4940
rect 27860 4915 27865 4935
rect 27865 4915 27885 4935
rect 27885 4915 27890 4935
rect 27860 4910 27890 4915
rect 26660 4285 26690 4290
rect 26660 4265 26665 4285
rect 26665 4265 26685 4285
rect 26685 4265 26690 4285
rect 26660 4260 26690 4265
rect 25460 3635 25490 3640
rect 25460 3615 25465 3635
rect 25465 3615 25485 3635
rect 25485 3615 25490 3635
rect 25460 3610 25490 3615
rect 25610 3610 25640 3640
rect 25760 3635 25790 3640
rect 25760 3615 25765 3635
rect 25765 3615 25785 3635
rect 25785 3615 25790 3635
rect 25760 3610 25790 3615
rect 26660 4135 26690 4140
rect 26660 4115 26665 4135
rect 26665 4115 26685 4135
rect 26685 4115 26690 4135
rect 26660 4110 26690 4115
rect 26660 4035 26690 4040
rect 26660 4015 26665 4035
rect 26665 4015 26685 4035
rect 26685 4015 26690 4035
rect 26660 4010 26690 4015
rect 26660 3935 26690 3940
rect 26660 3915 26665 3935
rect 26665 3915 26685 3935
rect 26685 3915 26690 3935
rect 26660 3910 26690 3915
rect 26660 3835 26690 3840
rect 26660 3815 26665 3835
rect 26665 3815 26685 3835
rect 26685 3815 26690 3835
rect 26660 3810 26690 3815
rect 26660 3735 26690 3740
rect 26660 3715 26665 3735
rect 26665 3715 26685 3735
rect 26685 3715 26690 3735
rect 26660 3710 26690 3715
rect 26210 3635 26240 3640
rect 26210 3615 26215 3635
rect 26215 3615 26235 3635
rect 26235 3615 26240 3635
rect 26210 3610 26240 3615
rect 26510 3635 26540 3640
rect 26510 3615 26515 3635
rect 26515 3615 26535 3635
rect 26535 3615 26540 3635
rect 26510 3610 26540 3615
rect 26810 3635 26840 3640
rect 26810 3615 26815 3635
rect 26815 3615 26835 3635
rect 26835 3615 26840 3635
rect 26810 3610 26840 3615
rect 27110 3635 27140 3640
rect 27110 3615 27115 3635
rect 27115 3615 27135 3635
rect 27135 3615 27140 3635
rect 27110 3610 27140 3615
rect 26660 3535 26690 3540
rect 26660 3515 26665 3535
rect 26665 3515 26685 3535
rect 26685 3515 26690 3535
rect 26660 3510 26690 3515
rect 26660 3435 26690 3440
rect 26660 3415 26665 3435
rect 26665 3415 26685 3435
rect 26685 3415 26690 3435
rect 26660 3410 26690 3415
rect 26660 3335 26690 3340
rect 26660 3315 26665 3335
rect 26665 3315 26685 3335
rect 26685 3315 26690 3335
rect 26660 3310 26690 3315
rect 26660 3235 26690 3240
rect 26660 3215 26665 3235
rect 26665 3215 26685 3235
rect 26685 3215 26690 3235
rect 26660 3210 26690 3215
rect 26660 3135 26690 3140
rect 26660 3115 26665 3135
rect 26665 3115 26685 3135
rect 26685 3115 26690 3135
rect 26660 3110 26690 3115
rect 27560 3635 27590 3640
rect 27560 3615 27565 3635
rect 27565 3615 27585 3635
rect 27585 3615 27590 3635
rect 27560 3610 27590 3615
rect 28760 5585 28790 5590
rect 28760 5565 28765 5585
rect 28765 5565 28785 5585
rect 28785 5565 28790 5585
rect 28760 5560 28790 5565
rect 32060 5585 32090 5590
rect 32060 5565 32065 5585
rect 32065 5565 32085 5585
rect 32085 5565 32090 5585
rect 32060 5560 32090 5565
rect 28760 5435 28790 5440
rect 28760 5415 28765 5435
rect 28765 5415 28785 5435
rect 28785 5415 28790 5435
rect 28760 5410 28790 5415
rect 28760 5335 28790 5340
rect 28760 5315 28765 5335
rect 28765 5315 28785 5335
rect 28785 5315 28790 5335
rect 28760 5310 28790 5315
rect 28760 5235 28790 5240
rect 28760 5215 28765 5235
rect 28765 5215 28785 5235
rect 28785 5215 28790 5235
rect 28760 5210 28790 5215
rect 28760 5135 28790 5140
rect 28760 5115 28765 5135
rect 28765 5115 28785 5135
rect 28785 5115 28790 5135
rect 28760 5110 28790 5115
rect 28760 5035 28790 5040
rect 28760 5015 28765 5035
rect 28765 5015 28785 5035
rect 28785 5015 28790 5035
rect 28760 5010 28790 5015
rect 28310 4935 28340 4940
rect 28310 4915 28315 4935
rect 28315 4915 28335 4935
rect 28335 4915 28340 4935
rect 28310 4910 28340 4915
rect 28610 4935 28640 4940
rect 28610 4915 28615 4935
rect 28615 4915 28635 4935
rect 28635 4915 28640 4935
rect 28610 4910 28640 4915
rect 28760 4910 28790 4940
rect 28160 4835 28190 4840
rect 28160 4815 28165 4835
rect 28165 4815 28185 4835
rect 28185 4815 28190 4835
rect 28160 4810 28190 4815
rect 28160 4735 28190 4740
rect 28160 4715 28165 4735
rect 28165 4715 28185 4735
rect 28185 4715 28190 4735
rect 28160 4710 28190 4715
rect 28160 4635 28190 4640
rect 28160 4615 28165 4635
rect 28165 4615 28185 4635
rect 28185 4615 28190 4635
rect 28160 4610 28190 4615
rect 28160 4535 28190 4540
rect 28160 4515 28165 4535
rect 28165 4515 28185 4535
rect 28185 4515 28190 4535
rect 28160 4510 28190 4515
rect 28160 4435 28190 4440
rect 28160 4415 28165 4435
rect 28165 4415 28185 4435
rect 28185 4415 28190 4435
rect 28160 4410 28190 4415
rect 28160 4285 28190 4290
rect 28160 4265 28165 4285
rect 28165 4265 28185 4285
rect 28185 4265 28190 4285
rect 28160 4260 28190 4265
rect 28160 4135 28190 4140
rect 28160 4115 28165 4135
rect 28165 4115 28185 4135
rect 28185 4115 28190 4135
rect 28160 4110 28190 4115
rect 28160 4035 28190 4040
rect 28160 4015 28165 4035
rect 28165 4015 28185 4035
rect 28185 4015 28190 4035
rect 28160 4010 28190 4015
rect 28160 3935 28190 3940
rect 28160 3915 28165 3935
rect 28165 3915 28185 3935
rect 28185 3915 28190 3935
rect 28160 3910 28190 3915
rect 28160 3835 28190 3840
rect 28160 3815 28165 3835
rect 28165 3815 28185 3835
rect 28185 3815 28190 3835
rect 28160 3810 28190 3815
rect 28160 3735 28190 3740
rect 28160 3715 28165 3735
rect 28165 3715 28185 3735
rect 28185 3715 28190 3735
rect 28160 3710 28190 3715
rect 27710 3610 27740 3640
rect 27860 3635 27890 3640
rect 27860 3615 27865 3635
rect 27865 3615 27885 3635
rect 27885 3615 27890 3635
rect 27860 3610 27890 3615
rect 28910 4935 28940 4940
rect 28910 4915 28915 4935
rect 28915 4915 28935 4935
rect 28935 4915 28940 4935
rect 28910 4910 28940 4915
rect 29210 4935 29240 4940
rect 29210 4915 29215 4935
rect 29215 4915 29235 4935
rect 29235 4915 29240 4935
rect 29210 4910 29240 4915
rect 29360 4910 29390 4940
rect 28760 4835 28790 4840
rect 28760 4815 28765 4835
rect 28765 4815 28785 4835
rect 28785 4815 28790 4835
rect 28760 4810 28790 4815
rect 28760 4735 28790 4740
rect 28760 4715 28765 4735
rect 28765 4715 28785 4735
rect 28785 4715 28790 4735
rect 28760 4710 28790 4715
rect 28760 4635 28790 4640
rect 28760 4615 28765 4635
rect 28765 4615 28785 4635
rect 28785 4615 28790 4635
rect 28760 4610 28790 4615
rect 28760 4535 28790 4540
rect 28760 4515 28765 4535
rect 28765 4515 28785 4535
rect 28785 4515 28790 4535
rect 28760 4510 28790 4515
rect 28760 4435 28790 4440
rect 28760 4415 28765 4435
rect 28765 4415 28785 4435
rect 28785 4415 28790 4435
rect 28760 4410 28790 4415
rect 28760 4285 28790 4290
rect 28760 4265 28765 4285
rect 28765 4265 28785 4285
rect 28785 4265 28790 4285
rect 28760 4260 28790 4265
rect 28760 4135 28790 4140
rect 28760 4115 28765 4135
rect 28765 4115 28785 4135
rect 28785 4115 28790 4135
rect 28760 4110 28790 4115
rect 28760 4035 28790 4040
rect 28760 4015 28765 4035
rect 28765 4015 28785 4035
rect 28785 4015 28790 4035
rect 28760 4010 28790 4015
rect 28760 3935 28790 3940
rect 28760 3915 28765 3935
rect 28765 3915 28785 3935
rect 28785 3915 28790 3935
rect 28760 3910 28790 3915
rect 28760 3835 28790 3840
rect 28760 3815 28765 3835
rect 28765 3815 28785 3835
rect 28785 3815 28790 3835
rect 28760 3810 28790 3815
rect 28760 3735 28790 3740
rect 28760 3715 28765 3735
rect 28765 3715 28785 3735
rect 28785 3715 28790 3735
rect 28760 3710 28790 3715
rect 28310 3635 28340 3640
rect 28310 3615 28315 3635
rect 28315 3615 28335 3635
rect 28335 3615 28340 3635
rect 28310 3610 28340 3615
rect 28610 3635 28640 3640
rect 28610 3615 28615 3635
rect 28615 3615 28635 3635
rect 28635 3615 28640 3635
rect 28610 3610 28640 3615
rect 29660 4935 29690 4940
rect 29660 4915 29665 4935
rect 29665 4915 29685 4935
rect 29685 4915 29690 4935
rect 29660 4910 29690 4915
rect 29960 4935 29990 4940
rect 29960 4915 29965 4935
rect 29965 4915 29985 4935
rect 29985 4915 29990 4935
rect 29960 4910 29990 4915
rect 30260 4935 30290 4940
rect 30260 4915 30265 4935
rect 30265 4915 30285 4935
rect 30285 4915 30290 4935
rect 30260 4910 30290 4915
rect 30560 4935 30590 4940
rect 30560 4915 30565 4935
rect 30565 4915 30585 4935
rect 30585 4915 30590 4935
rect 30560 4910 30590 4915
rect 30860 4935 30890 4940
rect 30860 4915 30865 4935
rect 30865 4915 30885 4935
rect 30885 4915 30890 4935
rect 30860 4910 30890 4915
rect 31160 4935 31190 4940
rect 31160 4915 31165 4935
rect 31165 4915 31185 4935
rect 31185 4915 31190 4935
rect 31160 4910 31190 4915
rect 32060 5435 32090 5440
rect 32060 5415 32065 5435
rect 32065 5415 32085 5435
rect 32085 5415 32090 5435
rect 32060 5410 32090 5415
rect 32060 5335 32090 5340
rect 32060 5315 32065 5335
rect 32065 5315 32085 5335
rect 32085 5315 32090 5335
rect 32060 5310 32090 5315
rect 32060 5235 32090 5240
rect 32060 5215 32065 5235
rect 32065 5215 32085 5235
rect 32085 5215 32090 5235
rect 32060 5210 32090 5215
rect 32060 5135 32090 5140
rect 32060 5115 32065 5135
rect 32065 5115 32085 5135
rect 32085 5115 32090 5135
rect 32060 5110 32090 5115
rect 32060 5035 32090 5040
rect 32060 5015 32065 5035
rect 32065 5015 32085 5035
rect 32085 5015 32090 5035
rect 32060 5010 32090 5015
rect 31460 4910 31490 4940
rect 28760 3610 28790 3640
rect 28160 3535 28190 3540
rect 28160 3515 28165 3535
rect 28165 3515 28185 3535
rect 28185 3515 28190 3535
rect 28160 3510 28190 3515
rect 28160 3435 28190 3440
rect 28160 3415 28165 3435
rect 28165 3415 28185 3435
rect 28185 3415 28190 3435
rect 28160 3410 28190 3415
rect 28160 3335 28190 3340
rect 28160 3315 28165 3335
rect 28165 3315 28185 3335
rect 28185 3315 28190 3335
rect 28160 3310 28190 3315
rect 28160 3235 28190 3240
rect 28160 3215 28165 3235
rect 28165 3215 28185 3235
rect 28185 3215 28190 3235
rect 28160 3210 28190 3215
rect 28160 3135 28190 3140
rect 28160 3115 28165 3135
rect 28165 3115 28185 3135
rect 28185 3115 28190 3135
rect 28160 3110 28190 3115
rect 24560 2985 24590 2990
rect 24560 2965 24565 2985
rect 24565 2965 24585 2985
rect 24585 2965 24590 2985
rect 24560 2960 24590 2965
rect 28160 2985 28190 2990
rect 28160 2965 28165 2985
rect 28165 2965 28185 2985
rect 28185 2965 28190 2985
rect 28160 2960 28190 2965
rect 28910 3635 28940 3640
rect 28910 3615 28915 3635
rect 28915 3615 28935 3635
rect 28935 3615 28940 3635
rect 28910 3610 28940 3615
rect 29210 3635 29240 3640
rect 29210 3615 29215 3635
rect 29215 3615 29235 3635
rect 29235 3615 29240 3635
rect 29210 3610 29240 3615
rect 31610 4935 31640 4940
rect 31610 4915 31615 4935
rect 31615 4915 31635 4935
rect 31635 4915 31640 4935
rect 31610 4910 31640 4915
rect 31910 4935 31940 4940
rect 31910 4915 31915 4935
rect 31915 4915 31935 4935
rect 31935 4915 31940 4935
rect 31910 4910 31940 4915
rect 32060 4910 32090 4940
rect 29360 3610 29390 3640
rect 28760 3535 28790 3540
rect 28760 3515 28765 3535
rect 28765 3515 28785 3535
rect 28785 3515 28790 3535
rect 28760 3510 28790 3515
rect 28760 3435 28790 3440
rect 28760 3415 28765 3435
rect 28765 3415 28785 3435
rect 28785 3415 28790 3435
rect 28760 3410 28790 3415
rect 28760 3335 28790 3340
rect 28760 3315 28765 3335
rect 28765 3315 28785 3335
rect 28785 3315 28790 3335
rect 28760 3310 28790 3315
rect 28760 3235 28790 3240
rect 28760 3215 28765 3235
rect 28765 3215 28785 3235
rect 28785 3215 28790 3235
rect 28760 3210 28790 3215
rect 28760 3135 28790 3140
rect 28760 3115 28765 3135
rect 28765 3115 28785 3135
rect 28785 3115 28790 3135
rect 28760 3110 28790 3115
rect 29660 3635 29690 3640
rect 29660 3615 29665 3635
rect 29665 3615 29685 3635
rect 29685 3615 29690 3635
rect 29660 3610 29690 3615
rect 29960 3635 29990 3640
rect 29960 3615 29965 3635
rect 29965 3615 29985 3635
rect 29985 3615 29990 3635
rect 29960 3610 29990 3615
rect 30260 3635 30290 3640
rect 30260 3615 30265 3635
rect 30265 3615 30285 3635
rect 30285 3615 30290 3635
rect 30260 3610 30290 3615
rect 30560 3635 30590 3640
rect 30560 3615 30565 3635
rect 30565 3615 30585 3635
rect 30585 3615 30590 3635
rect 30560 3610 30590 3615
rect 30860 3635 30890 3640
rect 30860 3615 30865 3635
rect 30865 3615 30885 3635
rect 30885 3615 30890 3635
rect 30860 3610 30890 3615
rect 31160 3635 31190 3640
rect 31160 3615 31165 3635
rect 31165 3615 31185 3635
rect 31185 3615 31190 3635
rect 31160 3610 31190 3615
rect 32060 4835 32090 4840
rect 32060 4815 32065 4835
rect 32065 4815 32085 4835
rect 32085 4815 32090 4835
rect 32060 4810 32090 4815
rect 32060 4735 32090 4740
rect 32060 4715 32065 4735
rect 32065 4715 32085 4735
rect 32085 4715 32090 4735
rect 32060 4710 32090 4715
rect 32060 4635 32090 4640
rect 32060 4615 32065 4635
rect 32065 4615 32085 4635
rect 32085 4615 32090 4635
rect 32060 4610 32090 4615
rect 32060 4535 32090 4540
rect 32060 4515 32065 4535
rect 32065 4515 32085 4535
rect 32085 4515 32090 4535
rect 32060 4510 32090 4515
rect 32060 4435 32090 4440
rect 32060 4415 32065 4435
rect 32065 4415 32085 4435
rect 32085 4415 32090 4435
rect 32060 4410 32090 4415
rect 32060 4285 32090 4290
rect 32060 4265 32065 4285
rect 32065 4265 32085 4285
rect 32085 4265 32090 4285
rect 32060 4260 32090 4265
rect 32060 4135 32090 4140
rect 32060 4115 32065 4135
rect 32065 4115 32085 4135
rect 32085 4115 32090 4135
rect 32060 4110 32090 4115
rect 32060 4035 32090 4040
rect 32060 4015 32065 4035
rect 32065 4015 32085 4035
rect 32085 4015 32090 4035
rect 32060 4010 32090 4015
rect 32060 3935 32090 3940
rect 32060 3915 32065 3935
rect 32065 3915 32085 3935
rect 32085 3915 32090 3935
rect 32060 3910 32090 3915
rect 32060 3835 32090 3840
rect 32060 3815 32065 3835
rect 32065 3815 32085 3835
rect 32085 3815 32090 3835
rect 32060 3810 32090 3815
rect 32060 3735 32090 3740
rect 32060 3715 32065 3735
rect 32065 3715 32085 3735
rect 32085 3715 32090 3735
rect 32060 3710 32090 3715
rect 31460 3610 31490 3640
rect 31610 3635 31640 3640
rect 31610 3615 31615 3635
rect 31615 3615 31635 3635
rect 31635 3615 31640 3635
rect 31610 3610 31640 3615
rect 31910 3635 31940 3640
rect 31910 3615 31915 3635
rect 31915 3615 31935 3635
rect 31935 3615 31940 3635
rect 31910 3610 31940 3615
rect 32060 3610 32090 3640
rect 32060 3535 32090 3540
rect 32060 3515 32065 3535
rect 32065 3515 32085 3535
rect 32085 3515 32090 3535
rect 32060 3510 32090 3515
rect 32060 3435 32090 3440
rect 32060 3415 32065 3435
rect 32065 3415 32085 3435
rect 32085 3415 32090 3435
rect 32060 3410 32090 3415
rect 32060 3335 32090 3340
rect 32060 3315 32065 3335
rect 32065 3315 32085 3335
rect 32085 3315 32090 3335
rect 32060 3310 32090 3315
rect 32060 3235 32090 3240
rect 32060 3215 32065 3235
rect 32065 3215 32085 3235
rect 32085 3215 32090 3235
rect 32060 3210 32090 3215
rect 32060 3135 32090 3140
rect 32060 3115 32065 3135
rect 32065 3115 32085 3135
rect 32085 3115 32090 3135
rect 32060 3110 32090 3115
rect 28760 2985 28790 2990
rect 28760 2965 28765 2985
rect 28765 2965 28785 2985
rect 28785 2965 28790 2985
rect 28760 2960 28790 2965
rect 32060 2985 32090 2990
rect 32060 2965 32065 2985
rect 32065 2965 32085 2985
rect 32085 2965 32090 2985
rect 32060 2960 32090 2965
rect -640 1685 -610 1690
rect -640 1665 -635 1685
rect -635 1665 -615 1685
rect -615 1665 -610 1685
rect -640 1660 -610 1665
rect -40 1685 -10 1690
rect -40 1665 -35 1685
rect -35 1665 -15 1685
rect -15 1665 -10 1685
rect -40 1660 -10 1665
rect -640 1535 -610 1540
rect -640 1515 -635 1535
rect -635 1515 -615 1535
rect -615 1515 -610 1535
rect -640 1510 -610 1515
rect -640 1435 -610 1440
rect -640 1415 -635 1435
rect -635 1415 -615 1435
rect -615 1415 -610 1435
rect -640 1410 -610 1415
rect -640 1335 -610 1340
rect -640 1315 -635 1335
rect -635 1315 -615 1335
rect -615 1315 -610 1335
rect -640 1310 -610 1315
rect -640 1235 -610 1240
rect -640 1215 -635 1235
rect -635 1215 -615 1235
rect -615 1215 -610 1235
rect -640 1210 -610 1215
rect -640 1135 -610 1140
rect -640 1115 -635 1135
rect -635 1115 -615 1135
rect -615 1115 -610 1135
rect -640 1110 -610 1115
rect -640 1035 -610 1040
rect -640 1015 -635 1035
rect -635 1015 -615 1035
rect -615 1015 -610 1035
rect -640 1010 -610 1015
rect -640 935 -610 940
rect -640 915 -635 935
rect -635 915 -615 935
rect -615 915 -610 935
rect -640 910 -610 915
rect -490 835 -460 840
rect -490 815 -485 835
rect -485 815 -465 835
rect -465 815 -460 835
rect -490 810 -460 815
rect 8360 1685 8390 1690
rect 8360 1665 8365 1685
rect 8365 1665 8385 1685
rect 8385 1665 8390 1685
rect 8360 1660 8390 1665
rect -40 1535 -10 1540
rect -40 1515 -35 1535
rect -35 1515 -15 1535
rect -15 1515 -10 1535
rect -40 1510 -10 1515
rect -40 1435 -10 1440
rect -40 1415 -35 1435
rect -35 1415 -15 1435
rect -15 1415 -10 1435
rect -40 1410 -10 1415
rect -40 1335 -10 1340
rect -40 1315 -35 1335
rect -35 1315 -15 1335
rect -15 1315 -10 1335
rect -40 1310 -10 1315
rect -40 1235 -10 1240
rect -40 1215 -35 1235
rect -35 1215 -15 1235
rect -15 1215 -10 1235
rect -40 1210 -10 1215
rect -40 1135 -10 1140
rect -40 1115 -35 1135
rect -35 1115 -15 1135
rect -15 1115 -10 1135
rect -40 1110 -10 1115
rect -40 1035 -10 1040
rect -40 1015 -35 1035
rect -35 1015 -15 1035
rect -15 1015 -10 1035
rect -40 1010 -10 1015
rect -40 935 -10 940
rect -40 915 -35 935
rect -35 915 -15 935
rect -15 915 -10 935
rect -40 910 -10 915
rect -340 810 -310 840
rect -640 735 -610 740
rect -640 715 -635 735
rect -635 715 -615 735
rect -615 715 -610 735
rect -640 710 -610 715
rect -640 635 -610 640
rect -640 615 -635 635
rect -635 615 -615 635
rect -615 615 -610 635
rect -640 610 -610 615
rect -640 535 -610 540
rect -640 515 -635 535
rect -635 515 -615 535
rect -615 515 -610 535
rect -640 510 -610 515
rect -640 435 -610 440
rect -640 415 -635 435
rect -635 415 -615 435
rect -615 415 -610 435
rect -640 410 -610 415
rect -640 335 -610 340
rect -640 315 -635 335
rect -635 315 -615 335
rect -615 315 -610 335
rect -640 310 -610 315
rect -640 235 -610 240
rect -640 215 -635 235
rect -635 215 -615 235
rect -615 215 -610 235
rect -640 210 -610 215
rect -640 135 -610 140
rect -640 115 -635 135
rect -635 115 -615 135
rect -615 115 -610 135
rect -640 110 -610 115
rect -190 835 -160 840
rect -190 815 -185 835
rect -185 815 -165 835
rect -165 815 -160 835
rect -190 810 -160 815
rect 10760 1685 10790 1690
rect 10760 1665 10765 1685
rect 10765 1665 10785 1685
rect 10785 1665 10790 1685
rect 10760 1660 10790 1665
rect 8360 1535 8390 1540
rect 8360 1515 8365 1535
rect 8365 1515 8385 1535
rect 8385 1515 8390 1535
rect 8360 1510 8390 1515
rect 8360 1435 8390 1440
rect 8360 1415 8365 1435
rect 8365 1415 8385 1435
rect 8385 1415 8390 1435
rect 8360 1410 8390 1415
rect 8360 1335 8390 1340
rect 8360 1315 8365 1335
rect 8365 1315 8385 1335
rect 8385 1315 8390 1335
rect 8360 1310 8390 1315
rect 8360 1235 8390 1240
rect 8360 1215 8365 1235
rect 8365 1215 8385 1235
rect 8385 1215 8390 1235
rect 8360 1210 8390 1215
rect 8360 1135 8390 1140
rect 8360 1115 8365 1135
rect 8365 1115 8385 1135
rect 8385 1115 8390 1135
rect 8360 1110 8390 1115
rect 8360 1035 8390 1040
rect 8360 1015 8365 1035
rect 8365 1015 8385 1035
rect 8385 1015 8390 1035
rect 8360 1010 8390 1015
rect 8360 935 8390 940
rect 8360 915 8365 935
rect 8365 915 8385 935
rect 8385 915 8390 935
rect 8360 910 8390 915
rect 110 835 140 840
rect 110 815 115 835
rect 115 815 135 835
rect 135 815 140 835
rect 110 810 140 815
rect 410 835 440 840
rect 410 815 415 835
rect 415 815 435 835
rect 435 815 440 835
rect 410 810 440 815
rect 710 835 740 840
rect 710 815 715 835
rect 715 815 735 835
rect 735 815 740 835
rect 710 810 740 815
rect 1010 835 1040 840
rect 1010 815 1015 835
rect 1015 815 1035 835
rect 1035 815 1040 835
rect 1010 810 1040 815
rect 1310 835 1340 840
rect 1310 815 1315 835
rect 1315 815 1335 835
rect 1335 815 1340 835
rect 1310 810 1340 815
rect 1610 835 1640 840
rect 1610 815 1615 835
rect 1615 815 1635 835
rect 1635 815 1640 835
rect 1610 810 1640 815
rect 1910 835 1940 840
rect 1910 815 1915 835
rect 1915 815 1935 835
rect 1935 815 1940 835
rect 1910 810 1940 815
rect 2210 835 2240 840
rect 2210 815 2215 835
rect 2215 815 2235 835
rect 2235 815 2240 835
rect 2210 810 2240 815
rect 2360 810 2390 840
rect 2510 835 2540 840
rect 2510 815 2515 835
rect 2515 815 2535 835
rect 2535 815 2540 835
rect 2510 810 2540 815
rect 2810 835 2840 840
rect 2810 815 2815 835
rect 2815 815 2835 835
rect 2835 815 2840 835
rect 2810 810 2840 815
rect 3110 835 3140 840
rect 3110 815 3115 835
rect 3115 815 3135 835
rect 3135 815 3140 835
rect 3110 810 3140 815
rect 3410 835 3440 840
rect 3410 815 3415 835
rect 3415 815 3435 835
rect 3435 815 3440 835
rect 3410 810 3440 815
rect 3710 835 3740 840
rect 3710 815 3715 835
rect 3715 815 3735 835
rect 3735 815 3740 835
rect 3710 810 3740 815
rect 3860 810 3890 840
rect 4010 835 4040 840
rect 4010 815 4015 835
rect 4015 815 4035 835
rect 4035 815 4040 835
rect 4010 810 4040 815
rect 4310 835 4340 840
rect 4310 815 4315 835
rect 4315 815 4335 835
rect 4335 815 4340 835
rect 4310 810 4340 815
rect 4460 810 4490 840
rect 4610 835 4640 840
rect 4610 815 4615 835
rect 4615 815 4635 835
rect 4635 815 4640 835
rect 4610 810 4640 815
rect 4910 835 4940 840
rect 4910 815 4915 835
rect 4915 815 4935 835
rect 4935 815 4940 835
rect 4910 810 4940 815
rect 5210 835 5240 840
rect 5210 815 5215 835
rect 5215 815 5235 835
rect 5235 815 5240 835
rect 5210 810 5240 815
rect 5510 835 5540 840
rect 5510 815 5515 835
rect 5515 815 5535 835
rect 5535 815 5540 835
rect 5510 810 5540 815
rect 5810 835 5840 840
rect 5810 815 5815 835
rect 5815 815 5835 835
rect 5835 815 5840 835
rect 5810 810 5840 815
rect 5960 810 5990 840
rect 6110 835 6140 840
rect 6110 815 6115 835
rect 6115 815 6135 835
rect 6135 815 6140 835
rect 6110 810 6140 815
rect 6410 835 6440 840
rect 6410 815 6415 835
rect 6415 815 6435 835
rect 6435 815 6440 835
rect 6410 810 6440 815
rect 6710 835 6740 840
rect 6710 815 6715 835
rect 6715 815 6735 835
rect 6735 815 6740 835
rect 6710 810 6740 815
rect 7010 835 7040 840
rect 7010 815 7015 835
rect 7015 815 7035 835
rect 7035 815 7040 835
rect 7010 810 7040 815
rect 7310 835 7340 840
rect 7310 815 7315 835
rect 7315 815 7335 835
rect 7335 815 7340 835
rect 7310 810 7340 815
rect 7610 835 7640 840
rect 7610 815 7615 835
rect 7615 815 7635 835
rect 7635 815 7640 835
rect 7610 810 7640 815
rect 7910 835 7940 840
rect 7910 815 7915 835
rect 7915 815 7935 835
rect 7935 815 7940 835
rect 7910 810 7940 815
rect 8210 835 8240 840
rect 8210 815 8215 835
rect 8215 815 8235 835
rect 8235 815 8240 835
rect 8210 810 8240 815
rect -40 735 -10 740
rect -40 715 -35 735
rect -35 715 -15 735
rect -15 715 -10 735
rect -40 710 -10 715
rect -40 635 -10 640
rect -40 615 -35 635
rect -35 615 -15 635
rect -15 615 -10 635
rect -40 610 -10 615
rect -40 535 -10 540
rect -40 515 -35 535
rect -35 515 -15 535
rect -15 515 -10 535
rect -40 510 -10 515
rect -40 435 -10 440
rect -40 415 -35 435
rect -35 415 -15 435
rect -15 415 -10 435
rect -40 410 -10 415
rect -40 335 -10 340
rect -40 315 -35 335
rect -35 315 -15 335
rect -15 315 -10 335
rect -40 310 -10 315
rect -40 235 -10 240
rect -40 215 -35 235
rect -35 215 -15 235
rect -15 215 -10 235
rect -40 210 -10 215
rect -40 135 -10 140
rect -40 115 -35 135
rect -35 115 -15 135
rect -15 115 -10 135
rect -40 110 -10 115
rect -640 -15 -610 -10
rect -640 -35 -635 -15
rect -635 -35 -615 -15
rect -615 -35 -610 -15
rect -640 -40 -610 -35
rect 8510 835 8540 840
rect 8510 815 8515 835
rect 8515 815 8535 835
rect 8535 815 8540 835
rect 8510 810 8540 815
rect 8810 835 8840 840
rect 8810 815 8815 835
rect 8815 815 8835 835
rect 8835 815 8840 835
rect 8810 810 8840 815
rect 9110 835 9140 840
rect 9110 815 9115 835
rect 9115 815 9135 835
rect 9135 815 9140 835
rect 9110 810 9140 815
rect 9410 835 9440 840
rect 9410 815 9415 835
rect 9415 815 9435 835
rect 9435 815 9440 835
rect 9410 810 9440 815
rect 15560 1685 15590 1690
rect 15560 1665 15565 1685
rect 15565 1665 15585 1685
rect 15585 1665 15590 1685
rect 15560 1660 15590 1665
rect 10760 1535 10790 1540
rect 10760 1515 10765 1535
rect 10765 1515 10785 1535
rect 10785 1515 10790 1535
rect 10760 1510 10790 1515
rect 10760 1435 10790 1440
rect 10760 1415 10765 1435
rect 10765 1415 10785 1435
rect 10785 1415 10790 1435
rect 10760 1410 10790 1415
rect 10760 1335 10790 1340
rect 10760 1315 10765 1335
rect 10765 1315 10785 1335
rect 10785 1315 10790 1335
rect 10760 1310 10790 1315
rect 10760 1235 10790 1240
rect 10760 1215 10765 1235
rect 10765 1215 10785 1235
rect 10785 1215 10790 1235
rect 10760 1210 10790 1215
rect 10760 1135 10790 1140
rect 10760 1115 10765 1135
rect 10765 1115 10785 1135
rect 10785 1115 10790 1135
rect 10760 1110 10790 1115
rect 10760 1035 10790 1040
rect 10760 1015 10765 1035
rect 10765 1015 10785 1035
rect 10785 1015 10790 1035
rect 10760 1010 10790 1015
rect 10760 935 10790 940
rect 10760 915 10765 935
rect 10765 915 10785 935
rect 10785 915 10790 935
rect 10760 910 10790 915
rect 9560 810 9590 840
rect 8360 735 8390 740
rect 8360 715 8365 735
rect 8365 715 8385 735
rect 8385 715 8390 735
rect 8360 710 8390 715
rect 8360 635 8390 640
rect 8360 615 8365 635
rect 8365 615 8385 635
rect 8385 615 8390 635
rect 8360 610 8390 615
rect 8360 535 8390 540
rect 8360 515 8365 535
rect 8365 515 8385 535
rect 8385 515 8390 535
rect 8360 510 8390 515
rect 8360 435 8390 440
rect 8360 415 8365 435
rect 8365 415 8385 435
rect 8385 415 8390 435
rect 8360 410 8390 415
rect 8360 335 8390 340
rect 8360 315 8365 335
rect 8365 315 8385 335
rect 8385 315 8390 335
rect 8360 310 8390 315
rect 8360 235 8390 240
rect 8360 215 8365 235
rect 8365 215 8385 235
rect 8385 215 8390 235
rect 8360 210 8390 215
rect 8360 135 8390 140
rect 8360 115 8365 135
rect 8365 115 8385 135
rect 8385 115 8390 135
rect 8360 110 8390 115
rect -40 -15 -10 -10
rect -40 -35 -35 -15
rect -35 -35 -15 -15
rect -15 -35 -10 -15
rect -40 -40 -10 -35
rect -640 -165 -610 -160
rect -640 -185 -635 -165
rect -635 -185 -615 -165
rect -615 -185 -610 -165
rect -640 -190 -610 -185
rect -640 -265 -610 -260
rect -640 -285 -635 -265
rect -635 -285 -615 -265
rect -615 -285 -610 -265
rect -640 -290 -610 -285
rect -640 -365 -610 -360
rect -640 -385 -635 -365
rect -635 -385 -615 -365
rect -615 -385 -610 -365
rect -640 -390 -610 -385
rect -640 -465 -610 -460
rect -640 -485 -635 -465
rect -635 -485 -615 -465
rect -615 -485 -610 -465
rect -640 -490 -610 -485
rect -640 -565 -610 -560
rect -640 -585 -635 -565
rect -635 -585 -615 -565
rect -615 -585 -610 -565
rect -640 -590 -610 -585
rect -640 -665 -610 -660
rect -640 -685 -635 -665
rect -635 -685 -615 -665
rect -615 -685 -610 -665
rect -640 -690 -610 -685
rect -640 -765 -610 -760
rect -640 -785 -635 -765
rect -635 -785 -615 -765
rect -615 -785 -610 -765
rect -640 -790 -610 -785
rect -490 -865 -460 -860
rect -490 -885 -485 -865
rect -485 -885 -465 -865
rect -465 -885 -460 -865
rect -490 -890 -460 -885
rect 9710 835 9740 840
rect 9710 815 9715 835
rect 9715 815 9735 835
rect 9735 815 9740 835
rect 9710 810 9740 815
rect 10010 835 10040 840
rect 10010 815 10015 835
rect 10015 815 10035 835
rect 10035 815 10040 835
rect 10010 810 10040 815
rect 10310 835 10340 840
rect 10310 815 10315 835
rect 10315 815 10335 835
rect 10335 815 10340 835
rect 10310 810 10340 815
rect 10610 835 10640 840
rect 10610 815 10615 835
rect 10615 815 10635 835
rect 10635 815 10640 835
rect 10610 810 10640 815
rect 10910 835 10940 840
rect 10910 815 10915 835
rect 10915 815 10935 835
rect 10935 815 10940 835
rect 10910 810 10940 815
rect 11210 835 11240 840
rect 11210 815 11215 835
rect 11215 815 11235 835
rect 11235 815 11240 835
rect 11210 810 11240 815
rect 11510 835 11540 840
rect 11510 815 11515 835
rect 11515 815 11535 835
rect 11535 815 11540 835
rect 11510 810 11540 815
rect 11810 835 11840 840
rect 11810 815 11815 835
rect 11815 815 11835 835
rect 11835 815 11840 835
rect 11810 810 11840 815
rect 10760 735 10790 740
rect 10760 715 10765 735
rect 10765 715 10785 735
rect 10785 715 10790 735
rect 10760 710 10790 715
rect 10760 635 10790 640
rect 10760 615 10765 635
rect 10765 615 10785 635
rect 10785 615 10790 635
rect 10760 610 10790 615
rect 10760 535 10790 540
rect 10760 515 10765 535
rect 10765 515 10785 535
rect 10785 515 10790 535
rect 10760 510 10790 515
rect 10760 435 10790 440
rect 10760 415 10765 435
rect 10765 415 10785 435
rect 10785 415 10790 435
rect 10760 410 10790 415
rect 10760 335 10790 340
rect 10760 315 10765 335
rect 10765 315 10785 335
rect 10785 315 10790 335
rect 10760 310 10790 315
rect 10760 235 10790 240
rect 10760 215 10765 235
rect 10765 215 10785 235
rect 10785 215 10790 235
rect 10760 210 10790 215
rect 10760 135 10790 140
rect 10760 115 10765 135
rect 10765 115 10785 135
rect 10785 115 10790 135
rect 10760 110 10790 115
rect 8360 -15 8390 -10
rect 8360 -35 8365 -15
rect 8365 -35 8385 -15
rect 8385 -35 8390 -15
rect 8360 -40 8390 -35
rect -40 -165 -10 -160
rect -40 -185 -35 -165
rect -35 -185 -15 -165
rect -15 -185 -10 -165
rect -40 -190 -10 -185
rect -40 -265 -10 -260
rect -40 -285 -35 -265
rect -35 -285 -15 -265
rect -15 -285 -10 -265
rect -40 -290 -10 -285
rect -40 -365 -10 -360
rect -40 -385 -35 -365
rect -35 -385 -15 -365
rect -15 -385 -10 -365
rect -40 -390 -10 -385
rect -40 -465 -10 -460
rect -40 -485 -35 -465
rect -35 -485 -15 -465
rect -15 -485 -10 -465
rect -40 -490 -10 -485
rect -40 -565 -10 -560
rect -40 -585 -35 -565
rect -35 -585 -15 -565
rect -15 -585 -10 -565
rect -40 -590 -10 -585
rect -40 -665 -10 -660
rect -40 -685 -35 -665
rect -35 -685 -15 -665
rect -15 -685 -10 -665
rect -40 -690 -10 -685
rect -40 -765 -10 -760
rect -40 -785 -35 -765
rect -35 -785 -15 -765
rect -15 -785 -10 -765
rect -40 -790 -10 -785
rect -340 -890 -310 -860
rect -640 -965 -610 -960
rect -640 -985 -635 -965
rect -635 -985 -615 -965
rect -615 -985 -610 -965
rect -640 -990 -610 -985
rect -640 -1065 -610 -1060
rect -640 -1085 -635 -1065
rect -635 -1085 -615 -1065
rect -615 -1085 -610 -1065
rect -640 -1090 -610 -1085
rect -640 -1165 -610 -1160
rect -640 -1185 -635 -1165
rect -635 -1185 -615 -1165
rect -615 -1185 -610 -1165
rect -640 -1190 -610 -1185
rect -640 -1265 -610 -1260
rect -640 -1285 -635 -1265
rect -635 -1285 -615 -1265
rect -615 -1285 -610 -1265
rect -640 -1290 -610 -1285
rect -640 -1365 -610 -1360
rect -640 -1385 -635 -1365
rect -635 -1385 -615 -1365
rect -615 -1385 -610 -1365
rect -640 -1390 -610 -1385
rect -640 -1465 -610 -1460
rect -640 -1485 -635 -1465
rect -635 -1485 -615 -1465
rect -615 -1485 -610 -1465
rect -640 -1490 -610 -1485
rect -640 -1565 -610 -1560
rect -640 -1585 -635 -1565
rect -635 -1585 -615 -1565
rect -615 -1585 -610 -1565
rect -640 -1590 -610 -1585
rect -190 -865 -160 -860
rect -190 -885 -185 -865
rect -185 -885 -165 -865
rect -165 -885 -160 -865
rect -190 -890 -160 -885
rect 10760 -15 10790 -10
rect 10760 -35 10765 -15
rect 10765 -35 10785 -15
rect 10785 -35 10790 -15
rect 10760 -40 10790 -35
rect 8360 -165 8390 -160
rect 8360 -185 8365 -165
rect 8365 -185 8385 -165
rect 8385 -185 8390 -165
rect 8360 -190 8390 -185
rect 8360 -265 8390 -260
rect 8360 -285 8365 -265
rect 8365 -285 8385 -265
rect 8385 -285 8390 -265
rect 8360 -290 8390 -285
rect 8360 -365 8390 -360
rect 8360 -385 8365 -365
rect 8365 -385 8385 -365
rect 8385 -385 8390 -365
rect 8360 -390 8390 -385
rect 8360 -465 8390 -460
rect 8360 -485 8365 -465
rect 8365 -485 8385 -465
rect 8385 -485 8390 -465
rect 8360 -490 8390 -485
rect 8360 -565 8390 -560
rect 8360 -585 8365 -565
rect 8365 -585 8385 -565
rect 8385 -585 8390 -565
rect 8360 -590 8390 -585
rect 8360 -665 8390 -660
rect 8360 -685 8365 -665
rect 8365 -685 8385 -665
rect 8385 -685 8390 -665
rect 8360 -690 8390 -685
rect 8360 -765 8390 -760
rect 8360 -785 8365 -765
rect 8365 -785 8385 -765
rect 8385 -785 8390 -765
rect 8360 -790 8390 -785
rect 110 -865 140 -860
rect 110 -885 115 -865
rect 115 -885 135 -865
rect 135 -885 140 -865
rect 110 -890 140 -885
rect 410 -865 440 -860
rect 410 -885 415 -865
rect 415 -885 435 -865
rect 435 -885 440 -865
rect 410 -890 440 -885
rect 710 -865 740 -860
rect 710 -885 715 -865
rect 715 -885 735 -865
rect 735 -885 740 -865
rect 710 -890 740 -885
rect 1010 -865 1040 -860
rect 1010 -885 1015 -865
rect 1015 -885 1035 -865
rect 1035 -885 1040 -865
rect 1010 -890 1040 -885
rect 1310 -865 1340 -860
rect 1310 -885 1315 -865
rect 1315 -885 1335 -865
rect 1335 -885 1340 -865
rect 1310 -890 1340 -885
rect 1610 -865 1640 -860
rect 1610 -885 1615 -865
rect 1615 -885 1635 -865
rect 1635 -885 1640 -865
rect 1610 -890 1640 -885
rect 1910 -865 1940 -860
rect 1910 -885 1915 -865
rect 1915 -885 1935 -865
rect 1935 -885 1940 -865
rect 1910 -890 1940 -885
rect 2210 -865 2240 -860
rect 2210 -885 2215 -865
rect 2215 -885 2235 -865
rect 2235 -885 2240 -865
rect 2210 -890 2240 -885
rect 2360 -890 2390 -860
rect 2510 -865 2540 -860
rect 2510 -885 2515 -865
rect 2515 -885 2535 -865
rect 2535 -885 2540 -865
rect 2510 -890 2540 -885
rect 2810 -865 2840 -860
rect 2810 -885 2815 -865
rect 2815 -885 2835 -865
rect 2835 -885 2840 -865
rect 2810 -890 2840 -885
rect 3110 -865 3140 -860
rect 3110 -885 3115 -865
rect 3115 -885 3135 -865
rect 3135 -885 3140 -865
rect 3110 -890 3140 -885
rect 3410 -865 3440 -860
rect 3410 -885 3415 -865
rect 3415 -885 3435 -865
rect 3435 -885 3440 -865
rect 3410 -890 3440 -885
rect 3710 -865 3740 -860
rect 3710 -885 3715 -865
rect 3715 -885 3735 -865
rect 3735 -885 3740 -865
rect 3710 -890 3740 -885
rect 3860 -890 3890 -860
rect 4010 -865 4040 -860
rect 4010 -885 4015 -865
rect 4015 -885 4035 -865
rect 4035 -885 4040 -865
rect 4010 -890 4040 -885
rect 4310 -865 4340 -860
rect 4310 -885 4315 -865
rect 4315 -885 4335 -865
rect 4335 -885 4340 -865
rect 4310 -890 4340 -885
rect 4460 -890 4490 -860
rect 4610 -865 4640 -860
rect 4610 -885 4615 -865
rect 4615 -885 4635 -865
rect 4635 -885 4640 -865
rect 4610 -890 4640 -885
rect 4910 -865 4940 -860
rect 4910 -885 4915 -865
rect 4915 -885 4935 -865
rect 4935 -885 4940 -865
rect 4910 -890 4940 -885
rect 5210 -865 5240 -860
rect 5210 -885 5215 -865
rect 5215 -885 5235 -865
rect 5235 -885 5240 -865
rect 5210 -890 5240 -885
rect 5510 -865 5540 -860
rect 5510 -885 5515 -865
rect 5515 -885 5535 -865
rect 5535 -885 5540 -865
rect 5510 -890 5540 -885
rect 5810 -865 5840 -860
rect 5810 -885 5815 -865
rect 5815 -885 5835 -865
rect 5835 -885 5840 -865
rect 5810 -890 5840 -885
rect 5960 -890 5990 -860
rect 6110 -865 6140 -860
rect 6110 -885 6115 -865
rect 6115 -885 6135 -865
rect 6135 -885 6140 -865
rect 6110 -890 6140 -885
rect 6410 -865 6440 -860
rect 6410 -885 6415 -865
rect 6415 -885 6435 -865
rect 6435 -885 6440 -865
rect 6410 -890 6440 -885
rect 6710 -865 6740 -860
rect 6710 -885 6715 -865
rect 6715 -885 6735 -865
rect 6735 -885 6740 -865
rect 6710 -890 6740 -885
rect 7010 -865 7040 -860
rect 7010 -885 7015 -865
rect 7015 -885 7035 -865
rect 7035 -885 7040 -865
rect 7010 -890 7040 -885
rect 7310 -865 7340 -860
rect 7310 -885 7315 -865
rect 7315 -885 7335 -865
rect 7335 -885 7340 -865
rect 7310 -890 7340 -885
rect 7610 -865 7640 -860
rect 7610 -885 7615 -865
rect 7615 -885 7635 -865
rect 7635 -885 7640 -865
rect 7610 -890 7640 -885
rect 7910 -865 7940 -860
rect 7910 -885 7915 -865
rect 7915 -885 7935 -865
rect 7935 -885 7940 -865
rect 7910 -890 7940 -885
rect 8210 -865 8240 -860
rect 8210 -885 8215 -865
rect 8215 -885 8235 -865
rect 8235 -885 8240 -865
rect 8210 -890 8240 -885
rect -40 -965 -10 -960
rect -40 -985 -35 -965
rect -35 -985 -15 -965
rect -15 -985 -10 -965
rect -40 -990 -10 -985
rect -40 -1065 -10 -1060
rect -40 -1085 -35 -1065
rect -35 -1085 -15 -1065
rect -15 -1085 -10 -1065
rect -40 -1090 -10 -1085
rect -40 -1165 -10 -1160
rect -40 -1185 -35 -1165
rect -35 -1185 -15 -1165
rect -15 -1185 -10 -1165
rect -40 -1190 -10 -1185
rect -40 -1265 -10 -1260
rect -40 -1285 -35 -1265
rect -35 -1285 -15 -1265
rect -15 -1285 -10 -1265
rect -40 -1290 -10 -1285
rect -40 -1365 -10 -1360
rect -40 -1385 -35 -1365
rect -35 -1385 -15 -1365
rect -15 -1385 -10 -1365
rect -40 -1390 -10 -1385
rect -40 -1465 -10 -1460
rect -40 -1485 -35 -1465
rect -35 -1485 -15 -1465
rect -15 -1485 -10 -1465
rect -40 -1490 -10 -1485
rect -40 -1565 -10 -1560
rect -40 -1585 -35 -1565
rect -35 -1585 -15 -1565
rect -15 -1585 -10 -1565
rect -40 -1590 -10 -1585
rect -640 -1715 -610 -1710
rect -640 -1735 -635 -1715
rect -635 -1735 -615 -1715
rect -615 -1735 -610 -1715
rect -640 -1740 -610 -1735
rect 8510 -865 8540 -860
rect 8510 -885 8515 -865
rect 8515 -885 8535 -865
rect 8535 -885 8540 -865
rect 8510 -890 8540 -885
rect 8810 -865 8840 -860
rect 8810 -885 8815 -865
rect 8815 -885 8835 -865
rect 8835 -885 8840 -865
rect 8810 -890 8840 -885
rect 9110 -865 9140 -860
rect 9110 -885 9115 -865
rect 9115 -885 9135 -865
rect 9135 -885 9140 -865
rect 9110 -890 9140 -885
rect 9410 -865 9440 -860
rect 9410 -885 9415 -865
rect 9415 -885 9435 -865
rect 9435 -885 9440 -865
rect 9410 -890 9440 -885
rect 10760 -165 10790 -160
rect 10760 -185 10765 -165
rect 10765 -185 10785 -165
rect 10785 -185 10790 -165
rect 10760 -190 10790 -185
rect 10760 -265 10790 -260
rect 10760 -285 10765 -265
rect 10765 -285 10785 -265
rect 10785 -285 10790 -265
rect 10760 -290 10790 -285
rect 10760 -365 10790 -360
rect 10760 -385 10765 -365
rect 10765 -385 10785 -365
rect 10785 -385 10790 -365
rect 10760 -390 10790 -385
rect 10760 -465 10790 -460
rect 10760 -485 10765 -465
rect 10765 -485 10785 -465
rect 10785 -485 10790 -465
rect 10760 -490 10790 -485
rect 10760 -565 10790 -560
rect 10760 -585 10765 -565
rect 10765 -585 10785 -565
rect 10785 -585 10790 -565
rect 10760 -590 10790 -585
rect 10760 -665 10790 -660
rect 10760 -685 10765 -665
rect 10765 -685 10785 -665
rect 10785 -685 10790 -665
rect 10760 -690 10790 -685
rect 10760 -765 10790 -760
rect 10760 -785 10765 -765
rect 10765 -785 10785 -765
rect 10785 -785 10790 -765
rect 10760 -790 10790 -785
rect 9560 -890 9590 -860
rect 8360 -965 8390 -960
rect 8360 -985 8365 -965
rect 8365 -985 8385 -965
rect 8385 -985 8390 -965
rect 8360 -990 8390 -985
rect 8360 -1065 8390 -1060
rect 8360 -1085 8365 -1065
rect 8365 -1085 8385 -1065
rect 8385 -1085 8390 -1065
rect 8360 -1090 8390 -1085
rect 8360 -1165 8390 -1160
rect 8360 -1185 8365 -1165
rect 8365 -1185 8385 -1165
rect 8385 -1185 8390 -1165
rect 8360 -1190 8390 -1185
rect 8360 -1265 8390 -1260
rect 8360 -1285 8365 -1265
rect 8365 -1285 8385 -1265
rect 8385 -1285 8390 -1265
rect 8360 -1290 8390 -1285
rect 8360 -1365 8390 -1360
rect 8360 -1385 8365 -1365
rect 8365 -1385 8385 -1365
rect 8385 -1385 8390 -1365
rect 8360 -1390 8390 -1385
rect 8360 -1465 8390 -1460
rect 8360 -1485 8365 -1465
rect 8365 -1485 8385 -1465
rect 8385 -1485 8390 -1465
rect 8360 -1490 8390 -1485
rect 8360 -1565 8390 -1560
rect 8360 -1585 8365 -1565
rect 8365 -1585 8385 -1565
rect 8385 -1585 8390 -1565
rect 8360 -1590 8390 -1585
rect -40 -1715 -10 -1710
rect -40 -1735 -35 -1715
rect -35 -1735 -15 -1715
rect -15 -1735 -10 -1715
rect -40 -1740 -10 -1735
rect 9710 -865 9740 -860
rect 9710 -885 9715 -865
rect 9715 -885 9735 -865
rect 9735 -885 9740 -865
rect 9710 -890 9740 -885
rect 10010 -865 10040 -860
rect 10010 -885 10015 -865
rect 10015 -885 10035 -865
rect 10035 -885 10040 -865
rect 10010 -890 10040 -885
rect 10310 -865 10340 -860
rect 10310 -885 10315 -865
rect 10315 -885 10335 -865
rect 10335 -885 10340 -865
rect 10310 -890 10340 -885
rect 10610 -865 10640 -860
rect 10610 -885 10615 -865
rect 10615 -885 10635 -865
rect 10635 -885 10640 -865
rect 10610 -890 10640 -885
rect 12110 835 12140 840
rect 12110 815 12115 835
rect 12115 815 12135 835
rect 12135 815 12140 835
rect 12110 810 12140 815
rect 12410 835 12440 840
rect 12410 815 12415 835
rect 12415 815 12435 835
rect 12435 815 12440 835
rect 12410 810 12440 815
rect 12560 810 12590 840
rect 12710 835 12740 840
rect 12710 815 12715 835
rect 12715 815 12735 835
rect 12735 815 12740 835
rect 12710 810 12740 815
rect 13010 835 13040 840
rect 13010 815 13015 835
rect 13015 815 13035 835
rect 13035 815 13040 835
rect 13010 810 13040 815
rect 13160 810 13190 840
rect 13310 835 13340 840
rect 13310 815 13315 835
rect 13315 815 13335 835
rect 13335 815 13340 835
rect 13310 810 13340 815
rect 13610 835 13640 840
rect 13610 815 13615 835
rect 13615 815 13635 835
rect 13635 815 13640 835
rect 13610 810 13640 815
rect 13760 810 13790 840
rect 13910 835 13940 840
rect 13910 815 13915 835
rect 13915 815 13935 835
rect 13935 815 13940 835
rect 13910 810 13940 815
rect 14210 835 14240 840
rect 14210 815 14215 835
rect 14215 815 14235 835
rect 14235 815 14240 835
rect 14210 810 14240 815
rect 17960 1685 17990 1690
rect 17960 1665 17965 1685
rect 17965 1665 17985 1685
rect 17985 1665 17990 1685
rect 17960 1660 17990 1665
rect 15560 1535 15590 1540
rect 15560 1515 15565 1535
rect 15565 1515 15585 1535
rect 15585 1515 15590 1535
rect 15560 1510 15590 1515
rect 15560 1435 15590 1440
rect 15560 1415 15565 1435
rect 15565 1415 15585 1435
rect 15585 1415 15590 1435
rect 15560 1410 15590 1415
rect 15560 1335 15590 1340
rect 15560 1315 15565 1335
rect 15565 1315 15585 1335
rect 15585 1315 15590 1335
rect 15560 1310 15590 1315
rect 15560 1235 15590 1240
rect 15560 1215 15565 1235
rect 15565 1215 15585 1235
rect 15585 1215 15590 1235
rect 15560 1210 15590 1215
rect 15560 1135 15590 1140
rect 15560 1115 15565 1135
rect 15565 1115 15585 1135
rect 15585 1115 15590 1135
rect 15560 1110 15590 1115
rect 15560 1035 15590 1040
rect 15560 1015 15565 1035
rect 15565 1015 15585 1035
rect 15585 1015 15590 1035
rect 15560 1010 15590 1015
rect 15560 935 15590 940
rect 15560 915 15565 935
rect 15565 915 15585 935
rect 15585 915 15590 935
rect 15560 910 15590 915
rect 14510 835 14540 840
rect 14510 815 14515 835
rect 14515 815 14535 835
rect 14535 815 14540 835
rect 14510 810 14540 815
rect 14810 835 14840 840
rect 14810 815 14815 835
rect 14815 815 14835 835
rect 14835 815 14840 835
rect 14810 810 14840 815
rect 15110 835 15140 840
rect 15110 815 15115 835
rect 15115 815 15135 835
rect 15135 815 15140 835
rect 15110 810 15140 815
rect 15410 835 15440 840
rect 15410 815 15415 835
rect 15415 815 15435 835
rect 15435 815 15440 835
rect 15410 810 15440 815
rect 10910 -865 10940 -860
rect 10910 -885 10915 -865
rect 10915 -885 10935 -865
rect 10935 -885 10940 -865
rect 10910 -890 10940 -885
rect 11210 -865 11240 -860
rect 11210 -885 11215 -865
rect 11215 -885 11235 -865
rect 11235 -885 11240 -865
rect 11210 -890 11240 -885
rect 11510 -865 11540 -860
rect 11510 -885 11515 -865
rect 11515 -885 11535 -865
rect 11535 -885 11540 -865
rect 11510 -890 11540 -885
rect 11810 -865 11840 -860
rect 11810 -885 11815 -865
rect 11815 -885 11835 -865
rect 11835 -885 11840 -865
rect 11810 -890 11840 -885
rect 10760 -965 10790 -960
rect 10760 -985 10765 -965
rect 10765 -985 10785 -965
rect 10785 -985 10790 -965
rect 10760 -990 10790 -985
rect 10760 -1065 10790 -1060
rect 10760 -1085 10765 -1065
rect 10765 -1085 10785 -1065
rect 10785 -1085 10790 -1065
rect 10760 -1090 10790 -1085
rect 10760 -1165 10790 -1160
rect 10760 -1185 10765 -1165
rect 10765 -1185 10785 -1165
rect 10785 -1185 10790 -1165
rect 10760 -1190 10790 -1185
rect 10760 -1265 10790 -1260
rect 10760 -1285 10765 -1265
rect 10765 -1285 10785 -1265
rect 10785 -1285 10790 -1265
rect 10760 -1290 10790 -1285
rect 10760 -1365 10790 -1360
rect 10760 -1385 10765 -1365
rect 10765 -1385 10785 -1365
rect 10785 -1385 10790 -1365
rect 10760 -1390 10790 -1385
rect 10760 -1465 10790 -1460
rect 10760 -1485 10765 -1465
rect 10765 -1485 10785 -1465
rect 10785 -1485 10790 -1465
rect 10760 -1490 10790 -1485
rect 10760 -1565 10790 -1560
rect 10760 -1585 10765 -1565
rect 10765 -1585 10785 -1565
rect 10785 -1585 10790 -1565
rect 10760 -1590 10790 -1585
rect 8360 -1715 8390 -1710
rect 8360 -1735 8365 -1715
rect 8365 -1735 8385 -1715
rect 8385 -1735 8390 -1715
rect 8360 -1740 8390 -1735
rect 12110 -865 12140 -860
rect 12110 -885 12115 -865
rect 12115 -885 12135 -865
rect 12135 -885 12140 -865
rect 12110 -890 12140 -885
rect 12410 -865 12440 -860
rect 12410 -885 12415 -865
rect 12415 -885 12435 -865
rect 12435 -885 12440 -865
rect 12410 -890 12440 -885
rect 12560 -890 12590 -860
rect 12710 -865 12740 -860
rect 12710 -885 12715 -865
rect 12715 -885 12735 -865
rect 12735 -885 12740 -865
rect 12710 -890 12740 -885
rect 13010 -865 13040 -860
rect 13010 -885 13015 -865
rect 13015 -885 13035 -865
rect 13035 -885 13040 -865
rect 13010 -890 13040 -885
rect 13160 -890 13190 -860
rect 13310 -865 13340 -860
rect 13310 -885 13315 -865
rect 13315 -885 13335 -865
rect 13335 -885 13340 -865
rect 13310 -890 13340 -885
rect 13610 -865 13640 -860
rect 13610 -885 13615 -865
rect 13615 -885 13635 -865
rect 13635 -885 13640 -865
rect 13610 -890 13640 -885
rect 13760 -890 13790 -860
rect 13910 -865 13940 -860
rect 13910 -885 13915 -865
rect 13915 -885 13935 -865
rect 13935 -885 13940 -865
rect 13910 -890 13940 -885
rect 14210 -865 14240 -860
rect 14210 -885 14215 -865
rect 14215 -885 14235 -865
rect 14235 -885 14240 -865
rect 14210 -890 14240 -885
rect 15710 835 15740 840
rect 15710 815 15715 835
rect 15715 815 15735 835
rect 15735 815 15740 835
rect 15710 810 15740 815
rect 16010 835 16040 840
rect 16010 815 16015 835
rect 16015 815 16035 835
rect 16035 815 16040 835
rect 16010 810 16040 815
rect 16310 835 16340 840
rect 16310 815 16315 835
rect 16315 815 16335 835
rect 16335 815 16340 835
rect 16310 810 16340 815
rect 16610 835 16640 840
rect 16610 815 16615 835
rect 16615 815 16635 835
rect 16635 815 16640 835
rect 16610 810 16640 815
rect 20360 1685 20390 1690
rect 20360 1665 20365 1685
rect 20365 1665 20385 1685
rect 20385 1665 20390 1685
rect 20360 1660 20390 1665
rect 17960 1535 17990 1540
rect 17960 1515 17965 1535
rect 17965 1515 17985 1535
rect 17985 1515 17990 1535
rect 17960 1510 17990 1515
rect 17960 1435 17990 1440
rect 17960 1415 17965 1435
rect 17965 1415 17985 1435
rect 17985 1415 17990 1435
rect 17960 1410 17990 1415
rect 17960 1335 17990 1340
rect 17960 1315 17965 1335
rect 17965 1315 17985 1335
rect 17985 1315 17990 1335
rect 17960 1310 17990 1315
rect 17960 1235 17990 1240
rect 17960 1215 17965 1235
rect 17965 1215 17985 1235
rect 17985 1215 17990 1235
rect 17960 1210 17990 1215
rect 17960 1135 17990 1140
rect 17960 1115 17965 1135
rect 17965 1115 17985 1135
rect 17985 1115 17990 1135
rect 17960 1110 17990 1115
rect 17960 1035 17990 1040
rect 17960 1015 17965 1035
rect 17965 1015 17985 1035
rect 17985 1015 17990 1035
rect 17960 1010 17990 1015
rect 17960 935 17990 940
rect 17960 915 17965 935
rect 17965 915 17985 935
rect 17985 915 17990 935
rect 17960 910 17990 915
rect 16760 810 16790 840
rect 15560 735 15590 740
rect 15560 715 15565 735
rect 15565 715 15585 735
rect 15585 715 15590 735
rect 15560 710 15590 715
rect 15560 635 15590 640
rect 15560 615 15565 635
rect 15565 615 15585 635
rect 15585 615 15590 635
rect 15560 610 15590 615
rect 15560 535 15590 540
rect 15560 515 15565 535
rect 15565 515 15585 535
rect 15585 515 15590 535
rect 15560 510 15590 515
rect 15560 435 15590 440
rect 15560 415 15565 435
rect 15565 415 15585 435
rect 15585 415 15590 435
rect 15560 410 15590 415
rect 15560 335 15590 340
rect 15560 315 15565 335
rect 15565 315 15585 335
rect 15585 315 15590 335
rect 15560 310 15590 315
rect 15560 235 15590 240
rect 15560 215 15565 235
rect 15565 215 15585 235
rect 15585 215 15590 235
rect 15560 210 15590 215
rect 15560 135 15590 140
rect 15560 115 15565 135
rect 15565 115 15585 135
rect 15585 115 15590 135
rect 15560 110 15590 115
rect 16910 835 16940 840
rect 16910 815 16915 835
rect 16915 815 16935 835
rect 16935 815 16940 835
rect 16910 810 16940 815
rect 17210 835 17240 840
rect 17210 815 17215 835
rect 17215 815 17235 835
rect 17235 815 17240 835
rect 17210 810 17240 815
rect 17510 835 17540 840
rect 17510 815 17515 835
rect 17515 815 17535 835
rect 17535 815 17540 835
rect 17510 810 17540 815
rect 17810 835 17840 840
rect 17810 815 17815 835
rect 17815 815 17835 835
rect 17835 815 17840 835
rect 17810 810 17840 815
rect 18110 835 18140 840
rect 18110 815 18115 835
rect 18115 815 18135 835
rect 18135 815 18140 835
rect 18110 810 18140 815
rect 18410 835 18440 840
rect 18410 815 18415 835
rect 18415 815 18435 835
rect 18435 815 18440 835
rect 18410 810 18440 815
rect 18710 835 18740 840
rect 18710 815 18715 835
rect 18715 815 18735 835
rect 18735 815 18740 835
rect 18710 810 18740 815
rect 19010 835 19040 840
rect 19010 815 19015 835
rect 19015 815 19035 835
rect 19035 815 19040 835
rect 19010 810 19040 815
rect 24560 1685 24590 1690
rect 24560 1665 24565 1685
rect 24565 1665 24585 1685
rect 24585 1665 24590 1685
rect 24560 1660 24590 1665
rect 20360 1535 20390 1540
rect 20360 1515 20365 1535
rect 20365 1515 20385 1535
rect 20385 1515 20390 1535
rect 20360 1510 20390 1515
rect 20360 1435 20390 1440
rect 20360 1415 20365 1435
rect 20365 1415 20385 1435
rect 20385 1415 20390 1435
rect 20360 1410 20390 1415
rect 20360 1335 20390 1340
rect 20360 1315 20365 1335
rect 20365 1315 20385 1335
rect 20385 1315 20390 1335
rect 20360 1310 20390 1315
rect 20360 1235 20390 1240
rect 20360 1215 20365 1235
rect 20365 1215 20385 1235
rect 20385 1215 20390 1235
rect 20360 1210 20390 1215
rect 20360 1135 20390 1140
rect 20360 1115 20365 1135
rect 20365 1115 20385 1135
rect 20385 1115 20390 1135
rect 20360 1110 20390 1115
rect 20360 1035 20390 1040
rect 20360 1015 20365 1035
rect 20365 1015 20385 1035
rect 20385 1015 20390 1035
rect 20360 1010 20390 1015
rect 20360 935 20390 940
rect 20360 915 20365 935
rect 20365 915 20385 935
rect 20385 915 20390 935
rect 20360 910 20390 915
rect 19160 810 19190 840
rect 17960 735 17990 740
rect 17960 715 17965 735
rect 17965 715 17985 735
rect 17985 715 17990 735
rect 17960 710 17990 715
rect 17960 635 17990 640
rect 17960 615 17965 635
rect 17965 615 17985 635
rect 17985 615 17990 635
rect 17960 610 17990 615
rect 17960 535 17990 540
rect 17960 515 17965 535
rect 17965 515 17985 535
rect 17985 515 17990 535
rect 17960 510 17990 515
rect 17960 435 17990 440
rect 17960 415 17965 435
rect 17965 415 17985 435
rect 17985 415 17990 435
rect 17960 410 17990 415
rect 17960 335 17990 340
rect 17960 315 17965 335
rect 17965 315 17985 335
rect 17985 315 17990 335
rect 17960 310 17990 315
rect 17960 235 17990 240
rect 17960 215 17965 235
rect 17965 215 17985 235
rect 17985 215 17990 235
rect 17960 210 17990 215
rect 17960 135 17990 140
rect 17960 115 17965 135
rect 17965 115 17985 135
rect 17985 115 17990 135
rect 17960 110 17990 115
rect 15560 -15 15590 -10
rect 15560 -35 15565 -15
rect 15565 -35 15585 -15
rect 15585 -35 15590 -15
rect 15560 -40 15590 -35
rect 19310 835 19340 840
rect 19310 815 19315 835
rect 19315 815 19335 835
rect 19335 815 19340 835
rect 19310 810 19340 815
rect 19610 835 19640 840
rect 19610 815 19615 835
rect 19615 815 19635 835
rect 19635 815 19640 835
rect 19610 810 19640 815
rect 19910 835 19940 840
rect 19910 815 19915 835
rect 19915 815 19935 835
rect 19935 815 19940 835
rect 19910 810 19940 815
rect 20210 835 20240 840
rect 20210 815 20215 835
rect 20215 815 20235 835
rect 20235 815 20240 835
rect 20210 810 20240 815
rect 20510 835 20540 840
rect 20510 815 20515 835
rect 20515 815 20535 835
rect 20535 815 20540 835
rect 20510 810 20540 815
rect 20810 835 20840 840
rect 20810 815 20815 835
rect 20815 815 20835 835
rect 20835 815 20840 835
rect 20810 810 20840 815
rect 21110 835 21140 840
rect 21110 815 21115 835
rect 21115 815 21135 835
rect 21135 815 21140 835
rect 21110 810 21140 815
rect 21410 835 21440 840
rect 21410 815 21415 835
rect 21415 815 21435 835
rect 21435 815 21440 835
rect 21410 810 21440 815
rect 20360 735 20390 740
rect 20360 715 20365 735
rect 20365 715 20385 735
rect 20385 715 20390 735
rect 20360 710 20390 715
rect 20360 635 20390 640
rect 20360 615 20365 635
rect 20365 615 20385 635
rect 20385 615 20390 635
rect 20360 610 20390 615
rect 20360 535 20390 540
rect 20360 515 20365 535
rect 20365 515 20385 535
rect 20385 515 20390 535
rect 20360 510 20390 515
rect 20360 435 20390 440
rect 20360 415 20365 435
rect 20365 415 20385 435
rect 20385 415 20390 435
rect 20360 410 20390 415
rect 20360 335 20390 340
rect 20360 315 20365 335
rect 20365 315 20385 335
rect 20385 315 20390 335
rect 20360 310 20390 315
rect 20360 235 20390 240
rect 20360 215 20365 235
rect 20365 215 20385 235
rect 20385 215 20390 235
rect 20360 210 20390 215
rect 20360 135 20390 140
rect 20360 115 20365 135
rect 20365 115 20385 135
rect 20385 115 20390 135
rect 20360 110 20390 115
rect 17960 -15 17990 -10
rect 17960 -35 17965 -15
rect 17965 -35 17985 -15
rect 17985 -35 17990 -15
rect 17960 -40 17990 -35
rect 15560 -165 15590 -160
rect 15560 -185 15565 -165
rect 15565 -185 15585 -165
rect 15585 -185 15590 -165
rect 15560 -190 15590 -185
rect 15560 -265 15590 -260
rect 15560 -285 15565 -265
rect 15565 -285 15585 -265
rect 15585 -285 15590 -265
rect 15560 -290 15590 -285
rect 15560 -365 15590 -360
rect 15560 -385 15565 -365
rect 15565 -385 15585 -365
rect 15585 -385 15590 -365
rect 15560 -390 15590 -385
rect 15560 -465 15590 -460
rect 15560 -485 15565 -465
rect 15565 -485 15585 -465
rect 15585 -485 15590 -465
rect 15560 -490 15590 -485
rect 15560 -565 15590 -560
rect 15560 -585 15565 -565
rect 15565 -585 15585 -565
rect 15585 -585 15590 -565
rect 15560 -590 15590 -585
rect 15560 -665 15590 -660
rect 15560 -685 15565 -665
rect 15565 -685 15585 -665
rect 15585 -685 15590 -665
rect 15560 -690 15590 -685
rect 15560 -765 15590 -760
rect 15560 -785 15565 -765
rect 15565 -785 15585 -765
rect 15585 -785 15590 -765
rect 15560 -790 15590 -785
rect 14510 -865 14540 -860
rect 14510 -885 14515 -865
rect 14515 -885 14535 -865
rect 14535 -885 14540 -865
rect 14510 -890 14540 -885
rect 14810 -865 14840 -860
rect 14810 -885 14815 -865
rect 14815 -885 14835 -865
rect 14835 -885 14840 -865
rect 14810 -890 14840 -885
rect 15110 -865 15140 -860
rect 15110 -885 15115 -865
rect 15115 -885 15135 -865
rect 15135 -885 15140 -865
rect 15110 -890 15140 -885
rect 15410 -865 15440 -860
rect 15410 -885 15415 -865
rect 15415 -885 15435 -865
rect 15435 -885 15440 -865
rect 15410 -890 15440 -885
rect 15710 -865 15740 -860
rect 15710 -885 15715 -865
rect 15715 -885 15735 -865
rect 15735 -885 15740 -865
rect 15710 -890 15740 -885
rect 16010 -865 16040 -860
rect 16010 -885 16015 -865
rect 16015 -885 16035 -865
rect 16035 -885 16040 -865
rect 16010 -890 16040 -885
rect 16310 -865 16340 -860
rect 16310 -885 16315 -865
rect 16315 -885 16335 -865
rect 16335 -885 16340 -865
rect 16310 -890 16340 -885
rect 16610 -865 16640 -860
rect 16610 -885 16615 -865
rect 16615 -885 16635 -865
rect 16635 -885 16640 -865
rect 16610 -890 16640 -885
rect 20360 -15 20390 -10
rect 20360 -35 20365 -15
rect 20365 -35 20385 -15
rect 20385 -35 20390 -15
rect 20360 -40 20390 -35
rect 17960 -165 17990 -160
rect 17960 -185 17965 -165
rect 17965 -185 17985 -165
rect 17985 -185 17990 -165
rect 17960 -190 17990 -185
rect 17960 -265 17990 -260
rect 17960 -285 17965 -265
rect 17965 -285 17985 -265
rect 17985 -285 17990 -265
rect 17960 -290 17990 -285
rect 17960 -365 17990 -360
rect 17960 -385 17965 -365
rect 17965 -385 17985 -365
rect 17985 -385 17990 -365
rect 17960 -390 17990 -385
rect 17960 -465 17990 -460
rect 17960 -485 17965 -465
rect 17965 -485 17985 -465
rect 17985 -485 17990 -465
rect 17960 -490 17990 -485
rect 17960 -565 17990 -560
rect 17960 -585 17965 -565
rect 17965 -585 17985 -565
rect 17985 -585 17990 -565
rect 17960 -590 17990 -585
rect 17960 -665 17990 -660
rect 17960 -685 17965 -665
rect 17965 -685 17985 -665
rect 17985 -685 17990 -665
rect 17960 -690 17990 -685
rect 17960 -765 17990 -760
rect 17960 -785 17965 -765
rect 17965 -785 17985 -765
rect 17985 -785 17990 -765
rect 17960 -790 17990 -785
rect 16760 -890 16790 -860
rect 15560 -965 15590 -960
rect 15560 -985 15565 -965
rect 15565 -985 15585 -965
rect 15585 -985 15590 -965
rect 15560 -990 15590 -985
rect 15560 -1065 15590 -1060
rect 15560 -1085 15565 -1065
rect 15565 -1085 15585 -1065
rect 15585 -1085 15590 -1065
rect 15560 -1090 15590 -1085
rect 15560 -1165 15590 -1160
rect 15560 -1185 15565 -1165
rect 15565 -1185 15585 -1165
rect 15585 -1185 15590 -1165
rect 15560 -1190 15590 -1185
rect 15560 -1265 15590 -1260
rect 15560 -1285 15565 -1265
rect 15565 -1285 15585 -1265
rect 15585 -1285 15590 -1265
rect 15560 -1290 15590 -1285
rect 15560 -1365 15590 -1360
rect 15560 -1385 15565 -1365
rect 15565 -1385 15585 -1365
rect 15585 -1385 15590 -1365
rect 15560 -1390 15590 -1385
rect 15560 -1465 15590 -1460
rect 15560 -1485 15565 -1465
rect 15565 -1485 15585 -1465
rect 15585 -1485 15590 -1465
rect 15560 -1490 15590 -1485
rect 15560 -1565 15590 -1560
rect 15560 -1585 15565 -1565
rect 15565 -1585 15585 -1565
rect 15585 -1585 15590 -1565
rect 15560 -1590 15590 -1585
rect 10760 -1715 10790 -1710
rect 10760 -1735 10765 -1715
rect 10765 -1735 10785 -1715
rect 10785 -1735 10790 -1715
rect 10760 -1740 10790 -1735
rect 16910 -865 16940 -860
rect 16910 -885 16915 -865
rect 16915 -885 16935 -865
rect 16935 -885 16940 -865
rect 16910 -890 16940 -885
rect 17210 -865 17240 -860
rect 17210 -885 17215 -865
rect 17215 -885 17235 -865
rect 17235 -885 17240 -865
rect 17210 -890 17240 -885
rect 17510 -865 17540 -860
rect 17510 -885 17515 -865
rect 17515 -885 17535 -865
rect 17535 -885 17540 -865
rect 17510 -890 17540 -885
rect 17810 -865 17840 -860
rect 17810 -885 17815 -865
rect 17815 -885 17835 -865
rect 17835 -885 17840 -865
rect 17810 -890 17840 -885
rect 18110 -865 18140 -860
rect 18110 -885 18115 -865
rect 18115 -885 18135 -865
rect 18135 -885 18140 -865
rect 18110 -890 18140 -885
rect 18410 -865 18440 -860
rect 18410 -885 18415 -865
rect 18415 -885 18435 -865
rect 18435 -885 18440 -865
rect 18410 -890 18440 -885
rect 18710 -865 18740 -860
rect 18710 -885 18715 -865
rect 18715 -885 18735 -865
rect 18735 -885 18740 -865
rect 18710 -890 18740 -885
rect 19010 -865 19040 -860
rect 19010 -885 19015 -865
rect 19015 -885 19035 -865
rect 19035 -885 19040 -865
rect 19010 -890 19040 -885
rect 20360 -165 20390 -160
rect 20360 -185 20365 -165
rect 20365 -185 20385 -165
rect 20385 -185 20390 -165
rect 20360 -190 20390 -185
rect 20360 -265 20390 -260
rect 20360 -285 20365 -265
rect 20365 -285 20385 -265
rect 20385 -285 20390 -265
rect 20360 -290 20390 -285
rect 20360 -365 20390 -360
rect 20360 -385 20365 -365
rect 20365 -385 20385 -365
rect 20385 -385 20390 -365
rect 20360 -390 20390 -385
rect 20360 -465 20390 -460
rect 20360 -485 20365 -465
rect 20365 -485 20385 -465
rect 20385 -485 20390 -465
rect 20360 -490 20390 -485
rect 20360 -565 20390 -560
rect 20360 -585 20365 -565
rect 20365 -585 20385 -565
rect 20385 -585 20390 -565
rect 20360 -590 20390 -585
rect 20360 -665 20390 -660
rect 20360 -685 20365 -665
rect 20365 -685 20385 -665
rect 20385 -685 20390 -665
rect 20360 -690 20390 -685
rect 20360 -765 20390 -760
rect 20360 -785 20365 -765
rect 20365 -785 20385 -765
rect 20385 -785 20390 -765
rect 20360 -790 20390 -785
rect 19160 -890 19190 -860
rect 17960 -965 17990 -960
rect 17960 -985 17965 -965
rect 17965 -985 17985 -965
rect 17985 -985 17990 -965
rect 17960 -990 17990 -985
rect 17960 -1065 17990 -1060
rect 17960 -1085 17965 -1065
rect 17965 -1085 17985 -1065
rect 17985 -1085 17990 -1065
rect 17960 -1090 17990 -1085
rect 17960 -1165 17990 -1160
rect 17960 -1185 17965 -1165
rect 17965 -1185 17985 -1165
rect 17985 -1185 17990 -1165
rect 17960 -1190 17990 -1185
rect 17960 -1265 17990 -1260
rect 17960 -1285 17965 -1265
rect 17965 -1285 17985 -1265
rect 17985 -1285 17990 -1265
rect 17960 -1290 17990 -1285
rect 17960 -1365 17990 -1360
rect 17960 -1385 17965 -1365
rect 17965 -1385 17985 -1365
rect 17985 -1385 17990 -1365
rect 17960 -1390 17990 -1385
rect 17960 -1465 17990 -1460
rect 17960 -1485 17965 -1465
rect 17965 -1485 17985 -1465
rect 17985 -1485 17990 -1465
rect 17960 -1490 17990 -1485
rect 17960 -1565 17990 -1560
rect 17960 -1585 17965 -1565
rect 17965 -1585 17985 -1565
rect 17985 -1585 17990 -1565
rect 17960 -1590 17990 -1585
rect 15560 -1715 15590 -1710
rect 15560 -1735 15565 -1715
rect 15565 -1735 15585 -1715
rect 15585 -1735 15590 -1715
rect 15560 -1740 15590 -1735
rect 19310 -865 19340 -860
rect 19310 -885 19315 -865
rect 19315 -885 19335 -865
rect 19335 -885 19340 -865
rect 19310 -890 19340 -885
rect 19610 -865 19640 -860
rect 19610 -885 19615 -865
rect 19615 -885 19635 -865
rect 19635 -885 19640 -865
rect 19610 -890 19640 -885
rect 19910 -865 19940 -860
rect 19910 -885 19915 -865
rect 19915 -885 19935 -865
rect 19935 -885 19940 -865
rect 19910 -890 19940 -885
rect 20210 -865 20240 -860
rect 20210 -885 20215 -865
rect 20215 -885 20235 -865
rect 20235 -885 20240 -865
rect 20210 -890 20240 -885
rect 21710 835 21740 840
rect 21710 815 21715 835
rect 21715 815 21735 835
rect 21735 815 21740 835
rect 21710 810 21740 815
rect 22010 835 22040 840
rect 22010 815 22015 835
rect 22015 815 22035 835
rect 22035 815 22040 835
rect 22010 810 22040 815
rect 22310 835 22340 840
rect 22310 815 22315 835
rect 22315 815 22335 835
rect 22335 815 22340 835
rect 22310 810 22340 815
rect 22460 810 22490 840
rect 22610 835 22640 840
rect 22610 815 22615 835
rect 22615 815 22635 835
rect 22635 815 22640 835
rect 22610 810 22640 815
rect 22910 835 22940 840
rect 22910 815 22915 835
rect 22915 815 22935 835
rect 22935 815 22940 835
rect 22910 810 22940 815
rect 23210 835 23240 840
rect 23210 815 23215 835
rect 23215 815 23235 835
rect 23235 815 23240 835
rect 23210 810 23240 815
rect 28760 1685 28790 1690
rect 28760 1665 28765 1685
rect 28765 1665 28785 1685
rect 28785 1665 28790 1685
rect 28760 1660 28790 1665
rect 24560 1535 24590 1540
rect 24560 1515 24565 1535
rect 24565 1515 24585 1535
rect 24585 1515 24590 1535
rect 24560 1510 24590 1515
rect 24560 1435 24590 1440
rect 24560 1415 24565 1435
rect 24565 1415 24585 1435
rect 24585 1415 24590 1435
rect 24560 1410 24590 1415
rect 24560 1335 24590 1340
rect 24560 1315 24565 1335
rect 24565 1315 24585 1335
rect 24585 1315 24590 1335
rect 24560 1310 24590 1315
rect 24560 1235 24590 1240
rect 24560 1215 24565 1235
rect 24565 1215 24585 1235
rect 24585 1215 24590 1235
rect 24560 1210 24590 1215
rect 24560 1135 24590 1140
rect 24560 1115 24565 1135
rect 24565 1115 24585 1135
rect 24585 1115 24590 1135
rect 24560 1110 24590 1115
rect 24560 1035 24590 1040
rect 24560 1015 24565 1035
rect 24565 1015 24585 1035
rect 24585 1015 24590 1035
rect 24560 1010 24590 1015
rect 24560 935 24590 940
rect 24560 915 24565 935
rect 24565 915 24585 935
rect 24585 915 24590 935
rect 24560 910 24590 915
rect 23510 835 23540 840
rect 23510 815 23515 835
rect 23515 815 23535 835
rect 23535 815 23540 835
rect 23510 810 23540 815
rect 23810 835 23840 840
rect 23810 815 23815 835
rect 23815 815 23835 835
rect 23835 815 23840 835
rect 23810 810 23840 815
rect 24110 835 24140 840
rect 24110 815 24115 835
rect 24115 815 24135 835
rect 24135 815 24140 835
rect 24110 810 24140 815
rect 24410 835 24440 840
rect 24410 815 24415 835
rect 24415 815 24435 835
rect 24435 815 24440 835
rect 24410 810 24440 815
rect 20510 -865 20540 -860
rect 20510 -885 20515 -865
rect 20515 -885 20535 -865
rect 20535 -885 20540 -865
rect 20510 -890 20540 -885
rect 20810 -865 20840 -860
rect 20810 -885 20815 -865
rect 20815 -885 20835 -865
rect 20835 -885 20840 -865
rect 20810 -890 20840 -885
rect 21110 -865 21140 -860
rect 21110 -885 21115 -865
rect 21115 -885 21135 -865
rect 21135 -885 21140 -865
rect 21110 -890 21140 -885
rect 21410 -865 21440 -860
rect 21410 -885 21415 -865
rect 21415 -885 21435 -865
rect 21435 -885 21440 -865
rect 21410 -890 21440 -885
rect 20360 -965 20390 -960
rect 20360 -985 20365 -965
rect 20365 -985 20385 -965
rect 20385 -985 20390 -965
rect 20360 -990 20390 -985
rect 20360 -1065 20390 -1060
rect 20360 -1085 20365 -1065
rect 20365 -1085 20385 -1065
rect 20385 -1085 20390 -1065
rect 20360 -1090 20390 -1085
rect 20360 -1165 20390 -1160
rect 20360 -1185 20365 -1165
rect 20365 -1185 20385 -1165
rect 20385 -1185 20390 -1165
rect 20360 -1190 20390 -1185
rect 20360 -1265 20390 -1260
rect 20360 -1285 20365 -1265
rect 20365 -1285 20385 -1265
rect 20385 -1285 20390 -1265
rect 20360 -1290 20390 -1285
rect 20360 -1365 20390 -1360
rect 20360 -1385 20365 -1365
rect 20365 -1385 20385 -1365
rect 20385 -1385 20390 -1365
rect 20360 -1390 20390 -1385
rect 20360 -1465 20390 -1460
rect 20360 -1485 20365 -1465
rect 20365 -1485 20385 -1465
rect 20385 -1485 20390 -1465
rect 20360 -1490 20390 -1485
rect 20360 -1565 20390 -1560
rect 20360 -1585 20365 -1565
rect 20365 -1585 20385 -1565
rect 20385 -1585 20390 -1565
rect 20360 -1590 20390 -1585
rect 17960 -1715 17990 -1710
rect 17960 -1735 17965 -1715
rect 17965 -1735 17985 -1715
rect 17985 -1735 17990 -1715
rect 17960 -1740 17990 -1735
rect 21710 -865 21740 -860
rect 21710 -885 21715 -865
rect 21715 -885 21735 -865
rect 21735 -885 21740 -865
rect 21710 -890 21740 -885
rect 22010 -865 22040 -860
rect 22010 -885 22015 -865
rect 22015 -885 22035 -865
rect 22035 -885 22040 -865
rect 22010 -890 22040 -885
rect 22310 -865 22340 -860
rect 22310 -885 22315 -865
rect 22315 -885 22335 -865
rect 22335 -885 22340 -865
rect 22310 -890 22340 -885
rect 22460 -890 22490 -860
rect 22610 -865 22640 -860
rect 22610 -885 22615 -865
rect 22615 -885 22635 -865
rect 22635 -885 22640 -865
rect 22610 -890 22640 -885
rect 22910 -865 22940 -860
rect 22910 -885 22915 -865
rect 22915 -885 22935 -865
rect 22935 -885 22940 -865
rect 22910 -890 22940 -885
rect 23210 -865 23240 -860
rect 23210 -885 23215 -865
rect 23215 -885 23235 -865
rect 23235 -885 23240 -865
rect 23210 -890 23240 -885
rect 24710 835 24740 840
rect 24710 815 24715 835
rect 24715 815 24735 835
rect 24735 815 24740 835
rect 24710 810 24740 815
rect 25010 835 25040 840
rect 25010 815 25015 835
rect 25015 815 25035 835
rect 25035 815 25040 835
rect 25010 810 25040 815
rect 25310 835 25340 840
rect 25310 815 25315 835
rect 25315 815 25335 835
rect 25335 815 25340 835
rect 25310 810 25340 815
rect 25610 835 25640 840
rect 25610 815 25615 835
rect 25615 815 25635 835
rect 25635 815 25640 835
rect 25610 810 25640 815
rect 25760 810 25790 840
rect 24560 735 24590 740
rect 24560 715 24565 735
rect 24565 715 24585 735
rect 24585 715 24590 735
rect 24560 710 24590 715
rect 24560 635 24590 640
rect 24560 615 24565 635
rect 24565 615 24585 635
rect 24585 615 24590 635
rect 24560 610 24590 615
rect 24560 535 24590 540
rect 24560 515 24565 535
rect 24565 515 24585 535
rect 24585 515 24590 535
rect 24560 510 24590 515
rect 24560 435 24590 440
rect 24560 415 24565 435
rect 24565 415 24585 435
rect 24585 415 24590 435
rect 24560 410 24590 415
rect 24560 335 24590 340
rect 24560 315 24565 335
rect 24565 315 24585 335
rect 24585 315 24590 335
rect 24560 310 24590 315
rect 24560 235 24590 240
rect 24560 215 24565 235
rect 24565 215 24585 235
rect 24585 215 24590 235
rect 24560 210 24590 215
rect 24560 135 24590 140
rect 24560 115 24565 135
rect 24565 115 24585 135
rect 24585 115 24590 135
rect 24560 110 24590 115
rect 25910 835 25940 840
rect 25910 815 25915 835
rect 25915 815 25935 835
rect 25935 815 25940 835
rect 25910 810 25940 815
rect 26210 835 26240 840
rect 26210 815 26215 835
rect 26215 815 26235 835
rect 26235 815 26240 835
rect 26210 810 26240 815
rect 26510 835 26540 840
rect 26510 815 26515 835
rect 26515 815 26535 835
rect 26535 815 26540 835
rect 26510 810 26540 815
rect 26660 810 26690 840
rect 26810 835 26840 840
rect 26810 815 26815 835
rect 26815 815 26835 835
rect 26835 815 26840 835
rect 26810 810 26840 815
rect 27110 835 27140 840
rect 27110 815 27115 835
rect 27115 815 27135 835
rect 27135 815 27140 835
rect 27110 810 27140 815
rect 27410 835 27440 840
rect 27410 815 27415 835
rect 27415 815 27435 835
rect 27435 815 27440 835
rect 27410 810 27440 815
rect 28760 1535 28790 1540
rect 28760 1515 28765 1535
rect 28765 1515 28785 1535
rect 28785 1515 28790 1535
rect 28760 1510 28790 1515
rect 28760 1435 28790 1440
rect 28760 1415 28765 1435
rect 28765 1415 28785 1435
rect 28785 1415 28790 1435
rect 28760 1410 28790 1415
rect 28760 1335 28790 1340
rect 28760 1315 28765 1335
rect 28765 1315 28785 1335
rect 28785 1315 28790 1335
rect 28760 1310 28790 1315
rect 28760 1235 28790 1240
rect 28760 1215 28765 1235
rect 28765 1215 28785 1235
rect 28785 1215 28790 1235
rect 28760 1210 28790 1215
rect 28760 1135 28790 1140
rect 28760 1115 28765 1135
rect 28765 1115 28785 1135
rect 28785 1115 28790 1135
rect 28760 1110 28790 1115
rect 28760 1035 28790 1040
rect 28760 1015 28765 1035
rect 28765 1015 28785 1035
rect 28785 1015 28790 1035
rect 28760 1010 28790 1015
rect 28760 935 28790 940
rect 28760 915 28765 935
rect 28765 915 28785 935
rect 28785 915 28790 935
rect 28760 910 28790 915
rect 27560 810 27590 840
rect 27710 835 27740 840
rect 27710 815 27715 835
rect 27715 815 27735 835
rect 27735 815 27740 835
rect 27710 810 27740 815
rect 28010 835 28040 840
rect 28010 815 28015 835
rect 28015 815 28035 835
rect 28035 815 28040 835
rect 28010 810 28040 815
rect 28310 835 28340 840
rect 28310 815 28315 835
rect 28315 815 28335 835
rect 28335 815 28340 835
rect 28310 810 28340 815
rect 28610 835 28640 840
rect 28610 815 28615 835
rect 28615 815 28635 835
rect 28635 815 28640 835
rect 28610 810 28640 815
rect 28760 735 28790 740
rect 28760 715 28765 735
rect 28765 715 28785 735
rect 28785 715 28790 735
rect 28760 710 28790 715
rect 28760 635 28790 640
rect 28760 615 28765 635
rect 28765 615 28785 635
rect 28785 615 28790 635
rect 28760 610 28790 615
rect 28760 535 28790 540
rect 28760 515 28765 535
rect 28765 515 28785 535
rect 28785 515 28790 535
rect 28760 510 28790 515
rect 28760 435 28790 440
rect 28760 415 28765 435
rect 28765 415 28785 435
rect 28785 415 28790 435
rect 28760 410 28790 415
rect 28760 335 28790 340
rect 28760 315 28765 335
rect 28765 315 28785 335
rect 28785 315 28790 335
rect 28760 310 28790 315
rect 28760 235 28790 240
rect 28760 215 28765 235
rect 28765 215 28785 235
rect 28785 215 28790 235
rect 28760 210 28790 215
rect 28760 135 28790 140
rect 28760 115 28765 135
rect 28765 115 28785 135
rect 28785 115 28790 135
rect 28760 110 28790 115
rect 24560 -15 24590 -10
rect 24560 -35 24565 -15
rect 24565 -35 24585 -15
rect 24585 -35 24590 -15
rect 24560 -40 24590 -35
rect 28760 -15 28790 -10
rect 28760 -35 28765 -15
rect 28765 -35 28785 -15
rect 28785 -35 28790 -15
rect 28760 -40 28790 -35
rect 24560 -165 24590 -160
rect 24560 -185 24565 -165
rect 24565 -185 24585 -165
rect 24585 -185 24590 -165
rect 24560 -190 24590 -185
rect 24560 -265 24590 -260
rect 24560 -285 24565 -265
rect 24565 -285 24585 -265
rect 24585 -285 24590 -265
rect 24560 -290 24590 -285
rect 24560 -365 24590 -360
rect 24560 -385 24565 -365
rect 24565 -385 24585 -365
rect 24585 -385 24590 -365
rect 24560 -390 24590 -385
rect 24560 -465 24590 -460
rect 24560 -485 24565 -465
rect 24565 -485 24585 -465
rect 24585 -485 24590 -465
rect 24560 -490 24590 -485
rect 24560 -565 24590 -560
rect 24560 -585 24565 -565
rect 24565 -585 24585 -565
rect 24585 -585 24590 -565
rect 24560 -590 24590 -585
rect 24560 -665 24590 -660
rect 24560 -685 24565 -665
rect 24565 -685 24585 -665
rect 24585 -685 24590 -665
rect 24560 -690 24590 -685
rect 24560 -765 24590 -760
rect 24560 -785 24565 -765
rect 24565 -785 24585 -765
rect 24585 -785 24590 -765
rect 24560 -790 24590 -785
rect 23510 -865 23540 -860
rect 23510 -885 23515 -865
rect 23515 -885 23535 -865
rect 23535 -885 23540 -865
rect 23510 -890 23540 -885
rect 23810 -865 23840 -860
rect 23810 -885 23815 -865
rect 23815 -885 23835 -865
rect 23835 -885 23840 -865
rect 23810 -890 23840 -885
rect 24110 -865 24140 -860
rect 24110 -885 24115 -865
rect 24115 -885 24135 -865
rect 24135 -885 24140 -865
rect 24110 -890 24140 -885
rect 24410 -865 24440 -860
rect 24410 -885 24415 -865
rect 24415 -885 24435 -865
rect 24435 -885 24440 -865
rect 24410 -890 24440 -885
rect 24710 -865 24740 -860
rect 24710 -885 24715 -865
rect 24715 -885 24735 -865
rect 24735 -885 24740 -865
rect 24710 -890 24740 -885
rect 25010 -865 25040 -860
rect 25010 -885 25015 -865
rect 25015 -885 25035 -865
rect 25035 -885 25040 -865
rect 25010 -890 25040 -885
rect 25310 -865 25340 -860
rect 25310 -885 25315 -865
rect 25315 -885 25335 -865
rect 25335 -885 25340 -865
rect 25310 -890 25340 -885
rect 25610 -865 25640 -860
rect 25610 -885 25615 -865
rect 25615 -885 25635 -865
rect 25635 -885 25640 -865
rect 25610 -890 25640 -885
rect 25760 -890 25790 -860
rect 24560 -965 24590 -960
rect 24560 -985 24565 -965
rect 24565 -985 24585 -965
rect 24585 -985 24590 -965
rect 24560 -990 24590 -985
rect 24560 -1065 24590 -1060
rect 24560 -1085 24565 -1065
rect 24565 -1085 24585 -1065
rect 24585 -1085 24590 -1065
rect 24560 -1090 24590 -1085
rect 24560 -1165 24590 -1160
rect 24560 -1185 24565 -1165
rect 24565 -1185 24585 -1165
rect 24585 -1185 24590 -1165
rect 24560 -1190 24590 -1185
rect 24560 -1265 24590 -1260
rect 24560 -1285 24565 -1265
rect 24565 -1285 24585 -1265
rect 24585 -1285 24590 -1265
rect 24560 -1290 24590 -1285
rect 24560 -1365 24590 -1360
rect 24560 -1385 24565 -1365
rect 24565 -1385 24585 -1365
rect 24585 -1385 24590 -1365
rect 24560 -1390 24590 -1385
rect 24560 -1465 24590 -1460
rect 24560 -1485 24565 -1465
rect 24565 -1485 24585 -1465
rect 24585 -1485 24590 -1465
rect 24560 -1490 24590 -1485
rect 24560 -1565 24590 -1560
rect 24560 -1585 24565 -1565
rect 24565 -1585 24585 -1565
rect 24585 -1585 24590 -1565
rect 24560 -1590 24590 -1585
rect 20360 -1715 20390 -1710
rect 20360 -1735 20365 -1715
rect 20365 -1735 20385 -1715
rect 20385 -1735 20390 -1715
rect 20360 -1740 20390 -1735
rect 25910 -865 25940 -860
rect 25910 -885 25915 -865
rect 25915 -885 25935 -865
rect 25935 -885 25940 -865
rect 25910 -890 25940 -885
rect 26210 -865 26240 -860
rect 26210 -885 26215 -865
rect 26215 -885 26235 -865
rect 26235 -885 26240 -865
rect 26210 -890 26240 -885
rect 26510 -865 26540 -860
rect 26510 -885 26515 -865
rect 26515 -885 26535 -865
rect 26535 -885 26540 -865
rect 26510 -890 26540 -885
rect 26660 -890 26690 -860
rect 26810 -865 26840 -860
rect 26810 -885 26815 -865
rect 26815 -885 26835 -865
rect 26835 -885 26840 -865
rect 26810 -890 26840 -885
rect 27110 -865 27140 -860
rect 27110 -885 27115 -865
rect 27115 -885 27135 -865
rect 27135 -885 27140 -865
rect 27110 -890 27140 -885
rect 27410 -865 27440 -860
rect 27410 -885 27415 -865
rect 27415 -885 27435 -865
rect 27435 -885 27440 -865
rect 27410 -890 27440 -885
rect 28760 -165 28790 -160
rect 28760 -185 28765 -165
rect 28765 -185 28785 -165
rect 28785 -185 28790 -165
rect 28760 -190 28790 -185
rect 28760 -265 28790 -260
rect 28760 -285 28765 -265
rect 28765 -285 28785 -265
rect 28785 -285 28790 -265
rect 28760 -290 28790 -285
rect 28760 -365 28790 -360
rect 28760 -385 28765 -365
rect 28765 -385 28785 -365
rect 28785 -385 28790 -365
rect 28760 -390 28790 -385
rect 28760 -465 28790 -460
rect 28760 -485 28765 -465
rect 28765 -485 28785 -465
rect 28785 -485 28790 -465
rect 28760 -490 28790 -485
rect 28760 -565 28790 -560
rect 28760 -585 28765 -565
rect 28765 -585 28785 -565
rect 28785 -585 28790 -565
rect 28760 -590 28790 -585
rect 28760 -665 28790 -660
rect 28760 -685 28765 -665
rect 28765 -685 28785 -665
rect 28785 -685 28790 -665
rect 28760 -690 28790 -685
rect 28760 -765 28790 -760
rect 28760 -785 28765 -765
rect 28765 -785 28785 -765
rect 28785 -785 28790 -765
rect 28760 -790 28790 -785
rect 27560 -890 27590 -860
rect 27710 -865 27740 -860
rect 27710 -885 27715 -865
rect 27715 -885 27735 -865
rect 27735 -885 27740 -865
rect 27710 -890 27740 -885
rect 28010 -865 28040 -860
rect 28010 -885 28015 -865
rect 28015 -885 28035 -865
rect 28035 -885 28040 -865
rect 28010 -890 28040 -885
rect 28310 -865 28340 -860
rect 28310 -885 28315 -865
rect 28315 -885 28335 -865
rect 28335 -885 28340 -865
rect 28310 -890 28340 -885
rect 28610 -865 28640 -860
rect 28610 -885 28615 -865
rect 28615 -885 28635 -865
rect 28635 -885 28640 -865
rect 28610 -890 28640 -885
rect 28760 -965 28790 -960
rect 28760 -985 28765 -965
rect 28765 -985 28785 -965
rect 28785 -985 28790 -965
rect 28760 -990 28790 -985
rect 28760 -1065 28790 -1060
rect 28760 -1085 28765 -1065
rect 28765 -1085 28785 -1065
rect 28785 -1085 28790 -1065
rect 28760 -1090 28790 -1085
rect 28760 -1165 28790 -1160
rect 28760 -1185 28765 -1165
rect 28765 -1185 28785 -1165
rect 28785 -1185 28790 -1165
rect 28760 -1190 28790 -1185
rect 28760 -1265 28790 -1260
rect 28760 -1285 28765 -1265
rect 28765 -1285 28785 -1265
rect 28785 -1285 28790 -1265
rect 28760 -1290 28790 -1285
rect 28760 -1365 28790 -1360
rect 28760 -1385 28765 -1365
rect 28765 -1385 28785 -1365
rect 28785 -1385 28790 -1365
rect 28760 -1390 28790 -1385
rect 28760 -1465 28790 -1460
rect 28760 -1485 28765 -1465
rect 28765 -1485 28785 -1465
rect 28785 -1485 28790 -1465
rect 28760 -1490 28790 -1485
rect 28760 -1565 28790 -1560
rect 28760 -1585 28765 -1565
rect 28765 -1585 28785 -1565
rect 28785 -1585 28790 -1565
rect 28760 -1590 28790 -1585
rect 24560 -1715 24590 -1710
rect 24560 -1735 24565 -1715
rect 24565 -1735 24585 -1715
rect 24585 -1735 24590 -1715
rect 24560 -1740 24590 -1735
rect 28760 -1715 28790 -1710
rect 28760 -1735 28765 -1715
rect 28765 -1735 28785 -1715
rect 28785 -1735 28790 -1715
rect 28760 -1740 28790 -1735
<< metal2 >>
rect -650 5590 17950 5600
rect -650 5560 -640 5590
rect -610 5560 -40 5590
rect -10 5560 4160 5590
rect 4190 5560 8360 5590
rect 8390 5560 8660 5590
rect 8690 5560 8960 5590
rect 8990 5560 9260 5590
rect 9290 5560 9560 5590
rect 9590 5560 9860 5590
rect 9890 5560 10160 5590
rect 10190 5560 10460 5590
rect 10490 5560 10760 5590
rect 10790 5560 11960 5590
rect 11990 5560 13160 5590
rect 13190 5560 14360 5590
rect 14390 5560 15560 5590
rect 15590 5560 17950 5590
rect -650 5500 17950 5560
rect 18000 5590 32100 5600
rect 18000 5560 20360 5590
rect 20390 5560 22460 5590
rect 22490 5560 24560 5590
rect 24590 5560 26660 5590
rect 26690 5560 28160 5590
rect 28190 5560 28760 5590
rect 28790 5560 32060 5590
rect 32090 5560 32100 5590
rect 18000 5500 32100 5560
rect -650 5440 32100 5450
rect -650 5410 -640 5440
rect -610 5410 8360 5440
rect 8390 5410 8660 5440
rect 8690 5410 8960 5440
rect 8990 5410 9260 5440
rect 9290 5410 9560 5440
rect 9590 5410 9860 5440
rect 9890 5410 10160 5440
rect 10190 5410 10460 5440
rect 10490 5410 10760 5440
rect 10790 5410 11960 5440
rect 11990 5410 13160 5440
rect 13190 5410 14360 5440
rect 14390 5410 15560 5440
rect 15590 5410 20360 5440
rect 20390 5410 22460 5440
rect 22490 5410 24560 5440
rect 24590 5410 26660 5440
rect 26690 5410 28160 5440
rect 28190 5410 28760 5440
rect 28790 5410 32060 5440
rect 32090 5410 32100 5440
rect -650 5400 32100 5410
rect -650 5340 32100 5350
rect -650 5310 -640 5340
rect -610 5310 8360 5340
rect 8390 5310 8660 5340
rect 8690 5310 8960 5340
rect 8990 5310 9260 5340
rect 9290 5310 9560 5340
rect 9590 5310 9860 5340
rect 9890 5310 10160 5340
rect 10190 5310 10460 5340
rect 10490 5310 10760 5340
rect 10790 5310 11960 5340
rect 11990 5310 13160 5340
rect 13190 5310 14360 5340
rect 14390 5310 15560 5340
rect 15590 5310 17960 5340
rect 17990 5310 20360 5340
rect 20390 5310 22460 5340
rect 22490 5310 24560 5340
rect 24590 5310 26660 5340
rect 26690 5310 28160 5340
rect 28190 5310 28760 5340
rect 28790 5310 32060 5340
rect 32090 5310 32100 5340
rect -650 5300 32100 5310
rect -650 5240 32100 5250
rect -650 5210 -640 5240
rect -610 5210 8360 5240
rect 8390 5210 8660 5240
rect 8690 5210 8960 5240
rect 8990 5210 9260 5240
rect 9290 5210 9560 5240
rect 9590 5210 9860 5240
rect 9890 5210 10160 5240
rect 10190 5210 10460 5240
rect 10490 5210 10760 5240
rect 10790 5210 11960 5240
rect 11990 5210 13160 5240
rect 13190 5210 14360 5240
rect 14390 5210 15560 5240
rect 15590 5210 17960 5240
rect 17990 5210 20360 5240
rect 20390 5210 22460 5240
rect 22490 5210 24560 5240
rect 24590 5210 26660 5240
rect 26690 5210 28160 5240
rect 28190 5210 28760 5240
rect 28790 5210 32060 5240
rect 32090 5210 32100 5240
rect -650 5200 32100 5210
rect -650 5140 32100 5150
rect -650 5110 -640 5140
rect -610 5110 8360 5140
rect 8390 5110 8660 5140
rect 8690 5110 8960 5140
rect 8990 5110 9260 5140
rect 9290 5110 9560 5140
rect 9590 5110 9860 5140
rect 9890 5110 10160 5140
rect 10190 5110 10460 5140
rect 10490 5110 10760 5140
rect 10790 5110 11960 5140
rect 11990 5110 13160 5140
rect 13190 5110 14360 5140
rect 14390 5110 15560 5140
rect 15590 5110 17960 5140
rect 17990 5110 20360 5140
rect 20390 5110 22460 5140
rect 22490 5110 24560 5140
rect 24590 5110 26660 5140
rect 26690 5110 28160 5140
rect 28190 5110 28760 5140
rect 28790 5110 32060 5140
rect 32090 5110 32100 5140
rect -650 5100 32100 5110
rect -650 5040 32100 5050
rect -650 5010 -640 5040
rect -610 5010 8360 5040
rect 8390 5010 8660 5040
rect 8690 5010 8960 5040
rect 8990 5010 9260 5040
rect 9290 5010 9560 5040
rect 9590 5010 9860 5040
rect 9890 5010 10160 5040
rect 10190 5010 10460 5040
rect 10490 5010 10760 5040
rect 10790 5010 11960 5040
rect 11990 5010 13160 5040
rect 13190 5010 14360 5040
rect 14390 5010 15560 5040
rect 15590 5010 17960 5040
rect 17990 5010 20360 5040
rect 20390 5010 22460 5040
rect 22490 5010 24560 5040
rect 24590 5010 26660 5040
rect 26690 5010 28160 5040
rect 28190 5010 28760 5040
rect 28790 5010 32060 5040
rect 32090 5010 32100 5040
rect -650 5000 32100 5010
rect -500 4940 -450 4950
rect -500 4910 -490 4940
rect -460 4910 -450 4940
rect -500 4900 -450 4910
rect -350 4940 -300 4950
rect -350 4910 -340 4940
rect -310 4910 -300 4940
rect -350 4900 -300 4910
rect -200 4940 -150 4950
rect -200 4910 -190 4940
rect -160 4910 -150 4940
rect -200 4900 -150 4910
rect 100 4940 150 4950
rect 100 4910 110 4940
rect 140 4910 150 4940
rect 100 4900 150 4910
rect 400 4940 450 4950
rect 400 4910 410 4940
rect 440 4910 450 4940
rect 400 4900 450 4910
rect 700 4940 750 4950
rect 700 4910 710 4940
rect 740 4910 750 4940
rect 700 4900 750 4910
rect 1000 4940 1050 4950
rect 1000 4910 1010 4940
rect 1040 4910 1050 4940
rect 1000 4900 1050 4910
rect 1150 4940 1200 4950
rect 1150 4910 1160 4940
rect 1190 4910 1200 4940
rect 1150 4900 1200 4910
rect 1300 4940 1350 4950
rect 1300 4910 1310 4940
rect 1340 4910 1350 4940
rect 1300 4900 1350 4910
rect 1600 4940 1650 4950
rect 1600 4910 1610 4940
rect 1640 4910 1650 4940
rect 1600 4900 1650 4910
rect 1900 4940 1950 4950
rect 1900 4910 1910 4940
rect 1940 4910 1950 4940
rect 1900 4900 1950 4910
rect 2050 4940 2100 4950
rect 2050 4910 2060 4940
rect 2090 4910 2100 4940
rect 2050 4900 2100 4910
rect 2200 4940 2250 4950
rect 2200 4910 2210 4940
rect 2240 4910 2250 4940
rect 2200 4900 2250 4910
rect 2500 4940 2550 4950
rect 2500 4910 2510 4940
rect 2540 4910 2550 4940
rect 2500 4900 2550 4910
rect 2800 4940 2850 4950
rect 2800 4910 2810 4940
rect 2840 4910 2850 4940
rect 2800 4900 2850 4910
rect 2950 4940 3000 4950
rect 2950 4910 2960 4940
rect 2990 4910 3000 4940
rect 2950 4900 3000 4910
rect 3100 4940 3150 4950
rect 3100 4910 3110 4940
rect 3140 4910 3150 4940
rect 3100 4900 3150 4910
rect 3400 4940 3450 4950
rect 3400 4910 3410 4940
rect 3440 4910 3450 4940
rect 3400 4900 3450 4910
rect 3700 4940 3750 4950
rect 3700 4910 3710 4940
rect 3740 4910 3750 4940
rect 3700 4900 3750 4910
rect 4000 4940 4050 4950
rect 4000 4910 4010 4940
rect 4040 4910 4050 4940
rect 4000 4900 4050 4910
rect 4300 4940 4350 4950
rect 4300 4910 4310 4940
rect 4340 4910 4350 4940
rect 4300 4900 4350 4910
rect 4600 4940 4650 4950
rect 4600 4910 4610 4940
rect 4640 4910 4650 4940
rect 4600 4900 4650 4910
rect 4900 4940 4950 4950
rect 4900 4910 4910 4940
rect 4940 4910 4950 4940
rect 4900 4900 4950 4910
rect 5200 4940 5250 4950
rect 5200 4910 5210 4940
rect 5240 4910 5250 4940
rect 5200 4900 5250 4910
rect 5350 4940 5400 4950
rect 5350 4910 5360 4940
rect 5390 4910 5400 4940
rect 5350 4900 5400 4910
rect 5500 4940 5550 4950
rect 5500 4910 5510 4940
rect 5540 4910 5550 4940
rect 5500 4900 5550 4910
rect 5800 4940 5850 4950
rect 5800 4910 5810 4940
rect 5840 4910 5850 4940
rect 5800 4900 5850 4910
rect 6100 4940 6150 4950
rect 6100 4910 6110 4940
rect 6140 4910 6150 4940
rect 6100 4900 6150 4910
rect 6250 4940 6300 4950
rect 6250 4910 6260 4940
rect 6290 4910 6300 4940
rect 6250 4900 6300 4910
rect 6400 4940 6450 4950
rect 6400 4910 6410 4940
rect 6440 4910 6450 4940
rect 6400 4900 6450 4910
rect 6700 4940 6750 4950
rect 6700 4910 6710 4940
rect 6740 4910 6750 4940
rect 6700 4900 6750 4910
rect 7000 4940 7050 4950
rect 7000 4910 7010 4940
rect 7040 4910 7050 4940
rect 7000 4900 7050 4910
rect 7150 4940 7200 4950
rect 7150 4910 7160 4940
rect 7190 4910 7200 4940
rect 7150 4900 7200 4910
rect 7300 4940 7350 4950
rect 7300 4910 7310 4940
rect 7340 4910 7350 4940
rect 7300 4900 7350 4910
rect 7600 4940 7650 4950
rect 7600 4910 7610 4940
rect 7640 4910 7650 4940
rect 7600 4900 7650 4910
rect 7900 4940 7950 4950
rect 7900 4910 7910 4940
rect 7940 4910 7950 4940
rect 7900 4900 7950 4910
rect 8200 4940 8250 4950
rect 8200 4910 8210 4940
rect 8240 4910 8250 4940
rect 8200 4900 8250 4910
rect 8500 4940 8550 4950
rect 8500 4910 8510 4940
rect 8540 4910 8550 4940
rect 8500 4900 8550 4910
rect 8800 4940 8850 4950
rect 8800 4910 8810 4940
rect 8840 4910 8850 4940
rect 8800 4900 8850 4910
rect 9100 4940 9150 4950
rect 9100 4910 9110 4940
rect 9140 4910 9150 4940
rect 9100 4900 9150 4910
rect 9400 4940 9450 4950
rect 9400 4910 9410 4940
rect 9440 4910 9450 4940
rect 9400 4900 9450 4910
rect 9700 4940 9750 4950
rect 9700 4910 9710 4940
rect 9740 4910 9750 4940
rect 9700 4900 9750 4910
rect 10000 4940 10050 4950
rect 10000 4910 10010 4940
rect 10040 4910 10050 4940
rect 10000 4900 10050 4910
rect 10300 4940 10350 4950
rect 10300 4910 10310 4940
rect 10340 4910 10350 4940
rect 10300 4900 10350 4910
rect 10600 4940 10650 4950
rect 10600 4910 10610 4940
rect 10640 4910 10650 4940
rect 10600 4900 10650 4910
rect 10900 4940 10950 4950
rect 10900 4910 10910 4940
rect 10940 4910 10950 4940
rect 10900 4900 10950 4910
rect 11200 4940 11250 4950
rect 11200 4910 11210 4940
rect 11240 4910 11250 4940
rect 11200 4900 11250 4910
rect 11350 4940 11400 4950
rect 11350 4910 11360 4940
rect 11390 4910 11400 4940
rect 11350 4900 11400 4910
rect 11500 4940 11550 4950
rect 11500 4910 11510 4940
rect 11540 4910 11550 4940
rect 11500 4900 11550 4910
rect 11800 4940 11850 4950
rect 11800 4910 11810 4940
rect 11840 4910 11850 4940
rect 11800 4900 11850 4910
rect 12100 4940 12150 4950
rect 12100 4910 12110 4940
rect 12140 4910 12150 4940
rect 12100 4900 12150 4910
rect 12400 4940 12450 4950
rect 12400 4910 12410 4940
rect 12440 4910 12450 4940
rect 12400 4900 12450 4910
rect 12550 4940 12600 4950
rect 12550 4910 12560 4940
rect 12590 4910 12600 4940
rect 12550 4900 12600 4910
rect 12700 4940 12750 4950
rect 12700 4910 12710 4940
rect 12740 4910 12750 4940
rect 12700 4900 12750 4910
rect 13000 4940 13050 4950
rect 13000 4910 13010 4940
rect 13040 4910 13050 4940
rect 13000 4900 13050 4910
rect 13300 4940 13350 4950
rect 13300 4910 13310 4940
rect 13340 4910 13350 4940
rect 13300 4900 13350 4910
rect 13600 4940 13650 4950
rect 13600 4910 13610 4940
rect 13640 4910 13650 4940
rect 13600 4900 13650 4910
rect 13750 4940 13800 4950
rect 13750 4910 13760 4940
rect 13790 4910 13800 4940
rect 13750 4900 13800 4910
rect 13900 4940 13950 4950
rect 13900 4910 13910 4940
rect 13940 4910 13950 4940
rect 13900 4900 13950 4910
rect 14200 4940 14250 4950
rect 14200 4910 14210 4940
rect 14240 4910 14250 4940
rect 14200 4900 14250 4910
rect 14500 4940 14550 4950
rect 14500 4910 14510 4940
rect 14540 4910 14550 4940
rect 14500 4900 14550 4910
rect 14800 4940 14850 4950
rect 14800 4910 14810 4940
rect 14840 4910 14850 4940
rect 14800 4900 14850 4910
rect 14950 4940 15000 4950
rect 14950 4910 14960 4940
rect 14990 4910 15000 4940
rect 14950 4900 15000 4910
rect 15100 4940 15150 4950
rect 15100 4910 15110 4940
rect 15140 4910 15150 4940
rect 15100 4900 15150 4910
rect 15400 4940 15450 4950
rect 15400 4910 15410 4940
rect 15440 4910 15450 4940
rect 15400 4900 15450 4910
rect 15700 4940 15750 4950
rect 15700 4910 15710 4940
rect 15740 4910 15750 4940
rect 15700 4900 15750 4910
rect 16000 4940 16050 4950
rect 16000 4910 16010 4940
rect 16040 4910 16050 4940
rect 16000 4900 16050 4910
rect 16300 4940 16350 4950
rect 16300 4910 16310 4940
rect 16340 4910 16350 4940
rect 16300 4900 16350 4910
rect 16600 4940 16650 4950
rect 16600 4910 16610 4940
rect 16640 4910 16650 4940
rect 16600 4900 16650 4910
rect 16750 4940 16800 4950
rect 16750 4910 16760 4940
rect 16790 4910 16800 4940
rect 16750 4900 16800 4910
rect 16900 4940 16950 4950
rect 16900 4910 16910 4940
rect 16940 4910 16950 4940
rect 16900 4900 16950 4910
rect 17200 4940 17250 4950
rect 17200 4910 17210 4940
rect 17240 4910 17250 4940
rect 17200 4900 17250 4910
rect 17500 4940 17550 4950
rect 17500 4910 17510 4940
rect 17540 4910 17550 4940
rect 17500 4900 17550 4910
rect 17800 4940 17850 4950
rect 17800 4910 17810 4940
rect 17840 4910 17850 4940
rect 17800 4900 17850 4910
rect 18100 4940 18150 4950
rect 18100 4910 18110 4940
rect 18140 4910 18150 4940
rect 18100 4900 18150 4910
rect 18400 4940 18450 4950
rect 18400 4910 18410 4940
rect 18440 4910 18450 4940
rect 18400 4900 18450 4910
rect 18700 4940 18750 4950
rect 18700 4910 18710 4940
rect 18740 4910 18750 4940
rect 18700 4900 18750 4910
rect 19000 4940 19050 4950
rect 19000 4910 19010 4940
rect 19040 4910 19050 4940
rect 19000 4900 19050 4910
rect 19150 4940 19200 4950
rect 19150 4910 19160 4940
rect 19190 4910 19200 4940
rect 19150 4900 19200 4910
rect 19300 4940 19350 4950
rect 19300 4910 19310 4940
rect 19340 4910 19350 4940
rect 19300 4900 19350 4910
rect 19600 4940 19650 4950
rect 19600 4910 19610 4940
rect 19640 4910 19650 4940
rect 19600 4900 19650 4910
rect 19900 4940 19950 4950
rect 19900 4910 19910 4940
rect 19940 4910 19950 4940
rect 19900 4900 19950 4910
rect 20200 4940 20250 4950
rect 20200 4910 20210 4940
rect 20240 4910 20250 4940
rect 20200 4900 20250 4910
rect 20500 4940 20550 4950
rect 20500 4910 20510 4940
rect 20540 4910 20550 4940
rect 20500 4900 20550 4910
rect 20800 4940 20850 4950
rect 20800 4910 20810 4940
rect 20840 4910 20850 4940
rect 20800 4900 20850 4910
rect 20950 4940 21000 4950
rect 20950 4910 20960 4940
rect 20990 4910 21000 4940
rect 20950 4900 21000 4910
rect 21100 4940 21150 4950
rect 21100 4910 21110 4940
rect 21140 4910 21150 4940
rect 21100 4900 21150 4910
rect 21400 4940 21450 4950
rect 21400 4910 21410 4940
rect 21440 4910 21450 4940
rect 21400 4900 21450 4910
rect 21700 4940 21750 4950
rect 21700 4910 21710 4940
rect 21740 4910 21750 4940
rect 21700 4900 21750 4910
rect 21850 4940 21900 4950
rect 21850 4910 21860 4940
rect 21890 4910 21900 4940
rect 21850 4900 21900 4910
rect 22000 4940 22050 4950
rect 22000 4910 22010 4940
rect 22040 4910 22050 4940
rect 22000 4900 22050 4910
rect 22300 4940 22350 4950
rect 22300 4910 22310 4940
rect 22340 4910 22350 4940
rect 22300 4900 22350 4910
rect 22600 4940 22650 4950
rect 22600 4910 22610 4940
rect 22640 4910 22650 4940
rect 22600 4900 22650 4910
rect 22900 4940 22950 4950
rect 22900 4910 22910 4940
rect 22940 4910 22950 4940
rect 22900 4900 22950 4910
rect 23050 4940 23100 4950
rect 23050 4910 23060 4940
rect 23090 4910 23100 4940
rect 23050 4900 23100 4910
rect 23200 4940 23250 4950
rect 23200 4910 23210 4940
rect 23240 4910 23250 4940
rect 23200 4900 23250 4910
rect 23350 4940 23400 4950
rect 23350 4910 23360 4940
rect 23390 4910 23400 4940
rect 23350 4900 23400 4910
rect 23500 4940 23550 4950
rect 23500 4910 23510 4940
rect 23540 4910 23550 4940
rect 23500 4900 23550 4910
rect 23650 4940 23700 4950
rect 23650 4910 23660 4940
rect 23690 4910 23700 4940
rect 23650 4900 23700 4910
rect 23800 4940 23850 4950
rect 23800 4910 23810 4940
rect 23840 4910 23850 4940
rect 23800 4900 23850 4910
rect 23950 4940 24000 4950
rect 23950 4910 23960 4940
rect 23990 4910 24000 4940
rect 23950 4900 24000 4910
rect 24100 4940 24150 4950
rect 24100 4910 24110 4940
rect 24140 4910 24150 4940
rect 24100 4900 24150 4910
rect 24400 4940 24450 4950
rect 24400 4910 24410 4940
rect 24440 4910 24450 4940
rect 24400 4900 24450 4910
rect 24700 4940 24750 4950
rect 24700 4910 24710 4940
rect 24740 4910 24750 4940
rect 24700 4900 24750 4910
rect 25000 4940 25050 4950
rect 25000 4910 25010 4940
rect 25040 4910 25050 4940
rect 25000 4900 25050 4910
rect 25450 4940 25500 4950
rect 25450 4910 25460 4940
rect 25490 4910 25500 4940
rect 25450 4900 25500 4910
rect 25600 4940 25650 4950
rect 25600 4910 25610 4940
rect 25640 4910 25650 4940
rect 25600 4900 25650 4910
rect 25750 4940 25800 4950
rect 25750 4910 25760 4940
rect 25790 4910 25800 4940
rect 25750 4900 25800 4910
rect 26200 4940 26250 4950
rect 26200 4910 26210 4940
rect 26240 4910 26250 4940
rect 26200 4900 26250 4910
rect 26500 4940 26550 4950
rect 26500 4910 26510 4940
rect 26540 4910 26550 4940
rect 26500 4900 26550 4910
rect 26800 4940 26850 4950
rect 26800 4910 26810 4940
rect 26840 4910 26850 4940
rect 26800 4900 26850 4910
rect 27100 4940 27150 4950
rect 27100 4910 27110 4940
rect 27140 4910 27150 4940
rect 27100 4900 27150 4910
rect 27550 4940 27600 4950
rect 27550 4910 27560 4940
rect 27590 4910 27600 4940
rect 27550 4900 27600 4910
rect 27700 4940 27750 4950
rect 27700 4910 27710 4940
rect 27740 4910 27750 4940
rect 27700 4900 27750 4910
rect 27850 4940 27900 4950
rect 27850 4910 27860 4940
rect 27890 4910 27900 4940
rect 27850 4900 27900 4910
rect 28300 4940 28350 4950
rect 28300 4910 28310 4940
rect 28340 4910 28350 4940
rect 28300 4900 28350 4910
rect 28600 4940 28650 4950
rect 28600 4910 28610 4940
rect 28640 4910 28650 4940
rect 28600 4900 28650 4910
rect 28750 4940 28800 4950
rect 28750 4910 28760 4940
rect 28790 4910 28800 4940
rect 28750 4900 28800 4910
rect 28900 4940 28950 4950
rect 28900 4910 28910 4940
rect 28940 4910 28950 4940
rect 28900 4900 28950 4910
rect 29200 4940 29250 4950
rect 29200 4910 29210 4940
rect 29240 4910 29250 4940
rect 29200 4900 29250 4910
rect 29350 4940 29400 4950
rect 29350 4910 29360 4940
rect 29390 4910 29400 4940
rect 29350 4900 29400 4910
rect 29650 4940 29700 4950
rect 29650 4910 29660 4940
rect 29690 4910 29700 4940
rect 29650 4900 29700 4910
rect 29800 4940 29850 4950
rect 29800 4910 29810 4940
rect 29840 4910 29850 4940
rect 29800 4900 29850 4910
rect 29950 4940 30000 4950
rect 29950 4910 29960 4940
rect 29990 4910 30000 4940
rect 29950 4900 30000 4910
rect 30250 4940 30300 4950
rect 30250 4910 30260 4940
rect 30290 4910 30300 4940
rect 30250 4900 30300 4910
rect 30400 4940 30450 4950
rect 30400 4910 30410 4940
rect 30440 4910 30450 4940
rect 30400 4900 30450 4910
rect 30550 4940 30600 4950
rect 30550 4910 30560 4940
rect 30590 4910 30600 4940
rect 30550 4900 30600 4910
rect 30850 4940 30900 4950
rect 30850 4910 30860 4940
rect 30890 4910 30900 4940
rect 30850 4900 30900 4910
rect 31000 4940 31050 4950
rect 31000 4910 31010 4940
rect 31040 4910 31050 4940
rect 31000 4900 31050 4910
rect 31150 4940 31200 4950
rect 31150 4910 31160 4940
rect 31190 4910 31200 4940
rect 31150 4900 31200 4910
rect 31450 4940 31500 4950
rect 31450 4910 31460 4940
rect 31490 4910 31500 4940
rect 31450 4900 31500 4910
rect 31600 4940 31650 4950
rect 31600 4910 31610 4940
rect 31640 4910 31650 4940
rect 31600 4900 31650 4910
rect 31900 4940 31950 4950
rect 31900 4910 31910 4940
rect 31940 4910 31950 4940
rect 31900 4900 31950 4910
rect 32050 4940 32100 4950
rect 32050 4910 32060 4940
rect 32090 4910 32100 4940
rect 32050 4900 32100 4910
rect -650 4840 32100 4850
rect -650 4810 -640 4840
rect -610 4810 -40 4840
rect -10 4810 4160 4840
rect 4190 4810 8360 4840
rect 8390 4810 8660 4840
rect 8690 4810 8960 4840
rect 8990 4810 9260 4840
rect 9290 4810 9560 4840
rect 9590 4810 9860 4840
rect 9890 4810 10160 4840
rect 10190 4810 10460 4840
rect 10490 4810 10760 4840
rect 10790 4810 11960 4840
rect 11990 4810 13160 4840
rect 13190 4810 14360 4840
rect 14390 4810 15560 4840
rect 15590 4810 17960 4840
rect 17990 4810 20360 4840
rect 20390 4810 22460 4840
rect 22490 4810 24560 4840
rect 24590 4810 26660 4840
rect 26690 4810 28160 4840
rect 28190 4810 28760 4840
rect 28790 4810 32060 4840
rect 32090 4810 32100 4840
rect -650 4800 32100 4810
rect -650 4740 32100 4750
rect -650 4710 -640 4740
rect -610 4710 -40 4740
rect -10 4710 4160 4740
rect 4190 4710 8360 4740
rect 8390 4710 8660 4740
rect 8690 4710 8960 4740
rect 8990 4710 9260 4740
rect 9290 4710 9560 4740
rect 9590 4710 9860 4740
rect 9890 4710 10160 4740
rect 10190 4710 10460 4740
rect 10490 4710 10760 4740
rect 10790 4710 11960 4740
rect 11990 4710 13160 4740
rect 13190 4710 14360 4740
rect 14390 4710 15560 4740
rect 15590 4710 17960 4740
rect 17990 4710 20360 4740
rect 20390 4710 22460 4740
rect 22490 4710 24560 4740
rect 24590 4710 26660 4740
rect 26690 4710 28160 4740
rect 28190 4710 28760 4740
rect 28790 4710 32060 4740
rect 32090 4710 32100 4740
rect -650 4700 32100 4710
rect -650 4640 32100 4650
rect -650 4610 -640 4640
rect -610 4610 -40 4640
rect -10 4610 4160 4640
rect 4190 4610 8360 4640
rect 8390 4610 8660 4640
rect 8690 4610 8960 4640
rect 8990 4610 9260 4640
rect 9290 4610 9560 4640
rect 9590 4610 9860 4640
rect 9890 4610 10160 4640
rect 10190 4610 10460 4640
rect 10490 4610 10760 4640
rect 10790 4610 11960 4640
rect 11990 4610 13160 4640
rect 13190 4610 14360 4640
rect 14390 4610 15560 4640
rect 15590 4610 17960 4640
rect 17990 4610 20360 4640
rect 20390 4610 22460 4640
rect 22490 4610 24560 4640
rect 24590 4610 26660 4640
rect 26690 4610 28160 4640
rect 28190 4610 28760 4640
rect 28790 4610 32060 4640
rect 32090 4610 32100 4640
rect -650 4600 32100 4610
rect -650 4540 32100 4550
rect -650 4510 -640 4540
rect -610 4510 -40 4540
rect -10 4510 4160 4540
rect 4190 4510 8360 4540
rect 8390 4510 8660 4540
rect 8690 4510 8960 4540
rect 8990 4510 9260 4540
rect 9290 4510 9560 4540
rect 9590 4510 9860 4540
rect 9890 4510 10160 4540
rect 10190 4510 10460 4540
rect 10490 4510 10760 4540
rect 10790 4510 11960 4540
rect 11990 4510 13160 4540
rect 13190 4510 14360 4540
rect 14390 4510 15560 4540
rect 15590 4510 17960 4540
rect 17990 4510 20360 4540
rect 20390 4510 22460 4540
rect 22490 4510 24560 4540
rect 24590 4510 26660 4540
rect 26690 4510 28160 4540
rect 28190 4510 28760 4540
rect 28790 4510 32060 4540
rect 32090 4510 32100 4540
rect -650 4500 32100 4510
rect -650 4440 32100 4450
rect -650 4410 -640 4440
rect -610 4410 -40 4440
rect -10 4410 4160 4440
rect 4190 4410 8360 4440
rect 8390 4410 8660 4440
rect 8690 4410 8960 4440
rect 8990 4410 9260 4440
rect 9290 4410 9560 4440
rect 9590 4410 9860 4440
rect 9890 4410 10160 4440
rect 10190 4410 10460 4440
rect 10490 4410 10760 4440
rect 10790 4410 11960 4440
rect 11990 4410 13160 4440
rect 13190 4410 14360 4440
rect 14390 4410 15560 4440
rect 15590 4410 20360 4440
rect 20390 4410 22460 4440
rect 22490 4410 24560 4440
rect 24590 4410 26660 4440
rect 26690 4410 28160 4440
rect 28190 4410 28760 4440
rect 28790 4410 32060 4440
rect 32090 4410 32100 4440
rect -650 4400 32100 4410
rect -650 4290 32100 4350
rect -650 4260 -640 4290
rect -610 4260 -40 4290
rect -10 4260 4160 4290
rect 4190 4260 8360 4290
rect 8390 4260 8660 4290
rect 8690 4260 8960 4290
rect 8990 4260 9260 4290
rect 9290 4260 9560 4290
rect 9590 4260 9860 4290
rect 9890 4260 10160 4290
rect 10190 4260 10460 4290
rect 10490 4260 10760 4290
rect 10790 4260 11960 4290
rect 11990 4260 13160 4290
rect 13190 4260 14360 4290
rect 14390 4260 15560 4290
rect 15590 4260 20360 4290
rect 20390 4260 22460 4290
rect 22490 4260 24560 4290
rect 24590 4260 26660 4290
rect 26690 4260 28160 4290
rect 28190 4260 28760 4290
rect 28790 4260 32060 4290
rect 32090 4260 32100 4290
rect -650 4200 32100 4260
rect -650 4140 32100 4150
rect -650 4110 -640 4140
rect -610 4110 8360 4140
rect 8390 4110 8660 4140
rect 8690 4110 8960 4140
rect 8990 4110 9260 4140
rect 9290 4110 9560 4140
rect 9590 4110 9860 4140
rect 9890 4110 10160 4140
rect 10190 4110 10460 4140
rect 10490 4110 10760 4140
rect 10790 4110 11960 4140
rect 11990 4110 13160 4140
rect 13190 4110 14360 4140
rect 14390 4110 15560 4140
rect 15590 4110 20360 4140
rect 20390 4110 22460 4140
rect 22490 4110 24560 4140
rect 24590 4110 26660 4140
rect 26690 4110 28160 4140
rect 28190 4110 28760 4140
rect 28790 4110 32060 4140
rect 32090 4110 32100 4140
rect -650 4100 32100 4110
rect -650 4040 32100 4050
rect -650 4010 -640 4040
rect -610 4010 8360 4040
rect 8390 4010 8660 4040
rect 8690 4010 8960 4040
rect 8990 4010 9260 4040
rect 9290 4010 9560 4040
rect 9590 4010 9860 4040
rect 9890 4010 10160 4040
rect 10190 4010 10460 4040
rect 10490 4010 10760 4040
rect 10790 4010 11960 4040
rect 11990 4010 13160 4040
rect 13190 4010 14360 4040
rect 14390 4010 15560 4040
rect 15590 4010 17960 4040
rect 17990 4010 20360 4040
rect 20390 4010 22460 4040
rect 22490 4010 24560 4040
rect 24590 4010 26660 4040
rect 26690 4010 28160 4040
rect 28190 4010 28760 4040
rect 28790 4010 32060 4040
rect 32090 4010 32100 4040
rect -650 4000 32100 4010
rect -650 3940 32100 3950
rect -650 3910 -640 3940
rect -610 3910 8360 3940
rect 8390 3910 8660 3940
rect 8690 3910 8960 3940
rect 8990 3910 9260 3940
rect 9290 3910 9560 3940
rect 9590 3910 9860 3940
rect 9890 3910 10160 3940
rect 10190 3910 10460 3940
rect 10490 3910 10760 3940
rect 10790 3910 11960 3940
rect 11990 3910 13160 3940
rect 13190 3910 14360 3940
rect 14390 3910 15560 3940
rect 15590 3910 17960 3940
rect 17990 3910 20360 3940
rect 20390 3910 22460 3940
rect 22490 3910 24560 3940
rect 24590 3910 26660 3940
rect 26690 3910 28160 3940
rect 28190 3910 28760 3940
rect 28790 3910 32060 3940
rect 32090 3910 32100 3940
rect -650 3900 32100 3910
rect -650 3840 32100 3850
rect -650 3810 -640 3840
rect -610 3810 8360 3840
rect 8390 3810 8660 3840
rect 8690 3810 8960 3840
rect 8990 3810 9260 3840
rect 9290 3810 9560 3840
rect 9590 3810 9860 3840
rect 9890 3810 10160 3840
rect 10190 3810 10460 3840
rect 10490 3810 10760 3840
rect 10790 3810 11960 3840
rect 11990 3810 13160 3840
rect 13190 3810 14360 3840
rect 14390 3810 15560 3840
rect 15590 3810 17960 3840
rect 17990 3810 20360 3840
rect 20390 3810 22460 3840
rect 22490 3810 24560 3840
rect 24590 3810 26660 3840
rect 26690 3810 28160 3840
rect 28190 3810 28760 3840
rect 28790 3810 32060 3840
rect 32090 3810 32100 3840
rect -650 3800 32100 3810
rect -650 3740 32100 3750
rect -650 3710 -640 3740
rect -610 3710 8360 3740
rect 8390 3710 8660 3740
rect 8690 3710 8960 3740
rect 8990 3710 9260 3740
rect 9290 3710 9560 3740
rect 9590 3710 9860 3740
rect 9890 3710 10160 3740
rect 10190 3710 10460 3740
rect 10490 3710 10760 3740
rect 10790 3710 11960 3740
rect 11990 3710 13160 3740
rect 13190 3710 14360 3740
rect 14390 3710 15560 3740
rect 15590 3710 17960 3740
rect 17990 3710 20360 3740
rect 20390 3710 22460 3740
rect 22490 3710 24560 3740
rect 24590 3710 26660 3740
rect 26690 3710 28160 3740
rect 28190 3710 28760 3740
rect 28790 3710 32060 3740
rect 32090 3710 32100 3740
rect -650 3700 32100 3710
rect -500 3640 -450 3650
rect -500 3610 -490 3640
rect -460 3610 -450 3640
rect -500 3600 -450 3610
rect -350 3640 -300 3650
rect -350 3610 -340 3640
rect -310 3610 -300 3640
rect -350 3600 -300 3610
rect -200 3640 -150 3650
rect -200 3610 -190 3640
rect -160 3610 -150 3640
rect -200 3600 -150 3610
rect 100 3640 150 3650
rect 100 3610 110 3640
rect 140 3610 150 3640
rect 100 3600 150 3610
rect 400 3640 450 3650
rect 400 3610 410 3640
rect 440 3610 450 3640
rect 400 3600 450 3610
rect 700 3640 750 3650
rect 700 3610 710 3640
rect 740 3610 750 3640
rect 700 3600 750 3610
rect 1000 3640 1050 3650
rect 1000 3610 1010 3640
rect 1040 3610 1050 3640
rect 1000 3600 1050 3610
rect 1150 3640 1200 3650
rect 1150 3610 1160 3640
rect 1190 3610 1200 3640
rect 1150 3600 1200 3610
rect 1300 3640 1350 3650
rect 1300 3610 1310 3640
rect 1340 3610 1350 3640
rect 1300 3600 1350 3610
rect 1600 3640 1650 3650
rect 1600 3610 1610 3640
rect 1640 3610 1650 3640
rect 1600 3600 1650 3610
rect 1900 3640 1950 3650
rect 1900 3610 1910 3640
rect 1940 3610 1950 3640
rect 1900 3600 1950 3610
rect 2050 3640 2100 3650
rect 2050 3610 2060 3640
rect 2090 3610 2100 3640
rect 2050 3600 2100 3610
rect 2200 3640 2250 3650
rect 2200 3610 2210 3640
rect 2240 3610 2250 3640
rect 2200 3600 2250 3610
rect 2500 3640 2550 3650
rect 2500 3610 2510 3640
rect 2540 3610 2550 3640
rect 2500 3600 2550 3610
rect 2800 3640 2850 3650
rect 2800 3610 2810 3640
rect 2840 3610 2850 3640
rect 2800 3600 2850 3610
rect 2950 3640 3000 3650
rect 2950 3610 2960 3640
rect 2990 3610 3000 3640
rect 2950 3600 3000 3610
rect 3100 3640 3150 3650
rect 3100 3610 3110 3640
rect 3140 3610 3150 3640
rect 3100 3600 3150 3610
rect 3400 3640 3450 3650
rect 3400 3610 3410 3640
rect 3440 3610 3450 3640
rect 3400 3600 3450 3610
rect 3700 3640 3750 3650
rect 3700 3610 3710 3640
rect 3740 3610 3750 3640
rect 3700 3600 3750 3610
rect 4000 3640 4050 3650
rect 4000 3610 4010 3640
rect 4040 3610 4050 3640
rect 4000 3600 4050 3610
rect 4300 3640 4350 3650
rect 4300 3610 4310 3640
rect 4340 3610 4350 3640
rect 4300 3600 4350 3610
rect 4600 3640 4650 3650
rect 4600 3610 4610 3640
rect 4640 3610 4650 3640
rect 4600 3600 4650 3610
rect 4900 3640 4950 3650
rect 4900 3610 4910 3640
rect 4940 3610 4950 3640
rect 4900 3600 4950 3610
rect 5200 3640 5250 3650
rect 5200 3610 5210 3640
rect 5240 3610 5250 3640
rect 5200 3600 5250 3610
rect 5350 3640 5400 3650
rect 5350 3610 5360 3640
rect 5390 3610 5400 3640
rect 5350 3600 5400 3610
rect 5500 3640 5550 3650
rect 5500 3610 5510 3640
rect 5540 3610 5550 3640
rect 5500 3600 5550 3610
rect 5800 3640 5850 3650
rect 5800 3610 5810 3640
rect 5840 3610 5850 3640
rect 5800 3600 5850 3610
rect 6100 3640 6150 3650
rect 6100 3610 6110 3640
rect 6140 3610 6150 3640
rect 6100 3600 6150 3610
rect 6250 3640 6300 3650
rect 6250 3610 6260 3640
rect 6290 3610 6300 3640
rect 6250 3600 6300 3610
rect 6400 3640 6450 3650
rect 6400 3610 6410 3640
rect 6440 3610 6450 3640
rect 6400 3600 6450 3610
rect 6700 3640 6750 3650
rect 6700 3610 6710 3640
rect 6740 3610 6750 3640
rect 6700 3600 6750 3610
rect 7000 3640 7050 3650
rect 7000 3610 7010 3640
rect 7040 3610 7050 3640
rect 7000 3600 7050 3610
rect 7150 3640 7200 3650
rect 7150 3610 7160 3640
rect 7190 3610 7200 3640
rect 7150 3600 7200 3610
rect 7300 3640 7350 3650
rect 7300 3610 7310 3640
rect 7340 3610 7350 3640
rect 7300 3600 7350 3610
rect 7600 3640 7650 3650
rect 7600 3610 7610 3640
rect 7640 3610 7650 3640
rect 7600 3600 7650 3610
rect 7900 3640 7950 3650
rect 7900 3610 7910 3640
rect 7940 3610 7950 3640
rect 7900 3600 7950 3610
rect 8200 3640 8250 3650
rect 8200 3610 8210 3640
rect 8240 3610 8250 3640
rect 8200 3600 8250 3610
rect 8500 3640 8550 3650
rect 8500 3610 8510 3640
rect 8540 3610 8550 3640
rect 8500 3600 8550 3610
rect 8800 3640 8850 3650
rect 8800 3610 8810 3640
rect 8840 3610 8850 3640
rect 8800 3600 8850 3610
rect 9100 3640 9150 3650
rect 9100 3610 9110 3640
rect 9140 3610 9150 3640
rect 9100 3600 9150 3610
rect 9400 3640 9450 3650
rect 9400 3610 9410 3640
rect 9440 3610 9450 3640
rect 9400 3600 9450 3610
rect 9700 3640 9750 3650
rect 9700 3610 9710 3640
rect 9740 3610 9750 3640
rect 9700 3600 9750 3610
rect 10000 3640 10050 3650
rect 10000 3610 10010 3640
rect 10040 3610 10050 3640
rect 10000 3600 10050 3610
rect 10300 3640 10350 3650
rect 10300 3610 10310 3640
rect 10340 3610 10350 3640
rect 10300 3600 10350 3610
rect 10600 3640 10650 3650
rect 10600 3610 10610 3640
rect 10640 3610 10650 3640
rect 10600 3600 10650 3610
rect 10900 3640 10950 3650
rect 10900 3610 10910 3640
rect 10940 3610 10950 3640
rect 10900 3600 10950 3610
rect 11200 3640 11250 3650
rect 11200 3610 11210 3640
rect 11240 3610 11250 3640
rect 11200 3600 11250 3610
rect 11350 3640 11400 3650
rect 11350 3610 11360 3640
rect 11390 3610 11400 3640
rect 11350 3600 11400 3610
rect 11500 3640 11550 3650
rect 11500 3610 11510 3640
rect 11540 3610 11550 3640
rect 11500 3600 11550 3610
rect 11800 3640 11850 3650
rect 11800 3610 11810 3640
rect 11840 3610 11850 3640
rect 11800 3600 11850 3610
rect 12100 3640 12150 3650
rect 12100 3610 12110 3640
rect 12140 3610 12150 3640
rect 12100 3600 12150 3610
rect 12400 3640 12450 3650
rect 12400 3610 12410 3640
rect 12440 3610 12450 3640
rect 12400 3600 12450 3610
rect 12550 3640 12600 3650
rect 12550 3610 12560 3640
rect 12590 3610 12600 3640
rect 12550 3600 12600 3610
rect 12700 3640 12750 3650
rect 12700 3610 12710 3640
rect 12740 3610 12750 3640
rect 12700 3600 12750 3610
rect 13000 3640 13050 3650
rect 13000 3610 13010 3640
rect 13040 3610 13050 3640
rect 13000 3600 13050 3610
rect 13300 3640 13350 3650
rect 13300 3610 13310 3640
rect 13340 3610 13350 3640
rect 13300 3600 13350 3610
rect 13600 3640 13650 3650
rect 13600 3610 13610 3640
rect 13640 3610 13650 3640
rect 13600 3600 13650 3610
rect 13750 3640 13800 3650
rect 13750 3610 13760 3640
rect 13790 3610 13800 3640
rect 13750 3600 13800 3610
rect 13900 3640 13950 3650
rect 13900 3610 13910 3640
rect 13940 3610 13950 3640
rect 13900 3600 13950 3610
rect 14200 3640 14250 3650
rect 14200 3610 14210 3640
rect 14240 3610 14250 3640
rect 14200 3600 14250 3610
rect 14500 3640 14550 3650
rect 14500 3610 14510 3640
rect 14540 3610 14550 3640
rect 14500 3600 14550 3610
rect 14800 3640 14850 3650
rect 14800 3610 14810 3640
rect 14840 3610 14850 3640
rect 14800 3600 14850 3610
rect 14950 3640 15000 3650
rect 14950 3610 14960 3640
rect 14990 3610 15000 3640
rect 14950 3600 15000 3610
rect 15100 3640 15150 3650
rect 15100 3610 15110 3640
rect 15140 3610 15150 3640
rect 15100 3600 15150 3610
rect 15400 3640 15450 3650
rect 15400 3610 15410 3640
rect 15440 3610 15450 3640
rect 15400 3600 15450 3610
rect 15700 3640 15750 3650
rect 15700 3610 15710 3640
rect 15740 3610 15750 3640
rect 15700 3600 15750 3610
rect 16000 3640 16050 3650
rect 16000 3610 16010 3640
rect 16040 3610 16050 3640
rect 16000 3600 16050 3610
rect 16300 3640 16350 3650
rect 16300 3610 16310 3640
rect 16340 3610 16350 3640
rect 16300 3600 16350 3610
rect 16600 3640 16650 3650
rect 16600 3610 16610 3640
rect 16640 3610 16650 3640
rect 16600 3600 16650 3610
rect 16750 3640 16800 3650
rect 16750 3610 16760 3640
rect 16790 3610 16800 3640
rect 16750 3600 16800 3610
rect 16900 3640 16950 3650
rect 16900 3610 16910 3640
rect 16940 3610 16950 3640
rect 16900 3600 16950 3610
rect 17200 3640 17250 3650
rect 17200 3610 17210 3640
rect 17240 3610 17250 3640
rect 17200 3600 17250 3610
rect 17500 3640 17550 3650
rect 17500 3610 17510 3640
rect 17540 3610 17550 3640
rect 17500 3600 17550 3610
rect 17800 3640 17850 3650
rect 17800 3610 17810 3640
rect 17840 3610 17850 3640
rect 17800 3600 17850 3610
rect 18100 3640 18150 3650
rect 18100 3610 18110 3640
rect 18140 3610 18150 3640
rect 18100 3600 18150 3610
rect 18400 3640 18450 3650
rect 18400 3610 18410 3640
rect 18440 3610 18450 3640
rect 18400 3600 18450 3610
rect 18700 3640 18750 3650
rect 18700 3610 18710 3640
rect 18740 3610 18750 3640
rect 18700 3600 18750 3610
rect 19000 3640 19050 3650
rect 19000 3610 19010 3640
rect 19040 3610 19050 3640
rect 19000 3600 19050 3610
rect 19150 3640 19200 3650
rect 19150 3610 19160 3640
rect 19190 3610 19200 3640
rect 19150 3600 19200 3610
rect 19300 3640 19350 3650
rect 19300 3610 19310 3640
rect 19340 3610 19350 3640
rect 19300 3600 19350 3610
rect 19600 3640 19650 3650
rect 19600 3610 19610 3640
rect 19640 3610 19650 3640
rect 19600 3600 19650 3610
rect 19900 3640 19950 3650
rect 19900 3610 19910 3640
rect 19940 3610 19950 3640
rect 19900 3600 19950 3610
rect 20200 3640 20250 3650
rect 20200 3610 20210 3640
rect 20240 3610 20250 3640
rect 20200 3600 20250 3610
rect 20500 3640 20550 3650
rect 20500 3610 20510 3640
rect 20540 3610 20550 3640
rect 20500 3600 20550 3610
rect 20800 3640 20850 3650
rect 20800 3610 20810 3640
rect 20840 3610 20850 3640
rect 20800 3600 20850 3610
rect 20950 3640 21000 3650
rect 20950 3610 20960 3640
rect 20990 3610 21000 3640
rect 20950 3600 21000 3610
rect 21100 3640 21150 3650
rect 21100 3610 21110 3640
rect 21140 3610 21150 3640
rect 21100 3600 21150 3610
rect 21400 3640 21450 3650
rect 21400 3610 21410 3640
rect 21440 3610 21450 3640
rect 21400 3600 21450 3610
rect 21700 3640 21750 3650
rect 21700 3610 21710 3640
rect 21740 3610 21750 3640
rect 21700 3600 21750 3610
rect 21850 3640 21900 3650
rect 21850 3610 21860 3640
rect 21890 3610 21900 3640
rect 21850 3600 21900 3610
rect 22000 3640 22050 3650
rect 22000 3610 22010 3640
rect 22040 3610 22050 3640
rect 22000 3600 22050 3610
rect 22300 3640 22350 3650
rect 22300 3610 22310 3640
rect 22340 3610 22350 3640
rect 22300 3600 22350 3610
rect 22600 3640 22650 3650
rect 22600 3610 22610 3640
rect 22640 3610 22650 3640
rect 22600 3600 22650 3610
rect 22900 3640 22950 3650
rect 22900 3610 22910 3640
rect 22940 3610 22950 3640
rect 22900 3600 22950 3610
rect 23050 3640 23100 3650
rect 23050 3610 23060 3640
rect 23090 3610 23100 3640
rect 23050 3600 23100 3610
rect 23200 3640 23250 3650
rect 23200 3610 23210 3640
rect 23240 3610 23250 3640
rect 23200 3600 23250 3610
rect 23350 3640 23400 3650
rect 23350 3610 23360 3640
rect 23390 3610 23400 3640
rect 23350 3600 23400 3610
rect 23500 3640 23550 3650
rect 23500 3610 23510 3640
rect 23540 3610 23550 3640
rect 23500 3600 23550 3610
rect 23650 3640 23700 3650
rect 23650 3610 23660 3640
rect 23690 3610 23700 3640
rect 23650 3600 23700 3610
rect 23800 3640 23850 3650
rect 23800 3610 23810 3640
rect 23840 3610 23850 3640
rect 23800 3600 23850 3610
rect 23950 3640 24000 3650
rect 23950 3610 23960 3640
rect 23990 3610 24000 3640
rect 23950 3600 24000 3610
rect 24100 3640 24150 3650
rect 24100 3610 24110 3640
rect 24140 3610 24150 3640
rect 24100 3600 24150 3610
rect 24400 3640 24450 3650
rect 24400 3610 24410 3640
rect 24440 3610 24450 3640
rect 24400 3600 24450 3610
rect 24700 3640 24750 3650
rect 24700 3610 24710 3640
rect 24740 3610 24750 3640
rect 24700 3600 24750 3610
rect 25000 3640 25050 3650
rect 25000 3610 25010 3640
rect 25040 3610 25050 3640
rect 25000 3600 25050 3610
rect 25450 3640 25500 3650
rect 25450 3610 25460 3640
rect 25490 3610 25500 3640
rect 25450 3600 25500 3610
rect 25600 3640 25650 3650
rect 25600 3610 25610 3640
rect 25640 3610 25650 3640
rect 25600 3600 25650 3610
rect 25750 3640 25800 3650
rect 25750 3610 25760 3640
rect 25790 3610 25800 3640
rect 25750 3600 25800 3610
rect 26200 3640 26250 3650
rect 26200 3610 26210 3640
rect 26240 3610 26250 3640
rect 26200 3600 26250 3610
rect 26500 3640 26550 3650
rect 26500 3610 26510 3640
rect 26540 3610 26550 3640
rect 26500 3600 26550 3610
rect 26800 3640 26850 3650
rect 26800 3610 26810 3640
rect 26840 3610 26850 3640
rect 26800 3600 26850 3610
rect 27100 3640 27150 3650
rect 27100 3610 27110 3640
rect 27140 3610 27150 3640
rect 27100 3600 27150 3610
rect 27550 3640 27600 3650
rect 27550 3610 27560 3640
rect 27590 3610 27600 3640
rect 27550 3600 27600 3610
rect 27700 3640 27750 3650
rect 27700 3610 27710 3640
rect 27740 3610 27750 3640
rect 27700 3600 27750 3610
rect 27850 3640 27900 3650
rect 27850 3610 27860 3640
rect 27890 3610 27900 3640
rect 27850 3600 27900 3610
rect 28300 3640 28350 3650
rect 28300 3610 28310 3640
rect 28340 3610 28350 3640
rect 28300 3600 28350 3610
rect 28600 3640 28650 3650
rect 28600 3610 28610 3640
rect 28640 3610 28650 3640
rect 28600 3600 28650 3610
rect 28750 3640 28800 3650
rect 28750 3610 28760 3640
rect 28790 3610 28800 3640
rect 28750 3600 28800 3610
rect 28900 3640 28950 3650
rect 28900 3610 28910 3640
rect 28940 3610 28950 3640
rect 28900 3600 28950 3610
rect 29200 3640 29250 3650
rect 29200 3610 29210 3640
rect 29240 3610 29250 3640
rect 29200 3600 29250 3610
rect 29350 3640 29400 3650
rect 29350 3610 29360 3640
rect 29390 3610 29400 3640
rect 29350 3600 29400 3610
rect 29650 3640 29700 3650
rect 29650 3610 29660 3640
rect 29690 3610 29700 3640
rect 29650 3600 29700 3610
rect 29800 3640 29850 3650
rect 29800 3610 29810 3640
rect 29840 3610 29850 3640
rect 29800 3600 29850 3610
rect 29950 3640 30000 3650
rect 29950 3610 29960 3640
rect 29990 3610 30000 3640
rect 29950 3600 30000 3610
rect 30250 3640 30300 3650
rect 30250 3610 30260 3640
rect 30290 3610 30300 3640
rect 30250 3600 30300 3610
rect 30400 3640 30450 3650
rect 30400 3610 30410 3640
rect 30440 3610 30450 3640
rect 30400 3600 30450 3610
rect 30550 3640 30600 3650
rect 30550 3610 30560 3640
rect 30590 3610 30600 3640
rect 30550 3600 30600 3610
rect 30850 3640 30900 3650
rect 30850 3610 30860 3640
rect 30890 3610 30900 3640
rect 30850 3600 30900 3610
rect 31000 3640 31050 3650
rect 31000 3610 31010 3640
rect 31040 3610 31050 3640
rect 31000 3600 31050 3610
rect 31150 3640 31200 3650
rect 31150 3610 31160 3640
rect 31190 3610 31200 3640
rect 31150 3600 31200 3610
rect 31450 3640 31500 3650
rect 31450 3610 31460 3640
rect 31490 3610 31500 3640
rect 31450 3600 31500 3610
rect 31600 3640 31650 3650
rect 31600 3610 31610 3640
rect 31640 3610 31650 3640
rect 31600 3600 31650 3610
rect 31900 3640 31950 3650
rect 31900 3610 31910 3640
rect 31940 3610 31950 3640
rect 31900 3600 31950 3610
rect 32050 3640 32100 3650
rect 32050 3610 32060 3640
rect 32090 3610 32100 3640
rect 32050 3600 32100 3610
rect -650 3540 32100 3550
rect -650 3510 -640 3540
rect -610 3510 -40 3540
rect -10 3510 4160 3540
rect 4190 3510 8360 3540
rect 8390 3510 8660 3540
rect 8690 3510 8960 3540
rect 8990 3510 9260 3540
rect 9290 3510 9560 3540
rect 9590 3510 9860 3540
rect 9890 3510 10160 3540
rect 10190 3510 10460 3540
rect 10490 3510 10760 3540
rect 10790 3510 11960 3540
rect 11990 3510 13160 3540
rect 13190 3510 14360 3540
rect 14390 3510 15560 3540
rect 15590 3510 17960 3540
rect 17990 3510 20360 3540
rect 20390 3510 22460 3540
rect 22490 3510 24560 3540
rect 24590 3510 26660 3540
rect 26690 3510 28160 3540
rect 28190 3510 28760 3540
rect 28790 3510 32060 3540
rect 32090 3510 32100 3540
rect -650 3500 32100 3510
rect -650 3440 32100 3450
rect -650 3410 -640 3440
rect -610 3410 -40 3440
rect -10 3410 4160 3440
rect 4190 3410 8360 3440
rect 8390 3410 8660 3440
rect 8690 3410 8960 3440
rect 8990 3410 9260 3440
rect 9290 3410 9560 3440
rect 9590 3410 9860 3440
rect 9890 3410 10160 3440
rect 10190 3410 10460 3440
rect 10490 3410 10760 3440
rect 10790 3410 11960 3440
rect 11990 3410 13160 3440
rect 13190 3410 14360 3440
rect 14390 3410 15560 3440
rect 15590 3410 17960 3440
rect 17990 3410 20360 3440
rect 20390 3410 22460 3440
rect 22490 3410 24560 3440
rect 24590 3410 26660 3440
rect 26690 3410 28160 3440
rect 28190 3410 28760 3440
rect 28790 3410 32060 3440
rect 32090 3410 32100 3440
rect -650 3400 32100 3410
rect -650 3340 32100 3350
rect -650 3310 -640 3340
rect -610 3310 -40 3340
rect -10 3310 4160 3340
rect 4190 3310 8360 3340
rect 8390 3310 8660 3340
rect 8690 3310 8960 3340
rect 8990 3310 9260 3340
rect 9290 3310 9560 3340
rect 9590 3310 9860 3340
rect 9890 3310 10160 3340
rect 10190 3310 10460 3340
rect 10490 3310 10760 3340
rect 10790 3310 11960 3340
rect 11990 3310 13160 3340
rect 13190 3310 14360 3340
rect 14390 3310 15560 3340
rect 15590 3310 17960 3340
rect 17990 3310 20360 3340
rect 20390 3310 22460 3340
rect 22490 3310 24560 3340
rect 24590 3310 26660 3340
rect 26690 3310 28160 3340
rect 28190 3310 28760 3340
rect 28790 3310 32060 3340
rect 32090 3310 32100 3340
rect -650 3300 32100 3310
rect -650 3240 32100 3250
rect -650 3210 -640 3240
rect -610 3210 -40 3240
rect -10 3210 4160 3240
rect 4190 3210 8360 3240
rect 8390 3210 8660 3240
rect 8690 3210 8960 3240
rect 8990 3210 9260 3240
rect 9290 3210 9560 3240
rect 9590 3210 9860 3240
rect 9890 3210 10160 3240
rect 10190 3210 10460 3240
rect 10490 3210 10760 3240
rect 10790 3210 11960 3240
rect 11990 3210 13160 3240
rect 13190 3210 14360 3240
rect 14390 3210 15560 3240
rect 15590 3210 17960 3240
rect 17990 3210 20360 3240
rect 20390 3210 22460 3240
rect 22490 3210 24560 3240
rect 24590 3210 26660 3240
rect 26690 3210 28160 3240
rect 28190 3210 28760 3240
rect 28790 3210 32060 3240
rect 32090 3210 32100 3240
rect -650 3200 32100 3210
rect -650 3140 32100 3150
rect -650 3110 -640 3140
rect -610 3110 -40 3140
rect -10 3110 4160 3140
rect 4190 3110 8360 3140
rect 8390 3110 8660 3140
rect 8690 3110 8960 3140
rect 8990 3110 9260 3140
rect 9290 3110 9560 3140
rect 9590 3110 9860 3140
rect 9890 3110 10160 3140
rect 10190 3110 10460 3140
rect 10490 3110 10760 3140
rect 10790 3110 11960 3140
rect 11990 3110 13160 3140
rect 13190 3110 14360 3140
rect 14390 3110 15560 3140
rect 15590 3110 20360 3140
rect 20390 3110 22460 3140
rect 22490 3110 24560 3140
rect 24590 3110 26660 3140
rect 26690 3110 28160 3140
rect 28190 3110 28760 3140
rect 28790 3110 32060 3140
rect 32090 3110 32100 3140
rect -650 3100 32100 3110
rect -650 3000 32100 3050
rect -650 2990 17950 3000
rect -650 2960 -640 2990
rect -610 2960 -40 2990
rect -10 2960 4160 2990
rect 4190 2960 8360 2990
rect 8390 2960 8660 2990
rect 8690 2960 8960 2990
rect 8990 2960 9260 2990
rect 9290 2960 9560 2990
rect 9590 2960 9860 2990
rect 9890 2960 10160 2990
rect 10190 2960 10460 2990
rect 10490 2960 10760 2990
rect 10790 2960 11960 2990
rect 11990 2960 13160 2990
rect 13190 2960 14360 2990
rect 14390 2960 15560 2990
rect 15590 2960 17950 2990
rect -650 2950 17950 2960
rect 18000 2990 32100 3000
rect 18000 2960 20360 2990
rect 20390 2960 24560 2990
rect 24590 2960 26660 2990
rect 26690 2960 28160 2990
rect 28190 2960 28760 2990
rect 28790 2960 32060 2990
rect 32090 2960 32100 2990
rect 18000 2950 32100 2960
rect -900 2800 32100 2850
rect -900 2700 28800 2750
rect -900 2600 28800 2650
rect -900 2300 28800 2550
rect -900 2200 28800 2250
rect -900 2100 28800 2150
rect -900 2000 28800 2050
rect -900 1690 28800 1700
rect -900 1660 -640 1690
rect -610 1660 -40 1690
rect -10 1660 8360 1690
rect 8390 1660 10760 1690
rect 10790 1660 15560 1690
rect 15590 1660 17960 1690
rect 17990 1660 20360 1690
rect 20390 1660 24560 1690
rect 24590 1660 28760 1690
rect 28790 1660 28800 1690
rect -900 1640 28800 1660
rect -900 1610 -640 1640
rect -610 1610 -40 1640
rect -10 1610 8360 1640
rect 8390 1610 10760 1640
rect 10790 1610 15560 1640
rect 15590 1610 17960 1640
rect 17990 1610 20360 1640
rect 20390 1610 24560 1640
rect 24590 1610 28760 1640
rect 28790 1610 28800 1640
rect -900 1600 28800 1610
rect -900 1540 28800 1550
rect -900 1510 -640 1540
rect -610 1510 -40 1540
rect -10 1510 8360 1540
rect 8390 1510 10760 1540
rect 10790 1510 15560 1540
rect 15590 1510 17960 1540
rect 17990 1510 20360 1540
rect 20390 1510 24560 1540
rect 24590 1510 28760 1540
rect 28790 1510 28800 1540
rect -900 1500 28800 1510
rect -900 1440 28800 1450
rect -900 1410 -640 1440
rect -610 1410 -40 1440
rect -10 1410 8360 1440
rect 8390 1410 10760 1440
rect 10790 1410 15560 1440
rect 15590 1410 17960 1440
rect 17990 1410 20360 1440
rect 20390 1410 24560 1440
rect 24590 1410 28760 1440
rect 28790 1410 28800 1440
rect -900 1400 28800 1410
rect -900 1340 28800 1350
rect -900 1310 -640 1340
rect -610 1310 -40 1340
rect -10 1310 8360 1340
rect 8390 1310 10760 1340
rect 10790 1310 15560 1340
rect 15590 1310 17960 1340
rect 17990 1310 20360 1340
rect 20390 1310 24560 1340
rect 24590 1310 28760 1340
rect 28790 1310 28800 1340
rect -900 1300 28800 1310
rect -900 1240 28800 1250
rect -900 1210 -640 1240
rect -610 1210 -40 1240
rect -10 1210 8360 1240
rect 8390 1210 10760 1240
rect 10790 1210 15560 1240
rect 15590 1210 17960 1240
rect 17990 1210 20360 1240
rect 20390 1210 24560 1240
rect 24590 1210 28760 1240
rect 28790 1210 28800 1240
rect -900 1200 28800 1210
rect -900 1140 28800 1150
rect -900 1110 -640 1140
rect -610 1110 -40 1140
rect -10 1110 8360 1140
rect 8390 1110 10760 1140
rect 10790 1110 15560 1140
rect 15590 1110 17960 1140
rect 17990 1110 20360 1140
rect 20390 1110 24560 1140
rect 24590 1110 28760 1140
rect 28790 1110 28800 1140
rect -900 1100 28800 1110
rect -900 1040 28800 1050
rect -900 1010 -640 1040
rect -610 1010 -40 1040
rect -10 1010 8360 1040
rect 8390 1010 10760 1040
rect 10790 1010 15560 1040
rect 15590 1010 17960 1040
rect 17990 1010 20360 1040
rect 20390 1010 24560 1040
rect 24590 1010 28760 1040
rect 28790 1010 28800 1040
rect -900 1000 28800 1010
rect -900 940 28800 950
rect -900 910 -640 940
rect -610 910 -40 940
rect -10 910 8360 940
rect 8390 910 10760 940
rect 10790 910 15560 940
rect 15590 910 17960 940
rect 17990 910 20360 940
rect 20390 910 24560 940
rect 24590 910 28760 940
rect 28790 910 28800 940
rect -900 900 28800 910
rect -500 840 -450 850
rect -500 810 -490 840
rect -460 810 -450 840
rect -500 800 -450 810
rect -350 840 -300 850
rect -350 810 -340 840
rect -310 810 -300 840
rect -350 800 -300 810
rect -200 840 -150 850
rect -200 810 -190 840
rect -160 810 -150 840
rect -200 800 -150 810
rect 100 840 150 850
rect 100 810 110 840
rect 140 810 150 840
rect 100 800 150 810
rect 400 840 450 850
rect 400 810 410 840
rect 440 810 450 840
rect 400 800 450 810
rect 700 840 750 850
rect 700 810 710 840
rect 740 810 750 840
rect 700 800 750 810
rect 1000 840 1050 850
rect 1000 810 1010 840
rect 1040 810 1050 840
rect 1000 800 1050 810
rect 1300 840 1350 850
rect 1300 810 1310 840
rect 1340 810 1350 840
rect 1300 800 1350 810
rect 1600 840 1650 850
rect 1600 810 1610 840
rect 1640 810 1650 840
rect 1600 800 1650 810
rect 1900 840 1950 850
rect 1900 810 1910 840
rect 1940 810 1950 840
rect 1900 800 1950 810
rect 2200 840 2250 850
rect 2200 810 2210 840
rect 2240 810 2250 840
rect 2200 800 2250 810
rect 2350 840 2400 850
rect 2350 810 2360 840
rect 2390 810 2400 840
rect 2350 800 2400 810
rect 2500 840 2550 850
rect 2500 810 2510 840
rect 2540 810 2550 840
rect 2500 800 2550 810
rect 2800 840 2850 850
rect 2800 810 2810 840
rect 2840 810 2850 840
rect 2800 800 2850 810
rect 3100 840 3150 850
rect 3100 810 3110 840
rect 3140 810 3150 840
rect 3100 800 3150 810
rect 3400 840 3450 850
rect 3400 810 3410 840
rect 3440 810 3450 840
rect 3400 800 3450 810
rect 3700 840 3750 850
rect 3700 810 3710 840
rect 3740 810 3750 840
rect 3700 800 3750 810
rect 3850 840 3900 850
rect 3850 810 3860 840
rect 3890 810 3900 840
rect 3850 800 3900 810
rect 4000 840 4050 850
rect 4000 810 4010 840
rect 4040 810 4050 840
rect 4000 800 4050 810
rect 4300 840 4350 850
rect 4300 810 4310 840
rect 4340 810 4350 840
rect 4300 800 4350 810
rect 4450 840 4500 850
rect 4450 810 4460 840
rect 4490 810 4500 840
rect 4450 800 4500 810
rect 4600 840 4650 850
rect 4600 810 4610 840
rect 4640 810 4650 840
rect 4600 800 4650 810
rect 4900 840 4950 850
rect 4900 810 4910 840
rect 4940 810 4950 840
rect 4900 800 4950 810
rect 5200 840 5250 850
rect 5200 810 5210 840
rect 5240 810 5250 840
rect 5200 800 5250 810
rect 5500 840 5550 850
rect 5500 810 5510 840
rect 5540 810 5550 840
rect 5500 800 5550 810
rect 5800 840 5850 850
rect 5800 810 5810 840
rect 5840 810 5850 840
rect 5800 800 5850 810
rect 5950 840 6000 850
rect 5950 810 5960 840
rect 5990 810 6000 840
rect 5950 800 6000 810
rect 6100 840 6150 850
rect 6100 810 6110 840
rect 6140 810 6150 840
rect 6100 800 6150 810
rect 6400 840 6450 850
rect 6400 810 6410 840
rect 6440 810 6450 840
rect 6400 800 6450 810
rect 6700 840 6750 850
rect 6700 810 6710 840
rect 6740 810 6750 840
rect 6700 800 6750 810
rect 7000 840 7050 850
rect 7000 810 7010 840
rect 7040 810 7050 840
rect 7000 800 7050 810
rect 7300 840 7350 850
rect 7300 810 7310 840
rect 7340 810 7350 840
rect 7300 800 7350 810
rect 7600 840 7650 850
rect 7600 810 7610 840
rect 7640 810 7650 840
rect 7600 800 7650 810
rect 7900 840 7950 850
rect 7900 810 7910 840
rect 7940 810 7950 840
rect 7900 800 7950 810
rect 8200 840 8250 850
rect 8200 810 8210 840
rect 8240 810 8250 840
rect 8200 800 8250 810
rect 8500 840 8550 850
rect 8500 810 8510 840
rect 8540 810 8550 840
rect 8500 800 8550 810
rect 8800 840 8850 850
rect 8800 810 8810 840
rect 8840 810 8850 840
rect 8800 800 8850 810
rect 9100 840 9150 850
rect 9100 810 9110 840
rect 9140 810 9150 840
rect 9100 800 9150 810
rect 9400 840 9450 850
rect 9400 810 9410 840
rect 9440 810 9450 840
rect 9400 800 9450 810
rect 9550 840 9600 850
rect 9550 810 9560 840
rect 9590 810 9600 840
rect 9550 800 9600 810
rect 9700 840 9750 850
rect 9700 810 9710 840
rect 9740 810 9750 840
rect 9700 800 9750 810
rect 10000 840 10050 850
rect 10000 810 10010 840
rect 10040 810 10050 840
rect 10000 800 10050 810
rect 10300 840 10350 850
rect 10300 810 10310 840
rect 10340 810 10350 840
rect 10300 800 10350 810
rect 10600 840 10650 850
rect 10600 810 10610 840
rect 10640 810 10650 840
rect 10600 800 10650 810
rect 10900 840 10950 850
rect 10900 810 10910 840
rect 10940 810 10950 840
rect 10900 800 10950 810
rect 11200 840 11250 850
rect 11200 810 11210 840
rect 11240 810 11250 840
rect 11200 800 11250 810
rect 11500 840 11550 850
rect 11500 810 11510 840
rect 11540 810 11550 840
rect 11500 800 11550 810
rect 11800 840 11850 850
rect 11800 810 11810 840
rect 11840 810 11850 840
rect 11800 800 11850 810
rect 12100 840 12150 850
rect 12100 810 12110 840
rect 12140 810 12150 840
rect 12100 800 12150 810
rect 12400 840 12450 850
rect 12400 810 12410 840
rect 12440 810 12450 840
rect 12400 800 12450 810
rect 12550 840 12600 850
rect 12550 810 12560 840
rect 12590 810 12600 840
rect 12550 800 12600 810
rect 12700 840 12750 850
rect 12700 810 12710 840
rect 12740 810 12750 840
rect 12700 800 12750 810
rect 13000 840 13050 850
rect 13000 810 13010 840
rect 13040 810 13050 840
rect 13000 800 13050 810
rect 13150 840 13200 850
rect 13150 810 13160 840
rect 13190 810 13200 840
rect 13150 800 13200 810
rect 13300 840 13350 850
rect 13300 810 13310 840
rect 13340 810 13350 840
rect 13300 800 13350 810
rect 13600 840 13650 850
rect 13600 810 13610 840
rect 13640 810 13650 840
rect 13600 800 13650 810
rect 13750 840 13800 850
rect 13750 810 13760 840
rect 13790 810 13800 840
rect 13750 800 13800 810
rect 13900 840 13950 850
rect 13900 810 13910 840
rect 13940 810 13950 840
rect 13900 800 13950 810
rect 14200 840 14250 850
rect 14200 810 14210 840
rect 14240 810 14250 840
rect 14200 800 14250 810
rect 14500 840 14550 850
rect 14500 810 14510 840
rect 14540 810 14550 840
rect 14500 800 14550 810
rect 14800 840 14850 850
rect 14800 810 14810 840
rect 14840 810 14850 840
rect 14800 800 14850 810
rect 15100 840 15150 850
rect 15100 810 15110 840
rect 15140 810 15150 840
rect 15100 800 15150 810
rect 15400 840 15450 850
rect 15400 810 15410 840
rect 15440 810 15450 840
rect 15400 800 15450 810
rect 15700 840 15750 850
rect 15700 810 15710 840
rect 15740 810 15750 840
rect 15700 800 15750 810
rect 16000 840 16050 850
rect 16000 810 16010 840
rect 16040 810 16050 840
rect 16000 800 16050 810
rect 16300 840 16350 850
rect 16300 810 16310 840
rect 16340 810 16350 840
rect 16300 800 16350 810
rect 16600 840 16650 850
rect 16600 810 16610 840
rect 16640 810 16650 840
rect 16600 800 16650 810
rect 16750 840 16800 850
rect 16750 810 16760 840
rect 16790 810 16800 840
rect 16750 800 16800 810
rect 16900 840 16950 850
rect 16900 810 16910 840
rect 16940 810 16950 840
rect 16900 800 16950 810
rect 17200 840 17250 850
rect 17200 810 17210 840
rect 17240 810 17250 840
rect 17200 800 17250 810
rect 17500 840 17550 850
rect 17500 810 17510 840
rect 17540 810 17550 840
rect 17500 800 17550 810
rect 17800 840 17850 850
rect 17800 810 17810 840
rect 17840 810 17850 840
rect 17800 800 17850 810
rect 18100 840 18150 850
rect 18100 810 18110 840
rect 18140 810 18150 840
rect 18100 800 18150 810
rect 18400 840 18450 850
rect 18400 810 18410 840
rect 18440 810 18450 840
rect 18400 800 18450 810
rect 18700 840 18750 850
rect 18700 810 18710 840
rect 18740 810 18750 840
rect 18700 800 18750 810
rect 19000 840 19050 850
rect 19000 810 19010 840
rect 19040 810 19050 840
rect 19000 800 19050 810
rect 19150 840 19200 850
rect 19150 810 19160 840
rect 19190 810 19200 840
rect 19150 800 19200 810
rect 19300 840 19350 850
rect 19300 810 19310 840
rect 19340 810 19350 840
rect 19300 800 19350 810
rect 19600 840 19650 850
rect 19600 810 19610 840
rect 19640 810 19650 840
rect 19600 800 19650 810
rect 19900 840 19950 850
rect 19900 810 19910 840
rect 19940 810 19950 840
rect 19900 800 19950 810
rect 20200 840 20250 850
rect 20200 810 20210 840
rect 20240 810 20250 840
rect 20200 800 20250 810
rect 20500 840 20550 850
rect 20500 810 20510 840
rect 20540 810 20550 840
rect 20500 800 20550 810
rect 20800 840 20850 850
rect 20800 810 20810 840
rect 20840 810 20850 840
rect 20800 800 20850 810
rect 21100 840 21150 850
rect 21100 810 21110 840
rect 21140 810 21150 840
rect 21100 800 21150 810
rect 21400 840 21450 850
rect 21400 810 21410 840
rect 21440 810 21450 840
rect 21400 800 21450 810
rect 21700 840 21750 850
rect 21700 810 21710 840
rect 21740 810 21750 840
rect 21700 800 21750 810
rect 22000 840 22050 850
rect 22000 810 22010 840
rect 22040 810 22050 840
rect 22000 800 22050 810
rect 22300 840 22350 850
rect 22300 810 22310 840
rect 22340 810 22350 840
rect 22300 800 22350 810
rect 22450 840 22500 850
rect 22450 810 22460 840
rect 22490 810 22500 840
rect 22450 800 22500 810
rect 22600 840 22650 850
rect 22600 810 22610 840
rect 22640 810 22650 840
rect 22600 800 22650 810
rect 22900 840 22950 850
rect 22900 810 22910 840
rect 22940 810 22950 840
rect 22900 800 22950 810
rect 23200 840 23250 850
rect 23200 810 23210 840
rect 23240 810 23250 840
rect 23200 800 23250 810
rect 23500 840 23550 850
rect 23500 810 23510 840
rect 23540 810 23550 840
rect 23500 800 23550 810
rect 23800 840 23850 850
rect 23800 810 23810 840
rect 23840 810 23850 840
rect 23800 800 23850 810
rect 24100 840 24150 850
rect 24100 810 24110 840
rect 24140 810 24150 840
rect 24100 800 24150 810
rect 24400 840 24450 850
rect 24400 810 24410 840
rect 24440 810 24450 840
rect 24400 800 24450 810
rect 24700 840 24750 850
rect 24700 810 24710 840
rect 24740 810 24750 840
rect 24700 800 24750 810
rect 25000 840 25050 850
rect 25000 810 25010 840
rect 25040 810 25050 840
rect 25000 800 25050 810
rect 25300 840 25350 850
rect 25300 810 25310 840
rect 25340 810 25350 840
rect 25300 800 25350 810
rect 25600 840 25650 850
rect 25600 810 25610 840
rect 25640 810 25650 840
rect 25600 800 25650 810
rect 25750 840 25800 850
rect 25750 810 25760 840
rect 25790 810 25800 840
rect 25750 800 25800 810
rect 25900 840 25950 850
rect 25900 810 25910 840
rect 25940 810 25950 840
rect 25900 800 25950 810
rect 26200 840 26250 850
rect 26200 810 26210 840
rect 26240 810 26250 840
rect 26200 800 26250 810
rect 26500 840 26550 850
rect 26500 810 26510 840
rect 26540 810 26550 840
rect 26500 800 26550 810
rect 26650 840 26700 850
rect 26650 810 26660 840
rect 26690 810 26700 840
rect 26650 800 26700 810
rect 26800 840 26850 850
rect 26800 810 26810 840
rect 26840 810 26850 840
rect 26800 800 26850 810
rect 27100 840 27150 850
rect 27100 810 27110 840
rect 27140 810 27150 840
rect 27100 800 27150 810
rect 27400 840 27450 850
rect 27400 810 27410 840
rect 27440 810 27450 840
rect 27400 800 27450 810
rect 27550 840 27600 850
rect 27550 810 27560 840
rect 27590 810 27600 840
rect 27550 800 27600 810
rect 27700 840 27750 850
rect 27700 810 27710 840
rect 27740 810 27750 840
rect 27700 800 27750 810
rect 28000 840 28050 850
rect 28000 810 28010 840
rect 28040 810 28050 840
rect 28000 800 28050 810
rect 28300 840 28350 850
rect 28300 810 28310 840
rect 28340 810 28350 840
rect 28300 800 28350 810
rect 28600 840 28650 850
rect 28600 810 28610 840
rect 28640 810 28650 840
rect 28600 800 28650 810
rect -900 740 28800 750
rect -900 710 -640 740
rect -610 710 -40 740
rect -10 710 8360 740
rect 8390 710 10760 740
rect 10790 710 15560 740
rect 15590 710 17960 740
rect 17990 710 20360 740
rect 20390 710 24560 740
rect 24590 710 28760 740
rect 28790 710 28800 740
rect -900 700 28800 710
rect -900 640 28800 650
rect -900 610 -640 640
rect -610 610 -40 640
rect -10 610 8360 640
rect 8390 610 10760 640
rect 10790 610 15560 640
rect 15590 610 17960 640
rect 17990 610 20360 640
rect 20390 610 24560 640
rect 24590 610 28760 640
rect 28790 610 28800 640
rect -900 600 28800 610
rect -900 540 28800 550
rect -900 510 -640 540
rect -610 510 -40 540
rect -10 510 8360 540
rect 8390 510 10760 540
rect 10790 510 15560 540
rect 15590 510 17960 540
rect 17990 510 20360 540
rect 20390 510 24560 540
rect 24590 510 28760 540
rect 28790 510 28800 540
rect -900 500 28800 510
rect -900 440 28800 450
rect -900 410 -640 440
rect -610 410 -40 440
rect -10 410 8360 440
rect 8390 410 10760 440
rect 10790 410 15560 440
rect 15590 410 17960 440
rect 17990 410 20360 440
rect 20390 410 24560 440
rect 24590 410 28760 440
rect 28790 410 28800 440
rect -900 400 28800 410
rect -900 340 28800 350
rect -900 310 -640 340
rect -610 310 -40 340
rect -10 310 8360 340
rect 8390 310 10760 340
rect 10790 310 15560 340
rect 15590 310 17960 340
rect 17990 310 20360 340
rect 20390 310 24560 340
rect 24590 310 28760 340
rect 28790 310 28800 340
rect -900 300 28800 310
rect -900 240 28800 250
rect -900 210 -640 240
rect -610 210 -40 240
rect -10 210 8360 240
rect 8390 210 10760 240
rect 10790 210 15560 240
rect 15590 210 17960 240
rect 17990 210 20360 240
rect 20390 210 24560 240
rect 24590 210 28760 240
rect 28790 210 28800 240
rect -900 200 28800 210
rect -900 140 28800 150
rect -900 110 -640 140
rect -610 110 -40 140
rect -10 110 8360 140
rect 8390 110 10760 140
rect 10790 110 15560 140
rect 15590 110 17960 140
rect 17990 110 20360 140
rect 20390 110 24560 140
rect 24590 110 28760 140
rect 28790 110 28800 140
rect -900 100 28800 110
rect -900 40 28800 50
rect -900 10 -640 40
rect -610 10 -40 40
rect -10 10 8360 40
rect 8390 10 10760 40
rect 10790 10 15560 40
rect 15590 10 17960 40
rect 17990 10 20360 40
rect 20390 10 24560 40
rect 24590 10 28760 40
rect 28790 10 28800 40
rect -900 -10 28800 10
rect -900 -40 -640 -10
rect -610 -40 -40 -10
rect -10 -40 8360 -10
rect 8390 -40 10760 -10
rect 10790 -40 15560 -10
rect 15590 -40 17960 -10
rect 17990 -40 20360 -10
rect 20390 -40 24560 -10
rect 24590 -40 28760 -10
rect 28790 -40 28800 -10
rect -900 -60 28800 -40
rect -900 -90 -640 -60
rect -610 -90 -40 -60
rect -10 -90 8360 -60
rect 8390 -90 10760 -60
rect 10790 -90 15560 -60
rect 15590 -90 17960 -60
rect 17990 -90 20360 -60
rect 20390 -90 24560 -60
rect 24590 -90 28760 -60
rect 28790 -90 28800 -60
rect -900 -100 28800 -90
rect -900 -160 28800 -150
rect -900 -190 -640 -160
rect -610 -190 -40 -160
rect -10 -190 8360 -160
rect 8390 -190 10760 -160
rect 10790 -190 15560 -160
rect 15590 -190 17960 -160
rect 17990 -190 20360 -160
rect 20390 -190 24560 -160
rect 24590 -190 28760 -160
rect 28790 -190 28800 -160
rect -900 -200 28800 -190
rect -900 -260 28800 -250
rect -900 -290 -640 -260
rect -610 -290 -40 -260
rect -10 -290 8360 -260
rect 8390 -290 10760 -260
rect 10790 -290 15560 -260
rect 15590 -290 17960 -260
rect 17990 -290 20360 -260
rect 20390 -290 24560 -260
rect 24590 -290 28760 -260
rect 28790 -290 28800 -260
rect -900 -300 28800 -290
rect -900 -360 28800 -350
rect -900 -390 -640 -360
rect -610 -390 -40 -360
rect -10 -390 8360 -360
rect 8390 -390 10760 -360
rect 10790 -390 15560 -360
rect 15590 -390 17960 -360
rect 17990 -390 20360 -360
rect 20390 -390 24560 -360
rect 24590 -390 28760 -360
rect 28790 -390 28800 -360
rect -900 -400 28800 -390
rect -900 -460 28800 -450
rect -900 -490 -640 -460
rect -610 -490 -40 -460
rect -10 -490 8360 -460
rect 8390 -490 10760 -460
rect 10790 -490 15560 -460
rect 15590 -490 17960 -460
rect 17990 -490 20360 -460
rect 20390 -490 24560 -460
rect 24590 -490 28760 -460
rect 28790 -490 28800 -460
rect -900 -500 28800 -490
rect -900 -560 28800 -550
rect -900 -590 -640 -560
rect -610 -590 -40 -560
rect -10 -590 8360 -560
rect 8390 -590 10760 -560
rect 10790 -590 15560 -560
rect 15590 -590 17960 -560
rect 17990 -590 20360 -560
rect 20390 -590 24560 -560
rect 24590 -590 28760 -560
rect 28790 -590 28800 -560
rect -900 -600 28800 -590
rect -900 -660 28800 -650
rect -900 -690 -640 -660
rect -610 -690 -40 -660
rect -10 -690 8360 -660
rect 8390 -690 10760 -660
rect 10790 -690 15560 -660
rect 15590 -690 17960 -660
rect 17990 -690 20360 -660
rect 20390 -690 24560 -660
rect 24590 -690 28760 -660
rect 28790 -690 28800 -660
rect -900 -700 28800 -690
rect -900 -760 28800 -750
rect -900 -790 -640 -760
rect -610 -790 -40 -760
rect -10 -790 8360 -760
rect 8390 -790 10760 -760
rect 10790 -790 15560 -760
rect 15590 -790 17960 -760
rect 17990 -790 20360 -760
rect 20390 -790 24560 -760
rect 24590 -790 28760 -760
rect 28790 -790 28800 -760
rect -900 -800 28800 -790
rect -500 -860 -450 -850
rect -500 -890 -490 -860
rect -460 -890 -450 -860
rect -500 -900 -450 -890
rect -350 -860 -300 -850
rect -350 -890 -340 -860
rect -310 -890 -300 -860
rect -350 -900 -300 -890
rect -200 -860 -150 -850
rect -200 -890 -190 -860
rect -160 -890 -150 -860
rect -200 -900 -150 -890
rect 100 -860 150 -850
rect 100 -890 110 -860
rect 140 -890 150 -860
rect 100 -900 150 -890
rect 400 -860 450 -850
rect 400 -890 410 -860
rect 440 -890 450 -860
rect 400 -900 450 -890
rect 700 -860 750 -850
rect 700 -890 710 -860
rect 740 -890 750 -860
rect 700 -900 750 -890
rect 1000 -860 1050 -850
rect 1000 -890 1010 -860
rect 1040 -890 1050 -860
rect 1000 -900 1050 -890
rect 1300 -860 1350 -850
rect 1300 -890 1310 -860
rect 1340 -890 1350 -860
rect 1300 -900 1350 -890
rect 1600 -860 1650 -850
rect 1600 -890 1610 -860
rect 1640 -890 1650 -860
rect 1600 -900 1650 -890
rect 1900 -860 1950 -850
rect 1900 -890 1910 -860
rect 1940 -890 1950 -860
rect 1900 -900 1950 -890
rect 2200 -860 2250 -850
rect 2200 -890 2210 -860
rect 2240 -890 2250 -860
rect 2200 -900 2250 -890
rect 2350 -860 2400 -850
rect 2350 -890 2360 -860
rect 2390 -890 2400 -860
rect 2350 -900 2400 -890
rect 2500 -860 2550 -850
rect 2500 -890 2510 -860
rect 2540 -890 2550 -860
rect 2500 -900 2550 -890
rect 2800 -860 2850 -850
rect 2800 -890 2810 -860
rect 2840 -890 2850 -860
rect 2800 -900 2850 -890
rect 3100 -860 3150 -850
rect 3100 -890 3110 -860
rect 3140 -890 3150 -860
rect 3100 -900 3150 -890
rect 3400 -860 3450 -850
rect 3400 -890 3410 -860
rect 3440 -890 3450 -860
rect 3400 -900 3450 -890
rect 3700 -860 3750 -850
rect 3700 -890 3710 -860
rect 3740 -890 3750 -860
rect 3700 -900 3750 -890
rect 3850 -860 3900 -850
rect 3850 -890 3860 -860
rect 3890 -890 3900 -860
rect 3850 -900 3900 -890
rect 4000 -860 4050 -850
rect 4000 -890 4010 -860
rect 4040 -890 4050 -860
rect 4000 -900 4050 -890
rect 4300 -860 4350 -850
rect 4300 -890 4310 -860
rect 4340 -890 4350 -860
rect 4300 -900 4350 -890
rect 4450 -860 4500 -850
rect 4450 -890 4460 -860
rect 4490 -890 4500 -860
rect 4450 -900 4500 -890
rect 4600 -860 4650 -850
rect 4600 -890 4610 -860
rect 4640 -890 4650 -860
rect 4600 -900 4650 -890
rect 4900 -860 4950 -850
rect 4900 -890 4910 -860
rect 4940 -890 4950 -860
rect 4900 -900 4950 -890
rect 5200 -860 5250 -850
rect 5200 -890 5210 -860
rect 5240 -890 5250 -860
rect 5200 -900 5250 -890
rect 5500 -860 5550 -850
rect 5500 -890 5510 -860
rect 5540 -890 5550 -860
rect 5500 -900 5550 -890
rect 5800 -860 5850 -850
rect 5800 -890 5810 -860
rect 5840 -890 5850 -860
rect 5800 -900 5850 -890
rect 5950 -860 6000 -850
rect 5950 -890 5960 -860
rect 5990 -890 6000 -860
rect 5950 -900 6000 -890
rect 6100 -860 6150 -850
rect 6100 -890 6110 -860
rect 6140 -890 6150 -860
rect 6100 -900 6150 -890
rect 6400 -860 6450 -850
rect 6400 -890 6410 -860
rect 6440 -890 6450 -860
rect 6400 -900 6450 -890
rect 6700 -860 6750 -850
rect 6700 -890 6710 -860
rect 6740 -890 6750 -860
rect 6700 -900 6750 -890
rect 7000 -860 7050 -850
rect 7000 -890 7010 -860
rect 7040 -890 7050 -860
rect 7000 -900 7050 -890
rect 7300 -860 7350 -850
rect 7300 -890 7310 -860
rect 7340 -890 7350 -860
rect 7300 -900 7350 -890
rect 7600 -860 7650 -850
rect 7600 -890 7610 -860
rect 7640 -890 7650 -860
rect 7600 -900 7650 -890
rect 7900 -860 7950 -850
rect 7900 -890 7910 -860
rect 7940 -890 7950 -860
rect 7900 -900 7950 -890
rect 8200 -860 8250 -850
rect 8200 -890 8210 -860
rect 8240 -890 8250 -860
rect 8200 -900 8250 -890
rect 8500 -860 8550 -850
rect 8500 -890 8510 -860
rect 8540 -890 8550 -860
rect 8500 -900 8550 -890
rect 8800 -860 8850 -850
rect 8800 -890 8810 -860
rect 8840 -890 8850 -860
rect 8800 -900 8850 -890
rect 9100 -860 9150 -850
rect 9100 -890 9110 -860
rect 9140 -890 9150 -860
rect 9100 -900 9150 -890
rect 9400 -860 9450 -850
rect 9400 -890 9410 -860
rect 9440 -890 9450 -860
rect 9400 -900 9450 -890
rect 9550 -860 9600 -850
rect 9550 -890 9560 -860
rect 9590 -890 9600 -860
rect 9550 -900 9600 -890
rect 9700 -860 9750 -850
rect 9700 -890 9710 -860
rect 9740 -890 9750 -860
rect 9700 -900 9750 -890
rect 10000 -860 10050 -850
rect 10000 -890 10010 -860
rect 10040 -890 10050 -860
rect 10000 -900 10050 -890
rect 10300 -860 10350 -850
rect 10300 -890 10310 -860
rect 10340 -890 10350 -860
rect 10300 -900 10350 -890
rect 10600 -860 10650 -850
rect 10600 -890 10610 -860
rect 10640 -890 10650 -860
rect 10600 -900 10650 -890
rect 10900 -860 10950 -850
rect 10900 -890 10910 -860
rect 10940 -890 10950 -860
rect 10900 -900 10950 -890
rect 11200 -860 11250 -850
rect 11200 -890 11210 -860
rect 11240 -890 11250 -860
rect 11200 -900 11250 -890
rect 11500 -860 11550 -850
rect 11500 -890 11510 -860
rect 11540 -890 11550 -860
rect 11500 -900 11550 -890
rect 11800 -860 11850 -850
rect 11800 -890 11810 -860
rect 11840 -890 11850 -860
rect 11800 -900 11850 -890
rect 12100 -860 12150 -850
rect 12100 -890 12110 -860
rect 12140 -890 12150 -860
rect 12100 -900 12150 -890
rect 12400 -860 12450 -850
rect 12400 -890 12410 -860
rect 12440 -890 12450 -860
rect 12400 -900 12450 -890
rect 12550 -860 12600 -850
rect 12550 -890 12560 -860
rect 12590 -890 12600 -860
rect 12550 -900 12600 -890
rect 12700 -860 12750 -850
rect 12700 -890 12710 -860
rect 12740 -890 12750 -860
rect 12700 -900 12750 -890
rect 13000 -860 13050 -850
rect 13000 -890 13010 -860
rect 13040 -890 13050 -860
rect 13000 -900 13050 -890
rect 13150 -860 13200 -850
rect 13150 -890 13160 -860
rect 13190 -890 13200 -860
rect 13150 -900 13200 -890
rect 13300 -860 13350 -850
rect 13300 -890 13310 -860
rect 13340 -890 13350 -860
rect 13300 -900 13350 -890
rect 13600 -860 13650 -850
rect 13600 -890 13610 -860
rect 13640 -890 13650 -860
rect 13600 -900 13650 -890
rect 13750 -860 13800 -850
rect 13750 -890 13760 -860
rect 13790 -890 13800 -860
rect 13750 -900 13800 -890
rect 13900 -860 13950 -850
rect 13900 -890 13910 -860
rect 13940 -890 13950 -860
rect 13900 -900 13950 -890
rect 14200 -860 14250 -850
rect 14200 -890 14210 -860
rect 14240 -890 14250 -860
rect 14200 -900 14250 -890
rect 14500 -860 14550 -850
rect 14500 -890 14510 -860
rect 14540 -890 14550 -860
rect 14500 -900 14550 -890
rect 14800 -860 14850 -850
rect 14800 -890 14810 -860
rect 14840 -890 14850 -860
rect 14800 -900 14850 -890
rect 15100 -860 15150 -850
rect 15100 -890 15110 -860
rect 15140 -890 15150 -860
rect 15100 -900 15150 -890
rect 15400 -860 15450 -850
rect 15400 -890 15410 -860
rect 15440 -890 15450 -860
rect 15400 -900 15450 -890
rect 15700 -860 15750 -850
rect 15700 -890 15710 -860
rect 15740 -890 15750 -860
rect 15700 -900 15750 -890
rect 16000 -860 16050 -850
rect 16000 -890 16010 -860
rect 16040 -890 16050 -860
rect 16000 -900 16050 -890
rect 16300 -860 16350 -850
rect 16300 -890 16310 -860
rect 16340 -890 16350 -860
rect 16300 -900 16350 -890
rect 16600 -860 16650 -850
rect 16600 -890 16610 -860
rect 16640 -890 16650 -860
rect 16600 -900 16650 -890
rect 16750 -860 16800 -850
rect 16750 -890 16760 -860
rect 16790 -890 16800 -860
rect 16750 -900 16800 -890
rect 16900 -860 16950 -850
rect 16900 -890 16910 -860
rect 16940 -890 16950 -860
rect 16900 -900 16950 -890
rect 17200 -860 17250 -850
rect 17200 -890 17210 -860
rect 17240 -890 17250 -860
rect 17200 -900 17250 -890
rect 17500 -860 17550 -850
rect 17500 -890 17510 -860
rect 17540 -890 17550 -860
rect 17500 -900 17550 -890
rect 17800 -860 17850 -850
rect 17800 -890 17810 -860
rect 17840 -890 17850 -860
rect 17800 -900 17850 -890
rect 18100 -860 18150 -850
rect 18100 -890 18110 -860
rect 18140 -890 18150 -860
rect 18100 -900 18150 -890
rect 18400 -860 18450 -850
rect 18400 -890 18410 -860
rect 18440 -890 18450 -860
rect 18400 -900 18450 -890
rect 18700 -860 18750 -850
rect 18700 -890 18710 -860
rect 18740 -890 18750 -860
rect 18700 -900 18750 -890
rect 19000 -860 19050 -850
rect 19000 -890 19010 -860
rect 19040 -890 19050 -860
rect 19000 -900 19050 -890
rect 19150 -860 19200 -850
rect 19150 -890 19160 -860
rect 19190 -890 19200 -860
rect 19150 -900 19200 -890
rect 19300 -860 19350 -850
rect 19300 -890 19310 -860
rect 19340 -890 19350 -860
rect 19300 -900 19350 -890
rect 19600 -860 19650 -850
rect 19600 -890 19610 -860
rect 19640 -890 19650 -860
rect 19600 -900 19650 -890
rect 19900 -860 19950 -850
rect 19900 -890 19910 -860
rect 19940 -890 19950 -860
rect 19900 -900 19950 -890
rect 20200 -860 20250 -850
rect 20200 -890 20210 -860
rect 20240 -890 20250 -860
rect 20200 -900 20250 -890
rect 20500 -860 20550 -850
rect 20500 -890 20510 -860
rect 20540 -890 20550 -860
rect 20500 -900 20550 -890
rect 20800 -860 20850 -850
rect 20800 -890 20810 -860
rect 20840 -890 20850 -860
rect 20800 -900 20850 -890
rect 21100 -860 21150 -850
rect 21100 -890 21110 -860
rect 21140 -890 21150 -860
rect 21100 -900 21150 -890
rect 21400 -860 21450 -850
rect 21400 -890 21410 -860
rect 21440 -890 21450 -860
rect 21400 -900 21450 -890
rect 21700 -860 21750 -850
rect 21700 -890 21710 -860
rect 21740 -890 21750 -860
rect 21700 -900 21750 -890
rect 22000 -860 22050 -850
rect 22000 -890 22010 -860
rect 22040 -890 22050 -860
rect 22000 -900 22050 -890
rect 22300 -860 22350 -850
rect 22300 -890 22310 -860
rect 22340 -890 22350 -860
rect 22300 -900 22350 -890
rect 22450 -860 22500 -850
rect 22450 -890 22460 -860
rect 22490 -890 22500 -860
rect 22450 -900 22500 -890
rect 22600 -860 22650 -850
rect 22600 -890 22610 -860
rect 22640 -890 22650 -860
rect 22600 -900 22650 -890
rect 22900 -860 22950 -850
rect 22900 -890 22910 -860
rect 22940 -890 22950 -860
rect 22900 -900 22950 -890
rect 23200 -860 23250 -850
rect 23200 -890 23210 -860
rect 23240 -890 23250 -860
rect 23200 -900 23250 -890
rect 23500 -860 23550 -850
rect 23500 -890 23510 -860
rect 23540 -890 23550 -860
rect 23500 -900 23550 -890
rect 23800 -860 23850 -850
rect 23800 -890 23810 -860
rect 23840 -890 23850 -860
rect 23800 -900 23850 -890
rect 24100 -860 24150 -850
rect 24100 -890 24110 -860
rect 24140 -890 24150 -860
rect 24100 -900 24150 -890
rect 24400 -860 24450 -850
rect 24400 -890 24410 -860
rect 24440 -890 24450 -860
rect 24400 -900 24450 -890
rect 24700 -860 24750 -850
rect 24700 -890 24710 -860
rect 24740 -890 24750 -860
rect 24700 -900 24750 -890
rect 25000 -860 25050 -850
rect 25000 -890 25010 -860
rect 25040 -890 25050 -860
rect 25000 -900 25050 -890
rect 25300 -860 25350 -850
rect 25300 -890 25310 -860
rect 25340 -890 25350 -860
rect 25300 -900 25350 -890
rect 25600 -860 25650 -850
rect 25600 -890 25610 -860
rect 25640 -890 25650 -860
rect 25600 -900 25650 -890
rect 25750 -860 25800 -850
rect 25750 -890 25760 -860
rect 25790 -890 25800 -860
rect 25750 -900 25800 -890
rect 25900 -860 25950 -850
rect 25900 -890 25910 -860
rect 25940 -890 25950 -860
rect 25900 -900 25950 -890
rect 26200 -860 26250 -850
rect 26200 -890 26210 -860
rect 26240 -890 26250 -860
rect 26200 -900 26250 -890
rect 26500 -860 26550 -850
rect 26500 -890 26510 -860
rect 26540 -890 26550 -860
rect 26500 -900 26550 -890
rect 26650 -860 26700 -850
rect 26650 -890 26660 -860
rect 26690 -890 26700 -860
rect 26650 -900 26700 -890
rect 26800 -860 26850 -850
rect 26800 -890 26810 -860
rect 26840 -890 26850 -860
rect 26800 -900 26850 -890
rect 27100 -860 27150 -850
rect 27100 -890 27110 -860
rect 27140 -890 27150 -860
rect 27100 -900 27150 -890
rect 27400 -860 27450 -850
rect 27400 -890 27410 -860
rect 27440 -890 27450 -860
rect 27400 -900 27450 -890
rect 27550 -860 27600 -850
rect 27550 -890 27560 -860
rect 27590 -890 27600 -860
rect 27550 -900 27600 -890
rect 27700 -860 27750 -850
rect 27700 -890 27710 -860
rect 27740 -890 27750 -860
rect 27700 -900 27750 -890
rect 28000 -860 28050 -850
rect 28000 -890 28010 -860
rect 28040 -890 28050 -860
rect 28000 -900 28050 -890
rect 28300 -860 28350 -850
rect 28300 -890 28310 -860
rect 28340 -890 28350 -860
rect 28300 -900 28350 -890
rect 28600 -860 28650 -850
rect 28600 -890 28610 -860
rect 28640 -890 28650 -860
rect 28600 -900 28650 -890
rect -900 -960 28800 -950
rect -900 -990 -640 -960
rect -610 -990 -40 -960
rect -10 -990 8360 -960
rect 8390 -990 10760 -960
rect 10790 -990 15560 -960
rect 15590 -990 17960 -960
rect 17990 -990 20360 -960
rect 20390 -990 24560 -960
rect 24590 -990 28760 -960
rect 28790 -990 28800 -960
rect -900 -1000 28800 -990
rect -900 -1060 28800 -1050
rect -900 -1090 -640 -1060
rect -610 -1090 -40 -1060
rect -10 -1090 8360 -1060
rect 8390 -1090 10760 -1060
rect 10790 -1090 15560 -1060
rect 15590 -1090 17960 -1060
rect 17990 -1090 20360 -1060
rect 20390 -1090 24560 -1060
rect 24590 -1090 28760 -1060
rect 28790 -1090 28800 -1060
rect -900 -1100 28800 -1090
rect -900 -1160 28800 -1150
rect -900 -1190 -640 -1160
rect -610 -1190 -40 -1160
rect -10 -1190 8360 -1160
rect 8390 -1190 10760 -1160
rect 10790 -1190 15560 -1160
rect 15590 -1190 17960 -1160
rect 17990 -1190 20360 -1160
rect 20390 -1190 24560 -1160
rect 24590 -1190 28760 -1160
rect 28790 -1190 28800 -1160
rect -900 -1200 28800 -1190
rect -900 -1260 28800 -1250
rect -900 -1290 -640 -1260
rect -610 -1290 -40 -1260
rect -10 -1290 8360 -1260
rect 8390 -1290 10760 -1260
rect 10790 -1290 15560 -1260
rect 15590 -1290 17960 -1260
rect 17990 -1290 20360 -1260
rect 20390 -1290 24560 -1260
rect 24590 -1290 28760 -1260
rect 28790 -1290 28800 -1260
rect -900 -1300 28800 -1290
rect -900 -1360 28800 -1350
rect -900 -1390 -640 -1360
rect -610 -1390 -40 -1360
rect -10 -1390 8360 -1360
rect 8390 -1390 10760 -1360
rect 10790 -1390 15560 -1360
rect 15590 -1390 17960 -1360
rect 17990 -1390 20360 -1360
rect 20390 -1390 24560 -1360
rect 24590 -1390 28760 -1360
rect 28790 -1390 28800 -1360
rect -900 -1400 28800 -1390
rect -900 -1460 28800 -1450
rect -900 -1490 -640 -1460
rect -610 -1490 -40 -1460
rect -10 -1490 8360 -1460
rect 8390 -1490 10760 -1460
rect 10790 -1490 15560 -1460
rect 15590 -1490 17960 -1460
rect 17990 -1490 20360 -1460
rect 20390 -1490 24560 -1460
rect 24590 -1490 28760 -1460
rect 28790 -1490 28800 -1460
rect -900 -1500 28800 -1490
rect -900 -1560 28800 -1550
rect -900 -1590 -640 -1560
rect -610 -1590 -40 -1560
rect -10 -1590 8360 -1560
rect 8390 -1590 10760 -1560
rect 10790 -1590 15560 -1560
rect 15590 -1590 17960 -1560
rect 17990 -1590 20360 -1560
rect 20390 -1590 24560 -1560
rect 24590 -1590 28760 -1560
rect 28790 -1590 28800 -1560
rect -900 -1600 28800 -1590
rect -900 -1660 28800 -1650
rect -900 -1690 -640 -1660
rect -610 -1690 -40 -1660
rect -10 -1690 8360 -1660
rect 8390 -1690 10760 -1660
rect 10790 -1690 15560 -1660
rect 15590 -1690 17960 -1660
rect 17990 -1690 20360 -1660
rect 20390 -1690 24560 -1660
rect 24590 -1690 28760 -1660
rect 28790 -1690 28800 -1660
rect -900 -1710 28800 -1690
rect -900 -1740 -640 -1710
rect -610 -1740 -40 -1710
rect -10 -1740 8360 -1710
rect 8390 -1740 10760 -1710
rect 10790 -1740 15560 -1710
rect 15590 -1740 17960 -1710
rect 17990 -1740 20360 -1710
rect 20390 -1740 24560 -1710
rect 24590 -1740 28760 -1710
rect 28790 -1740 28800 -1710
rect -900 -1750 28800 -1740
<< via2 >>
rect -640 5560 -610 5590
rect 8360 5560 8390 5590
rect 8660 5560 8690 5590
rect 8960 5560 8990 5590
rect 9260 5560 9290 5590
rect 9560 5560 9590 5590
rect 9860 5560 9890 5590
rect 10160 5560 10190 5590
rect 10460 5560 10490 5590
rect 10760 5560 10790 5590
rect 11960 5560 11990 5590
rect 13160 5560 13190 5590
rect 14360 5560 14390 5590
rect 15560 5560 15590 5590
rect 20360 5560 20390 5590
rect 22460 5560 22490 5590
rect 24560 5560 24590 5590
rect 26660 5560 26690 5590
rect 28160 5560 28190 5590
rect 28760 5560 28790 5590
rect 32060 5560 32090 5590
rect -490 4910 -460 4940
rect -340 4910 -310 4940
rect -190 4910 -160 4940
rect 110 4910 140 4940
rect 410 4910 440 4940
rect 710 4910 740 4940
rect 1010 4910 1040 4940
rect 1160 4910 1190 4940
rect 1310 4910 1340 4940
rect 1610 4910 1640 4940
rect 1910 4910 1940 4940
rect 2060 4910 2090 4940
rect 2210 4910 2240 4940
rect 2510 4910 2540 4940
rect 2810 4910 2840 4940
rect 2960 4910 2990 4940
rect 3110 4910 3140 4940
rect 3410 4910 3440 4940
rect 3710 4910 3740 4940
rect 4010 4910 4040 4940
rect 4310 4910 4340 4940
rect 4610 4910 4640 4940
rect 4910 4910 4940 4940
rect 5210 4910 5240 4940
rect 5360 4910 5390 4940
rect 5510 4910 5540 4940
rect 5810 4910 5840 4940
rect 6110 4910 6140 4940
rect 6260 4910 6290 4940
rect 6410 4910 6440 4940
rect 6710 4910 6740 4940
rect 7010 4910 7040 4940
rect 7160 4910 7190 4940
rect 7310 4910 7340 4940
rect 7610 4910 7640 4940
rect 7910 4910 7940 4940
rect 8210 4910 8240 4940
rect 8510 4910 8540 4940
rect 8810 4910 8840 4940
rect 9110 4910 9140 4940
rect 9410 4910 9440 4940
rect 9710 4910 9740 4940
rect 10010 4910 10040 4940
rect 10310 4910 10340 4940
rect 10610 4910 10640 4940
rect 10910 4910 10940 4940
rect 11210 4910 11240 4940
rect 11360 4910 11390 4940
rect 11510 4910 11540 4940
rect 11810 4910 11840 4940
rect 12110 4910 12140 4940
rect 12410 4910 12440 4940
rect 12560 4910 12590 4940
rect 12710 4910 12740 4940
rect 13010 4910 13040 4940
rect 13310 4910 13340 4940
rect 13610 4910 13640 4940
rect 13760 4910 13790 4940
rect 13910 4910 13940 4940
rect 14210 4910 14240 4940
rect 14510 4910 14540 4940
rect 14810 4910 14840 4940
rect 14960 4910 14990 4940
rect 15110 4910 15140 4940
rect 15410 4910 15440 4940
rect 15710 4910 15740 4940
rect 16010 4910 16040 4940
rect 16310 4910 16340 4940
rect 16610 4910 16640 4940
rect 16760 4910 16790 4940
rect 16910 4910 16940 4940
rect 17210 4910 17240 4940
rect 17510 4910 17540 4940
rect 17810 4910 17840 4940
rect 18110 4910 18140 4940
rect 18410 4910 18440 4940
rect 18710 4910 18740 4940
rect 19010 4910 19040 4940
rect 19160 4910 19190 4940
rect 19310 4910 19340 4940
rect 19610 4910 19640 4940
rect 19910 4910 19940 4940
rect 20210 4910 20240 4940
rect 20510 4910 20540 4940
rect 20810 4910 20840 4940
rect 20960 4910 20990 4940
rect 21110 4910 21140 4940
rect 21410 4910 21440 4940
rect 21710 4910 21740 4940
rect 21860 4910 21890 4940
rect 22010 4910 22040 4940
rect 22310 4910 22340 4940
rect 22610 4910 22640 4940
rect 22910 4910 22940 4940
rect 23060 4910 23090 4940
rect 23210 4910 23240 4940
rect 23360 4910 23390 4940
rect 23510 4910 23540 4940
rect 23660 4910 23690 4940
rect 23810 4910 23840 4940
rect 23960 4910 23990 4940
rect 24110 4910 24140 4940
rect 24410 4910 24440 4940
rect 24710 4910 24740 4940
rect 25010 4910 25040 4940
rect 25460 4910 25490 4940
rect 25610 4910 25640 4940
rect 25760 4910 25790 4940
rect 26210 4910 26240 4940
rect 26510 4910 26540 4940
rect 26810 4910 26840 4940
rect 27110 4910 27140 4940
rect 27560 4910 27590 4940
rect 27710 4910 27740 4940
rect 27860 4910 27890 4940
rect 28310 4910 28340 4940
rect 28610 4910 28640 4940
rect 28760 4910 28790 4940
rect 28910 4910 28940 4940
rect 29210 4910 29240 4940
rect 29360 4910 29390 4940
rect 29660 4910 29690 4940
rect 29810 4910 29840 4940
rect 29960 4910 29990 4940
rect 30260 4910 30290 4940
rect 30410 4910 30440 4940
rect 30560 4910 30590 4940
rect 30860 4910 30890 4940
rect 31010 4910 31040 4940
rect 31160 4910 31190 4940
rect 31460 4910 31490 4940
rect 31610 4910 31640 4940
rect 31910 4910 31940 4940
rect 32060 4910 32090 4940
rect -640 4260 -610 4290
rect -40 4260 -10 4290
rect 4160 4260 4190 4290
rect 8360 4260 8390 4290
rect 8660 4260 8690 4290
rect 8960 4260 8990 4290
rect 9260 4260 9290 4290
rect 9560 4260 9590 4290
rect 9860 4260 9890 4290
rect 10160 4260 10190 4290
rect 10460 4260 10490 4290
rect 10760 4260 10790 4290
rect 11960 4260 11990 4290
rect 13160 4260 13190 4290
rect 14360 4260 14390 4290
rect 15560 4260 15590 4290
rect 20360 4260 20390 4290
rect 22460 4260 22490 4290
rect 24560 4260 24590 4290
rect 26660 4260 26690 4290
rect 28160 4260 28190 4290
rect 28760 4260 28790 4290
rect 32060 4260 32090 4290
rect -490 3610 -460 3640
rect -340 3610 -310 3640
rect -190 3610 -160 3640
rect 110 3610 140 3640
rect 410 3610 440 3640
rect 710 3610 740 3640
rect 1010 3610 1040 3640
rect 1160 3610 1190 3640
rect 1310 3610 1340 3640
rect 1610 3610 1640 3640
rect 1910 3610 1940 3640
rect 2060 3610 2090 3640
rect 2210 3610 2240 3640
rect 2510 3610 2540 3640
rect 2810 3610 2840 3640
rect 2960 3610 2990 3640
rect 3110 3610 3140 3640
rect 3410 3610 3440 3640
rect 3710 3610 3740 3640
rect 4010 3610 4040 3640
rect 4310 3610 4340 3640
rect 4610 3610 4640 3640
rect 4910 3610 4940 3640
rect 5210 3610 5240 3640
rect 5360 3610 5390 3640
rect 5510 3610 5540 3640
rect 5810 3610 5840 3640
rect 6110 3610 6140 3640
rect 6260 3610 6290 3640
rect 6410 3610 6440 3640
rect 6710 3610 6740 3640
rect 7010 3610 7040 3640
rect 7160 3610 7190 3640
rect 7310 3610 7340 3640
rect 7610 3610 7640 3640
rect 7910 3610 7940 3640
rect 8210 3610 8240 3640
rect 8510 3610 8540 3640
rect 8810 3610 8840 3640
rect 9110 3610 9140 3640
rect 9410 3610 9440 3640
rect 9710 3610 9740 3640
rect 10010 3610 10040 3640
rect 10310 3610 10340 3640
rect 10610 3610 10640 3640
rect 10910 3610 10940 3640
rect 11210 3610 11240 3640
rect 11360 3610 11390 3640
rect 11510 3610 11540 3640
rect 11810 3610 11840 3640
rect 12110 3610 12140 3640
rect 12410 3610 12440 3640
rect 12560 3610 12590 3640
rect 12710 3610 12740 3640
rect 13010 3610 13040 3640
rect 13310 3610 13340 3640
rect 13610 3610 13640 3640
rect 13760 3610 13790 3640
rect 13910 3610 13940 3640
rect 14210 3610 14240 3640
rect 14510 3610 14540 3640
rect 14810 3610 14840 3640
rect 14960 3610 14990 3640
rect 15110 3610 15140 3640
rect 15410 3610 15440 3640
rect 15710 3610 15740 3640
rect 16010 3610 16040 3640
rect 16310 3610 16340 3640
rect 16610 3610 16640 3640
rect 16760 3610 16790 3640
rect 16910 3610 16940 3640
rect 17210 3610 17240 3640
rect 17510 3610 17540 3640
rect 17810 3610 17840 3640
rect 18110 3610 18140 3640
rect 18410 3610 18440 3640
rect 18710 3610 18740 3640
rect 19010 3610 19040 3640
rect 19160 3610 19190 3640
rect 19310 3610 19340 3640
rect 19610 3610 19640 3640
rect 19910 3610 19940 3640
rect 20210 3610 20240 3640
rect 20510 3610 20540 3640
rect 20810 3610 20840 3640
rect 20960 3610 20990 3640
rect 21110 3610 21140 3640
rect 21410 3610 21440 3640
rect 21710 3610 21740 3640
rect 21860 3610 21890 3640
rect 22010 3610 22040 3640
rect 22310 3610 22340 3640
rect 22610 3610 22640 3640
rect 22910 3610 22940 3640
rect 23060 3610 23090 3640
rect 23210 3610 23240 3640
rect 23360 3610 23390 3640
rect 23510 3610 23540 3640
rect 23660 3610 23690 3640
rect 23810 3610 23840 3640
rect 23960 3610 23990 3640
rect 24110 3610 24140 3640
rect 24410 3610 24440 3640
rect 24710 3610 24740 3640
rect 25010 3610 25040 3640
rect 25460 3610 25490 3640
rect 25610 3610 25640 3640
rect 25760 3610 25790 3640
rect 26210 3610 26240 3640
rect 26510 3610 26540 3640
rect 26810 3610 26840 3640
rect 27110 3610 27140 3640
rect 27560 3610 27590 3640
rect 27710 3610 27740 3640
rect 27860 3610 27890 3640
rect 28310 3610 28340 3640
rect 28610 3610 28640 3640
rect 28760 3610 28790 3640
rect 28910 3610 28940 3640
rect 29210 3610 29240 3640
rect 29360 3610 29390 3640
rect 29660 3610 29690 3640
rect 29810 3610 29840 3640
rect 29960 3610 29990 3640
rect 30260 3610 30290 3640
rect 30410 3610 30440 3640
rect 30560 3610 30590 3640
rect 30860 3610 30890 3640
rect 31010 3610 31040 3640
rect 31160 3610 31190 3640
rect 31460 3610 31490 3640
rect 31610 3610 31640 3640
rect 31910 3610 31940 3640
rect 32060 3610 32090 3640
rect -640 2960 -610 2990
rect -40 2960 -10 2990
rect 4160 2960 4190 2990
rect 8360 2960 8390 2990
rect 8660 2960 8690 2990
rect 8960 2960 8990 2990
rect 9260 2960 9290 2990
rect 9560 2960 9590 2990
rect 9860 2960 9890 2990
rect 10160 2960 10190 2990
rect 10460 2960 10490 2990
rect 10760 2960 10790 2990
rect 11960 2960 11990 2990
rect 13160 2960 13190 2990
rect 14360 2960 14390 2990
rect 15560 2960 15590 2990
rect 20360 2960 20390 2990
rect 24560 2960 24590 2990
rect 26660 2960 26690 2990
rect 28160 2960 28190 2990
rect 28760 2960 28790 2990
rect 32060 2960 32090 2990
rect -640 1660 -610 1690
rect -40 1660 -10 1690
rect 8360 1660 8390 1690
rect 10760 1660 10790 1690
rect 15560 1660 15590 1690
rect 17960 1660 17990 1690
rect 20360 1660 20390 1690
rect 24560 1660 24590 1690
rect 28760 1660 28790 1690
rect -640 1610 -610 1640
rect -40 1610 -10 1640
rect 8360 1610 8390 1640
rect 10760 1610 10790 1640
rect 15560 1610 15590 1640
rect 17960 1610 17990 1640
rect 20360 1610 20390 1640
rect 24560 1610 24590 1640
rect 28760 1610 28790 1640
rect -490 810 -460 840
rect -340 810 -310 840
rect -190 810 -160 840
rect 110 810 140 840
rect 410 810 440 840
rect 710 810 740 840
rect 1010 810 1040 840
rect 1310 810 1340 840
rect 1610 810 1640 840
rect 1910 810 1940 840
rect 2210 810 2240 840
rect 2360 810 2390 840
rect 2510 810 2540 840
rect 2810 810 2840 840
rect 3110 810 3140 840
rect 3410 810 3440 840
rect 3710 810 3740 840
rect 3860 810 3890 840
rect 4010 810 4040 840
rect 4310 810 4340 840
rect 4460 810 4490 840
rect 4610 810 4640 840
rect 4910 810 4940 840
rect 5210 810 5240 840
rect 5510 810 5540 840
rect 5810 810 5840 840
rect 5960 810 5990 840
rect 6110 810 6140 840
rect 6410 810 6440 840
rect 6710 810 6740 840
rect 7010 810 7040 840
rect 7310 810 7340 840
rect 7610 810 7640 840
rect 7910 810 7940 840
rect 8210 810 8240 840
rect 8510 810 8540 840
rect 8810 810 8840 840
rect 9110 810 9140 840
rect 9410 810 9440 840
rect 9560 810 9590 840
rect 9710 810 9740 840
rect 10010 810 10040 840
rect 10310 810 10340 840
rect 10610 810 10640 840
rect 10910 810 10940 840
rect 11210 810 11240 840
rect 11510 810 11540 840
rect 11810 810 11840 840
rect 12110 810 12140 840
rect 12410 810 12440 840
rect 12560 810 12590 840
rect 12710 810 12740 840
rect 13010 810 13040 840
rect 13160 810 13190 840
rect 13310 810 13340 840
rect 13610 810 13640 840
rect 13760 810 13790 840
rect 13910 810 13940 840
rect 14210 810 14240 840
rect 14510 810 14540 840
rect 14810 810 14840 840
rect 15110 810 15140 840
rect 15410 810 15440 840
rect 15710 810 15740 840
rect 16010 810 16040 840
rect 16310 810 16340 840
rect 16610 810 16640 840
rect 16760 810 16790 840
rect 16910 810 16940 840
rect 17210 810 17240 840
rect 17510 810 17540 840
rect 17810 810 17840 840
rect 18110 810 18140 840
rect 18410 810 18440 840
rect 18710 810 18740 840
rect 19010 810 19040 840
rect 19160 810 19190 840
rect 19310 810 19340 840
rect 19610 810 19640 840
rect 19910 810 19940 840
rect 20210 810 20240 840
rect 20510 810 20540 840
rect 20810 810 20840 840
rect 21110 810 21140 840
rect 21410 810 21440 840
rect 21710 810 21740 840
rect 22010 810 22040 840
rect 22310 810 22340 840
rect 22460 810 22490 840
rect 22610 810 22640 840
rect 22910 810 22940 840
rect 23210 810 23240 840
rect 23510 810 23540 840
rect 23810 810 23840 840
rect 24110 810 24140 840
rect 24410 810 24440 840
rect 24710 810 24740 840
rect 25010 810 25040 840
rect 25310 810 25340 840
rect 25610 810 25640 840
rect 25760 810 25790 840
rect 25910 810 25940 840
rect 26210 810 26240 840
rect 26510 810 26540 840
rect 26660 810 26690 840
rect 26810 810 26840 840
rect 27110 810 27140 840
rect 27410 810 27440 840
rect 27560 810 27590 840
rect 27710 810 27740 840
rect 28010 810 28040 840
rect 28310 810 28340 840
rect 28610 810 28640 840
rect -640 10 -610 40
rect -40 10 -10 40
rect 8360 10 8390 40
rect 10760 10 10790 40
rect 15560 10 15590 40
rect 17960 10 17990 40
rect 20360 10 20390 40
rect 24560 10 24590 40
rect 28760 10 28790 40
rect -640 -40 -610 -10
rect -40 -40 -10 -10
rect 8360 -40 8390 -10
rect 10760 -40 10790 -10
rect 15560 -40 15590 -10
rect 17960 -40 17990 -10
rect 20360 -40 20390 -10
rect 24560 -40 24590 -10
rect 28760 -40 28790 -10
rect -640 -90 -610 -60
rect -40 -90 -10 -60
rect 8360 -90 8390 -60
rect 10760 -90 10790 -60
rect 15560 -90 15590 -60
rect 17960 -90 17990 -60
rect 20360 -90 20390 -60
rect 24560 -90 24590 -60
rect 28760 -90 28790 -60
rect -490 -890 -460 -860
rect -340 -890 -310 -860
rect -190 -890 -160 -860
rect 110 -890 140 -860
rect 410 -890 440 -860
rect 710 -890 740 -860
rect 1010 -890 1040 -860
rect 1310 -890 1340 -860
rect 1610 -890 1640 -860
rect 1910 -890 1940 -860
rect 2210 -890 2240 -860
rect 2360 -890 2390 -860
rect 2510 -890 2540 -860
rect 2810 -890 2840 -860
rect 3110 -890 3140 -860
rect 3410 -890 3440 -860
rect 3710 -890 3740 -860
rect 3860 -890 3890 -860
rect 4010 -890 4040 -860
rect 4310 -890 4340 -860
rect 4460 -890 4490 -860
rect 4610 -890 4640 -860
rect 4910 -890 4940 -860
rect 5210 -890 5240 -860
rect 5510 -890 5540 -860
rect 5810 -890 5840 -860
rect 5960 -890 5990 -860
rect 6110 -890 6140 -860
rect 6410 -890 6440 -860
rect 6710 -890 6740 -860
rect 7010 -890 7040 -860
rect 7310 -890 7340 -860
rect 7610 -890 7640 -860
rect 7910 -890 7940 -860
rect 8210 -890 8240 -860
rect 8510 -890 8540 -860
rect 8810 -890 8840 -860
rect 9110 -890 9140 -860
rect 9410 -890 9440 -860
rect 9560 -890 9590 -860
rect 9710 -890 9740 -860
rect 10010 -890 10040 -860
rect 10310 -890 10340 -860
rect 10610 -890 10640 -860
rect 10910 -890 10940 -860
rect 11210 -890 11240 -860
rect 11510 -890 11540 -860
rect 11810 -890 11840 -860
rect 12110 -890 12140 -860
rect 12410 -890 12440 -860
rect 12560 -890 12590 -860
rect 12710 -890 12740 -860
rect 13010 -890 13040 -860
rect 13160 -890 13190 -860
rect 13310 -890 13340 -860
rect 13610 -890 13640 -860
rect 13760 -890 13790 -860
rect 13910 -890 13940 -860
rect 14210 -890 14240 -860
rect 14510 -890 14540 -860
rect 14810 -890 14840 -860
rect 15110 -890 15140 -860
rect 15410 -890 15440 -860
rect 15710 -890 15740 -860
rect 16010 -890 16040 -860
rect 16310 -890 16340 -860
rect 16610 -890 16640 -860
rect 16760 -890 16790 -860
rect 16910 -890 16940 -860
rect 17210 -890 17240 -860
rect 17510 -890 17540 -860
rect 17810 -890 17840 -860
rect 18110 -890 18140 -860
rect 18410 -890 18440 -860
rect 18710 -890 18740 -860
rect 19010 -890 19040 -860
rect 19160 -890 19190 -860
rect 19310 -890 19340 -860
rect 19610 -890 19640 -860
rect 19910 -890 19940 -860
rect 20210 -890 20240 -860
rect 20510 -890 20540 -860
rect 20810 -890 20840 -860
rect 21110 -890 21140 -860
rect 21410 -890 21440 -860
rect 21710 -890 21740 -860
rect 22010 -890 22040 -860
rect 22310 -890 22340 -860
rect 22460 -890 22490 -860
rect 22610 -890 22640 -860
rect 22910 -890 22940 -860
rect 23210 -890 23240 -860
rect 23510 -890 23540 -860
rect 23810 -890 23840 -860
rect 24110 -890 24140 -860
rect 24410 -890 24440 -860
rect 24710 -890 24740 -860
rect 25010 -890 25040 -860
rect 25310 -890 25340 -860
rect 25610 -890 25640 -860
rect 25760 -890 25790 -860
rect 25910 -890 25940 -860
rect 26210 -890 26240 -860
rect 26510 -890 26540 -860
rect 26660 -890 26690 -860
rect 26810 -890 26840 -860
rect 27110 -890 27140 -860
rect 27410 -890 27440 -860
rect 27560 -890 27590 -860
rect 27710 -890 27740 -860
rect 28010 -890 28040 -860
rect 28310 -890 28340 -860
rect 28610 -890 28640 -860
rect -640 -1690 -610 -1660
rect -40 -1690 -10 -1660
rect 8360 -1690 8390 -1660
rect 10760 -1690 10790 -1660
rect 15560 -1690 15590 -1660
rect 17960 -1690 17990 -1660
rect 20360 -1690 20390 -1660
rect 24560 -1690 24590 -1660
rect 28760 -1690 28790 -1660
rect -640 -1740 -610 -1710
rect -40 -1740 -10 -1710
rect 8360 -1740 8390 -1710
rect 10760 -1740 10790 -1710
rect 15560 -1740 15590 -1710
rect 17960 -1740 17990 -1710
rect 20360 -1740 20390 -1710
rect 24560 -1740 24590 -1710
rect 28760 -1740 28790 -1710
<< metal3 >>
rect -650 5590 17950 5600
rect -650 5560 -640 5590
rect -610 5560 8360 5590
rect 8390 5560 8660 5590
rect 8690 5560 8960 5590
rect 8990 5560 9260 5590
rect 9290 5560 9560 5590
rect 9590 5560 9860 5590
rect 9890 5560 10160 5590
rect 10190 5560 10460 5590
rect 10490 5560 10760 5590
rect 10790 5560 11960 5590
rect 11990 5560 13160 5590
rect 13190 5560 14360 5590
rect 14390 5560 15560 5590
rect 15590 5560 17950 5590
rect -650 5500 17950 5560
rect 18000 5590 32100 5600
rect 18000 5560 20360 5590
rect 20390 5560 22460 5590
rect 22490 5560 24560 5590
rect 24590 5560 26660 5590
rect 26690 5560 28160 5590
rect 28190 5560 28760 5590
rect 28790 5560 32060 5590
rect 32090 5560 32100 5590
rect 18000 5500 32100 5560
rect -650 5400 32100 5450
rect -650 5300 32100 5350
rect -650 5200 32100 5250
rect -650 5100 32100 5150
rect -650 5000 32100 5050
rect -500 4945 -450 4950
rect -500 4905 -495 4945
rect -455 4905 -450 4945
rect -500 4900 -450 4905
rect -350 4945 -300 4950
rect -350 4905 -345 4945
rect -305 4905 -300 4945
rect -350 4900 -300 4905
rect -200 4945 -150 4950
rect -200 4905 -195 4945
rect -155 4905 -150 4945
rect -200 4900 -150 4905
rect 100 4945 150 4950
rect 100 4905 105 4945
rect 145 4905 150 4945
rect 100 4900 150 4905
rect 400 4945 450 4950
rect 400 4905 405 4945
rect 445 4905 450 4945
rect 400 4900 450 4905
rect 700 4945 750 4950
rect 700 4905 705 4945
rect 745 4905 750 4945
rect 700 4900 750 4905
rect 1000 4945 1050 4950
rect 1000 4905 1005 4945
rect 1045 4905 1050 4945
rect 1000 4900 1050 4905
rect 1150 4945 1200 4950
rect 1150 4905 1155 4945
rect 1195 4905 1200 4945
rect 1150 4900 1200 4905
rect 1300 4945 1350 4950
rect 1300 4905 1305 4945
rect 1345 4905 1350 4945
rect 1300 4900 1350 4905
rect 1600 4945 1650 4950
rect 1600 4905 1605 4945
rect 1645 4905 1650 4945
rect 1600 4900 1650 4905
rect 1900 4945 1950 4950
rect 1900 4905 1905 4945
rect 1945 4905 1950 4945
rect 1900 4900 1950 4905
rect 2050 4945 2100 4950
rect 2050 4905 2055 4945
rect 2095 4905 2100 4945
rect 2050 4900 2100 4905
rect 2200 4945 2250 4950
rect 2200 4905 2205 4945
rect 2245 4905 2250 4945
rect 2200 4900 2250 4905
rect 2500 4945 2550 4950
rect 2500 4905 2505 4945
rect 2545 4905 2550 4945
rect 2500 4900 2550 4905
rect 2800 4945 2850 4950
rect 2800 4905 2805 4945
rect 2845 4905 2850 4945
rect 2800 4900 2850 4905
rect 2950 4945 3000 4950
rect 2950 4905 2955 4945
rect 2995 4905 3000 4945
rect 2950 4900 3000 4905
rect 3100 4945 3150 4950
rect 3100 4905 3105 4945
rect 3145 4905 3150 4945
rect 3100 4900 3150 4905
rect 3400 4945 3450 4950
rect 3400 4905 3405 4945
rect 3445 4905 3450 4945
rect 3400 4900 3450 4905
rect 3700 4945 3750 4950
rect 3700 4905 3705 4945
rect 3745 4905 3750 4945
rect 3700 4900 3750 4905
rect 4000 4945 4050 4950
rect 4000 4905 4005 4945
rect 4045 4905 4050 4945
rect 4000 4900 4050 4905
rect 4300 4945 4350 4950
rect 4300 4905 4305 4945
rect 4345 4905 4350 4945
rect 4300 4900 4350 4905
rect 4600 4945 4650 4950
rect 4600 4905 4605 4945
rect 4645 4905 4650 4945
rect 4600 4900 4650 4905
rect 4900 4945 4950 4950
rect 4900 4905 4905 4945
rect 4945 4905 4950 4945
rect 4900 4900 4950 4905
rect 5200 4945 5250 4950
rect 5200 4905 5205 4945
rect 5245 4905 5250 4945
rect 5200 4900 5250 4905
rect 5350 4945 5400 4950
rect 5350 4905 5355 4945
rect 5395 4905 5400 4945
rect 5350 4900 5400 4905
rect 5500 4945 5550 4950
rect 5500 4905 5505 4945
rect 5545 4905 5550 4945
rect 5500 4900 5550 4905
rect 5800 4945 5850 4950
rect 5800 4905 5805 4945
rect 5845 4905 5850 4945
rect 5800 4900 5850 4905
rect 6100 4945 6150 4950
rect 6100 4905 6105 4945
rect 6145 4905 6150 4945
rect 6100 4900 6150 4905
rect 6250 4945 6300 4950
rect 6250 4905 6255 4945
rect 6295 4905 6300 4945
rect 6250 4900 6300 4905
rect 6400 4945 6450 4950
rect 6400 4905 6405 4945
rect 6445 4905 6450 4945
rect 6400 4900 6450 4905
rect 6700 4945 6750 4950
rect 6700 4905 6705 4945
rect 6745 4905 6750 4945
rect 6700 4900 6750 4905
rect 7000 4945 7050 4950
rect 7000 4905 7005 4945
rect 7045 4905 7050 4945
rect 7000 4900 7050 4905
rect 7150 4945 7200 4950
rect 7150 4905 7155 4945
rect 7195 4905 7200 4945
rect 7150 4900 7200 4905
rect 7300 4945 7350 4950
rect 7300 4905 7305 4945
rect 7345 4905 7350 4945
rect 7300 4900 7350 4905
rect 7600 4945 7650 4950
rect 7600 4905 7605 4945
rect 7645 4905 7650 4945
rect 7600 4900 7650 4905
rect 7900 4945 7950 4950
rect 7900 4905 7905 4945
rect 7945 4905 7950 4945
rect 7900 4900 7950 4905
rect 8200 4945 8250 4950
rect 8200 4905 8205 4945
rect 8245 4905 8250 4945
rect 8200 4900 8250 4905
rect 8500 4945 8550 4950
rect 8500 4905 8505 4945
rect 8545 4905 8550 4945
rect 8500 4900 8550 4905
rect 8800 4945 8850 4950
rect 8800 4905 8805 4945
rect 8845 4905 8850 4945
rect 8800 4900 8850 4905
rect 9100 4945 9150 4950
rect 9100 4905 9105 4945
rect 9145 4905 9150 4945
rect 9100 4900 9150 4905
rect 9400 4945 9450 4950
rect 9400 4905 9405 4945
rect 9445 4905 9450 4945
rect 9400 4900 9450 4905
rect 9700 4945 9750 4950
rect 9700 4905 9705 4945
rect 9745 4905 9750 4945
rect 9700 4900 9750 4905
rect 10000 4945 10050 4950
rect 10000 4905 10005 4945
rect 10045 4905 10050 4945
rect 10000 4900 10050 4905
rect 10300 4945 10350 4950
rect 10300 4905 10305 4945
rect 10345 4905 10350 4945
rect 10300 4900 10350 4905
rect 10600 4945 10650 4950
rect 10600 4905 10605 4945
rect 10645 4905 10650 4945
rect 10600 4900 10650 4905
rect 10900 4945 10950 4950
rect 10900 4905 10905 4945
rect 10945 4905 10950 4945
rect 10900 4900 10950 4905
rect 11200 4945 11250 4950
rect 11200 4905 11205 4945
rect 11245 4905 11250 4945
rect 11200 4900 11250 4905
rect 11350 4945 11400 4950
rect 11350 4905 11355 4945
rect 11395 4905 11400 4945
rect 11350 4900 11400 4905
rect 11500 4945 11550 4950
rect 11500 4905 11505 4945
rect 11545 4905 11550 4945
rect 11500 4900 11550 4905
rect 11800 4945 11850 4950
rect 11800 4905 11805 4945
rect 11845 4905 11850 4945
rect 11800 4900 11850 4905
rect 12100 4945 12150 4950
rect 12100 4905 12105 4945
rect 12145 4905 12150 4945
rect 12100 4900 12150 4905
rect 12400 4945 12450 4950
rect 12400 4905 12405 4945
rect 12445 4905 12450 4945
rect 12400 4900 12450 4905
rect 12550 4945 12600 4950
rect 12550 4905 12555 4945
rect 12595 4905 12600 4945
rect 12550 4900 12600 4905
rect 12700 4945 12750 4950
rect 12700 4905 12705 4945
rect 12745 4905 12750 4945
rect 12700 4900 12750 4905
rect 13000 4945 13050 4950
rect 13000 4905 13005 4945
rect 13045 4905 13050 4945
rect 13000 4900 13050 4905
rect 13300 4945 13350 4950
rect 13300 4905 13305 4945
rect 13345 4905 13350 4945
rect 13300 4900 13350 4905
rect 13600 4945 13650 4950
rect 13600 4905 13605 4945
rect 13645 4905 13650 4945
rect 13600 4900 13650 4905
rect 13750 4945 13800 4950
rect 13750 4905 13755 4945
rect 13795 4905 13800 4945
rect 13750 4900 13800 4905
rect 13900 4945 13950 4950
rect 13900 4905 13905 4945
rect 13945 4905 13950 4945
rect 13900 4900 13950 4905
rect 14200 4945 14250 4950
rect 14200 4905 14205 4945
rect 14245 4905 14250 4945
rect 14200 4900 14250 4905
rect 14500 4945 14550 4950
rect 14500 4905 14505 4945
rect 14545 4905 14550 4945
rect 14500 4900 14550 4905
rect 14800 4945 14850 4950
rect 14800 4905 14805 4945
rect 14845 4905 14850 4945
rect 14800 4900 14850 4905
rect 14950 4945 15000 4950
rect 14950 4905 14955 4945
rect 14995 4905 15000 4945
rect 14950 4900 15000 4905
rect 15100 4945 15150 4950
rect 15100 4905 15105 4945
rect 15145 4905 15150 4945
rect 15100 4900 15150 4905
rect 15400 4945 15450 4950
rect 15400 4905 15405 4945
rect 15445 4905 15450 4945
rect 15400 4900 15450 4905
rect 15700 4945 15750 4950
rect 15700 4905 15705 4945
rect 15745 4905 15750 4945
rect 15700 4900 15750 4905
rect 16000 4945 16050 4950
rect 16000 4905 16005 4945
rect 16045 4905 16050 4945
rect 16000 4900 16050 4905
rect 16300 4945 16350 4950
rect 16300 4905 16305 4945
rect 16345 4905 16350 4945
rect 16300 4900 16350 4905
rect 16600 4945 16650 4950
rect 16600 4905 16605 4945
rect 16645 4905 16650 4945
rect 16600 4900 16650 4905
rect 16750 4945 16800 4950
rect 16750 4905 16755 4945
rect 16795 4905 16800 4945
rect 16750 4900 16800 4905
rect 16900 4945 16950 4950
rect 16900 4905 16905 4945
rect 16945 4905 16950 4945
rect 16900 4900 16950 4905
rect 17200 4945 17250 4950
rect 17200 4905 17205 4945
rect 17245 4905 17250 4945
rect 17200 4900 17250 4905
rect 17500 4945 17550 4950
rect 17500 4905 17505 4945
rect 17545 4905 17550 4945
rect 17500 4900 17550 4905
rect 17800 4945 17850 4950
rect 17800 4905 17805 4945
rect 17845 4905 17850 4945
rect 17800 4900 17850 4905
rect 18100 4945 18150 4950
rect 18100 4905 18105 4945
rect 18145 4905 18150 4945
rect 18100 4900 18150 4905
rect 18400 4945 18450 4950
rect 18400 4905 18405 4945
rect 18445 4905 18450 4945
rect 18400 4900 18450 4905
rect 18700 4945 18750 4950
rect 18700 4905 18705 4945
rect 18745 4905 18750 4945
rect 18700 4900 18750 4905
rect 19000 4945 19050 4950
rect 19000 4905 19005 4945
rect 19045 4905 19050 4945
rect 19000 4900 19050 4905
rect 19150 4945 19200 4950
rect 19150 4905 19155 4945
rect 19195 4905 19200 4945
rect 19150 4900 19200 4905
rect 19300 4945 19350 4950
rect 19300 4905 19305 4945
rect 19345 4905 19350 4945
rect 19300 4900 19350 4905
rect 19600 4945 19650 4950
rect 19600 4905 19605 4945
rect 19645 4905 19650 4945
rect 19600 4900 19650 4905
rect 19900 4945 19950 4950
rect 19900 4905 19905 4945
rect 19945 4905 19950 4945
rect 19900 4900 19950 4905
rect 20200 4945 20250 4950
rect 20200 4905 20205 4945
rect 20245 4905 20250 4945
rect 20200 4900 20250 4905
rect 20500 4945 20550 4950
rect 20500 4905 20505 4945
rect 20545 4905 20550 4945
rect 20500 4900 20550 4905
rect 20800 4945 20850 4950
rect 20800 4905 20805 4945
rect 20845 4905 20850 4945
rect 20800 4900 20850 4905
rect 20950 4945 21000 4950
rect 20950 4905 20955 4945
rect 20995 4905 21000 4945
rect 20950 4900 21000 4905
rect 21100 4945 21150 4950
rect 21100 4905 21105 4945
rect 21145 4905 21150 4945
rect 21100 4900 21150 4905
rect 21400 4940 21450 4950
rect 21400 4910 21410 4940
rect 21440 4910 21450 4940
rect 21400 4900 21450 4910
rect 21700 4945 21750 4950
rect 21700 4905 21705 4945
rect 21745 4905 21750 4945
rect 21700 4900 21750 4905
rect 21850 4945 21900 4950
rect 21850 4905 21855 4945
rect 21895 4905 21900 4945
rect 21850 4900 21900 4905
rect 22000 4945 22050 4950
rect 22000 4905 22005 4945
rect 22045 4905 22050 4945
rect 22000 4900 22050 4905
rect 22300 4945 22350 4950
rect 22300 4905 22305 4945
rect 22345 4905 22350 4945
rect 22300 4900 22350 4905
rect 22600 4945 22650 4950
rect 22600 4905 22605 4945
rect 22645 4905 22650 4945
rect 22600 4900 22650 4905
rect 22900 4945 22950 4950
rect 22900 4905 22905 4945
rect 22945 4905 22950 4945
rect 22900 4900 22950 4905
rect 23050 4945 23100 4950
rect 23050 4905 23055 4945
rect 23095 4905 23100 4945
rect 23050 4900 23100 4905
rect 23200 4945 23250 4950
rect 23200 4905 23205 4945
rect 23245 4905 23250 4945
rect 23200 4900 23250 4905
rect 23350 4945 23400 4950
rect 23350 4905 23355 4945
rect 23395 4905 23400 4945
rect 23350 4900 23400 4905
rect 23500 4940 23550 4950
rect 23500 4910 23510 4940
rect 23540 4910 23550 4940
rect 23500 4900 23550 4910
rect 23650 4945 23700 4950
rect 23650 4905 23655 4945
rect 23695 4905 23700 4945
rect 23650 4900 23700 4905
rect 23800 4945 23850 4950
rect 23800 4905 23805 4945
rect 23845 4905 23850 4945
rect 23800 4900 23850 4905
rect 23950 4945 24000 4950
rect 23950 4905 23955 4945
rect 23995 4905 24000 4945
rect 23950 4900 24000 4905
rect 24100 4945 24150 4950
rect 24100 4905 24105 4945
rect 24145 4905 24150 4945
rect 24100 4900 24150 4905
rect 24400 4945 24450 4950
rect 24400 4905 24405 4945
rect 24445 4905 24450 4945
rect 24400 4900 24450 4905
rect 24700 4945 24750 4950
rect 24700 4905 24705 4945
rect 24745 4905 24750 4945
rect 24700 4900 24750 4905
rect 25000 4945 25050 4950
rect 25000 4905 25005 4945
rect 25045 4905 25050 4945
rect 25000 4900 25050 4905
rect 25450 4945 25500 4950
rect 25450 4905 25455 4945
rect 25495 4905 25500 4945
rect 25450 4900 25500 4905
rect 25600 4945 25650 4950
rect 25600 4905 25605 4945
rect 25645 4905 25650 4945
rect 25600 4900 25650 4905
rect 25750 4945 25800 4950
rect 25750 4905 25755 4945
rect 25795 4905 25800 4945
rect 25750 4900 25800 4905
rect 26200 4945 26250 4950
rect 26200 4905 26205 4945
rect 26245 4905 26250 4945
rect 26200 4900 26250 4905
rect 26500 4945 26550 4950
rect 26500 4905 26505 4945
rect 26545 4905 26550 4945
rect 26500 4900 26550 4905
rect 26800 4945 26850 4950
rect 26800 4905 26805 4945
rect 26845 4905 26850 4945
rect 26800 4900 26850 4905
rect 27100 4945 27150 4950
rect 27100 4905 27105 4945
rect 27145 4905 27150 4945
rect 27100 4900 27150 4905
rect 27550 4945 27600 4950
rect 27550 4905 27555 4945
rect 27595 4905 27600 4945
rect 27550 4900 27600 4905
rect 27700 4945 27750 4950
rect 27700 4905 27705 4945
rect 27745 4905 27750 4945
rect 27700 4900 27750 4905
rect 27850 4945 27900 4950
rect 27850 4905 27855 4945
rect 27895 4905 27900 4945
rect 27850 4900 27900 4905
rect 28300 4945 28350 4950
rect 28300 4905 28305 4945
rect 28345 4905 28350 4945
rect 28300 4900 28350 4905
rect 28600 4945 28650 4950
rect 28600 4905 28605 4945
rect 28645 4905 28650 4945
rect 28600 4900 28650 4905
rect 28750 4945 28800 4950
rect 28750 4905 28755 4945
rect 28795 4905 28800 4945
rect 28750 4900 28800 4905
rect 28900 4945 28950 4950
rect 28900 4905 28905 4945
rect 28945 4905 28950 4945
rect 28900 4900 28950 4905
rect 29200 4945 29250 4950
rect 29200 4905 29205 4945
rect 29245 4905 29250 4945
rect 29200 4900 29250 4905
rect 29350 4945 29400 4950
rect 29350 4905 29355 4945
rect 29395 4905 29400 4945
rect 29350 4900 29400 4905
rect 29650 4945 29700 4950
rect 29650 4905 29655 4945
rect 29695 4905 29700 4945
rect 29650 4900 29700 4905
rect 29800 4940 29850 4950
rect 29800 4910 29810 4940
rect 29840 4910 29850 4940
rect 29800 4900 29850 4910
rect 29950 4945 30000 4950
rect 29950 4905 29955 4945
rect 29995 4905 30000 4945
rect 29950 4900 30000 4905
rect 30250 4945 30300 4950
rect 30250 4905 30255 4945
rect 30295 4905 30300 4945
rect 30250 4900 30300 4905
rect 30400 4940 30450 4950
rect 30400 4910 30410 4940
rect 30440 4910 30450 4940
rect 30400 4900 30450 4910
rect 30550 4945 30600 4950
rect 30550 4905 30555 4945
rect 30595 4905 30600 4945
rect 30550 4900 30600 4905
rect 30850 4945 30900 4950
rect 30850 4905 30855 4945
rect 30895 4905 30900 4945
rect 30850 4900 30900 4905
rect 31000 4945 31050 4950
rect 31000 4905 31005 4945
rect 31045 4905 31050 4945
rect 31000 4900 31050 4905
rect 31150 4940 31200 4950
rect 31150 4910 31160 4940
rect 31190 4910 31200 4940
rect 31150 4900 31200 4910
rect 31450 4945 31500 4950
rect 31450 4905 31455 4945
rect 31495 4905 31500 4945
rect 31450 4900 31500 4905
rect 31600 4945 31650 4950
rect 31600 4905 31605 4945
rect 31645 4905 31650 4945
rect 31600 4900 31650 4905
rect 31900 4945 31950 4950
rect 31900 4905 31905 4945
rect 31945 4905 31950 4945
rect 31900 4900 31950 4905
rect 32050 4945 32100 4950
rect 32050 4905 32055 4945
rect 32095 4905 32100 4945
rect 32050 4900 32100 4905
rect -650 4800 32100 4850
rect -650 4745 32100 4750
rect -650 4705 13755 4745
rect 13795 4705 14955 4745
rect 14995 4705 29355 4745
rect 29395 4705 31455 4745
rect 31495 4705 32100 4745
rect -650 4700 32100 4705
rect -650 4600 32100 4650
rect -650 4545 32100 4550
rect -650 4505 11355 4545
rect 11395 4505 12555 4545
rect 12595 4505 20955 4545
rect 20995 4505 21855 4545
rect 21895 4505 23055 4545
rect 23095 4505 23955 4545
rect 23995 4505 28755 4545
rect 28795 4505 32055 4545
rect 32095 4505 32100 4545
rect -650 4500 32100 4505
rect -650 4400 32100 4450
rect -650 4290 32100 4350
rect -650 4260 -640 4290
rect -610 4260 -40 4290
rect -10 4260 4160 4290
rect 4190 4260 8360 4290
rect 8390 4260 8660 4290
rect 8690 4260 8960 4290
rect 8990 4260 9260 4290
rect 9290 4260 9560 4290
rect 9590 4260 9860 4290
rect 9890 4260 10160 4290
rect 10190 4260 10460 4290
rect 10490 4260 10760 4290
rect 10790 4260 11960 4290
rect 11990 4260 13160 4290
rect 13190 4260 14360 4290
rect 14390 4260 15560 4290
rect 15590 4260 20360 4290
rect 20390 4260 22460 4290
rect 22490 4260 24560 4290
rect 24590 4260 26660 4290
rect 26690 4260 28160 4290
rect 28190 4260 28760 4290
rect 28790 4260 32060 4290
rect 32090 4260 32100 4290
rect -650 4200 32100 4260
rect -650 4100 32100 4150
rect -650 4045 32100 4050
rect -650 4005 31005 4045
rect 31045 4005 32100 4045
rect -650 4000 32100 4005
rect -650 3900 32100 3950
rect -650 3845 32100 3850
rect -650 3805 10905 3845
rect 10945 3805 11205 3845
rect 11245 3805 11505 3845
rect 11545 3805 11805 3845
rect 11845 3805 12105 3845
rect 12145 3805 12405 3845
rect 12445 3805 12705 3845
rect 12745 3805 13005 3845
rect 13045 3805 13305 3845
rect 13345 3805 13605 3845
rect 13645 3805 13905 3845
rect 13945 3805 14205 3845
rect 14245 3805 14505 3845
rect 14545 3805 14805 3845
rect 14845 3805 20505 3845
rect 20545 3805 20805 3845
rect 20845 3805 21105 3845
rect 21145 3805 21405 3845
rect 21445 3805 21705 3845
rect 21745 3805 22005 3845
rect 22045 3805 22305 3845
rect 22345 3805 22455 3845
rect 22495 3805 22605 3845
rect 22645 3805 22905 3845
rect 22945 3805 23205 3845
rect 23245 3805 23505 3845
rect 23545 3805 23805 3845
rect 23845 3805 24105 3845
rect 24145 3805 24405 3845
rect 24445 3805 28305 3845
rect 28345 3805 28605 3845
rect 28645 3805 28905 3845
rect 28945 3805 29205 3845
rect 29245 3805 29655 3845
rect 29695 3805 31605 3845
rect 31645 3805 31905 3845
rect 31945 3805 32100 3845
rect -650 3800 32100 3805
rect -650 3700 32100 3750
rect -500 3645 -450 3650
rect -500 3605 -495 3645
rect -455 3605 -450 3645
rect -500 3600 -450 3605
rect -350 3645 -300 3650
rect -350 3605 -345 3645
rect -305 3605 -300 3645
rect -350 3600 -300 3605
rect -200 3645 -150 3650
rect -200 3605 -195 3645
rect -155 3605 -150 3645
rect -200 3600 -150 3605
rect 100 3645 150 3650
rect 100 3605 105 3645
rect 145 3605 150 3645
rect 100 3600 150 3605
rect 400 3645 450 3650
rect 400 3605 405 3645
rect 445 3605 450 3645
rect 400 3600 450 3605
rect 700 3645 750 3650
rect 700 3605 705 3645
rect 745 3605 750 3645
rect 700 3600 750 3605
rect 1000 3645 1050 3650
rect 1000 3605 1005 3645
rect 1045 3605 1050 3645
rect 1000 3600 1050 3605
rect 1150 3645 1200 3650
rect 1150 3605 1155 3645
rect 1195 3605 1200 3645
rect 1150 3600 1200 3605
rect 1300 3645 1350 3650
rect 1300 3605 1305 3645
rect 1345 3605 1350 3645
rect 1300 3600 1350 3605
rect 1600 3645 1650 3650
rect 1600 3605 1605 3645
rect 1645 3605 1650 3645
rect 1600 3600 1650 3605
rect 1900 3645 1950 3650
rect 1900 3605 1905 3645
rect 1945 3605 1950 3645
rect 1900 3600 1950 3605
rect 2050 3645 2100 3650
rect 2050 3605 2055 3645
rect 2095 3605 2100 3645
rect 2050 3600 2100 3605
rect 2200 3645 2250 3650
rect 2200 3605 2205 3645
rect 2245 3605 2250 3645
rect 2200 3600 2250 3605
rect 2500 3645 2550 3650
rect 2500 3605 2505 3645
rect 2545 3605 2550 3645
rect 2500 3600 2550 3605
rect 2800 3645 2850 3650
rect 2800 3605 2805 3645
rect 2845 3605 2850 3645
rect 2800 3600 2850 3605
rect 2950 3645 3000 3650
rect 2950 3605 2955 3645
rect 2995 3605 3000 3645
rect 2950 3600 3000 3605
rect 3100 3645 3150 3650
rect 3100 3605 3105 3645
rect 3145 3605 3150 3645
rect 3100 3600 3150 3605
rect 3400 3645 3450 3650
rect 3400 3605 3405 3645
rect 3445 3605 3450 3645
rect 3400 3600 3450 3605
rect 3700 3645 3750 3650
rect 3700 3605 3705 3645
rect 3745 3605 3750 3645
rect 3700 3600 3750 3605
rect 4000 3645 4050 3650
rect 4000 3605 4005 3645
rect 4045 3605 4050 3645
rect 4000 3600 4050 3605
rect 4300 3645 4350 3650
rect 4300 3605 4305 3645
rect 4345 3605 4350 3645
rect 4300 3600 4350 3605
rect 4600 3645 4650 3650
rect 4600 3605 4605 3645
rect 4645 3605 4650 3645
rect 4600 3600 4650 3605
rect 4900 3645 4950 3650
rect 4900 3605 4905 3645
rect 4945 3605 4950 3645
rect 4900 3600 4950 3605
rect 5200 3645 5250 3650
rect 5200 3605 5205 3645
rect 5245 3605 5250 3645
rect 5200 3600 5250 3605
rect 5350 3645 5400 3650
rect 5350 3605 5355 3645
rect 5395 3605 5400 3645
rect 5350 3600 5400 3605
rect 5500 3645 5550 3650
rect 5500 3605 5505 3645
rect 5545 3605 5550 3645
rect 5500 3600 5550 3605
rect 5800 3645 5850 3650
rect 5800 3605 5805 3645
rect 5845 3605 5850 3645
rect 5800 3600 5850 3605
rect 6100 3645 6150 3650
rect 6100 3605 6105 3645
rect 6145 3605 6150 3645
rect 6100 3600 6150 3605
rect 6250 3645 6300 3650
rect 6250 3605 6255 3645
rect 6295 3605 6300 3645
rect 6250 3600 6300 3605
rect 6400 3645 6450 3650
rect 6400 3605 6405 3645
rect 6445 3605 6450 3645
rect 6400 3600 6450 3605
rect 6700 3645 6750 3650
rect 6700 3605 6705 3645
rect 6745 3605 6750 3645
rect 6700 3600 6750 3605
rect 7000 3645 7050 3650
rect 7000 3605 7005 3645
rect 7045 3605 7050 3645
rect 7000 3600 7050 3605
rect 7150 3645 7200 3650
rect 7150 3605 7155 3645
rect 7195 3605 7200 3645
rect 7150 3600 7200 3605
rect 7300 3645 7350 3650
rect 7300 3605 7305 3645
rect 7345 3605 7350 3645
rect 7300 3600 7350 3605
rect 7600 3645 7650 3650
rect 7600 3605 7605 3645
rect 7645 3605 7650 3645
rect 7600 3600 7650 3605
rect 7900 3645 7950 3650
rect 7900 3605 7905 3645
rect 7945 3605 7950 3645
rect 7900 3600 7950 3605
rect 8200 3645 8250 3650
rect 8200 3605 8205 3645
rect 8245 3605 8250 3645
rect 8200 3600 8250 3605
rect 8500 3645 8550 3650
rect 8500 3605 8505 3645
rect 8545 3605 8550 3645
rect 8500 3600 8550 3605
rect 8800 3645 8850 3650
rect 8800 3605 8805 3645
rect 8845 3605 8850 3645
rect 8800 3600 8850 3605
rect 9100 3645 9150 3650
rect 9100 3605 9105 3645
rect 9145 3605 9150 3645
rect 9100 3600 9150 3605
rect 9400 3645 9450 3650
rect 9400 3605 9405 3645
rect 9445 3605 9450 3645
rect 9400 3600 9450 3605
rect 9700 3645 9750 3650
rect 9700 3605 9705 3645
rect 9745 3605 9750 3645
rect 9700 3600 9750 3605
rect 10000 3645 10050 3650
rect 10000 3605 10005 3645
rect 10045 3605 10050 3645
rect 10000 3600 10050 3605
rect 10300 3645 10350 3650
rect 10300 3605 10305 3645
rect 10345 3605 10350 3645
rect 10300 3600 10350 3605
rect 10600 3645 10650 3650
rect 10600 3605 10605 3645
rect 10645 3605 10650 3645
rect 10600 3600 10650 3605
rect 10900 3645 10950 3650
rect 10900 3605 10905 3645
rect 10945 3605 10950 3645
rect 10900 3600 10950 3605
rect 11200 3645 11250 3650
rect 11200 3605 11205 3645
rect 11245 3605 11250 3645
rect 11200 3600 11250 3605
rect 11350 3645 11400 3650
rect 11350 3605 11355 3645
rect 11395 3605 11400 3645
rect 11350 3600 11400 3605
rect 11500 3645 11550 3650
rect 11500 3605 11505 3645
rect 11545 3605 11550 3645
rect 11500 3600 11550 3605
rect 11800 3645 11850 3650
rect 11800 3605 11805 3645
rect 11845 3605 11850 3645
rect 11800 3600 11850 3605
rect 12100 3645 12150 3650
rect 12100 3605 12105 3645
rect 12145 3605 12150 3645
rect 12100 3600 12150 3605
rect 12400 3645 12450 3650
rect 12400 3605 12405 3645
rect 12445 3605 12450 3645
rect 12400 3600 12450 3605
rect 12550 3645 12600 3650
rect 12550 3605 12555 3645
rect 12595 3605 12600 3645
rect 12550 3600 12600 3605
rect 12700 3645 12750 3650
rect 12700 3605 12705 3645
rect 12745 3605 12750 3645
rect 12700 3600 12750 3605
rect 13000 3645 13050 3650
rect 13000 3605 13005 3645
rect 13045 3605 13050 3645
rect 13000 3600 13050 3605
rect 13300 3645 13350 3650
rect 13300 3605 13305 3645
rect 13345 3605 13350 3645
rect 13300 3600 13350 3605
rect 13600 3645 13650 3650
rect 13600 3605 13605 3645
rect 13645 3605 13650 3645
rect 13600 3600 13650 3605
rect 13750 3645 13800 3650
rect 13750 3605 13755 3645
rect 13795 3605 13800 3645
rect 13750 3600 13800 3605
rect 13900 3645 13950 3650
rect 13900 3605 13905 3645
rect 13945 3605 13950 3645
rect 13900 3600 13950 3605
rect 14200 3645 14250 3650
rect 14200 3605 14205 3645
rect 14245 3605 14250 3645
rect 14200 3600 14250 3605
rect 14500 3645 14550 3650
rect 14500 3605 14505 3645
rect 14545 3605 14550 3645
rect 14500 3600 14550 3605
rect 14800 3645 14850 3650
rect 14800 3605 14805 3645
rect 14845 3605 14850 3645
rect 14800 3600 14850 3605
rect 14950 3645 15000 3650
rect 14950 3605 14955 3645
rect 14995 3605 15000 3645
rect 14950 3600 15000 3605
rect 15100 3645 15150 3650
rect 15100 3605 15105 3645
rect 15145 3605 15150 3645
rect 15100 3600 15150 3605
rect 15400 3645 15450 3650
rect 15400 3605 15405 3645
rect 15445 3605 15450 3645
rect 15400 3600 15450 3605
rect 15700 3645 15750 3650
rect 15700 3605 15705 3645
rect 15745 3605 15750 3645
rect 15700 3600 15750 3605
rect 16000 3645 16050 3650
rect 16000 3605 16005 3645
rect 16045 3605 16050 3645
rect 16000 3600 16050 3605
rect 16300 3645 16350 3650
rect 16300 3605 16305 3645
rect 16345 3605 16350 3645
rect 16300 3600 16350 3605
rect 16600 3645 16650 3650
rect 16600 3605 16605 3645
rect 16645 3605 16650 3645
rect 16600 3600 16650 3605
rect 16750 3645 16800 3650
rect 16750 3605 16755 3645
rect 16795 3605 16800 3645
rect 16750 3600 16800 3605
rect 16900 3645 16950 3650
rect 16900 3605 16905 3645
rect 16945 3605 16950 3645
rect 16900 3600 16950 3605
rect 17200 3645 17250 3650
rect 17200 3605 17205 3645
rect 17245 3605 17250 3645
rect 17200 3600 17250 3605
rect 17500 3645 17550 3650
rect 17500 3605 17505 3645
rect 17545 3605 17550 3645
rect 17500 3600 17550 3605
rect 17800 3645 17850 3650
rect 17800 3605 17805 3645
rect 17845 3605 17850 3645
rect 17800 3600 17850 3605
rect 18100 3645 18150 3650
rect 18100 3605 18105 3645
rect 18145 3605 18150 3645
rect 18100 3600 18150 3605
rect 18400 3645 18450 3650
rect 18400 3605 18405 3645
rect 18445 3605 18450 3645
rect 18400 3600 18450 3605
rect 18700 3645 18750 3650
rect 18700 3605 18705 3645
rect 18745 3605 18750 3645
rect 18700 3600 18750 3605
rect 19000 3645 19050 3650
rect 19000 3605 19005 3645
rect 19045 3605 19050 3645
rect 19000 3600 19050 3605
rect 19150 3645 19200 3650
rect 19150 3605 19155 3645
rect 19195 3605 19200 3645
rect 19150 3600 19200 3605
rect 19300 3645 19350 3650
rect 19300 3605 19305 3645
rect 19345 3605 19350 3645
rect 19300 3600 19350 3605
rect 19600 3645 19650 3650
rect 19600 3605 19605 3645
rect 19645 3605 19650 3645
rect 19600 3600 19650 3605
rect 19900 3645 19950 3650
rect 19900 3605 19905 3645
rect 19945 3605 19950 3645
rect 19900 3600 19950 3605
rect 20200 3645 20250 3650
rect 20200 3605 20205 3645
rect 20245 3605 20250 3645
rect 20200 3600 20250 3605
rect 20500 3645 20550 3650
rect 20500 3605 20505 3645
rect 20545 3605 20550 3645
rect 20500 3600 20550 3605
rect 20800 3645 20850 3650
rect 20800 3605 20805 3645
rect 20845 3605 20850 3645
rect 20800 3600 20850 3605
rect 20950 3645 21000 3650
rect 20950 3605 20955 3645
rect 20995 3605 21000 3645
rect 20950 3600 21000 3605
rect 21100 3645 21150 3650
rect 21100 3605 21105 3645
rect 21145 3605 21150 3645
rect 21100 3600 21150 3605
rect 21400 3640 21450 3650
rect 21400 3610 21410 3640
rect 21440 3610 21450 3640
rect 21400 3600 21450 3610
rect 21700 3645 21750 3650
rect 21700 3605 21705 3645
rect 21745 3605 21750 3645
rect 21700 3600 21750 3605
rect 21850 3645 21900 3650
rect 21850 3605 21855 3645
rect 21895 3605 21900 3645
rect 21850 3600 21900 3605
rect 22000 3645 22050 3650
rect 22000 3605 22005 3645
rect 22045 3605 22050 3645
rect 22000 3600 22050 3605
rect 22300 3645 22350 3650
rect 22300 3605 22305 3645
rect 22345 3605 22350 3645
rect 22300 3600 22350 3605
rect 22600 3645 22650 3650
rect 22600 3605 22605 3645
rect 22645 3605 22650 3645
rect 22600 3600 22650 3605
rect 22900 3645 22950 3650
rect 22900 3605 22905 3645
rect 22945 3605 22950 3645
rect 22900 3600 22950 3605
rect 23050 3645 23100 3650
rect 23050 3605 23055 3645
rect 23095 3605 23100 3645
rect 23050 3600 23100 3605
rect 23200 3645 23250 3650
rect 23200 3605 23205 3645
rect 23245 3605 23250 3645
rect 23200 3600 23250 3605
rect 23350 3645 23400 3650
rect 23350 3605 23355 3645
rect 23395 3605 23400 3645
rect 23350 3600 23400 3605
rect 23500 3640 23550 3650
rect 23500 3610 23510 3640
rect 23540 3610 23550 3640
rect 23500 3600 23550 3610
rect 23650 3645 23700 3650
rect 23650 3605 23655 3645
rect 23695 3605 23700 3645
rect 23650 3600 23700 3605
rect 23800 3645 23850 3650
rect 23800 3605 23805 3645
rect 23845 3605 23850 3645
rect 23800 3600 23850 3605
rect 23950 3645 24000 3650
rect 23950 3605 23955 3645
rect 23995 3605 24000 3645
rect 23950 3600 24000 3605
rect 24100 3645 24150 3650
rect 24100 3605 24105 3645
rect 24145 3605 24150 3645
rect 24100 3600 24150 3605
rect 24400 3645 24450 3650
rect 24400 3605 24405 3645
rect 24445 3605 24450 3645
rect 24400 3600 24450 3605
rect 24700 3645 24750 3650
rect 24700 3605 24705 3645
rect 24745 3605 24750 3645
rect 24700 3600 24750 3605
rect 25000 3645 25050 3650
rect 25000 3605 25005 3645
rect 25045 3605 25050 3645
rect 25000 3600 25050 3605
rect 25450 3645 25500 3650
rect 25450 3605 25455 3645
rect 25495 3605 25500 3645
rect 25450 3600 25500 3605
rect 25600 3645 25650 3650
rect 25600 3605 25605 3645
rect 25645 3605 25650 3645
rect 25600 3600 25650 3605
rect 25750 3645 25800 3650
rect 25750 3605 25755 3645
rect 25795 3605 25800 3645
rect 25750 3600 25800 3605
rect 26200 3645 26250 3650
rect 26200 3605 26205 3645
rect 26245 3605 26250 3645
rect 26200 3600 26250 3605
rect 26500 3645 26550 3650
rect 26500 3605 26505 3645
rect 26545 3605 26550 3645
rect 26500 3600 26550 3605
rect 26800 3645 26850 3650
rect 26800 3605 26805 3645
rect 26845 3605 26850 3645
rect 26800 3600 26850 3605
rect 27100 3645 27150 3650
rect 27100 3605 27105 3645
rect 27145 3605 27150 3645
rect 27100 3600 27150 3605
rect 27550 3645 27600 3650
rect 27550 3605 27555 3645
rect 27595 3605 27600 3645
rect 27550 3600 27600 3605
rect 27700 3645 27750 3650
rect 27700 3605 27705 3645
rect 27745 3605 27750 3645
rect 27700 3600 27750 3605
rect 27850 3645 27900 3650
rect 27850 3605 27855 3645
rect 27895 3605 27900 3645
rect 27850 3600 27900 3605
rect 28300 3645 28350 3650
rect 28300 3605 28305 3645
rect 28345 3605 28350 3645
rect 28300 3600 28350 3605
rect 28600 3645 28650 3650
rect 28600 3605 28605 3645
rect 28645 3605 28650 3645
rect 28600 3600 28650 3605
rect 28750 3645 28800 3650
rect 28750 3605 28755 3645
rect 28795 3605 28800 3645
rect 28750 3600 28800 3605
rect 28900 3645 28950 3650
rect 28900 3605 28905 3645
rect 28945 3605 28950 3645
rect 28900 3600 28950 3605
rect 29200 3645 29250 3650
rect 29200 3605 29205 3645
rect 29245 3605 29250 3645
rect 29200 3600 29250 3605
rect 29350 3645 29400 3650
rect 29350 3605 29355 3645
rect 29395 3605 29400 3645
rect 29350 3600 29400 3605
rect 29650 3645 29700 3650
rect 29650 3605 29655 3645
rect 29695 3605 29700 3645
rect 29650 3600 29700 3605
rect 29800 3640 29850 3650
rect 29800 3610 29810 3640
rect 29840 3610 29850 3640
rect 29800 3600 29850 3610
rect 29950 3645 30000 3650
rect 29950 3605 29955 3645
rect 29995 3605 30000 3645
rect 29950 3600 30000 3605
rect 30250 3645 30300 3650
rect 30250 3605 30255 3645
rect 30295 3605 30300 3645
rect 30250 3600 30300 3605
rect 30400 3640 30450 3650
rect 30400 3610 30410 3640
rect 30440 3610 30450 3640
rect 30400 3600 30450 3610
rect 30550 3645 30600 3650
rect 30550 3605 30555 3645
rect 30595 3605 30600 3645
rect 30550 3600 30600 3605
rect 30850 3645 30900 3650
rect 30850 3605 30855 3645
rect 30895 3605 30900 3645
rect 30850 3600 30900 3605
rect 31000 3645 31050 3650
rect 31000 3605 31005 3645
rect 31045 3605 31050 3645
rect 31000 3600 31050 3605
rect 31150 3640 31200 3650
rect 31150 3610 31160 3640
rect 31190 3610 31200 3640
rect 31150 3600 31200 3610
rect 31450 3645 31500 3650
rect 31450 3605 31455 3645
rect 31495 3605 31500 3645
rect 31450 3600 31500 3605
rect 31600 3645 31650 3650
rect 31600 3605 31605 3645
rect 31645 3605 31650 3645
rect 31600 3600 31650 3605
rect 31900 3645 31950 3650
rect 31900 3605 31905 3645
rect 31945 3605 31950 3645
rect 31900 3600 31950 3605
rect 32050 3645 32100 3650
rect 32050 3605 32055 3645
rect 32095 3605 32100 3645
rect 32050 3600 32100 3605
rect -650 3500 32100 3550
rect -650 3445 32100 3450
rect -650 3405 -345 3445
rect -305 3405 105 3445
rect 145 3405 405 3445
rect 445 3405 2055 3445
rect 2095 3405 3705 3445
rect 3745 3405 4005 3445
rect 4045 3405 4305 3445
rect 4345 3405 4605 3445
rect 4645 3405 6255 3445
rect 6295 3405 7905 3445
rect 7945 3405 8205 3445
rect 8245 3405 18105 3445
rect 18145 3405 18405 3445
rect 18445 3405 19905 3445
rect 19945 3405 20205 3445
rect 20245 3405 24705 3445
rect 24745 3405 25005 3445
rect 25045 3405 26205 3445
rect 26245 3405 26505 3445
rect 26545 3405 26805 3445
rect 26845 3405 27105 3445
rect 27145 3405 32100 3445
rect -650 3400 32100 3405
rect -650 3345 32100 3350
rect -650 3305 705 3345
rect 745 3305 1005 3345
rect 1045 3305 1155 3345
rect 1195 3305 1305 3345
rect 1345 3305 1605 3345
rect 1645 3305 2505 3345
rect 2545 3305 2805 3345
rect 2845 3305 2955 3345
rect 2995 3305 3105 3345
rect 3145 3305 3405 3345
rect 3445 3305 4905 3345
rect 4945 3305 5205 3345
rect 5245 3305 5355 3345
rect 5395 3305 5505 3345
rect 5545 3305 5805 3345
rect 5845 3305 6705 3345
rect 6745 3305 7005 3345
rect 7045 3305 7155 3345
rect 7195 3305 7305 3345
rect 7345 3305 7605 3345
rect 7645 3305 9555 3345
rect 9595 3305 25455 3345
rect 25495 3305 25755 3345
rect 25795 3305 27555 3345
rect 27595 3305 27855 3345
rect 27895 3305 29955 3345
rect 29995 3305 30255 3345
rect 30295 3305 30555 3345
rect 30595 3305 30855 3345
rect 30895 3305 32100 3345
rect -650 3300 32100 3305
rect -650 3245 32100 3250
rect -650 3205 1905 3245
rect 1945 3205 2205 3245
rect 2245 3205 6105 3245
rect 6145 3205 6405 3245
rect 6445 3205 32100 3245
rect -650 3200 32100 3205
rect -650 3145 32100 3150
rect -650 3105 -495 3145
rect -455 3105 -195 3145
rect -155 3105 32100 3145
rect -650 3100 32100 3105
rect -650 3000 32100 3050
rect -650 2990 17950 3000
rect -650 2960 -640 2990
rect -610 2960 -40 2990
rect -10 2960 4160 2990
rect 4190 2960 8360 2990
rect 8390 2960 8660 2990
rect 8690 2960 8960 2990
rect 8990 2960 9260 2990
rect 9290 2960 9560 2990
rect 9590 2960 9860 2990
rect 9890 2960 10160 2990
rect 10190 2960 10460 2990
rect 10490 2960 10760 2990
rect 10790 2960 11960 2990
rect 11990 2960 13160 2990
rect 13190 2960 14360 2990
rect 14390 2960 15560 2990
rect 15590 2960 17950 2990
rect -650 2950 17950 2960
rect 18000 2990 32100 3000
rect 18000 2960 20360 2990
rect 20390 2960 24560 2990
rect 24590 2960 26660 2990
rect 26690 2960 28160 2990
rect 28190 2960 28760 2990
rect 28790 2960 32060 2990
rect 32090 2960 32100 2990
rect 18000 2950 32100 2960
rect -900 2800 32100 2850
rect -900 2745 28800 2750
rect -900 2705 13305 2745
rect 13345 2705 13605 2745
rect 13645 2705 13905 2745
rect 13945 2705 14205 2745
rect 14245 2705 18705 2745
rect 18745 2705 19005 2745
rect 19045 2705 19305 2745
rect 19345 2705 28800 2745
rect -900 2700 28800 2705
rect -900 2600 28800 2650
rect -900 2300 28800 2550
rect -900 2200 28800 2250
rect -900 2145 28800 2150
rect -900 2105 12105 2145
rect 12145 2105 12405 2145
rect 12445 2105 12705 2145
rect 12745 2105 13005 2145
rect 13045 2105 16305 2145
rect 16345 2105 16605 2145
rect 16645 2105 16905 2145
rect 16945 2105 17205 2145
rect 17245 2105 28800 2145
rect -900 2100 28800 2105
rect -900 2000 28800 2050
rect -900 1690 28800 1700
rect -900 1660 -640 1690
rect -610 1660 -40 1690
rect -10 1660 8360 1690
rect 8390 1660 10760 1690
rect 10790 1660 15560 1690
rect 15590 1660 17960 1690
rect 17990 1660 20360 1690
rect 20390 1660 24560 1690
rect 24590 1660 28760 1690
rect 28790 1660 28800 1690
rect -900 1640 28800 1660
rect -900 1610 -640 1640
rect -610 1610 -40 1640
rect -10 1610 8360 1640
rect 8390 1610 10760 1640
rect 10790 1610 15560 1640
rect 15590 1610 17960 1640
rect 17990 1610 20360 1640
rect 20390 1610 24560 1640
rect 24590 1610 28760 1640
rect 28790 1610 28800 1640
rect -900 1600 28800 1610
rect -900 1500 28800 1550
rect -900 1400 28800 1450
rect -900 1345 28800 1350
rect -900 1305 -495 1345
rect -455 1305 -195 1345
rect -155 1305 28800 1345
rect -900 1300 28800 1305
rect -900 1245 28800 1250
rect -900 1205 3705 1245
rect 3745 1205 4005 1245
rect 4045 1205 4305 1245
rect 4345 1205 4605 1245
rect 4645 1205 28800 1245
rect -900 1200 28800 1205
rect -900 1145 28800 1150
rect -900 1105 1305 1145
rect 1345 1105 1605 1145
rect 1645 1105 1905 1145
rect 1945 1105 2205 1145
rect 2245 1105 2355 1145
rect 2395 1105 2505 1145
rect 2545 1105 2805 1145
rect 2845 1105 3105 1145
rect 3145 1105 3405 1145
rect 3445 1105 4905 1145
rect 4945 1105 5205 1145
rect 5245 1105 5505 1145
rect 5545 1105 5805 1145
rect 5845 1105 5955 1145
rect 5995 1105 6105 1145
rect 6145 1105 6405 1145
rect 6445 1105 6705 1145
rect 6745 1105 7005 1145
rect 7045 1105 21705 1145
rect 21745 1105 22005 1145
rect 22045 1105 22305 1145
rect 22345 1105 22605 1145
rect 22645 1105 22905 1145
rect 22945 1105 23205 1145
rect 23245 1105 28800 1145
rect -900 1100 28800 1105
rect -900 1045 28800 1050
rect -900 1005 -345 1045
rect -305 1005 105 1045
rect 145 1005 405 1045
rect 445 1005 705 1045
rect 745 1005 1005 1045
rect 1045 1005 3855 1045
rect 3895 1005 4455 1045
rect 4495 1005 7305 1045
rect 7345 1005 7605 1045
rect 7645 1005 7905 1045
rect 7945 1005 8205 1045
rect 8245 1005 8505 1045
rect 8545 1005 8805 1045
rect 8845 1005 9105 1045
rect 9145 1005 9405 1045
rect 9445 1005 9705 1045
rect 9745 1005 10005 1045
rect 10045 1005 10305 1045
rect 10345 1005 10605 1045
rect 10645 1005 10905 1045
rect 10945 1005 11205 1045
rect 11245 1005 11505 1045
rect 11545 1005 11805 1045
rect 11845 1005 14505 1045
rect 14545 1005 14805 1045
rect 14845 1005 15105 1045
rect 15145 1005 15405 1045
rect 15445 1005 20505 1045
rect 20545 1005 20805 1045
rect 20845 1005 21105 1045
rect 21145 1005 21405 1045
rect 21445 1005 23505 1045
rect 23545 1005 23805 1045
rect 23845 1005 24105 1045
rect 24145 1005 24405 1045
rect 24445 1005 28800 1045
rect -900 1000 28800 1005
rect -900 900 28800 950
rect -500 845 -450 850
rect -500 805 -495 845
rect -455 805 -450 845
rect -500 800 -450 805
rect -350 845 -300 850
rect -350 805 -345 845
rect -305 805 -300 845
rect -350 800 -300 805
rect -200 845 -150 850
rect -200 805 -195 845
rect -155 805 -150 845
rect -200 800 -150 805
rect 100 845 150 850
rect 100 805 105 845
rect 145 805 150 845
rect 100 800 150 805
rect 400 845 450 850
rect 400 805 405 845
rect 445 805 450 845
rect 400 800 450 805
rect 700 845 750 850
rect 700 805 705 845
rect 745 805 750 845
rect 700 800 750 805
rect 1000 845 1050 850
rect 1000 805 1005 845
rect 1045 805 1050 845
rect 1000 800 1050 805
rect 1300 845 1350 850
rect 1300 805 1305 845
rect 1345 805 1350 845
rect 1300 800 1350 805
rect 1600 845 1650 850
rect 1600 805 1605 845
rect 1645 805 1650 845
rect 1600 800 1650 805
rect 1900 845 1950 850
rect 1900 805 1905 845
rect 1945 805 1950 845
rect 1900 800 1950 805
rect 2200 845 2250 850
rect 2200 805 2205 845
rect 2245 805 2250 845
rect 2200 800 2250 805
rect 2350 845 2400 850
rect 2350 805 2355 845
rect 2395 805 2400 845
rect 2350 800 2400 805
rect 2500 845 2550 850
rect 2500 805 2505 845
rect 2545 805 2550 845
rect 2500 800 2550 805
rect 2800 845 2850 850
rect 2800 805 2805 845
rect 2845 805 2850 845
rect 2800 800 2850 805
rect 3100 845 3150 850
rect 3100 805 3105 845
rect 3145 805 3150 845
rect 3100 800 3150 805
rect 3400 845 3450 850
rect 3400 805 3405 845
rect 3445 805 3450 845
rect 3400 800 3450 805
rect 3700 845 3750 850
rect 3700 805 3705 845
rect 3745 805 3750 845
rect 3700 800 3750 805
rect 3850 845 3900 850
rect 3850 805 3855 845
rect 3895 805 3900 845
rect 3850 800 3900 805
rect 4000 845 4050 850
rect 4000 805 4005 845
rect 4045 805 4050 845
rect 4000 800 4050 805
rect 4300 845 4350 850
rect 4300 805 4305 845
rect 4345 805 4350 845
rect 4300 800 4350 805
rect 4450 845 4500 850
rect 4450 805 4455 845
rect 4495 805 4500 845
rect 4450 800 4500 805
rect 4600 845 4650 850
rect 4600 805 4605 845
rect 4645 805 4650 845
rect 4600 800 4650 805
rect 4900 845 4950 850
rect 4900 805 4905 845
rect 4945 805 4950 845
rect 4900 800 4950 805
rect 5200 845 5250 850
rect 5200 805 5205 845
rect 5245 805 5250 845
rect 5200 800 5250 805
rect 5500 845 5550 850
rect 5500 805 5505 845
rect 5545 805 5550 845
rect 5500 800 5550 805
rect 5800 845 5850 850
rect 5800 805 5805 845
rect 5845 805 5850 845
rect 5800 800 5850 805
rect 5950 845 6000 850
rect 5950 805 5955 845
rect 5995 805 6000 845
rect 5950 800 6000 805
rect 6100 845 6150 850
rect 6100 805 6105 845
rect 6145 805 6150 845
rect 6100 800 6150 805
rect 6400 845 6450 850
rect 6400 805 6405 845
rect 6445 805 6450 845
rect 6400 800 6450 805
rect 6700 845 6750 850
rect 6700 805 6705 845
rect 6745 805 6750 845
rect 6700 800 6750 805
rect 7000 845 7050 850
rect 7000 805 7005 845
rect 7045 805 7050 845
rect 7000 800 7050 805
rect 7300 845 7350 850
rect 7300 805 7305 845
rect 7345 805 7350 845
rect 7300 800 7350 805
rect 7600 845 7650 850
rect 7600 805 7605 845
rect 7645 805 7650 845
rect 7600 800 7650 805
rect 7900 845 7950 850
rect 7900 805 7905 845
rect 7945 805 7950 845
rect 7900 800 7950 805
rect 8200 845 8250 850
rect 8200 805 8205 845
rect 8245 805 8250 845
rect 8200 800 8250 805
rect 8500 845 8550 850
rect 8500 805 8505 845
rect 8545 805 8550 845
rect 8500 800 8550 805
rect 8800 845 8850 850
rect 8800 805 8805 845
rect 8845 805 8850 845
rect 8800 800 8850 805
rect 9100 845 9150 850
rect 9100 805 9105 845
rect 9145 805 9150 845
rect 9100 800 9150 805
rect 9400 845 9450 850
rect 9400 805 9405 845
rect 9445 805 9450 845
rect 9400 800 9450 805
rect 9550 845 9600 850
rect 9550 805 9555 845
rect 9595 805 9600 845
rect 9550 800 9600 805
rect 9700 845 9750 850
rect 9700 805 9705 845
rect 9745 805 9750 845
rect 9700 800 9750 805
rect 10000 845 10050 850
rect 10000 805 10005 845
rect 10045 805 10050 845
rect 10000 800 10050 805
rect 10300 845 10350 850
rect 10300 805 10305 845
rect 10345 805 10350 845
rect 10300 800 10350 805
rect 10600 845 10650 850
rect 10600 805 10605 845
rect 10645 805 10650 845
rect 10600 800 10650 805
rect 10900 845 10950 850
rect 10900 805 10905 845
rect 10945 805 10950 845
rect 10900 800 10950 805
rect 11200 845 11250 850
rect 11200 805 11205 845
rect 11245 805 11250 845
rect 11200 800 11250 805
rect 11500 845 11550 850
rect 11500 805 11505 845
rect 11545 805 11550 845
rect 11500 800 11550 805
rect 11800 845 11850 850
rect 11800 805 11805 845
rect 11845 805 11850 845
rect 11800 800 11850 805
rect 12100 845 12150 850
rect 12100 805 12105 845
rect 12145 805 12150 845
rect 12100 800 12150 805
rect 12400 845 12450 850
rect 12400 805 12405 845
rect 12445 805 12450 845
rect 12400 800 12450 805
rect 12550 845 12600 850
rect 12550 805 12555 845
rect 12595 805 12600 845
rect 12550 800 12600 805
rect 12700 845 12750 850
rect 12700 805 12705 845
rect 12745 805 12750 845
rect 12700 800 12750 805
rect 13000 845 13050 850
rect 13000 805 13005 845
rect 13045 805 13050 845
rect 13000 800 13050 805
rect 13150 840 13200 850
rect 13150 810 13160 840
rect 13190 810 13200 840
rect 13150 800 13200 810
rect 13300 845 13350 850
rect 13300 805 13305 845
rect 13345 805 13350 845
rect 13300 800 13350 805
rect 13600 845 13650 850
rect 13600 805 13605 845
rect 13645 805 13650 845
rect 13600 800 13650 805
rect 13750 845 13800 850
rect 13750 805 13755 845
rect 13795 805 13800 845
rect 13750 800 13800 805
rect 13900 845 13950 850
rect 13900 805 13905 845
rect 13945 805 13950 845
rect 13900 800 13950 805
rect 14200 845 14250 850
rect 14200 805 14205 845
rect 14245 805 14250 845
rect 14200 800 14250 805
rect 14500 845 14550 850
rect 14500 805 14505 845
rect 14545 805 14550 845
rect 14500 800 14550 805
rect 14800 845 14850 850
rect 14800 805 14805 845
rect 14845 805 14850 845
rect 14800 800 14850 805
rect 15100 845 15150 850
rect 15100 805 15105 845
rect 15145 805 15150 845
rect 15100 800 15150 805
rect 15400 845 15450 850
rect 15400 805 15405 845
rect 15445 805 15450 845
rect 15400 800 15450 805
rect 15700 845 15750 850
rect 15700 805 15705 845
rect 15745 805 15750 845
rect 15700 800 15750 805
rect 16000 845 16050 850
rect 16000 805 16005 845
rect 16045 805 16050 845
rect 16000 800 16050 805
rect 16300 845 16350 850
rect 16300 805 16305 845
rect 16345 805 16350 845
rect 16300 800 16350 805
rect 16600 845 16650 850
rect 16600 805 16605 845
rect 16645 805 16650 845
rect 16600 800 16650 805
rect 16750 845 16800 850
rect 16750 805 16755 845
rect 16795 805 16800 845
rect 16750 800 16800 805
rect 16900 845 16950 850
rect 16900 805 16905 845
rect 16945 805 16950 845
rect 16900 800 16950 805
rect 17200 845 17250 850
rect 17200 805 17205 845
rect 17245 805 17250 845
rect 17200 800 17250 805
rect 17500 845 17550 850
rect 17500 805 17505 845
rect 17545 805 17550 845
rect 17500 800 17550 805
rect 17800 845 17850 850
rect 17800 805 17805 845
rect 17845 805 17850 845
rect 17800 800 17850 805
rect 18100 845 18150 850
rect 18100 805 18105 845
rect 18145 805 18150 845
rect 18100 800 18150 805
rect 18400 845 18450 850
rect 18400 805 18405 845
rect 18445 805 18450 845
rect 18400 800 18450 805
rect 18700 845 18750 850
rect 18700 805 18705 845
rect 18745 805 18750 845
rect 18700 800 18750 805
rect 19000 845 19050 850
rect 19000 805 19005 845
rect 19045 805 19050 845
rect 19000 800 19050 805
rect 19150 845 19200 850
rect 19150 805 19155 845
rect 19195 805 19200 845
rect 19150 800 19200 805
rect 19300 845 19350 850
rect 19300 805 19305 845
rect 19345 805 19350 845
rect 19300 800 19350 805
rect 19600 845 19650 850
rect 19600 805 19605 845
rect 19645 805 19650 845
rect 19600 800 19650 805
rect 19900 845 19950 850
rect 19900 805 19905 845
rect 19945 805 19950 845
rect 19900 800 19950 805
rect 20200 845 20250 850
rect 20200 805 20205 845
rect 20245 805 20250 845
rect 20200 800 20250 805
rect 20500 845 20550 850
rect 20500 805 20505 845
rect 20545 805 20550 845
rect 20500 800 20550 805
rect 20800 845 20850 850
rect 20800 805 20805 845
rect 20845 805 20850 845
rect 20800 800 20850 805
rect 21100 845 21150 850
rect 21100 805 21105 845
rect 21145 805 21150 845
rect 21100 800 21150 805
rect 21400 845 21450 850
rect 21400 805 21405 845
rect 21445 805 21450 845
rect 21400 800 21450 805
rect 21700 845 21750 850
rect 21700 805 21705 845
rect 21745 805 21750 845
rect 21700 800 21750 805
rect 22000 845 22050 850
rect 22000 805 22005 845
rect 22045 805 22050 845
rect 22000 800 22050 805
rect 22300 845 22350 850
rect 22300 805 22305 845
rect 22345 805 22350 845
rect 22300 800 22350 805
rect 22450 845 22500 850
rect 22450 805 22455 845
rect 22495 805 22500 845
rect 22450 800 22500 805
rect 22600 845 22650 850
rect 22600 805 22605 845
rect 22645 805 22650 845
rect 22600 800 22650 805
rect 22900 845 22950 850
rect 22900 805 22905 845
rect 22945 805 22950 845
rect 22900 800 22950 805
rect 23200 845 23250 850
rect 23200 805 23205 845
rect 23245 805 23250 845
rect 23200 800 23250 805
rect 23500 845 23550 850
rect 23500 805 23505 845
rect 23545 805 23550 845
rect 23500 800 23550 805
rect 23800 845 23850 850
rect 23800 805 23805 845
rect 23845 805 23850 845
rect 23800 800 23850 805
rect 24100 845 24150 850
rect 24100 805 24105 845
rect 24145 805 24150 845
rect 24100 800 24150 805
rect 24400 845 24450 850
rect 24400 805 24405 845
rect 24445 805 24450 845
rect 24400 800 24450 805
rect 24700 845 24750 850
rect 24700 805 24705 845
rect 24745 805 24750 845
rect 24700 800 24750 805
rect 25000 845 25050 850
rect 25000 805 25005 845
rect 25045 805 25050 845
rect 25000 800 25050 805
rect 25300 845 25350 850
rect 25300 805 25305 845
rect 25345 805 25350 845
rect 25300 800 25350 805
rect 25600 845 25650 850
rect 25600 805 25605 845
rect 25645 805 25650 845
rect 25600 800 25650 805
rect 25750 845 25800 850
rect 25750 805 25755 845
rect 25795 805 25800 845
rect 25750 800 25800 805
rect 25900 845 25950 850
rect 25900 805 25905 845
rect 25945 805 25950 845
rect 25900 800 25950 805
rect 26200 845 26250 850
rect 26200 805 26205 845
rect 26245 805 26250 845
rect 26200 800 26250 805
rect 26500 845 26550 850
rect 26500 805 26505 845
rect 26545 805 26550 845
rect 26500 800 26550 805
rect 26650 845 26700 850
rect 26650 805 26655 845
rect 26695 805 26700 845
rect 26650 800 26700 805
rect 26800 845 26850 850
rect 26800 805 26805 845
rect 26845 805 26850 845
rect 26800 800 26850 805
rect 27100 845 27150 850
rect 27100 805 27105 845
rect 27145 805 27150 845
rect 27100 800 27150 805
rect 27400 845 27450 850
rect 27400 805 27405 845
rect 27445 805 27450 845
rect 27400 800 27450 805
rect 27550 845 27600 850
rect 27550 805 27555 845
rect 27595 805 27600 845
rect 27550 800 27600 805
rect 27700 845 27750 850
rect 27700 805 27705 845
rect 27745 805 27750 845
rect 27700 800 27750 805
rect 28000 845 28050 850
rect 28000 805 28005 845
rect 28045 805 28050 845
rect 28000 800 28050 805
rect 28300 845 28350 850
rect 28300 805 28305 845
rect 28345 805 28350 845
rect 28300 800 28350 805
rect 28600 845 28650 850
rect 28600 805 28605 845
rect 28645 805 28650 845
rect 28600 800 28650 805
rect -900 700 28800 750
rect -900 645 28800 650
rect -900 605 15705 645
rect 15745 605 16005 645
rect 16045 605 16305 645
rect 16345 605 16605 645
rect 16645 605 16905 645
rect 16945 605 17205 645
rect 17245 605 17505 645
rect 17545 605 17805 645
rect 17845 605 18105 645
rect 18145 605 18405 645
rect 18445 605 18705 645
rect 18745 605 19005 645
rect 19045 605 19305 645
rect 19345 605 19605 645
rect 19645 605 19905 645
rect 19945 605 20205 645
rect 20245 605 24705 645
rect 24745 605 25005 645
rect 25045 605 25305 645
rect 25345 605 25605 645
rect 25645 605 25905 645
rect 25945 605 26205 645
rect 26245 605 26505 645
rect 26545 605 26655 645
rect 26695 605 26805 645
rect 26845 605 27105 645
rect 27145 605 27405 645
rect 27445 605 27705 645
rect 27745 605 28005 645
rect 28045 605 28305 645
rect 28345 605 28605 645
rect 28645 605 28800 645
rect -900 600 28800 605
rect -900 500 28800 550
rect -900 400 24700 450
rect 26550 400 26800 450
rect 28650 400 28800 450
rect -900 300 28800 350
rect -900 200 28800 250
rect -900 100 28800 150
rect -900 40 28800 50
rect -900 10 -640 40
rect -610 10 -40 40
rect -10 10 8360 40
rect 8390 10 10760 40
rect 10790 10 15560 40
rect 15590 10 17960 40
rect 17990 10 20360 40
rect 20390 10 24560 40
rect 24590 10 28760 40
rect 28790 10 28800 40
rect -900 -10 28800 10
rect -900 -40 -640 -10
rect -610 -40 -40 -10
rect -10 -40 8360 -10
rect 8390 -40 10760 -10
rect 10790 -40 15560 -10
rect 15590 -40 17960 -10
rect 17990 -40 20360 -10
rect 20390 -40 24560 -10
rect 24590 -40 28760 -10
rect 28790 -40 28800 -10
rect -900 -60 28800 -40
rect -900 -90 -640 -60
rect -610 -90 -40 -60
rect -10 -90 8360 -60
rect 8390 -90 10760 -60
rect 10790 -90 15560 -60
rect 15590 -90 17960 -60
rect 17990 -90 20360 -60
rect 20390 -90 24560 -60
rect 24590 -90 28760 -60
rect 28790 -90 28800 -60
rect -900 -100 28800 -90
rect -900 -200 28800 -150
rect -900 -300 28800 -250
rect -900 -400 28800 -350
rect -900 -455 28800 -450
rect -900 -495 16755 -455
rect 16795 -495 25755 -455
rect 25795 -495 27555 -455
rect 27595 -495 28800 -455
rect -900 -500 28800 -495
rect -900 -600 28800 -550
rect -900 -700 28800 -650
rect -900 -800 28800 -750
rect -500 -855 -450 -850
rect -500 -895 -495 -855
rect -455 -895 -450 -855
rect -500 -900 -450 -895
rect -350 -855 -300 -850
rect -350 -895 -345 -855
rect -305 -895 -300 -855
rect -350 -900 -300 -895
rect -200 -855 -150 -850
rect -200 -895 -195 -855
rect -155 -895 -150 -855
rect -200 -900 -150 -895
rect 100 -855 150 -850
rect 100 -895 105 -855
rect 145 -895 150 -855
rect 100 -900 150 -895
rect 400 -855 450 -850
rect 400 -895 405 -855
rect 445 -895 450 -855
rect 400 -900 450 -895
rect 700 -855 750 -850
rect 700 -895 705 -855
rect 745 -895 750 -855
rect 700 -900 750 -895
rect 1000 -855 1050 -850
rect 1000 -895 1005 -855
rect 1045 -895 1050 -855
rect 1000 -900 1050 -895
rect 1300 -855 1350 -850
rect 1300 -895 1305 -855
rect 1345 -895 1350 -855
rect 1300 -900 1350 -895
rect 1600 -855 1650 -850
rect 1600 -895 1605 -855
rect 1645 -895 1650 -855
rect 1600 -900 1650 -895
rect 1900 -855 1950 -850
rect 1900 -895 1905 -855
rect 1945 -895 1950 -855
rect 1900 -900 1950 -895
rect 2200 -855 2250 -850
rect 2200 -895 2205 -855
rect 2245 -895 2250 -855
rect 2200 -900 2250 -895
rect 2350 -855 2400 -850
rect 2350 -895 2355 -855
rect 2395 -895 2400 -855
rect 2350 -900 2400 -895
rect 2500 -855 2550 -850
rect 2500 -895 2505 -855
rect 2545 -895 2550 -855
rect 2500 -900 2550 -895
rect 2800 -855 2850 -850
rect 2800 -895 2805 -855
rect 2845 -895 2850 -855
rect 2800 -900 2850 -895
rect 3100 -855 3150 -850
rect 3100 -895 3105 -855
rect 3145 -895 3150 -855
rect 3100 -900 3150 -895
rect 3400 -855 3450 -850
rect 3400 -895 3405 -855
rect 3445 -895 3450 -855
rect 3400 -900 3450 -895
rect 3700 -855 3750 -850
rect 3700 -895 3705 -855
rect 3745 -895 3750 -855
rect 3700 -900 3750 -895
rect 3850 -855 3900 -850
rect 3850 -895 3855 -855
rect 3895 -895 3900 -855
rect 3850 -900 3900 -895
rect 4000 -855 4050 -850
rect 4000 -895 4005 -855
rect 4045 -895 4050 -855
rect 4000 -900 4050 -895
rect 4300 -855 4350 -850
rect 4300 -895 4305 -855
rect 4345 -895 4350 -855
rect 4300 -900 4350 -895
rect 4450 -855 4500 -850
rect 4450 -895 4455 -855
rect 4495 -895 4500 -855
rect 4450 -900 4500 -895
rect 4600 -855 4650 -850
rect 4600 -895 4605 -855
rect 4645 -895 4650 -855
rect 4600 -900 4650 -895
rect 4900 -855 4950 -850
rect 4900 -895 4905 -855
rect 4945 -895 4950 -855
rect 4900 -900 4950 -895
rect 5200 -855 5250 -850
rect 5200 -895 5205 -855
rect 5245 -895 5250 -855
rect 5200 -900 5250 -895
rect 5500 -855 5550 -850
rect 5500 -895 5505 -855
rect 5545 -895 5550 -855
rect 5500 -900 5550 -895
rect 5800 -855 5850 -850
rect 5800 -895 5805 -855
rect 5845 -895 5850 -855
rect 5800 -900 5850 -895
rect 5950 -855 6000 -850
rect 5950 -895 5955 -855
rect 5995 -895 6000 -855
rect 5950 -900 6000 -895
rect 6100 -855 6150 -850
rect 6100 -895 6105 -855
rect 6145 -895 6150 -855
rect 6100 -900 6150 -895
rect 6400 -855 6450 -850
rect 6400 -895 6405 -855
rect 6445 -895 6450 -855
rect 6400 -900 6450 -895
rect 6700 -855 6750 -850
rect 6700 -895 6705 -855
rect 6745 -895 6750 -855
rect 6700 -900 6750 -895
rect 7000 -855 7050 -850
rect 7000 -895 7005 -855
rect 7045 -895 7050 -855
rect 7000 -900 7050 -895
rect 7300 -855 7350 -850
rect 7300 -895 7305 -855
rect 7345 -895 7350 -855
rect 7300 -900 7350 -895
rect 7600 -855 7650 -850
rect 7600 -895 7605 -855
rect 7645 -895 7650 -855
rect 7600 -900 7650 -895
rect 7900 -855 7950 -850
rect 7900 -895 7905 -855
rect 7945 -895 7950 -855
rect 7900 -900 7950 -895
rect 8200 -855 8250 -850
rect 8200 -895 8205 -855
rect 8245 -895 8250 -855
rect 8200 -900 8250 -895
rect 8500 -855 8550 -850
rect 8500 -895 8505 -855
rect 8545 -895 8550 -855
rect 8500 -900 8550 -895
rect 8800 -855 8850 -850
rect 8800 -895 8805 -855
rect 8845 -895 8850 -855
rect 8800 -900 8850 -895
rect 9100 -855 9150 -850
rect 9100 -895 9105 -855
rect 9145 -895 9150 -855
rect 9100 -900 9150 -895
rect 9400 -855 9450 -850
rect 9400 -895 9405 -855
rect 9445 -895 9450 -855
rect 9400 -900 9450 -895
rect 9550 -855 9600 -850
rect 9550 -895 9555 -855
rect 9595 -895 9600 -855
rect 9550 -900 9600 -895
rect 9700 -855 9750 -850
rect 9700 -895 9705 -855
rect 9745 -895 9750 -855
rect 9700 -900 9750 -895
rect 10000 -855 10050 -850
rect 10000 -895 10005 -855
rect 10045 -895 10050 -855
rect 10000 -900 10050 -895
rect 10300 -855 10350 -850
rect 10300 -895 10305 -855
rect 10345 -895 10350 -855
rect 10300 -900 10350 -895
rect 10600 -855 10650 -850
rect 10600 -895 10605 -855
rect 10645 -895 10650 -855
rect 10600 -900 10650 -895
rect 10900 -855 10950 -850
rect 10900 -895 10905 -855
rect 10945 -895 10950 -855
rect 10900 -900 10950 -895
rect 11200 -855 11250 -850
rect 11200 -895 11205 -855
rect 11245 -895 11250 -855
rect 11200 -900 11250 -895
rect 11500 -855 11550 -850
rect 11500 -895 11505 -855
rect 11545 -895 11550 -855
rect 11500 -900 11550 -895
rect 11800 -855 11850 -850
rect 11800 -895 11805 -855
rect 11845 -895 11850 -855
rect 11800 -900 11850 -895
rect 12100 -855 12150 -850
rect 12100 -895 12105 -855
rect 12145 -895 12150 -855
rect 12100 -900 12150 -895
rect 12400 -855 12450 -850
rect 12400 -895 12405 -855
rect 12445 -895 12450 -855
rect 12400 -900 12450 -895
rect 12550 -855 12600 -850
rect 12550 -895 12555 -855
rect 12595 -895 12600 -855
rect 12550 -900 12600 -895
rect 12700 -855 12750 -850
rect 12700 -895 12705 -855
rect 12745 -895 12750 -855
rect 12700 -900 12750 -895
rect 13000 -855 13050 -850
rect 13000 -895 13005 -855
rect 13045 -895 13050 -855
rect 13000 -900 13050 -895
rect 13150 -860 13200 -850
rect 13150 -890 13160 -860
rect 13190 -890 13200 -860
rect 13150 -900 13200 -890
rect 13300 -855 13350 -850
rect 13300 -895 13305 -855
rect 13345 -895 13350 -855
rect 13300 -900 13350 -895
rect 13600 -855 13650 -850
rect 13600 -895 13605 -855
rect 13645 -895 13650 -855
rect 13600 -900 13650 -895
rect 13750 -855 13800 -850
rect 13750 -895 13755 -855
rect 13795 -895 13800 -855
rect 13750 -900 13800 -895
rect 13900 -855 13950 -850
rect 13900 -895 13905 -855
rect 13945 -895 13950 -855
rect 13900 -900 13950 -895
rect 14200 -855 14250 -850
rect 14200 -895 14205 -855
rect 14245 -895 14250 -855
rect 14200 -900 14250 -895
rect 14500 -855 14550 -850
rect 14500 -895 14505 -855
rect 14545 -895 14550 -855
rect 14500 -900 14550 -895
rect 14800 -855 14850 -850
rect 14800 -895 14805 -855
rect 14845 -895 14850 -855
rect 14800 -900 14850 -895
rect 15100 -855 15150 -850
rect 15100 -895 15105 -855
rect 15145 -895 15150 -855
rect 15100 -900 15150 -895
rect 15400 -855 15450 -850
rect 15400 -895 15405 -855
rect 15445 -895 15450 -855
rect 15400 -900 15450 -895
rect 15700 -855 15750 -850
rect 15700 -895 15705 -855
rect 15745 -895 15750 -855
rect 15700 -900 15750 -895
rect 16000 -855 16050 -850
rect 16000 -895 16005 -855
rect 16045 -895 16050 -855
rect 16000 -900 16050 -895
rect 16300 -855 16350 -850
rect 16300 -895 16305 -855
rect 16345 -895 16350 -855
rect 16300 -900 16350 -895
rect 16600 -855 16650 -850
rect 16600 -895 16605 -855
rect 16645 -895 16650 -855
rect 16600 -900 16650 -895
rect 16750 -855 16800 -850
rect 16750 -895 16755 -855
rect 16795 -895 16800 -855
rect 16750 -900 16800 -895
rect 16900 -855 16950 -850
rect 16900 -895 16905 -855
rect 16945 -895 16950 -855
rect 16900 -900 16950 -895
rect 17200 -855 17250 -850
rect 17200 -895 17205 -855
rect 17245 -895 17250 -855
rect 17200 -900 17250 -895
rect 17500 -855 17550 -850
rect 17500 -895 17505 -855
rect 17545 -895 17550 -855
rect 17500 -900 17550 -895
rect 17800 -855 17850 -850
rect 17800 -895 17805 -855
rect 17845 -895 17850 -855
rect 17800 -900 17850 -895
rect 18100 -855 18150 -850
rect 18100 -895 18105 -855
rect 18145 -895 18150 -855
rect 18100 -900 18150 -895
rect 18400 -855 18450 -850
rect 18400 -895 18405 -855
rect 18445 -895 18450 -855
rect 18400 -900 18450 -895
rect 18700 -855 18750 -850
rect 18700 -895 18705 -855
rect 18745 -895 18750 -855
rect 18700 -900 18750 -895
rect 19000 -855 19050 -850
rect 19000 -895 19005 -855
rect 19045 -895 19050 -855
rect 19000 -900 19050 -895
rect 19150 -855 19200 -850
rect 19150 -895 19155 -855
rect 19195 -895 19200 -855
rect 19150 -900 19200 -895
rect 19300 -855 19350 -850
rect 19300 -895 19305 -855
rect 19345 -895 19350 -855
rect 19300 -900 19350 -895
rect 19600 -855 19650 -850
rect 19600 -895 19605 -855
rect 19645 -895 19650 -855
rect 19600 -900 19650 -895
rect 19900 -855 19950 -850
rect 19900 -895 19905 -855
rect 19945 -895 19950 -855
rect 19900 -900 19950 -895
rect 20200 -855 20250 -850
rect 20200 -895 20205 -855
rect 20245 -895 20250 -855
rect 20200 -900 20250 -895
rect 20500 -855 20550 -850
rect 20500 -895 20505 -855
rect 20545 -895 20550 -855
rect 20500 -900 20550 -895
rect 20800 -855 20850 -850
rect 20800 -895 20805 -855
rect 20845 -895 20850 -855
rect 20800 -900 20850 -895
rect 21100 -855 21150 -850
rect 21100 -895 21105 -855
rect 21145 -895 21150 -855
rect 21100 -900 21150 -895
rect 21400 -855 21450 -850
rect 21400 -895 21405 -855
rect 21445 -895 21450 -855
rect 21400 -900 21450 -895
rect 21700 -855 21750 -850
rect 21700 -895 21705 -855
rect 21745 -895 21750 -855
rect 21700 -900 21750 -895
rect 22000 -855 22050 -850
rect 22000 -895 22005 -855
rect 22045 -895 22050 -855
rect 22000 -900 22050 -895
rect 22300 -855 22350 -850
rect 22300 -895 22305 -855
rect 22345 -895 22350 -855
rect 22300 -900 22350 -895
rect 22450 -855 22500 -850
rect 22450 -895 22455 -855
rect 22495 -895 22500 -855
rect 22450 -900 22500 -895
rect 22600 -855 22650 -850
rect 22600 -895 22605 -855
rect 22645 -895 22650 -855
rect 22600 -900 22650 -895
rect 22900 -855 22950 -850
rect 22900 -895 22905 -855
rect 22945 -895 22950 -855
rect 22900 -900 22950 -895
rect 23200 -855 23250 -850
rect 23200 -895 23205 -855
rect 23245 -895 23250 -855
rect 23200 -900 23250 -895
rect 23500 -855 23550 -850
rect 23500 -895 23505 -855
rect 23545 -895 23550 -855
rect 23500 -900 23550 -895
rect 23800 -855 23850 -850
rect 23800 -895 23805 -855
rect 23845 -895 23850 -855
rect 23800 -900 23850 -895
rect 24100 -855 24150 -850
rect 24100 -895 24105 -855
rect 24145 -895 24150 -855
rect 24100 -900 24150 -895
rect 24400 -855 24450 -850
rect 24400 -895 24405 -855
rect 24445 -895 24450 -855
rect 24400 -900 24450 -895
rect 24700 -855 24750 -850
rect 24700 -895 24705 -855
rect 24745 -895 24750 -855
rect 24700 -900 24750 -895
rect 25000 -855 25050 -850
rect 25000 -895 25005 -855
rect 25045 -895 25050 -855
rect 25000 -900 25050 -895
rect 25300 -855 25350 -850
rect 25300 -895 25305 -855
rect 25345 -895 25350 -855
rect 25300 -900 25350 -895
rect 25600 -855 25650 -850
rect 25600 -895 25605 -855
rect 25645 -895 25650 -855
rect 25600 -900 25650 -895
rect 25750 -855 25800 -850
rect 25750 -895 25755 -855
rect 25795 -895 25800 -855
rect 25750 -900 25800 -895
rect 25900 -855 25950 -850
rect 25900 -895 25905 -855
rect 25945 -895 25950 -855
rect 25900 -900 25950 -895
rect 26200 -855 26250 -850
rect 26200 -895 26205 -855
rect 26245 -895 26250 -855
rect 26200 -900 26250 -895
rect 26500 -855 26550 -850
rect 26500 -895 26505 -855
rect 26545 -895 26550 -855
rect 26500 -900 26550 -895
rect 26650 -855 26700 -850
rect 26650 -895 26655 -855
rect 26695 -895 26700 -855
rect 26650 -900 26700 -895
rect 26800 -855 26850 -850
rect 26800 -895 26805 -855
rect 26845 -895 26850 -855
rect 26800 -900 26850 -895
rect 27100 -855 27150 -850
rect 27100 -895 27105 -855
rect 27145 -895 27150 -855
rect 27100 -900 27150 -895
rect 27400 -855 27450 -850
rect 27400 -895 27405 -855
rect 27445 -895 27450 -855
rect 27400 -900 27450 -895
rect 27550 -855 27600 -850
rect 27550 -895 27555 -855
rect 27595 -895 27600 -855
rect 27550 -900 27600 -895
rect 27700 -855 27750 -850
rect 27700 -895 27705 -855
rect 27745 -895 27750 -855
rect 27700 -900 27750 -895
rect 28000 -855 28050 -850
rect 28000 -895 28005 -855
rect 28045 -895 28050 -855
rect 28000 -900 28050 -895
rect 28300 -855 28350 -850
rect 28300 -895 28305 -855
rect 28345 -895 28350 -855
rect 28300 -900 28350 -895
rect 28600 -855 28650 -850
rect 28600 -895 28605 -855
rect 28645 -895 28650 -855
rect 28600 -900 28650 -895
rect -900 -1000 28800 -950
rect -900 -1100 28800 -1050
rect -900 -1200 28800 -1150
rect -900 -1300 28800 -1250
rect -900 -1400 28800 -1350
rect -900 -1500 28800 -1450
rect -900 -1600 28800 -1550
rect -900 -1660 28800 -1650
rect -900 -1690 -640 -1660
rect -610 -1690 -40 -1660
rect -10 -1690 8360 -1660
rect 8390 -1690 10760 -1660
rect 10790 -1690 15560 -1660
rect 15590 -1690 17960 -1660
rect 17990 -1690 20360 -1660
rect 20390 -1690 24560 -1660
rect 24590 -1690 28760 -1660
rect 28790 -1690 28800 -1660
rect -900 -1710 28800 -1690
rect -900 -1740 -640 -1710
rect -610 -1740 -40 -1710
rect -10 -1740 8360 -1710
rect 8390 -1740 10760 -1710
rect 10790 -1740 15560 -1710
rect 15590 -1740 17960 -1710
rect 17990 -1740 20360 -1710
rect 20390 -1740 24560 -1710
rect 24590 -1740 28760 -1710
rect 28790 -1740 28800 -1710
rect -900 -1750 28800 -1740
<< via3 >>
rect -495 4940 -455 4945
rect -495 4910 -490 4940
rect -490 4910 -460 4940
rect -460 4910 -455 4940
rect -495 4905 -455 4910
rect -345 4940 -305 4945
rect -345 4910 -340 4940
rect -340 4910 -310 4940
rect -310 4910 -305 4940
rect -345 4905 -305 4910
rect -195 4940 -155 4945
rect -195 4910 -190 4940
rect -190 4910 -160 4940
rect -160 4910 -155 4940
rect -195 4905 -155 4910
rect 105 4940 145 4945
rect 105 4910 110 4940
rect 110 4910 140 4940
rect 140 4910 145 4940
rect 105 4905 145 4910
rect 405 4940 445 4945
rect 405 4910 410 4940
rect 410 4910 440 4940
rect 440 4910 445 4940
rect 405 4905 445 4910
rect 705 4940 745 4945
rect 705 4910 710 4940
rect 710 4910 740 4940
rect 740 4910 745 4940
rect 705 4905 745 4910
rect 1005 4940 1045 4945
rect 1005 4910 1010 4940
rect 1010 4910 1040 4940
rect 1040 4910 1045 4940
rect 1005 4905 1045 4910
rect 1155 4940 1195 4945
rect 1155 4910 1160 4940
rect 1160 4910 1190 4940
rect 1190 4910 1195 4940
rect 1155 4905 1195 4910
rect 1305 4940 1345 4945
rect 1305 4910 1310 4940
rect 1310 4910 1340 4940
rect 1340 4910 1345 4940
rect 1305 4905 1345 4910
rect 1605 4940 1645 4945
rect 1605 4910 1610 4940
rect 1610 4910 1640 4940
rect 1640 4910 1645 4940
rect 1605 4905 1645 4910
rect 1905 4940 1945 4945
rect 1905 4910 1910 4940
rect 1910 4910 1940 4940
rect 1940 4910 1945 4940
rect 1905 4905 1945 4910
rect 2055 4940 2095 4945
rect 2055 4910 2060 4940
rect 2060 4910 2090 4940
rect 2090 4910 2095 4940
rect 2055 4905 2095 4910
rect 2205 4940 2245 4945
rect 2205 4910 2210 4940
rect 2210 4910 2240 4940
rect 2240 4910 2245 4940
rect 2205 4905 2245 4910
rect 2505 4940 2545 4945
rect 2505 4910 2510 4940
rect 2510 4910 2540 4940
rect 2540 4910 2545 4940
rect 2505 4905 2545 4910
rect 2805 4940 2845 4945
rect 2805 4910 2810 4940
rect 2810 4910 2840 4940
rect 2840 4910 2845 4940
rect 2805 4905 2845 4910
rect 2955 4940 2995 4945
rect 2955 4910 2960 4940
rect 2960 4910 2990 4940
rect 2990 4910 2995 4940
rect 2955 4905 2995 4910
rect 3105 4940 3145 4945
rect 3105 4910 3110 4940
rect 3110 4910 3140 4940
rect 3140 4910 3145 4940
rect 3105 4905 3145 4910
rect 3405 4940 3445 4945
rect 3405 4910 3410 4940
rect 3410 4910 3440 4940
rect 3440 4910 3445 4940
rect 3405 4905 3445 4910
rect 3705 4940 3745 4945
rect 3705 4910 3710 4940
rect 3710 4910 3740 4940
rect 3740 4910 3745 4940
rect 3705 4905 3745 4910
rect 4005 4940 4045 4945
rect 4005 4910 4010 4940
rect 4010 4910 4040 4940
rect 4040 4910 4045 4940
rect 4005 4905 4045 4910
rect 4305 4940 4345 4945
rect 4305 4910 4310 4940
rect 4310 4910 4340 4940
rect 4340 4910 4345 4940
rect 4305 4905 4345 4910
rect 4605 4940 4645 4945
rect 4605 4910 4610 4940
rect 4610 4910 4640 4940
rect 4640 4910 4645 4940
rect 4605 4905 4645 4910
rect 4905 4940 4945 4945
rect 4905 4910 4910 4940
rect 4910 4910 4940 4940
rect 4940 4910 4945 4940
rect 4905 4905 4945 4910
rect 5205 4940 5245 4945
rect 5205 4910 5210 4940
rect 5210 4910 5240 4940
rect 5240 4910 5245 4940
rect 5205 4905 5245 4910
rect 5355 4940 5395 4945
rect 5355 4910 5360 4940
rect 5360 4910 5390 4940
rect 5390 4910 5395 4940
rect 5355 4905 5395 4910
rect 5505 4940 5545 4945
rect 5505 4910 5510 4940
rect 5510 4910 5540 4940
rect 5540 4910 5545 4940
rect 5505 4905 5545 4910
rect 5805 4940 5845 4945
rect 5805 4910 5810 4940
rect 5810 4910 5840 4940
rect 5840 4910 5845 4940
rect 5805 4905 5845 4910
rect 6105 4940 6145 4945
rect 6105 4910 6110 4940
rect 6110 4910 6140 4940
rect 6140 4910 6145 4940
rect 6105 4905 6145 4910
rect 6255 4940 6295 4945
rect 6255 4910 6260 4940
rect 6260 4910 6290 4940
rect 6290 4910 6295 4940
rect 6255 4905 6295 4910
rect 6405 4940 6445 4945
rect 6405 4910 6410 4940
rect 6410 4910 6440 4940
rect 6440 4910 6445 4940
rect 6405 4905 6445 4910
rect 6705 4940 6745 4945
rect 6705 4910 6710 4940
rect 6710 4910 6740 4940
rect 6740 4910 6745 4940
rect 6705 4905 6745 4910
rect 7005 4940 7045 4945
rect 7005 4910 7010 4940
rect 7010 4910 7040 4940
rect 7040 4910 7045 4940
rect 7005 4905 7045 4910
rect 7155 4940 7195 4945
rect 7155 4910 7160 4940
rect 7160 4910 7190 4940
rect 7190 4910 7195 4940
rect 7155 4905 7195 4910
rect 7305 4940 7345 4945
rect 7305 4910 7310 4940
rect 7310 4910 7340 4940
rect 7340 4910 7345 4940
rect 7305 4905 7345 4910
rect 7605 4940 7645 4945
rect 7605 4910 7610 4940
rect 7610 4910 7640 4940
rect 7640 4910 7645 4940
rect 7605 4905 7645 4910
rect 7905 4940 7945 4945
rect 7905 4910 7910 4940
rect 7910 4910 7940 4940
rect 7940 4910 7945 4940
rect 7905 4905 7945 4910
rect 8205 4940 8245 4945
rect 8205 4910 8210 4940
rect 8210 4910 8240 4940
rect 8240 4910 8245 4940
rect 8205 4905 8245 4910
rect 8505 4940 8545 4945
rect 8505 4910 8510 4940
rect 8510 4910 8540 4940
rect 8540 4910 8545 4940
rect 8505 4905 8545 4910
rect 8805 4940 8845 4945
rect 8805 4910 8810 4940
rect 8810 4910 8840 4940
rect 8840 4910 8845 4940
rect 8805 4905 8845 4910
rect 9105 4940 9145 4945
rect 9105 4910 9110 4940
rect 9110 4910 9140 4940
rect 9140 4910 9145 4940
rect 9105 4905 9145 4910
rect 9405 4940 9445 4945
rect 9405 4910 9410 4940
rect 9410 4910 9440 4940
rect 9440 4910 9445 4940
rect 9405 4905 9445 4910
rect 9705 4940 9745 4945
rect 9705 4910 9710 4940
rect 9710 4910 9740 4940
rect 9740 4910 9745 4940
rect 9705 4905 9745 4910
rect 10005 4940 10045 4945
rect 10005 4910 10010 4940
rect 10010 4910 10040 4940
rect 10040 4910 10045 4940
rect 10005 4905 10045 4910
rect 10305 4940 10345 4945
rect 10305 4910 10310 4940
rect 10310 4910 10340 4940
rect 10340 4910 10345 4940
rect 10305 4905 10345 4910
rect 10605 4940 10645 4945
rect 10605 4910 10610 4940
rect 10610 4910 10640 4940
rect 10640 4910 10645 4940
rect 10605 4905 10645 4910
rect 10905 4940 10945 4945
rect 10905 4910 10910 4940
rect 10910 4910 10940 4940
rect 10940 4910 10945 4940
rect 10905 4905 10945 4910
rect 11205 4940 11245 4945
rect 11205 4910 11210 4940
rect 11210 4910 11240 4940
rect 11240 4910 11245 4940
rect 11205 4905 11245 4910
rect 11355 4940 11395 4945
rect 11355 4910 11360 4940
rect 11360 4910 11390 4940
rect 11390 4910 11395 4940
rect 11355 4905 11395 4910
rect 11505 4940 11545 4945
rect 11505 4910 11510 4940
rect 11510 4910 11540 4940
rect 11540 4910 11545 4940
rect 11505 4905 11545 4910
rect 11805 4940 11845 4945
rect 11805 4910 11810 4940
rect 11810 4910 11840 4940
rect 11840 4910 11845 4940
rect 11805 4905 11845 4910
rect 12105 4940 12145 4945
rect 12105 4910 12110 4940
rect 12110 4910 12140 4940
rect 12140 4910 12145 4940
rect 12105 4905 12145 4910
rect 12405 4940 12445 4945
rect 12405 4910 12410 4940
rect 12410 4910 12440 4940
rect 12440 4910 12445 4940
rect 12405 4905 12445 4910
rect 12555 4940 12595 4945
rect 12555 4910 12560 4940
rect 12560 4910 12590 4940
rect 12590 4910 12595 4940
rect 12555 4905 12595 4910
rect 12705 4940 12745 4945
rect 12705 4910 12710 4940
rect 12710 4910 12740 4940
rect 12740 4910 12745 4940
rect 12705 4905 12745 4910
rect 13005 4940 13045 4945
rect 13005 4910 13010 4940
rect 13010 4910 13040 4940
rect 13040 4910 13045 4940
rect 13005 4905 13045 4910
rect 13305 4940 13345 4945
rect 13305 4910 13310 4940
rect 13310 4910 13340 4940
rect 13340 4910 13345 4940
rect 13305 4905 13345 4910
rect 13605 4940 13645 4945
rect 13605 4910 13610 4940
rect 13610 4910 13640 4940
rect 13640 4910 13645 4940
rect 13605 4905 13645 4910
rect 13755 4940 13795 4945
rect 13755 4910 13760 4940
rect 13760 4910 13790 4940
rect 13790 4910 13795 4940
rect 13755 4905 13795 4910
rect 13905 4940 13945 4945
rect 13905 4910 13910 4940
rect 13910 4910 13940 4940
rect 13940 4910 13945 4940
rect 13905 4905 13945 4910
rect 14205 4940 14245 4945
rect 14205 4910 14210 4940
rect 14210 4910 14240 4940
rect 14240 4910 14245 4940
rect 14205 4905 14245 4910
rect 14505 4940 14545 4945
rect 14505 4910 14510 4940
rect 14510 4910 14540 4940
rect 14540 4910 14545 4940
rect 14505 4905 14545 4910
rect 14805 4940 14845 4945
rect 14805 4910 14810 4940
rect 14810 4910 14840 4940
rect 14840 4910 14845 4940
rect 14805 4905 14845 4910
rect 14955 4940 14995 4945
rect 14955 4910 14960 4940
rect 14960 4910 14990 4940
rect 14990 4910 14995 4940
rect 14955 4905 14995 4910
rect 15105 4940 15145 4945
rect 15105 4910 15110 4940
rect 15110 4910 15140 4940
rect 15140 4910 15145 4940
rect 15105 4905 15145 4910
rect 15405 4940 15445 4945
rect 15405 4910 15410 4940
rect 15410 4910 15440 4940
rect 15440 4910 15445 4940
rect 15405 4905 15445 4910
rect 15705 4940 15745 4945
rect 15705 4910 15710 4940
rect 15710 4910 15740 4940
rect 15740 4910 15745 4940
rect 15705 4905 15745 4910
rect 16005 4940 16045 4945
rect 16005 4910 16010 4940
rect 16010 4910 16040 4940
rect 16040 4910 16045 4940
rect 16005 4905 16045 4910
rect 16305 4940 16345 4945
rect 16305 4910 16310 4940
rect 16310 4910 16340 4940
rect 16340 4910 16345 4940
rect 16305 4905 16345 4910
rect 16605 4940 16645 4945
rect 16605 4910 16610 4940
rect 16610 4910 16640 4940
rect 16640 4910 16645 4940
rect 16605 4905 16645 4910
rect 16755 4940 16795 4945
rect 16755 4910 16760 4940
rect 16760 4910 16790 4940
rect 16790 4910 16795 4940
rect 16755 4905 16795 4910
rect 16905 4940 16945 4945
rect 16905 4910 16910 4940
rect 16910 4910 16940 4940
rect 16940 4910 16945 4940
rect 16905 4905 16945 4910
rect 17205 4940 17245 4945
rect 17205 4910 17210 4940
rect 17210 4910 17240 4940
rect 17240 4910 17245 4940
rect 17205 4905 17245 4910
rect 17505 4940 17545 4945
rect 17505 4910 17510 4940
rect 17510 4910 17540 4940
rect 17540 4910 17545 4940
rect 17505 4905 17545 4910
rect 17805 4940 17845 4945
rect 17805 4910 17810 4940
rect 17810 4910 17840 4940
rect 17840 4910 17845 4940
rect 17805 4905 17845 4910
rect 18105 4940 18145 4945
rect 18105 4910 18110 4940
rect 18110 4910 18140 4940
rect 18140 4910 18145 4940
rect 18105 4905 18145 4910
rect 18405 4940 18445 4945
rect 18405 4910 18410 4940
rect 18410 4910 18440 4940
rect 18440 4910 18445 4940
rect 18405 4905 18445 4910
rect 18705 4940 18745 4945
rect 18705 4910 18710 4940
rect 18710 4910 18740 4940
rect 18740 4910 18745 4940
rect 18705 4905 18745 4910
rect 19005 4940 19045 4945
rect 19005 4910 19010 4940
rect 19010 4910 19040 4940
rect 19040 4910 19045 4940
rect 19005 4905 19045 4910
rect 19155 4940 19195 4945
rect 19155 4910 19160 4940
rect 19160 4910 19190 4940
rect 19190 4910 19195 4940
rect 19155 4905 19195 4910
rect 19305 4940 19345 4945
rect 19305 4910 19310 4940
rect 19310 4910 19340 4940
rect 19340 4910 19345 4940
rect 19305 4905 19345 4910
rect 19605 4940 19645 4945
rect 19605 4910 19610 4940
rect 19610 4910 19640 4940
rect 19640 4910 19645 4940
rect 19605 4905 19645 4910
rect 19905 4940 19945 4945
rect 19905 4910 19910 4940
rect 19910 4910 19940 4940
rect 19940 4910 19945 4940
rect 19905 4905 19945 4910
rect 20205 4940 20245 4945
rect 20205 4910 20210 4940
rect 20210 4910 20240 4940
rect 20240 4910 20245 4940
rect 20205 4905 20245 4910
rect 20505 4940 20545 4945
rect 20505 4910 20510 4940
rect 20510 4910 20540 4940
rect 20540 4910 20545 4940
rect 20505 4905 20545 4910
rect 20805 4940 20845 4945
rect 20805 4910 20810 4940
rect 20810 4910 20840 4940
rect 20840 4910 20845 4940
rect 20805 4905 20845 4910
rect 20955 4940 20995 4945
rect 20955 4910 20960 4940
rect 20960 4910 20990 4940
rect 20990 4910 20995 4940
rect 20955 4905 20995 4910
rect 21105 4940 21145 4945
rect 21105 4910 21110 4940
rect 21110 4910 21140 4940
rect 21140 4910 21145 4940
rect 21105 4905 21145 4910
rect 21705 4940 21745 4945
rect 21705 4910 21710 4940
rect 21710 4910 21740 4940
rect 21740 4910 21745 4940
rect 21705 4905 21745 4910
rect 21855 4940 21895 4945
rect 21855 4910 21860 4940
rect 21860 4910 21890 4940
rect 21890 4910 21895 4940
rect 21855 4905 21895 4910
rect 22005 4940 22045 4945
rect 22005 4910 22010 4940
rect 22010 4910 22040 4940
rect 22040 4910 22045 4940
rect 22005 4905 22045 4910
rect 22305 4940 22345 4945
rect 22305 4910 22310 4940
rect 22310 4910 22340 4940
rect 22340 4910 22345 4940
rect 22305 4905 22345 4910
rect 22605 4940 22645 4945
rect 22605 4910 22610 4940
rect 22610 4910 22640 4940
rect 22640 4910 22645 4940
rect 22605 4905 22645 4910
rect 22905 4940 22945 4945
rect 22905 4910 22910 4940
rect 22910 4910 22940 4940
rect 22940 4910 22945 4940
rect 22905 4905 22945 4910
rect 23055 4940 23095 4945
rect 23055 4910 23060 4940
rect 23060 4910 23090 4940
rect 23090 4910 23095 4940
rect 23055 4905 23095 4910
rect 23205 4940 23245 4945
rect 23205 4910 23210 4940
rect 23210 4910 23240 4940
rect 23240 4910 23245 4940
rect 23205 4905 23245 4910
rect 23355 4940 23395 4945
rect 23355 4910 23360 4940
rect 23360 4910 23390 4940
rect 23390 4910 23395 4940
rect 23355 4905 23395 4910
rect 23655 4940 23695 4945
rect 23655 4910 23660 4940
rect 23660 4910 23690 4940
rect 23690 4910 23695 4940
rect 23655 4905 23695 4910
rect 23805 4940 23845 4945
rect 23805 4910 23810 4940
rect 23810 4910 23840 4940
rect 23840 4910 23845 4940
rect 23805 4905 23845 4910
rect 23955 4940 23995 4945
rect 23955 4910 23960 4940
rect 23960 4910 23990 4940
rect 23990 4910 23995 4940
rect 23955 4905 23995 4910
rect 24105 4940 24145 4945
rect 24105 4910 24110 4940
rect 24110 4910 24140 4940
rect 24140 4910 24145 4940
rect 24105 4905 24145 4910
rect 24405 4940 24445 4945
rect 24405 4910 24410 4940
rect 24410 4910 24440 4940
rect 24440 4910 24445 4940
rect 24405 4905 24445 4910
rect 24705 4940 24745 4945
rect 24705 4910 24710 4940
rect 24710 4910 24740 4940
rect 24740 4910 24745 4940
rect 24705 4905 24745 4910
rect 25005 4940 25045 4945
rect 25005 4910 25010 4940
rect 25010 4910 25040 4940
rect 25040 4910 25045 4940
rect 25005 4905 25045 4910
rect 25455 4940 25495 4945
rect 25455 4910 25460 4940
rect 25460 4910 25490 4940
rect 25490 4910 25495 4940
rect 25455 4905 25495 4910
rect 25605 4940 25645 4945
rect 25605 4910 25610 4940
rect 25610 4910 25640 4940
rect 25640 4910 25645 4940
rect 25605 4905 25645 4910
rect 25755 4940 25795 4945
rect 25755 4910 25760 4940
rect 25760 4910 25790 4940
rect 25790 4910 25795 4940
rect 25755 4905 25795 4910
rect 26205 4940 26245 4945
rect 26205 4910 26210 4940
rect 26210 4910 26240 4940
rect 26240 4910 26245 4940
rect 26205 4905 26245 4910
rect 26505 4940 26545 4945
rect 26505 4910 26510 4940
rect 26510 4910 26540 4940
rect 26540 4910 26545 4940
rect 26505 4905 26545 4910
rect 26805 4940 26845 4945
rect 26805 4910 26810 4940
rect 26810 4910 26840 4940
rect 26840 4910 26845 4940
rect 26805 4905 26845 4910
rect 27105 4940 27145 4945
rect 27105 4910 27110 4940
rect 27110 4910 27140 4940
rect 27140 4910 27145 4940
rect 27105 4905 27145 4910
rect 27555 4940 27595 4945
rect 27555 4910 27560 4940
rect 27560 4910 27590 4940
rect 27590 4910 27595 4940
rect 27555 4905 27595 4910
rect 27705 4940 27745 4945
rect 27705 4910 27710 4940
rect 27710 4910 27740 4940
rect 27740 4910 27745 4940
rect 27705 4905 27745 4910
rect 27855 4940 27895 4945
rect 27855 4910 27860 4940
rect 27860 4910 27890 4940
rect 27890 4910 27895 4940
rect 27855 4905 27895 4910
rect 28305 4940 28345 4945
rect 28305 4910 28310 4940
rect 28310 4910 28340 4940
rect 28340 4910 28345 4940
rect 28305 4905 28345 4910
rect 28605 4940 28645 4945
rect 28605 4910 28610 4940
rect 28610 4910 28640 4940
rect 28640 4910 28645 4940
rect 28605 4905 28645 4910
rect 28755 4940 28795 4945
rect 28755 4910 28760 4940
rect 28760 4910 28790 4940
rect 28790 4910 28795 4940
rect 28755 4905 28795 4910
rect 28905 4940 28945 4945
rect 28905 4910 28910 4940
rect 28910 4910 28940 4940
rect 28940 4910 28945 4940
rect 28905 4905 28945 4910
rect 29205 4940 29245 4945
rect 29205 4910 29210 4940
rect 29210 4910 29240 4940
rect 29240 4910 29245 4940
rect 29205 4905 29245 4910
rect 29355 4940 29395 4945
rect 29355 4910 29360 4940
rect 29360 4910 29390 4940
rect 29390 4910 29395 4940
rect 29355 4905 29395 4910
rect 29655 4940 29695 4945
rect 29655 4910 29660 4940
rect 29660 4910 29690 4940
rect 29690 4910 29695 4940
rect 29655 4905 29695 4910
rect 29955 4940 29995 4945
rect 29955 4910 29960 4940
rect 29960 4910 29990 4940
rect 29990 4910 29995 4940
rect 29955 4905 29995 4910
rect 30255 4940 30295 4945
rect 30255 4910 30260 4940
rect 30260 4910 30290 4940
rect 30290 4910 30295 4940
rect 30255 4905 30295 4910
rect 30555 4940 30595 4945
rect 30555 4910 30560 4940
rect 30560 4910 30590 4940
rect 30590 4910 30595 4940
rect 30555 4905 30595 4910
rect 30855 4940 30895 4945
rect 30855 4910 30860 4940
rect 30860 4910 30890 4940
rect 30890 4910 30895 4940
rect 30855 4905 30895 4910
rect 31005 4940 31045 4945
rect 31005 4910 31010 4940
rect 31010 4910 31040 4940
rect 31040 4910 31045 4940
rect 31005 4905 31045 4910
rect 31455 4940 31495 4945
rect 31455 4910 31460 4940
rect 31460 4910 31490 4940
rect 31490 4910 31495 4940
rect 31455 4905 31495 4910
rect 31605 4940 31645 4945
rect 31605 4910 31610 4940
rect 31610 4910 31640 4940
rect 31640 4910 31645 4940
rect 31605 4905 31645 4910
rect 31905 4940 31945 4945
rect 31905 4910 31910 4940
rect 31910 4910 31940 4940
rect 31940 4910 31945 4940
rect 31905 4905 31945 4910
rect 32055 4940 32095 4945
rect 32055 4910 32060 4940
rect 32060 4910 32090 4940
rect 32090 4910 32095 4940
rect 32055 4905 32095 4910
rect 13755 4705 13795 4745
rect 14955 4705 14995 4745
rect 29355 4705 29395 4745
rect 31455 4705 31495 4745
rect 11355 4505 11395 4545
rect 12555 4505 12595 4545
rect 20955 4505 20995 4545
rect 21855 4505 21895 4545
rect 23055 4505 23095 4545
rect 23955 4505 23995 4545
rect 28755 4505 28795 4545
rect 32055 4505 32095 4545
rect 31005 4005 31045 4045
rect 10905 3805 10945 3845
rect 11205 3805 11245 3845
rect 11505 3805 11545 3845
rect 11805 3805 11845 3845
rect 12105 3805 12145 3845
rect 12405 3805 12445 3845
rect 12705 3805 12745 3845
rect 13005 3805 13045 3845
rect 13305 3805 13345 3845
rect 13605 3805 13645 3845
rect 13905 3805 13945 3845
rect 14205 3805 14245 3845
rect 14505 3805 14545 3845
rect 14805 3805 14845 3845
rect 20505 3805 20545 3845
rect 20805 3805 20845 3845
rect 21105 3805 21145 3845
rect 21405 3805 21445 3845
rect 21705 3805 21745 3845
rect 22005 3805 22045 3845
rect 22305 3805 22345 3845
rect 22455 3805 22495 3845
rect 22605 3805 22645 3845
rect 22905 3805 22945 3845
rect 23205 3805 23245 3845
rect 23505 3805 23545 3845
rect 23805 3805 23845 3845
rect 24105 3805 24145 3845
rect 24405 3805 24445 3845
rect 28305 3805 28345 3845
rect 28605 3805 28645 3845
rect 28905 3805 28945 3845
rect 29205 3805 29245 3845
rect 29655 3805 29695 3845
rect 31605 3805 31645 3845
rect 31905 3805 31945 3845
rect -495 3640 -455 3645
rect -495 3610 -490 3640
rect -490 3610 -460 3640
rect -460 3610 -455 3640
rect -495 3605 -455 3610
rect -345 3640 -305 3645
rect -345 3610 -340 3640
rect -340 3610 -310 3640
rect -310 3610 -305 3640
rect -345 3605 -305 3610
rect -195 3640 -155 3645
rect -195 3610 -190 3640
rect -190 3610 -160 3640
rect -160 3610 -155 3640
rect -195 3605 -155 3610
rect 105 3640 145 3645
rect 105 3610 110 3640
rect 110 3610 140 3640
rect 140 3610 145 3640
rect 105 3605 145 3610
rect 405 3640 445 3645
rect 405 3610 410 3640
rect 410 3610 440 3640
rect 440 3610 445 3640
rect 405 3605 445 3610
rect 705 3640 745 3645
rect 705 3610 710 3640
rect 710 3610 740 3640
rect 740 3610 745 3640
rect 705 3605 745 3610
rect 1005 3640 1045 3645
rect 1005 3610 1010 3640
rect 1010 3610 1040 3640
rect 1040 3610 1045 3640
rect 1005 3605 1045 3610
rect 1155 3640 1195 3645
rect 1155 3610 1160 3640
rect 1160 3610 1190 3640
rect 1190 3610 1195 3640
rect 1155 3605 1195 3610
rect 1305 3640 1345 3645
rect 1305 3610 1310 3640
rect 1310 3610 1340 3640
rect 1340 3610 1345 3640
rect 1305 3605 1345 3610
rect 1605 3640 1645 3645
rect 1605 3610 1610 3640
rect 1610 3610 1640 3640
rect 1640 3610 1645 3640
rect 1605 3605 1645 3610
rect 1905 3640 1945 3645
rect 1905 3610 1910 3640
rect 1910 3610 1940 3640
rect 1940 3610 1945 3640
rect 1905 3605 1945 3610
rect 2055 3640 2095 3645
rect 2055 3610 2060 3640
rect 2060 3610 2090 3640
rect 2090 3610 2095 3640
rect 2055 3605 2095 3610
rect 2205 3640 2245 3645
rect 2205 3610 2210 3640
rect 2210 3610 2240 3640
rect 2240 3610 2245 3640
rect 2205 3605 2245 3610
rect 2505 3640 2545 3645
rect 2505 3610 2510 3640
rect 2510 3610 2540 3640
rect 2540 3610 2545 3640
rect 2505 3605 2545 3610
rect 2805 3640 2845 3645
rect 2805 3610 2810 3640
rect 2810 3610 2840 3640
rect 2840 3610 2845 3640
rect 2805 3605 2845 3610
rect 2955 3640 2995 3645
rect 2955 3610 2960 3640
rect 2960 3610 2990 3640
rect 2990 3610 2995 3640
rect 2955 3605 2995 3610
rect 3105 3640 3145 3645
rect 3105 3610 3110 3640
rect 3110 3610 3140 3640
rect 3140 3610 3145 3640
rect 3105 3605 3145 3610
rect 3405 3640 3445 3645
rect 3405 3610 3410 3640
rect 3410 3610 3440 3640
rect 3440 3610 3445 3640
rect 3405 3605 3445 3610
rect 3705 3640 3745 3645
rect 3705 3610 3710 3640
rect 3710 3610 3740 3640
rect 3740 3610 3745 3640
rect 3705 3605 3745 3610
rect 4005 3640 4045 3645
rect 4005 3610 4010 3640
rect 4010 3610 4040 3640
rect 4040 3610 4045 3640
rect 4005 3605 4045 3610
rect 4305 3640 4345 3645
rect 4305 3610 4310 3640
rect 4310 3610 4340 3640
rect 4340 3610 4345 3640
rect 4305 3605 4345 3610
rect 4605 3640 4645 3645
rect 4605 3610 4610 3640
rect 4610 3610 4640 3640
rect 4640 3610 4645 3640
rect 4605 3605 4645 3610
rect 4905 3640 4945 3645
rect 4905 3610 4910 3640
rect 4910 3610 4940 3640
rect 4940 3610 4945 3640
rect 4905 3605 4945 3610
rect 5205 3640 5245 3645
rect 5205 3610 5210 3640
rect 5210 3610 5240 3640
rect 5240 3610 5245 3640
rect 5205 3605 5245 3610
rect 5355 3640 5395 3645
rect 5355 3610 5360 3640
rect 5360 3610 5390 3640
rect 5390 3610 5395 3640
rect 5355 3605 5395 3610
rect 5505 3640 5545 3645
rect 5505 3610 5510 3640
rect 5510 3610 5540 3640
rect 5540 3610 5545 3640
rect 5505 3605 5545 3610
rect 5805 3640 5845 3645
rect 5805 3610 5810 3640
rect 5810 3610 5840 3640
rect 5840 3610 5845 3640
rect 5805 3605 5845 3610
rect 6105 3640 6145 3645
rect 6105 3610 6110 3640
rect 6110 3610 6140 3640
rect 6140 3610 6145 3640
rect 6105 3605 6145 3610
rect 6255 3640 6295 3645
rect 6255 3610 6260 3640
rect 6260 3610 6290 3640
rect 6290 3610 6295 3640
rect 6255 3605 6295 3610
rect 6405 3640 6445 3645
rect 6405 3610 6410 3640
rect 6410 3610 6440 3640
rect 6440 3610 6445 3640
rect 6405 3605 6445 3610
rect 6705 3640 6745 3645
rect 6705 3610 6710 3640
rect 6710 3610 6740 3640
rect 6740 3610 6745 3640
rect 6705 3605 6745 3610
rect 7005 3640 7045 3645
rect 7005 3610 7010 3640
rect 7010 3610 7040 3640
rect 7040 3610 7045 3640
rect 7005 3605 7045 3610
rect 7155 3640 7195 3645
rect 7155 3610 7160 3640
rect 7160 3610 7190 3640
rect 7190 3610 7195 3640
rect 7155 3605 7195 3610
rect 7305 3640 7345 3645
rect 7305 3610 7310 3640
rect 7310 3610 7340 3640
rect 7340 3610 7345 3640
rect 7305 3605 7345 3610
rect 7605 3640 7645 3645
rect 7605 3610 7610 3640
rect 7610 3610 7640 3640
rect 7640 3610 7645 3640
rect 7605 3605 7645 3610
rect 7905 3640 7945 3645
rect 7905 3610 7910 3640
rect 7910 3610 7940 3640
rect 7940 3610 7945 3640
rect 7905 3605 7945 3610
rect 8205 3640 8245 3645
rect 8205 3610 8210 3640
rect 8210 3610 8240 3640
rect 8240 3610 8245 3640
rect 8205 3605 8245 3610
rect 8505 3640 8545 3645
rect 8505 3610 8510 3640
rect 8510 3610 8540 3640
rect 8540 3610 8545 3640
rect 8505 3605 8545 3610
rect 8805 3640 8845 3645
rect 8805 3610 8810 3640
rect 8810 3610 8840 3640
rect 8840 3610 8845 3640
rect 8805 3605 8845 3610
rect 9105 3640 9145 3645
rect 9105 3610 9110 3640
rect 9110 3610 9140 3640
rect 9140 3610 9145 3640
rect 9105 3605 9145 3610
rect 9405 3640 9445 3645
rect 9405 3610 9410 3640
rect 9410 3610 9440 3640
rect 9440 3610 9445 3640
rect 9405 3605 9445 3610
rect 9705 3640 9745 3645
rect 9705 3610 9710 3640
rect 9710 3610 9740 3640
rect 9740 3610 9745 3640
rect 9705 3605 9745 3610
rect 10005 3640 10045 3645
rect 10005 3610 10010 3640
rect 10010 3610 10040 3640
rect 10040 3610 10045 3640
rect 10005 3605 10045 3610
rect 10305 3640 10345 3645
rect 10305 3610 10310 3640
rect 10310 3610 10340 3640
rect 10340 3610 10345 3640
rect 10305 3605 10345 3610
rect 10605 3640 10645 3645
rect 10605 3610 10610 3640
rect 10610 3610 10640 3640
rect 10640 3610 10645 3640
rect 10605 3605 10645 3610
rect 10905 3640 10945 3645
rect 10905 3610 10910 3640
rect 10910 3610 10940 3640
rect 10940 3610 10945 3640
rect 10905 3605 10945 3610
rect 11205 3640 11245 3645
rect 11205 3610 11210 3640
rect 11210 3610 11240 3640
rect 11240 3610 11245 3640
rect 11205 3605 11245 3610
rect 11355 3640 11395 3645
rect 11355 3610 11360 3640
rect 11360 3610 11390 3640
rect 11390 3610 11395 3640
rect 11355 3605 11395 3610
rect 11505 3640 11545 3645
rect 11505 3610 11510 3640
rect 11510 3610 11540 3640
rect 11540 3610 11545 3640
rect 11505 3605 11545 3610
rect 11805 3640 11845 3645
rect 11805 3610 11810 3640
rect 11810 3610 11840 3640
rect 11840 3610 11845 3640
rect 11805 3605 11845 3610
rect 12105 3640 12145 3645
rect 12105 3610 12110 3640
rect 12110 3610 12140 3640
rect 12140 3610 12145 3640
rect 12105 3605 12145 3610
rect 12405 3640 12445 3645
rect 12405 3610 12410 3640
rect 12410 3610 12440 3640
rect 12440 3610 12445 3640
rect 12405 3605 12445 3610
rect 12555 3640 12595 3645
rect 12555 3610 12560 3640
rect 12560 3610 12590 3640
rect 12590 3610 12595 3640
rect 12555 3605 12595 3610
rect 12705 3640 12745 3645
rect 12705 3610 12710 3640
rect 12710 3610 12740 3640
rect 12740 3610 12745 3640
rect 12705 3605 12745 3610
rect 13005 3640 13045 3645
rect 13005 3610 13010 3640
rect 13010 3610 13040 3640
rect 13040 3610 13045 3640
rect 13005 3605 13045 3610
rect 13305 3640 13345 3645
rect 13305 3610 13310 3640
rect 13310 3610 13340 3640
rect 13340 3610 13345 3640
rect 13305 3605 13345 3610
rect 13605 3640 13645 3645
rect 13605 3610 13610 3640
rect 13610 3610 13640 3640
rect 13640 3610 13645 3640
rect 13605 3605 13645 3610
rect 13755 3640 13795 3645
rect 13755 3610 13760 3640
rect 13760 3610 13790 3640
rect 13790 3610 13795 3640
rect 13755 3605 13795 3610
rect 13905 3640 13945 3645
rect 13905 3610 13910 3640
rect 13910 3610 13940 3640
rect 13940 3610 13945 3640
rect 13905 3605 13945 3610
rect 14205 3640 14245 3645
rect 14205 3610 14210 3640
rect 14210 3610 14240 3640
rect 14240 3610 14245 3640
rect 14205 3605 14245 3610
rect 14505 3640 14545 3645
rect 14505 3610 14510 3640
rect 14510 3610 14540 3640
rect 14540 3610 14545 3640
rect 14505 3605 14545 3610
rect 14805 3640 14845 3645
rect 14805 3610 14810 3640
rect 14810 3610 14840 3640
rect 14840 3610 14845 3640
rect 14805 3605 14845 3610
rect 14955 3640 14995 3645
rect 14955 3610 14960 3640
rect 14960 3610 14990 3640
rect 14990 3610 14995 3640
rect 14955 3605 14995 3610
rect 15105 3640 15145 3645
rect 15105 3610 15110 3640
rect 15110 3610 15140 3640
rect 15140 3610 15145 3640
rect 15105 3605 15145 3610
rect 15405 3640 15445 3645
rect 15405 3610 15410 3640
rect 15410 3610 15440 3640
rect 15440 3610 15445 3640
rect 15405 3605 15445 3610
rect 15705 3640 15745 3645
rect 15705 3610 15710 3640
rect 15710 3610 15740 3640
rect 15740 3610 15745 3640
rect 15705 3605 15745 3610
rect 16005 3640 16045 3645
rect 16005 3610 16010 3640
rect 16010 3610 16040 3640
rect 16040 3610 16045 3640
rect 16005 3605 16045 3610
rect 16305 3640 16345 3645
rect 16305 3610 16310 3640
rect 16310 3610 16340 3640
rect 16340 3610 16345 3640
rect 16305 3605 16345 3610
rect 16605 3640 16645 3645
rect 16605 3610 16610 3640
rect 16610 3610 16640 3640
rect 16640 3610 16645 3640
rect 16605 3605 16645 3610
rect 16755 3640 16795 3645
rect 16755 3610 16760 3640
rect 16760 3610 16790 3640
rect 16790 3610 16795 3640
rect 16755 3605 16795 3610
rect 16905 3640 16945 3645
rect 16905 3610 16910 3640
rect 16910 3610 16940 3640
rect 16940 3610 16945 3640
rect 16905 3605 16945 3610
rect 17205 3640 17245 3645
rect 17205 3610 17210 3640
rect 17210 3610 17240 3640
rect 17240 3610 17245 3640
rect 17205 3605 17245 3610
rect 17505 3640 17545 3645
rect 17505 3610 17510 3640
rect 17510 3610 17540 3640
rect 17540 3610 17545 3640
rect 17505 3605 17545 3610
rect 17805 3640 17845 3645
rect 17805 3610 17810 3640
rect 17810 3610 17840 3640
rect 17840 3610 17845 3640
rect 17805 3605 17845 3610
rect 18105 3640 18145 3645
rect 18105 3610 18110 3640
rect 18110 3610 18140 3640
rect 18140 3610 18145 3640
rect 18105 3605 18145 3610
rect 18405 3640 18445 3645
rect 18405 3610 18410 3640
rect 18410 3610 18440 3640
rect 18440 3610 18445 3640
rect 18405 3605 18445 3610
rect 18705 3640 18745 3645
rect 18705 3610 18710 3640
rect 18710 3610 18740 3640
rect 18740 3610 18745 3640
rect 18705 3605 18745 3610
rect 19005 3640 19045 3645
rect 19005 3610 19010 3640
rect 19010 3610 19040 3640
rect 19040 3610 19045 3640
rect 19005 3605 19045 3610
rect 19155 3640 19195 3645
rect 19155 3610 19160 3640
rect 19160 3610 19190 3640
rect 19190 3610 19195 3640
rect 19155 3605 19195 3610
rect 19305 3640 19345 3645
rect 19305 3610 19310 3640
rect 19310 3610 19340 3640
rect 19340 3610 19345 3640
rect 19305 3605 19345 3610
rect 19605 3640 19645 3645
rect 19605 3610 19610 3640
rect 19610 3610 19640 3640
rect 19640 3610 19645 3640
rect 19605 3605 19645 3610
rect 19905 3640 19945 3645
rect 19905 3610 19910 3640
rect 19910 3610 19940 3640
rect 19940 3610 19945 3640
rect 19905 3605 19945 3610
rect 20205 3640 20245 3645
rect 20205 3610 20210 3640
rect 20210 3610 20240 3640
rect 20240 3610 20245 3640
rect 20205 3605 20245 3610
rect 20505 3640 20545 3645
rect 20505 3610 20510 3640
rect 20510 3610 20540 3640
rect 20540 3610 20545 3640
rect 20505 3605 20545 3610
rect 20805 3640 20845 3645
rect 20805 3610 20810 3640
rect 20810 3610 20840 3640
rect 20840 3610 20845 3640
rect 20805 3605 20845 3610
rect 20955 3640 20995 3645
rect 20955 3610 20960 3640
rect 20960 3610 20990 3640
rect 20990 3610 20995 3640
rect 20955 3605 20995 3610
rect 21105 3640 21145 3645
rect 21105 3610 21110 3640
rect 21110 3610 21140 3640
rect 21140 3610 21145 3640
rect 21105 3605 21145 3610
rect 21705 3640 21745 3645
rect 21705 3610 21710 3640
rect 21710 3610 21740 3640
rect 21740 3610 21745 3640
rect 21705 3605 21745 3610
rect 21855 3640 21895 3645
rect 21855 3610 21860 3640
rect 21860 3610 21890 3640
rect 21890 3610 21895 3640
rect 21855 3605 21895 3610
rect 22005 3640 22045 3645
rect 22005 3610 22010 3640
rect 22010 3610 22040 3640
rect 22040 3610 22045 3640
rect 22005 3605 22045 3610
rect 22305 3640 22345 3645
rect 22305 3610 22310 3640
rect 22310 3610 22340 3640
rect 22340 3610 22345 3640
rect 22305 3605 22345 3610
rect 22605 3640 22645 3645
rect 22605 3610 22610 3640
rect 22610 3610 22640 3640
rect 22640 3610 22645 3640
rect 22605 3605 22645 3610
rect 22905 3640 22945 3645
rect 22905 3610 22910 3640
rect 22910 3610 22940 3640
rect 22940 3610 22945 3640
rect 22905 3605 22945 3610
rect 23055 3640 23095 3645
rect 23055 3610 23060 3640
rect 23060 3610 23090 3640
rect 23090 3610 23095 3640
rect 23055 3605 23095 3610
rect 23205 3640 23245 3645
rect 23205 3610 23210 3640
rect 23210 3610 23240 3640
rect 23240 3610 23245 3640
rect 23205 3605 23245 3610
rect 23355 3640 23395 3645
rect 23355 3610 23360 3640
rect 23360 3610 23390 3640
rect 23390 3610 23395 3640
rect 23355 3605 23395 3610
rect 23655 3640 23695 3645
rect 23655 3610 23660 3640
rect 23660 3610 23690 3640
rect 23690 3610 23695 3640
rect 23655 3605 23695 3610
rect 23805 3640 23845 3645
rect 23805 3610 23810 3640
rect 23810 3610 23840 3640
rect 23840 3610 23845 3640
rect 23805 3605 23845 3610
rect 23955 3640 23995 3645
rect 23955 3610 23960 3640
rect 23960 3610 23990 3640
rect 23990 3610 23995 3640
rect 23955 3605 23995 3610
rect 24105 3640 24145 3645
rect 24105 3610 24110 3640
rect 24110 3610 24140 3640
rect 24140 3610 24145 3640
rect 24105 3605 24145 3610
rect 24405 3640 24445 3645
rect 24405 3610 24410 3640
rect 24410 3610 24440 3640
rect 24440 3610 24445 3640
rect 24405 3605 24445 3610
rect 24705 3640 24745 3645
rect 24705 3610 24710 3640
rect 24710 3610 24740 3640
rect 24740 3610 24745 3640
rect 24705 3605 24745 3610
rect 25005 3640 25045 3645
rect 25005 3610 25010 3640
rect 25010 3610 25040 3640
rect 25040 3610 25045 3640
rect 25005 3605 25045 3610
rect 25455 3640 25495 3645
rect 25455 3610 25460 3640
rect 25460 3610 25490 3640
rect 25490 3610 25495 3640
rect 25455 3605 25495 3610
rect 25605 3640 25645 3645
rect 25605 3610 25610 3640
rect 25610 3610 25640 3640
rect 25640 3610 25645 3640
rect 25605 3605 25645 3610
rect 25755 3640 25795 3645
rect 25755 3610 25760 3640
rect 25760 3610 25790 3640
rect 25790 3610 25795 3640
rect 25755 3605 25795 3610
rect 26205 3640 26245 3645
rect 26205 3610 26210 3640
rect 26210 3610 26240 3640
rect 26240 3610 26245 3640
rect 26205 3605 26245 3610
rect 26505 3640 26545 3645
rect 26505 3610 26510 3640
rect 26510 3610 26540 3640
rect 26540 3610 26545 3640
rect 26505 3605 26545 3610
rect 26805 3640 26845 3645
rect 26805 3610 26810 3640
rect 26810 3610 26840 3640
rect 26840 3610 26845 3640
rect 26805 3605 26845 3610
rect 27105 3640 27145 3645
rect 27105 3610 27110 3640
rect 27110 3610 27140 3640
rect 27140 3610 27145 3640
rect 27105 3605 27145 3610
rect 27555 3640 27595 3645
rect 27555 3610 27560 3640
rect 27560 3610 27590 3640
rect 27590 3610 27595 3640
rect 27555 3605 27595 3610
rect 27705 3640 27745 3645
rect 27705 3610 27710 3640
rect 27710 3610 27740 3640
rect 27740 3610 27745 3640
rect 27705 3605 27745 3610
rect 27855 3640 27895 3645
rect 27855 3610 27860 3640
rect 27860 3610 27890 3640
rect 27890 3610 27895 3640
rect 27855 3605 27895 3610
rect 28305 3640 28345 3645
rect 28305 3610 28310 3640
rect 28310 3610 28340 3640
rect 28340 3610 28345 3640
rect 28305 3605 28345 3610
rect 28605 3640 28645 3645
rect 28605 3610 28610 3640
rect 28610 3610 28640 3640
rect 28640 3610 28645 3640
rect 28605 3605 28645 3610
rect 28755 3640 28795 3645
rect 28755 3610 28760 3640
rect 28760 3610 28790 3640
rect 28790 3610 28795 3640
rect 28755 3605 28795 3610
rect 28905 3640 28945 3645
rect 28905 3610 28910 3640
rect 28910 3610 28940 3640
rect 28940 3610 28945 3640
rect 28905 3605 28945 3610
rect 29205 3640 29245 3645
rect 29205 3610 29210 3640
rect 29210 3610 29240 3640
rect 29240 3610 29245 3640
rect 29205 3605 29245 3610
rect 29355 3640 29395 3645
rect 29355 3610 29360 3640
rect 29360 3610 29390 3640
rect 29390 3610 29395 3640
rect 29355 3605 29395 3610
rect 29655 3640 29695 3645
rect 29655 3610 29660 3640
rect 29660 3610 29690 3640
rect 29690 3610 29695 3640
rect 29655 3605 29695 3610
rect 29955 3640 29995 3645
rect 29955 3610 29960 3640
rect 29960 3610 29990 3640
rect 29990 3610 29995 3640
rect 29955 3605 29995 3610
rect 30255 3640 30295 3645
rect 30255 3610 30260 3640
rect 30260 3610 30290 3640
rect 30290 3610 30295 3640
rect 30255 3605 30295 3610
rect 30555 3640 30595 3645
rect 30555 3610 30560 3640
rect 30560 3610 30590 3640
rect 30590 3610 30595 3640
rect 30555 3605 30595 3610
rect 30855 3640 30895 3645
rect 30855 3610 30860 3640
rect 30860 3610 30890 3640
rect 30890 3610 30895 3640
rect 30855 3605 30895 3610
rect 31005 3640 31045 3645
rect 31005 3610 31010 3640
rect 31010 3610 31040 3640
rect 31040 3610 31045 3640
rect 31005 3605 31045 3610
rect 31455 3640 31495 3645
rect 31455 3610 31460 3640
rect 31460 3610 31490 3640
rect 31490 3610 31495 3640
rect 31455 3605 31495 3610
rect 31605 3640 31645 3645
rect 31605 3610 31610 3640
rect 31610 3610 31640 3640
rect 31640 3610 31645 3640
rect 31605 3605 31645 3610
rect 31905 3640 31945 3645
rect 31905 3610 31910 3640
rect 31910 3610 31940 3640
rect 31940 3610 31945 3640
rect 31905 3605 31945 3610
rect 32055 3640 32095 3645
rect 32055 3610 32060 3640
rect 32060 3610 32090 3640
rect 32090 3610 32095 3640
rect 32055 3605 32095 3610
rect -345 3405 -305 3445
rect 105 3405 145 3445
rect 405 3405 445 3445
rect 2055 3405 2095 3445
rect 3705 3405 3745 3445
rect 4005 3405 4045 3445
rect 4305 3405 4345 3445
rect 4605 3405 4645 3445
rect 6255 3405 6295 3445
rect 7905 3405 7945 3445
rect 8205 3405 8245 3445
rect 18105 3405 18145 3445
rect 18405 3405 18445 3445
rect 19905 3405 19945 3445
rect 20205 3405 20245 3445
rect 24705 3405 24745 3445
rect 25005 3405 25045 3445
rect 26205 3405 26245 3445
rect 26505 3405 26545 3445
rect 26805 3405 26845 3445
rect 27105 3405 27145 3445
rect 705 3305 745 3345
rect 1005 3305 1045 3345
rect 1155 3305 1195 3345
rect 1305 3305 1345 3345
rect 1605 3305 1645 3345
rect 2505 3305 2545 3345
rect 2805 3305 2845 3345
rect 2955 3305 2995 3345
rect 3105 3305 3145 3345
rect 3405 3305 3445 3345
rect 4905 3305 4945 3345
rect 5205 3305 5245 3345
rect 5355 3305 5395 3345
rect 5505 3305 5545 3345
rect 5805 3305 5845 3345
rect 6705 3305 6745 3345
rect 7005 3305 7045 3345
rect 7155 3305 7195 3345
rect 7305 3305 7345 3345
rect 7605 3305 7645 3345
rect 9555 3305 9595 3345
rect 25455 3305 25495 3345
rect 25755 3305 25795 3345
rect 27555 3305 27595 3345
rect 27855 3305 27895 3345
rect 29955 3305 29995 3345
rect 30255 3305 30295 3345
rect 30555 3305 30595 3345
rect 30855 3305 30895 3345
rect 1905 3205 1945 3245
rect 2205 3205 2245 3245
rect 6105 3205 6145 3245
rect 6405 3205 6445 3245
rect -495 3105 -455 3145
rect -195 3105 -155 3145
rect 13305 2705 13345 2745
rect 13605 2705 13645 2745
rect 13905 2705 13945 2745
rect 14205 2705 14245 2745
rect 18705 2705 18745 2745
rect 19005 2705 19045 2745
rect 19305 2705 19345 2745
rect 12105 2105 12145 2145
rect 12405 2105 12445 2145
rect 12705 2105 12745 2145
rect 13005 2105 13045 2145
rect 16305 2105 16345 2145
rect 16605 2105 16645 2145
rect 16905 2105 16945 2145
rect 17205 2105 17245 2145
rect -495 1305 -455 1345
rect -195 1305 -155 1345
rect 3705 1205 3745 1245
rect 4005 1205 4045 1245
rect 4305 1205 4345 1245
rect 4605 1205 4645 1245
rect 1305 1105 1345 1145
rect 1605 1105 1645 1145
rect 1905 1105 1945 1145
rect 2205 1105 2245 1145
rect 2355 1105 2395 1145
rect 2505 1105 2545 1145
rect 2805 1105 2845 1145
rect 3105 1105 3145 1145
rect 3405 1105 3445 1145
rect 4905 1105 4945 1145
rect 5205 1105 5245 1145
rect 5505 1105 5545 1145
rect 5805 1105 5845 1145
rect 5955 1105 5995 1145
rect 6105 1105 6145 1145
rect 6405 1105 6445 1145
rect 6705 1105 6745 1145
rect 7005 1105 7045 1145
rect 21705 1105 21745 1145
rect 22005 1105 22045 1145
rect 22305 1105 22345 1145
rect 22605 1105 22645 1145
rect 22905 1105 22945 1145
rect 23205 1105 23245 1145
rect -345 1005 -305 1045
rect 105 1005 145 1045
rect 405 1005 445 1045
rect 705 1005 745 1045
rect 1005 1005 1045 1045
rect 3855 1005 3895 1045
rect 4455 1005 4495 1045
rect 7305 1005 7345 1045
rect 7605 1005 7645 1045
rect 7905 1005 7945 1045
rect 8205 1005 8245 1045
rect 8505 1005 8545 1045
rect 8805 1005 8845 1045
rect 9105 1005 9145 1045
rect 9405 1005 9445 1045
rect 9705 1005 9745 1045
rect 10005 1005 10045 1045
rect 10305 1005 10345 1045
rect 10605 1005 10645 1045
rect 10905 1005 10945 1045
rect 11205 1005 11245 1045
rect 11505 1005 11545 1045
rect 11805 1005 11845 1045
rect 14505 1005 14545 1045
rect 14805 1005 14845 1045
rect 15105 1005 15145 1045
rect 15405 1005 15445 1045
rect 20505 1005 20545 1045
rect 20805 1005 20845 1045
rect 21105 1005 21145 1045
rect 21405 1005 21445 1045
rect 23505 1005 23545 1045
rect 23805 1005 23845 1045
rect 24105 1005 24145 1045
rect 24405 1005 24445 1045
rect -495 840 -455 845
rect -495 810 -490 840
rect -490 810 -460 840
rect -460 810 -455 840
rect -495 805 -455 810
rect -345 840 -305 845
rect -345 810 -340 840
rect -340 810 -310 840
rect -310 810 -305 840
rect -345 805 -305 810
rect -195 840 -155 845
rect -195 810 -190 840
rect -190 810 -160 840
rect -160 810 -155 840
rect -195 805 -155 810
rect 105 840 145 845
rect 105 810 110 840
rect 110 810 140 840
rect 140 810 145 840
rect 105 805 145 810
rect 405 840 445 845
rect 405 810 410 840
rect 410 810 440 840
rect 440 810 445 840
rect 405 805 445 810
rect 705 840 745 845
rect 705 810 710 840
rect 710 810 740 840
rect 740 810 745 840
rect 705 805 745 810
rect 1005 840 1045 845
rect 1005 810 1010 840
rect 1010 810 1040 840
rect 1040 810 1045 840
rect 1005 805 1045 810
rect 1305 840 1345 845
rect 1305 810 1310 840
rect 1310 810 1340 840
rect 1340 810 1345 840
rect 1305 805 1345 810
rect 1605 840 1645 845
rect 1605 810 1610 840
rect 1610 810 1640 840
rect 1640 810 1645 840
rect 1605 805 1645 810
rect 1905 840 1945 845
rect 1905 810 1910 840
rect 1910 810 1940 840
rect 1940 810 1945 840
rect 1905 805 1945 810
rect 2205 840 2245 845
rect 2205 810 2210 840
rect 2210 810 2240 840
rect 2240 810 2245 840
rect 2205 805 2245 810
rect 2355 840 2395 845
rect 2355 810 2360 840
rect 2360 810 2390 840
rect 2390 810 2395 840
rect 2355 805 2395 810
rect 2505 840 2545 845
rect 2505 810 2510 840
rect 2510 810 2540 840
rect 2540 810 2545 840
rect 2505 805 2545 810
rect 2805 840 2845 845
rect 2805 810 2810 840
rect 2810 810 2840 840
rect 2840 810 2845 840
rect 2805 805 2845 810
rect 3105 840 3145 845
rect 3105 810 3110 840
rect 3110 810 3140 840
rect 3140 810 3145 840
rect 3105 805 3145 810
rect 3405 840 3445 845
rect 3405 810 3410 840
rect 3410 810 3440 840
rect 3440 810 3445 840
rect 3405 805 3445 810
rect 3705 840 3745 845
rect 3705 810 3710 840
rect 3710 810 3740 840
rect 3740 810 3745 840
rect 3705 805 3745 810
rect 3855 840 3895 845
rect 3855 810 3860 840
rect 3860 810 3890 840
rect 3890 810 3895 840
rect 3855 805 3895 810
rect 4005 840 4045 845
rect 4005 810 4010 840
rect 4010 810 4040 840
rect 4040 810 4045 840
rect 4005 805 4045 810
rect 4305 840 4345 845
rect 4305 810 4310 840
rect 4310 810 4340 840
rect 4340 810 4345 840
rect 4305 805 4345 810
rect 4455 840 4495 845
rect 4455 810 4460 840
rect 4460 810 4490 840
rect 4490 810 4495 840
rect 4455 805 4495 810
rect 4605 840 4645 845
rect 4605 810 4610 840
rect 4610 810 4640 840
rect 4640 810 4645 840
rect 4605 805 4645 810
rect 4905 840 4945 845
rect 4905 810 4910 840
rect 4910 810 4940 840
rect 4940 810 4945 840
rect 4905 805 4945 810
rect 5205 840 5245 845
rect 5205 810 5210 840
rect 5210 810 5240 840
rect 5240 810 5245 840
rect 5205 805 5245 810
rect 5505 840 5545 845
rect 5505 810 5510 840
rect 5510 810 5540 840
rect 5540 810 5545 840
rect 5505 805 5545 810
rect 5805 840 5845 845
rect 5805 810 5810 840
rect 5810 810 5840 840
rect 5840 810 5845 840
rect 5805 805 5845 810
rect 5955 840 5995 845
rect 5955 810 5960 840
rect 5960 810 5990 840
rect 5990 810 5995 840
rect 5955 805 5995 810
rect 6105 840 6145 845
rect 6105 810 6110 840
rect 6110 810 6140 840
rect 6140 810 6145 840
rect 6105 805 6145 810
rect 6405 840 6445 845
rect 6405 810 6410 840
rect 6410 810 6440 840
rect 6440 810 6445 840
rect 6405 805 6445 810
rect 6705 840 6745 845
rect 6705 810 6710 840
rect 6710 810 6740 840
rect 6740 810 6745 840
rect 6705 805 6745 810
rect 7005 840 7045 845
rect 7005 810 7010 840
rect 7010 810 7040 840
rect 7040 810 7045 840
rect 7005 805 7045 810
rect 7305 840 7345 845
rect 7305 810 7310 840
rect 7310 810 7340 840
rect 7340 810 7345 840
rect 7305 805 7345 810
rect 7605 840 7645 845
rect 7605 810 7610 840
rect 7610 810 7640 840
rect 7640 810 7645 840
rect 7605 805 7645 810
rect 7905 840 7945 845
rect 7905 810 7910 840
rect 7910 810 7940 840
rect 7940 810 7945 840
rect 7905 805 7945 810
rect 8205 840 8245 845
rect 8205 810 8210 840
rect 8210 810 8240 840
rect 8240 810 8245 840
rect 8205 805 8245 810
rect 8505 840 8545 845
rect 8505 810 8510 840
rect 8510 810 8540 840
rect 8540 810 8545 840
rect 8505 805 8545 810
rect 8805 840 8845 845
rect 8805 810 8810 840
rect 8810 810 8840 840
rect 8840 810 8845 840
rect 8805 805 8845 810
rect 9105 840 9145 845
rect 9105 810 9110 840
rect 9110 810 9140 840
rect 9140 810 9145 840
rect 9105 805 9145 810
rect 9405 840 9445 845
rect 9405 810 9410 840
rect 9410 810 9440 840
rect 9440 810 9445 840
rect 9405 805 9445 810
rect 9555 840 9595 845
rect 9555 810 9560 840
rect 9560 810 9590 840
rect 9590 810 9595 840
rect 9555 805 9595 810
rect 9705 840 9745 845
rect 9705 810 9710 840
rect 9710 810 9740 840
rect 9740 810 9745 840
rect 9705 805 9745 810
rect 10005 840 10045 845
rect 10005 810 10010 840
rect 10010 810 10040 840
rect 10040 810 10045 840
rect 10005 805 10045 810
rect 10305 840 10345 845
rect 10305 810 10310 840
rect 10310 810 10340 840
rect 10340 810 10345 840
rect 10305 805 10345 810
rect 10605 840 10645 845
rect 10605 810 10610 840
rect 10610 810 10640 840
rect 10640 810 10645 840
rect 10605 805 10645 810
rect 10905 840 10945 845
rect 10905 810 10910 840
rect 10910 810 10940 840
rect 10940 810 10945 840
rect 10905 805 10945 810
rect 11205 840 11245 845
rect 11205 810 11210 840
rect 11210 810 11240 840
rect 11240 810 11245 840
rect 11205 805 11245 810
rect 11505 840 11545 845
rect 11505 810 11510 840
rect 11510 810 11540 840
rect 11540 810 11545 840
rect 11505 805 11545 810
rect 11805 840 11845 845
rect 11805 810 11810 840
rect 11810 810 11840 840
rect 11840 810 11845 840
rect 11805 805 11845 810
rect 12105 840 12145 845
rect 12105 810 12110 840
rect 12110 810 12140 840
rect 12140 810 12145 840
rect 12105 805 12145 810
rect 12405 840 12445 845
rect 12405 810 12410 840
rect 12410 810 12440 840
rect 12440 810 12445 840
rect 12405 805 12445 810
rect 12555 840 12595 845
rect 12555 810 12560 840
rect 12560 810 12590 840
rect 12590 810 12595 840
rect 12555 805 12595 810
rect 12705 840 12745 845
rect 12705 810 12710 840
rect 12710 810 12740 840
rect 12740 810 12745 840
rect 12705 805 12745 810
rect 13005 840 13045 845
rect 13005 810 13010 840
rect 13010 810 13040 840
rect 13040 810 13045 840
rect 13005 805 13045 810
rect 13305 840 13345 845
rect 13305 810 13310 840
rect 13310 810 13340 840
rect 13340 810 13345 840
rect 13305 805 13345 810
rect 13605 840 13645 845
rect 13605 810 13610 840
rect 13610 810 13640 840
rect 13640 810 13645 840
rect 13605 805 13645 810
rect 13755 840 13795 845
rect 13755 810 13760 840
rect 13760 810 13790 840
rect 13790 810 13795 840
rect 13755 805 13795 810
rect 13905 840 13945 845
rect 13905 810 13910 840
rect 13910 810 13940 840
rect 13940 810 13945 840
rect 13905 805 13945 810
rect 14205 840 14245 845
rect 14205 810 14210 840
rect 14210 810 14240 840
rect 14240 810 14245 840
rect 14205 805 14245 810
rect 14505 840 14545 845
rect 14505 810 14510 840
rect 14510 810 14540 840
rect 14540 810 14545 840
rect 14505 805 14545 810
rect 14805 840 14845 845
rect 14805 810 14810 840
rect 14810 810 14840 840
rect 14840 810 14845 840
rect 14805 805 14845 810
rect 15105 840 15145 845
rect 15105 810 15110 840
rect 15110 810 15140 840
rect 15140 810 15145 840
rect 15105 805 15145 810
rect 15405 840 15445 845
rect 15405 810 15410 840
rect 15410 810 15440 840
rect 15440 810 15445 840
rect 15405 805 15445 810
rect 15705 840 15745 845
rect 15705 810 15710 840
rect 15710 810 15740 840
rect 15740 810 15745 840
rect 15705 805 15745 810
rect 16005 840 16045 845
rect 16005 810 16010 840
rect 16010 810 16040 840
rect 16040 810 16045 840
rect 16005 805 16045 810
rect 16305 840 16345 845
rect 16305 810 16310 840
rect 16310 810 16340 840
rect 16340 810 16345 840
rect 16305 805 16345 810
rect 16605 840 16645 845
rect 16605 810 16610 840
rect 16610 810 16640 840
rect 16640 810 16645 840
rect 16605 805 16645 810
rect 16755 840 16795 845
rect 16755 810 16760 840
rect 16760 810 16790 840
rect 16790 810 16795 840
rect 16755 805 16795 810
rect 16905 840 16945 845
rect 16905 810 16910 840
rect 16910 810 16940 840
rect 16940 810 16945 840
rect 16905 805 16945 810
rect 17205 840 17245 845
rect 17205 810 17210 840
rect 17210 810 17240 840
rect 17240 810 17245 840
rect 17205 805 17245 810
rect 17505 840 17545 845
rect 17505 810 17510 840
rect 17510 810 17540 840
rect 17540 810 17545 840
rect 17505 805 17545 810
rect 17805 840 17845 845
rect 17805 810 17810 840
rect 17810 810 17840 840
rect 17840 810 17845 840
rect 17805 805 17845 810
rect 18105 840 18145 845
rect 18105 810 18110 840
rect 18110 810 18140 840
rect 18140 810 18145 840
rect 18105 805 18145 810
rect 18405 840 18445 845
rect 18405 810 18410 840
rect 18410 810 18440 840
rect 18440 810 18445 840
rect 18405 805 18445 810
rect 18705 840 18745 845
rect 18705 810 18710 840
rect 18710 810 18740 840
rect 18740 810 18745 840
rect 18705 805 18745 810
rect 19005 840 19045 845
rect 19005 810 19010 840
rect 19010 810 19040 840
rect 19040 810 19045 840
rect 19005 805 19045 810
rect 19155 840 19195 845
rect 19155 810 19160 840
rect 19160 810 19190 840
rect 19190 810 19195 840
rect 19155 805 19195 810
rect 19305 840 19345 845
rect 19305 810 19310 840
rect 19310 810 19340 840
rect 19340 810 19345 840
rect 19305 805 19345 810
rect 19605 840 19645 845
rect 19605 810 19610 840
rect 19610 810 19640 840
rect 19640 810 19645 840
rect 19605 805 19645 810
rect 19905 840 19945 845
rect 19905 810 19910 840
rect 19910 810 19940 840
rect 19940 810 19945 840
rect 19905 805 19945 810
rect 20205 840 20245 845
rect 20205 810 20210 840
rect 20210 810 20240 840
rect 20240 810 20245 840
rect 20205 805 20245 810
rect 20505 840 20545 845
rect 20505 810 20510 840
rect 20510 810 20540 840
rect 20540 810 20545 840
rect 20505 805 20545 810
rect 20805 840 20845 845
rect 20805 810 20810 840
rect 20810 810 20840 840
rect 20840 810 20845 840
rect 20805 805 20845 810
rect 21105 840 21145 845
rect 21105 810 21110 840
rect 21110 810 21140 840
rect 21140 810 21145 840
rect 21105 805 21145 810
rect 21405 840 21445 845
rect 21405 810 21410 840
rect 21410 810 21440 840
rect 21440 810 21445 840
rect 21405 805 21445 810
rect 21705 840 21745 845
rect 21705 810 21710 840
rect 21710 810 21740 840
rect 21740 810 21745 840
rect 21705 805 21745 810
rect 22005 840 22045 845
rect 22005 810 22010 840
rect 22010 810 22040 840
rect 22040 810 22045 840
rect 22005 805 22045 810
rect 22305 840 22345 845
rect 22305 810 22310 840
rect 22310 810 22340 840
rect 22340 810 22345 840
rect 22305 805 22345 810
rect 22455 840 22495 845
rect 22455 810 22460 840
rect 22460 810 22490 840
rect 22490 810 22495 840
rect 22455 805 22495 810
rect 22605 840 22645 845
rect 22605 810 22610 840
rect 22610 810 22640 840
rect 22640 810 22645 840
rect 22605 805 22645 810
rect 22905 840 22945 845
rect 22905 810 22910 840
rect 22910 810 22940 840
rect 22940 810 22945 840
rect 22905 805 22945 810
rect 23205 840 23245 845
rect 23205 810 23210 840
rect 23210 810 23240 840
rect 23240 810 23245 840
rect 23205 805 23245 810
rect 23505 840 23545 845
rect 23505 810 23510 840
rect 23510 810 23540 840
rect 23540 810 23545 840
rect 23505 805 23545 810
rect 23805 840 23845 845
rect 23805 810 23810 840
rect 23810 810 23840 840
rect 23840 810 23845 840
rect 23805 805 23845 810
rect 24105 840 24145 845
rect 24105 810 24110 840
rect 24110 810 24140 840
rect 24140 810 24145 840
rect 24105 805 24145 810
rect 24405 840 24445 845
rect 24405 810 24410 840
rect 24410 810 24440 840
rect 24440 810 24445 840
rect 24405 805 24445 810
rect 24705 840 24745 845
rect 24705 810 24710 840
rect 24710 810 24740 840
rect 24740 810 24745 840
rect 24705 805 24745 810
rect 25005 840 25045 845
rect 25005 810 25010 840
rect 25010 810 25040 840
rect 25040 810 25045 840
rect 25005 805 25045 810
rect 25305 840 25345 845
rect 25305 810 25310 840
rect 25310 810 25340 840
rect 25340 810 25345 840
rect 25305 805 25345 810
rect 25605 840 25645 845
rect 25605 810 25610 840
rect 25610 810 25640 840
rect 25640 810 25645 840
rect 25605 805 25645 810
rect 25755 840 25795 845
rect 25755 810 25760 840
rect 25760 810 25790 840
rect 25790 810 25795 840
rect 25755 805 25795 810
rect 25905 840 25945 845
rect 25905 810 25910 840
rect 25910 810 25940 840
rect 25940 810 25945 840
rect 25905 805 25945 810
rect 26205 840 26245 845
rect 26205 810 26210 840
rect 26210 810 26240 840
rect 26240 810 26245 840
rect 26205 805 26245 810
rect 26505 840 26545 845
rect 26505 810 26510 840
rect 26510 810 26540 840
rect 26540 810 26545 840
rect 26505 805 26545 810
rect 26655 840 26695 845
rect 26655 810 26660 840
rect 26660 810 26690 840
rect 26690 810 26695 840
rect 26655 805 26695 810
rect 26805 840 26845 845
rect 26805 810 26810 840
rect 26810 810 26840 840
rect 26840 810 26845 840
rect 26805 805 26845 810
rect 27105 840 27145 845
rect 27105 810 27110 840
rect 27110 810 27140 840
rect 27140 810 27145 840
rect 27105 805 27145 810
rect 27405 840 27445 845
rect 27405 810 27410 840
rect 27410 810 27440 840
rect 27440 810 27445 840
rect 27405 805 27445 810
rect 27555 840 27595 845
rect 27555 810 27560 840
rect 27560 810 27590 840
rect 27590 810 27595 840
rect 27555 805 27595 810
rect 27705 840 27745 845
rect 27705 810 27710 840
rect 27710 810 27740 840
rect 27740 810 27745 840
rect 27705 805 27745 810
rect 28005 840 28045 845
rect 28005 810 28010 840
rect 28010 810 28040 840
rect 28040 810 28045 840
rect 28005 805 28045 810
rect 28305 840 28345 845
rect 28305 810 28310 840
rect 28310 810 28340 840
rect 28340 810 28345 840
rect 28305 805 28345 810
rect 28605 840 28645 845
rect 28605 810 28610 840
rect 28610 810 28640 840
rect 28640 810 28645 840
rect 28605 805 28645 810
rect 15705 605 15745 645
rect 16005 605 16045 645
rect 16305 605 16345 645
rect 16605 605 16645 645
rect 16905 605 16945 645
rect 17205 605 17245 645
rect 17505 605 17545 645
rect 17805 605 17845 645
rect 18105 605 18145 645
rect 18405 605 18445 645
rect 18705 605 18745 645
rect 19005 605 19045 645
rect 19305 605 19345 645
rect 19605 605 19645 645
rect 19905 605 19945 645
rect 20205 605 20245 645
rect 24705 605 24745 645
rect 25005 605 25045 645
rect 25305 605 25345 645
rect 25605 605 25645 645
rect 25905 605 25945 645
rect 26205 605 26245 645
rect 26505 605 26545 645
rect 26655 605 26695 645
rect 26805 605 26845 645
rect 27105 605 27145 645
rect 27405 605 27445 645
rect 27705 605 27745 645
rect 28005 605 28045 645
rect 28305 605 28345 645
rect 28605 605 28645 645
rect 16755 -495 16795 -455
rect 25755 -495 25795 -455
rect 27555 -495 27595 -455
rect -495 -860 -455 -855
rect -495 -890 -490 -860
rect -490 -890 -460 -860
rect -460 -890 -455 -860
rect -495 -895 -455 -890
rect -345 -860 -305 -855
rect -345 -890 -340 -860
rect -340 -890 -310 -860
rect -310 -890 -305 -860
rect -345 -895 -305 -890
rect -195 -860 -155 -855
rect -195 -890 -190 -860
rect -190 -890 -160 -860
rect -160 -890 -155 -860
rect -195 -895 -155 -890
rect 105 -860 145 -855
rect 105 -890 110 -860
rect 110 -890 140 -860
rect 140 -890 145 -860
rect 105 -895 145 -890
rect 405 -860 445 -855
rect 405 -890 410 -860
rect 410 -890 440 -860
rect 440 -890 445 -860
rect 405 -895 445 -890
rect 705 -860 745 -855
rect 705 -890 710 -860
rect 710 -890 740 -860
rect 740 -890 745 -860
rect 705 -895 745 -890
rect 1005 -860 1045 -855
rect 1005 -890 1010 -860
rect 1010 -890 1040 -860
rect 1040 -890 1045 -860
rect 1005 -895 1045 -890
rect 1305 -860 1345 -855
rect 1305 -890 1310 -860
rect 1310 -890 1340 -860
rect 1340 -890 1345 -860
rect 1305 -895 1345 -890
rect 1605 -860 1645 -855
rect 1605 -890 1610 -860
rect 1610 -890 1640 -860
rect 1640 -890 1645 -860
rect 1605 -895 1645 -890
rect 1905 -860 1945 -855
rect 1905 -890 1910 -860
rect 1910 -890 1940 -860
rect 1940 -890 1945 -860
rect 1905 -895 1945 -890
rect 2205 -860 2245 -855
rect 2205 -890 2210 -860
rect 2210 -890 2240 -860
rect 2240 -890 2245 -860
rect 2205 -895 2245 -890
rect 2355 -860 2395 -855
rect 2355 -890 2360 -860
rect 2360 -890 2390 -860
rect 2390 -890 2395 -860
rect 2355 -895 2395 -890
rect 2505 -860 2545 -855
rect 2505 -890 2510 -860
rect 2510 -890 2540 -860
rect 2540 -890 2545 -860
rect 2505 -895 2545 -890
rect 2805 -860 2845 -855
rect 2805 -890 2810 -860
rect 2810 -890 2840 -860
rect 2840 -890 2845 -860
rect 2805 -895 2845 -890
rect 3105 -860 3145 -855
rect 3105 -890 3110 -860
rect 3110 -890 3140 -860
rect 3140 -890 3145 -860
rect 3105 -895 3145 -890
rect 3405 -860 3445 -855
rect 3405 -890 3410 -860
rect 3410 -890 3440 -860
rect 3440 -890 3445 -860
rect 3405 -895 3445 -890
rect 3705 -860 3745 -855
rect 3705 -890 3710 -860
rect 3710 -890 3740 -860
rect 3740 -890 3745 -860
rect 3705 -895 3745 -890
rect 3855 -860 3895 -855
rect 3855 -890 3860 -860
rect 3860 -890 3890 -860
rect 3890 -890 3895 -860
rect 3855 -895 3895 -890
rect 4005 -860 4045 -855
rect 4005 -890 4010 -860
rect 4010 -890 4040 -860
rect 4040 -890 4045 -860
rect 4005 -895 4045 -890
rect 4305 -860 4345 -855
rect 4305 -890 4310 -860
rect 4310 -890 4340 -860
rect 4340 -890 4345 -860
rect 4305 -895 4345 -890
rect 4455 -860 4495 -855
rect 4455 -890 4460 -860
rect 4460 -890 4490 -860
rect 4490 -890 4495 -860
rect 4455 -895 4495 -890
rect 4605 -860 4645 -855
rect 4605 -890 4610 -860
rect 4610 -890 4640 -860
rect 4640 -890 4645 -860
rect 4605 -895 4645 -890
rect 4905 -860 4945 -855
rect 4905 -890 4910 -860
rect 4910 -890 4940 -860
rect 4940 -890 4945 -860
rect 4905 -895 4945 -890
rect 5205 -860 5245 -855
rect 5205 -890 5210 -860
rect 5210 -890 5240 -860
rect 5240 -890 5245 -860
rect 5205 -895 5245 -890
rect 5505 -860 5545 -855
rect 5505 -890 5510 -860
rect 5510 -890 5540 -860
rect 5540 -890 5545 -860
rect 5505 -895 5545 -890
rect 5805 -860 5845 -855
rect 5805 -890 5810 -860
rect 5810 -890 5840 -860
rect 5840 -890 5845 -860
rect 5805 -895 5845 -890
rect 5955 -860 5995 -855
rect 5955 -890 5960 -860
rect 5960 -890 5990 -860
rect 5990 -890 5995 -860
rect 5955 -895 5995 -890
rect 6105 -860 6145 -855
rect 6105 -890 6110 -860
rect 6110 -890 6140 -860
rect 6140 -890 6145 -860
rect 6105 -895 6145 -890
rect 6405 -860 6445 -855
rect 6405 -890 6410 -860
rect 6410 -890 6440 -860
rect 6440 -890 6445 -860
rect 6405 -895 6445 -890
rect 6705 -860 6745 -855
rect 6705 -890 6710 -860
rect 6710 -890 6740 -860
rect 6740 -890 6745 -860
rect 6705 -895 6745 -890
rect 7005 -860 7045 -855
rect 7005 -890 7010 -860
rect 7010 -890 7040 -860
rect 7040 -890 7045 -860
rect 7005 -895 7045 -890
rect 7305 -860 7345 -855
rect 7305 -890 7310 -860
rect 7310 -890 7340 -860
rect 7340 -890 7345 -860
rect 7305 -895 7345 -890
rect 7605 -860 7645 -855
rect 7605 -890 7610 -860
rect 7610 -890 7640 -860
rect 7640 -890 7645 -860
rect 7605 -895 7645 -890
rect 7905 -860 7945 -855
rect 7905 -890 7910 -860
rect 7910 -890 7940 -860
rect 7940 -890 7945 -860
rect 7905 -895 7945 -890
rect 8205 -860 8245 -855
rect 8205 -890 8210 -860
rect 8210 -890 8240 -860
rect 8240 -890 8245 -860
rect 8205 -895 8245 -890
rect 8505 -860 8545 -855
rect 8505 -890 8510 -860
rect 8510 -890 8540 -860
rect 8540 -890 8545 -860
rect 8505 -895 8545 -890
rect 8805 -860 8845 -855
rect 8805 -890 8810 -860
rect 8810 -890 8840 -860
rect 8840 -890 8845 -860
rect 8805 -895 8845 -890
rect 9105 -860 9145 -855
rect 9105 -890 9110 -860
rect 9110 -890 9140 -860
rect 9140 -890 9145 -860
rect 9105 -895 9145 -890
rect 9405 -860 9445 -855
rect 9405 -890 9410 -860
rect 9410 -890 9440 -860
rect 9440 -890 9445 -860
rect 9405 -895 9445 -890
rect 9555 -860 9595 -855
rect 9555 -890 9560 -860
rect 9560 -890 9590 -860
rect 9590 -890 9595 -860
rect 9555 -895 9595 -890
rect 9705 -860 9745 -855
rect 9705 -890 9710 -860
rect 9710 -890 9740 -860
rect 9740 -890 9745 -860
rect 9705 -895 9745 -890
rect 10005 -860 10045 -855
rect 10005 -890 10010 -860
rect 10010 -890 10040 -860
rect 10040 -890 10045 -860
rect 10005 -895 10045 -890
rect 10305 -860 10345 -855
rect 10305 -890 10310 -860
rect 10310 -890 10340 -860
rect 10340 -890 10345 -860
rect 10305 -895 10345 -890
rect 10605 -860 10645 -855
rect 10605 -890 10610 -860
rect 10610 -890 10640 -860
rect 10640 -890 10645 -860
rect 10605 -895 10645 -890
rect 10905 -860 10945 -855
rect 10905 -890 10910 -860
rect 10910 -890 10940 -860
rect 10940 -890 10945 -860
rect 10905 -895 10945 -890
rect 11205 -860 11245 -855
rect 11205 -890 11210 -860
rect 11210 -890 11240 -860
rect 11240 -890 11245 -860
rect 11205 -895 11245 -890
rect 11505 -860 11545 -855
rect 11505 -890 11510 -860
rect 11510 -890 11540 -860
rect 11540 -890 11545 -860
rect 11505 -895 11545 -890
rect 11805 -860 11845 -855
rect 11805 -890 11810 -860
rect 11810 -890 11840 -860
rect 11840 -890 11845 -860
rect 11805 -895 11845 -890
rect 12105 -860 12145 -855
rect 12105 -890 12110 -860
rect 12110 -890 12140 -860
rect 12140 -890 12145 -860
rect 12105 -895 12145 -890
rect 12405 -860 12445 -855
rect 12405 -890 12410 -860
rect 12410 -890 12440 -860
rect 12440 -890 12445 -860
rect 12405 -895 12445 -890
rect 12555 -860 12595 -855
rect 12555 -890 12560 -860
rect 12560 -890 12590 -860
rect 12590 -890 12595 -860
rect 12555 -895 12595 -890
rect 12705 -860 12745 -855
rect 12705 -890 12710 -860
rect 12710 -890 12740 -860
rect 12740 -890 12745 -860
rect 12705 -895 12745 -890
rect 13005 -860 13045 -855
rect 13005 -890 13010 -860
rect 13010 -890 13040 -860
rect 13040 -890 13045 -860
rect 13005 -895 13045 -890
rect 13305 -860 13345 -855
rect 13305 -890 13310 -860
rect 13310 -890 13340 -860
rect 13340 -890 13345 -860
rect 13305 -895 13345 -890
rect 13605 -860 13645 -855
rect 13605 -890 13610 -860
rect 13610 -890 13640 -860
rect 13640 -890 13645 -860
rect 13605 -895 13645 -890
rect 13755 -860 13795 -855
rect 13755 -890 13760 -860
rect 13760 -890 13790 -860
rect 13790 -890 13795 -860
rect 13755 -895 13795 -890
rect 13905 -860 13945 -855
rect 13905 -890 13910 -860
rect 13910 -890 13940 -860
rect 13940 -890 13945 -860
rect 13905 -895 13945 -890
rect 14205 -860 14245 -855
rect 14205 -890 14210 -860
rect 14210 -890 14240 -860
rect 14240 -890 14245 -860
rect 14205 -895 14245 -890
rect 14505 -860 14545 -855
rect 14505 -890 14510 -860
rect 14510 -890 14540 -860
rect 14540 -890 14545 -860
rect 14505 -895 14545 -890
rect 14805 -860 14845 -855
rect 14805 -890 14810 -860
rect 14810 -890 14840 -860
rect 14840 -890 14845 -860
rect 14805 -895 14845 -890
rect 15105 -860 15145 -855
rect 15105 -890 15110 -860
rect 15110 -890 15140 -860
rect 15140 -890 15145 -860
rect 15105 -895 15145 -890
rect 15405 -860 15445 -855
rect 15405 -890 15410 -860
rect 15410 -890 15440 -860
rect 15440 -890 15445 -860
rect 15405 -895 15445 -890
rect 15705 -860 15745 -855
rect 15705 -890 15710 -860
rect 15710 -890 15740 -860
rect 15740 -890 15745 -860
rect 15705 -895 15745 -890
rect 16005 -860 16045 -855
rect 16005 -890 16010 -860
rect 16010 -890 16040 -860
rect 16040 -890 16045 -860
rect 16005 -895 16045 -890
rect 16305 -860 16345 -855
rect 16305 -890 16310 -860
rect 16310 -890 16340 -860
rect 16340 -890 16345 -860
rect 16305 -895 16345 -890
rect 16605 -860 16645 -855
rect 16605 -890 16610 -860
rect 16610 -890 16640 -860
rect 16640 -890 16645 -860
rect 16605 -895 16645 -890
rect 16755 -860 16795 -855
rect 16755 -890 16760 -860
rect 16760 -890 16790 -860
rect 16790 -890 16795 -860
rect 16755 -895 16795 -890
rect 16905 -860 16945 -855
rect 16905 -890 16910 -860
rect 16910 -890 16940 -860
rect 16940 -890 16945 -860
rect 16905 -895 16945 -890
rect 17205 -860 17245 -855
rect 17205 -890 17210 -860
rect 17210 -890 17240 -860
rect 17240 -890 17245 -860
rect 17205 -895 17245 -890
rect 17505 -860 17545 -855
rect 17505 -890 17510 -860
rect 17510 -890 17540 -860
rect 17540 -890 17545 -860
rect 17505 -895 17545 -890
rect 17805 -860 17845 -855
rect 17805 -890 17810 -860
rect 17810 -890 17840 -860
rect 17840 -890 17845 -860
rect 17805 -895 17845 -890
rect 18105 -860 18145 -855
rect 18105 -890 18110 -860
rect 18110 -890 18140 -860
rect 18140 -890 18145 -860
rect 18105 -895 18145 -890
rect 18405 -860 18445 -855
rect 18405 -890 18410 -860
rect 18410 -890 18440 -860
rect 18440 -890 18445 -860
rect 18405 -895 18445 -890
rect 18705 -860 18745 -855
rect 18705 -890 18710 -860
rect 18710 -890 18740 -860
rect 18740 -890 18745 -860
rect 18705 -895 18745 -890
rect 19005 -860 19045 -855
rect 19005 -890 19010 -860
rect 19010 -890 19040 -860
rect 19040 -890 19045 -860
rect 19005 -895 19045 -890
rect 19155 -860 19195 -855
rect 19155 -890 19160 -860
rect 19160 -890 19190 -860
rect 19190 -890 19195 -860
rect 19155 -895 19195 -890
rect 19305 -860 19345 -855
rect 19305 -890 19310 -860
rect 19310 -890 19340 -860
rect 19340 -890 19345 -860
rect 19305 -895 19345 -890
rect 19605 -860 19645 -855
rect 19605 -890 19610 -860
rect 19610 -890 19640 -860
rect 19640 -890 19645 -860
rect 19605 -895 19645 -890
rect 19905 -860 19945 -855
rect 19905 -890 19910 -860
rect 19910 -890 19940 -860
rect 19940 -890 19945 -860
rect 19905 -895 19945 -890
rect 20205 -860 20245 -855
rect 20205 -890 20210 -860
rect 20210 -890 20240 -860
rect 20240 -890 20245 -860
rect 20205 -895 20245 -890
rect 20505 -860 20545 -855
rect 20505 -890 20510 -860
rect 20510 -890 20540 -860
rect 20540 -890 20545 -860
rect 20505 -895 20545 -890
rect 20805 -860 20845 -855
rect 20805 -890 20810 -860
rect 20810 -890 20840 -860
rect 20840 -890 20845 -860
rect 20805 -895 20845 -890
rect 21105 -860 21145 -855
rect 21105 -890 21110 -860
rect 21110 -890 21140 -860
rect 21140 -890 21145 -860
rect 21105 -895 21145 -890
rect 21405 -860 21445 -855
rect 21405 -890 21410 -860
rect 21410 -890 21440 -860
rect 21440 -890 21445 -860
rect 21405 -895 21445 -890
rect 21705 -860 21745 -855
rect 21705 -890 21710 -860
rect 21710 -890 21740 -860
rect 21740 -890 21745 -860
rect 21705 -895 21745 -890
rect 22005 -860 22045 -855
rect 22005 -890 22010 -860
rect 22010 -890 22040 -860
rect 22040 -890 22045 -860
rect 22005 -895 22045 -890
rect 22305 -860 22345 -855
rect 22305 -890 22310 -860
rect 22310 -890 22340 -860
rect 22340 -890 22345 -860
rect 22305 -895 22345 -890
rect 22455 -860 22495 -855
rect 22455 -890 22460 -860
rect 22460 -890 22490 -860
rect 22490 -890 22495 -860
rect 22455 -895 22495 -890
rect 22605 -860 22645 -855
rect 22605 -890 22610 -860
rect 22610 -890 22640 -860
rect 22640 -890 22645 -860
rect 22605 -895 22645 -890
rect 22905 -860 22945 -855
rect 22905 -890 22910 -860
rect 22910 -890 22940 -860
rect 22940 -890 22945 -860
rect 22905 -895 22945 -890
rect 23205 -860 23245 -855
rect 23205 -890 23210 -860
rect 23210 -890 23240 -860
rect 23240 -890 23245 -860
rect 23205 -895 23245 -890
rect 23505 -860 23545 -855
rect 23505 -890 23510 -860
rect 23510 -890 23540 -860
rect 23540 -890 23545 -860
rect 23505 -895 23545 -890
rect 23805 -860 23845 -855
rect 23805 -890 23810 -860
rect 23810 -890 23840 -860
rect 23840 -890 23845 -860
rect 23805 -895 23845 -890
rect 24105 -860 24145 -855
rect 24105 -890 24110 -860
rect 24110 -890 24140 -860
rect 24140 -890 24145 -860
rect 24105 -895 24145 -890
rect 24405 -860 24445 -855
rect 24405 -890 24410 -860
rect 24410 -890 24440 -860
rect 24440 -890 24445 -860
rect 24405 -895 24445 -890
rect 24705 -860 24745 -855
rect 24705 -890 24710 -860
rect 24710 -890 24740 -860
rect 24740 -890 24745 -860
rect 24705 -895 24745 -890
rect 25005 -860 25045 -855
rect 25005 -890 25010 -860
rect 25010 -890 25040 -860
rect 25040 -890 25045 -860
rect 25005 -895 25045 -890
rect 25305 -860 25345 -855
rect 25305 -890 25310 -860
rect 25310 -890 25340 -860
rect 25340 -890 25345 -860
rect 25305 -895 25345 -890
rect 25605 -860 25645 -855
rect 25605 -890 25610 -860
rect 25610 -890 25640 -860
rect 25640 -890 25645 -860
rect 25605 -895 25645 -890
rect 25755 -860 25795 -855
rect 25755 -890 25760 -860
rect 25760 -890 25790 -860
rect 25790 -890 25795 -860
rect 25755 -895 25795 -890
rect 25905 -860 25945 -855
rect 25905 -890 25910 -860
rect 25910 -890 25940 -860
rect 25940 -890 25945 -860
rect 25905 -895 25945 -890
rect 26205 -860 26245 -855
rect 26205 -890 26210 -860
rect 26210 -890 26240 -860
rect 26240 -890 26245 -860
rect 26205 -895 26245 -890
rect 26505 -860 26545 -855
rect 26505 -890 26510 -860
rect 26510 -890 26540 -860
rect 26540 -890 26545 -860
rect 26505 -895 26545 -890
rect 26655 -860 26695 -855
rect 26655 -890 26660 -860
rect 26660 -890 26690 -860
rect 26690 -890 26695 -860
rect 26655 -895 26695 -890
rect 26805 -860 26845 -855
rect 26805 -890 26810 -860
rect 26810 -890 26840 -860
rect 26840 -890 26845 -860
rect 26805 -895 26845 -890
rect 27105 -860 27145 -855
rect 27105 -890 27110 -860
rect 27110 -890 27140 -860
rect 27140 -890 27145 -860
rect 27105 -895 27145 -890
rect 27405 -860 27445 -855
rect 27405 -890 27410 -860
rect 27410 -890 27440 -860
rect 27440 -890 27445 -860
rect 27405 -895 27445 -890
rect 27555 -860 27595 -855
rect 27555 -890 27560 -860
rect 27560 -890 27590 -860
rect 27590 -890 27595 -860
rect 27555 -895 27595 -890
rect 27705 -860 27745 -855
rect 27705 -890 27710 -860
rect 27710 -890 27740 -860
rect 27740 -890 27745 -860
rect 27705 -895 27745 -890
rect 28005 -860 28045 -855
rect 28005 -890 28010 -860
rect 28010 -890 28040 -860
rect 28040 -890 28045 -860
rect 28005 -895 28045 -890
rect 28305 -860 28345 -855
rect 28305 -890 28310 -860
rect 28310 -890 28340 -860
rect 28340 -890 28345 -860
rect 28305 -895 28345 -890
rect 28605 -860 28645 -855
rect 28605 -890 28610 -860
rect 28610 -890 28640 -860
rect 28640 -890 28645 -860
rect 28605 -895 28645 -890
<< metal4 >>
rect -500 4945 -450 4950
rect -500 4905 -495 4945
rect -455 4905 -450 4945
rect -500 3645 -450 4905
rect -500 3605 -495 3645
rect -455 3605 -450 3645
rect -500 3145 -450 3605
rect -350 4945 -300 5000
rect -350 4905 -345 4945
rect -305 4905 -300 4945
rect -350 3645 -300 4905
rect -350 3605 -345 3645
rect -305 3605 -300 3645
rect -350 3445 -300 3605
rect -350 3405 -345 3445
rect -305 3405 -300 3445
rect -350 3400 -300 3405
rect -200 4945 -150 4950
rect -200 4905 -195 4945
rect -155 4905 -150 4945
rect -200 3645 -150 4905
rect -200 3605 -195 3645
rect -155 3605 -150 3645
rect -500 3105 -495 3145
rect -455 3105 -450 3145
rect -500 3100 -450 3105
rect -200 3145 -150 3605
rect 100 4945 150 4950
rect 100 4905 105 4945
rect 145 4905 150 4945
rect 100 3645 150 4905
rect 100 3605 105 3645
rect 145 3605 150 3645
rect 100 3445 150 3605
rect 100 3405 105 3445
rect 145 3405 150 3445
rect 100 3400 150 3405
rect 400 4945 450 4950
rect 400 4905 405 4945
rect 445 4905 450 4945
rect 400 3645 450 4905
rect 400 3605 405 3645
rect 445 3605 450 3645
rect 400 3445 450 3605
rect 400 3405 405 3445
rect 445 3405 450 3445
rect 400 3400 450 3405
rect 700 4945 750 4950
rect 700 4905 705 4945
rect 745 4905 750 4945
rect 700 3645 750 4905
rect 700 3605 705 3645
rect 745 3605 750 3645
rect 700 3345 750 3605
rect 700 3305 705 3345
rect 745 3305 750 3345
rect 700 3300 750 3305
rect 1000 4945 1050 4950
rect 1000 4905 1005 4945
rect 1045 4905 1050 4945
rect 1000 3645 1050 4905
rect 1000 3605 1005 3645
rect 1045 3605 1050 3645
rect 1000 3345 1050 3605
rect 1000 3305 1005 3345
rect 1045 3305 1050 3345
rect 1000 3300 1050 3305
rect 1150 4945 1200 4950
rect 1150 4905 1155 4945
rect 1195 4905 1200 4945
rect 1150 3645 1200 4905
rect 1150 3605 1155 3645
rect 1195 3605 1200 3645
rect 1150 3345 1200 3605
rect 1150 3305 1155 3345
rect 1195 3305 1200 3345
rect 1150 3300 1200 3305
rect 1300 4945 1350 4950
rect 1300 4905 1305 4945
rect 1345 4905 1350 4945
rect 1300 3645 1350 4905
rect 1300 3605 1305 3645
rect 1345 3605 1350 3645
rect 1300 3345 1350 3605
rect 1300 3305 1305 3345
rect 1345 3305 1350 3345
rect 1300 3300 1350 3305
rect 1600 4945 1650 4950
rect 1600 4905 1605 4945
rect 1645 4905 1650 4945
rect 1600 3645 1650 4905
rect 1600 3605 1605 3645
rect 1645 3605 1650 3645
rect 1600 3345 1650 3605
rect 1600 3305 1605 3345
rect 1645 3305 1650 3345
rect 1600 3300 1650 3305
rect 1900 4945 1950 4950
rect 1900 4905 1905 4945
rect 1945 4905 1950 4945
rect 1900 3645 1950 4905
rect 1900 3605 1905 3645
rect 1945 3605 1950 3645
rect 1900 3245 1950 3605
rect 2050 4945 2100 4950
rect 2050 4905 2055 4945
rect 2095 4905 2100 4945
rect 2050 3645 2100 4905
rect 2050 3605 2055 3645
rect 2095 3605 2100 3645
rect 2050 3445 2100 3605
rect 2050 3405 2055 3445
rect 2095 3405 2100 3445
rect 2050 3400 2100 3405
rect 2200 4945 2250 4950
rect 2200 4905 2205 4945
rect 2245 4905 2250 4945
rect 2200 3645 2250 4905
rect 2200 3605 2205 3645
rect 2245 3605 2250 3645
rect 1900 3205 1905 3245
rect 1945 3205 1950 3245
rect 1900 3200 1950 3205
rect 2200 3245 2250 3605
rect 2500 4945 2550 4950
rect 2500 4905 2505 4945
rect 2545 4905 2550 4945
rect 2500 3645 2550 4905
rect 2500 3605 2505 3645
rect 2545 3605 2550 3645
rect 2500 3345 2550 3605
rect 2500 3305 2505 3345
rect 2545 3305 2550 3345
rect 2500 3300 2550 3305
rect 2800 4945 2850 4950
rect 2800 4905 2805 4945
rect 2845 4905 2850 4945
rect 2800 3645 2850 4905
rect 2800 3605 2805 3645
rect 2845 3605 2850 3645
rect 2800 3345 2850 3605
rect 2800 3305 2805 3345
rect 2845 3305 2850 3345
rect 2800 3300 2850 3305
rect 2950 4945 3000 4950
rect 2950 4905 2955 4945
rect 2995 4905 3000 4945
rect 2950 3645 3000 4905
rect 2950 3605 2955 3645
rect 2995 3605 3000 3645
rect 2950 3345 3000 3605
rect 2950 3305 2955 3345
rect 2995 3305 3000 3345
rect 2950 3300 3000 3305
rect 3100 4945 3150 4950
rect 3100 4905 3105 4945
rect 3145 4905 3150 4945
rect 3100 3645 3150 4905
rect 3100 3605 3105 3645
rect 3145 3605 3150 3645
rect 3100 3345 3150 3605
rect 3100 3305 3105 3345
rect 3145 3305 3150 3345
rect 3100 3300 3150 3305
rect 3400 4945 3450 4950
rect 3400 4905 3405 4945
rect 3445 4905 3450 4945
rect 3400 3645 3450 4905
rect 3400 3605 3405 3645
rect 3445 3605 3450 3645
rect 3400 3345 3450 3605
rect 3700 4945 3750 4950
rect 3700 4905 3705 4945
rect 3745 4905 3750 4945
rect 3700 3645 3750 4905
rect 3700 3605 3705 3645
rect 3745 3605 3750 3645
rect 3700 3445 3750 3605
rect 3700 3405 3705 3445
rect 3745 3405 3750 3445
rect 3700 3400 3750 3405
rect 4000 4945 4050 4950
rect 4000 4905 4005 4945
rect 4045 4905 4050 4945
rect 4000 3645 4050 4905
rect 4000 3605 4005 3645
rect 4045 3605 4050 3645
rect 4000 3445 4050 3605
rect 4000 3405 4005 3445
rect 4045 3405 4050 3445
rect 4000 3400 4050 3405
rect 4300 4945 4350 4950
rect 4300 4905 4305 4945
rect 4345 4905 4350 4945
rect 4300 3645 4350 4905
rect 4300 3605 4305 3645
rect 4345 3605 4350 3645
rect 4300 3445 4350 3605
rect 4300 3405 4305 3445
rect 4345 3405 4350 3445
rect 4300 3400 4350 3405
rect 4600 4945 4650 4950
rect 4600 4905 4605 4945
rect 4645 4905 4650 4945
rect 4600 3645 4650 4905
rect 4600 3605 4605 3645
rect 4645 3605 4650 3645
rect 4600 3445 4650 3605
rect 4600 3405 4605 3445
rect 4645 3405 4650 3445
rect 4600 3400 4650 3405
rect 4900 4945 4950 4950
rect 4900 4905 4905 4945
rect 4945 4905 4950 4945
rect 4900 3645 4950 4905
rect 4900 3605 4905 3645
rect 4945 3605 4950 3645
rect 3400 3305 3405 3345
rect 3445 3305 3450 3345
rect 3400 3300 3450 3305
rect 4900 3345 4950 3605
rect 4900 3305 4905 3345
rect 4945 3305 4950 3345
rect 4900 3300 4950 3305
rect 5200 4945 5250 4950
rect 5200 4905 5205 4945
rect 5245 4905 5250 4945
rect 5200 3645 5250 4905
rect 5200 3605 5205 3645
rect 5245 3605 5250 3645
rect 5200 3345 5250 3605
rect 5200 3305 5205 3345
rect 5245 3305 5250 3345
rect 5200 3300 5250 3305
rect 5350 4945 5400 4950
rect 5350 4905 5355 4945
rect 5395 4905 5400 4945
rect 5350 3645 5400 4905
rect 5350 3605 5355 3645
rect 5395 3605 5400 3645
rect 5350 3345 5400 3605
rect 5350 3305 5355 3345
rect 5395 3305 5400 3345
rect 5350 3300 5400 3305
rect 5500 4945 5550 4950
rect 5500 4905 5505 4945
rect 5545 4905 5550 4945
rect 5500 3645 5550 4905
rect 5500 3605 5505 3645
rect 5545 3605 5550 3645
rect 5500 3345 5550 3605
rect 5500 3305 5505 3345
rect 5545 3305 5550 3345
rect 5500 3300 5550 3305
rect 5800 4945 5850 4950
rect 5800 4905 5805 4945
rect 5845 4905 5850 4945
rect 5800 3645 5850 4905
rect 5800 3605 5805 3645
rect 5845 3605 5850 3645
rect 5800 3345 5850 3605
rect 5800 3305 5805 3345
rect 5845 3305 5850 3345
rect 5800 3300 5850 3305
rect 6100 4945 6150 4950
rect 6100 4905 6105 4945
rect 6145 4905 6150 4945
rect 6100 3645 6150 4905
rect 6100 3605 6105 3645
rect 6145 3605 6150 3645
rect 2200 3205 2205 3245
rect 2245 3205 2250 3245
rect 2200 3200 2250 3205
rect 6100 3245 6150 3605
rect 6250 4945 6300 4950
rect 6250 4905 6255 4945
rect 6295 4905 6300 4945
rect 6250 3645 6300 4905
rect 6250 3605 6255 3645
rect 6295 3605 6300 3645
rect 6250 3445 6300 3605
rect 6250 3405 6255 3445
rect 6295 3405 6300 3445
rect 6250 3400 6300 3405
rect 6400 4945 6450 4950
rect 6400 4905 6405 4945
rect 6445 4905 6450 4945
rect 6400 3645 6450 4905
rect 6400 3605 6405 3645
rect 6445 3605 6450 3645
rect 6100 3205 6105 3245
rect 6145 3205 6150 3245
rect 6100 3200 6150 3205
rect 6400 3245 6450 3605
rect 6700 4945 6750 4950
rect 6700 4905 6705 4945
rect 6745 4905 6750 4945
rect 6700 3645 6750 4905
rect 6700 3605 6705 3645
rect 6745 3605 6750 3645
rect 6700 3345 6750 3605
rect 6700 3305 6705 3345
rect 6745 3305 6750 3345
rect 6700 3300 6750 3305
rect 7000 4945 7050 4950
rect 7000 4905 7005 4945
rect 7045 4905 7050 4945
rect 7000 3645 7050 4905
rect 7000 3605 7005 3645
rect 7045 3605 7050 3645
rect 7000 3345 7050 3605
rect 7000 3305 7005 3345
rect 7045 3305 7050 3345
rect 7000 3300 7050 3305
rect 7150 4945 7200 4950
rect 7150 4905 7155 4945
rect 7195 4905 7200 4945
rect 7150 3645 7200 4905
rect 7150 3605 7155 3645
rect 7195 3605 7200 3645
rect 7150 3345 7200 3605
rect 7150 3305 7155 3345
rect 7195 3305 7200 3345
rect 7150 3300 7200 3305
rect 7300 4945 7350 4950
rect 7300 4905 7305 4945
rect 7345 4905 7350 4945
rect 7300 3645 7350 4905
rect 7300 3605 7305 3645
rect 7345 3605 7350 3645
rect 7300 3345 7350 3605
rect 7300 3305 7305 3345
rect 7345 3305 7350 3345
rect 7300 3300 7350 3305
rect 7600 4945 7650 4950
rect 7600 4905 7605 4945
rect 7645 4905 7650 4945
rect 7600 3645 7650 4905
rect 7600 3605 7605 3645
rect 7645 3605 7650 3645
rect 7600 3345 7650 3605
rect 7900 4945 7950 4950
rect 7900 4905 7905 4945
rect 7945 4905 7950 4945
rect 7900 3645 7950 4905
rect 7900 3605 7905 3645
rect 7945 3605 7950 3645
rect 7900 3445 7950 3605
rect 7900 3405 7905 3445
rect 7945 3405 7950 3445
rect 7900 3400 7950 3405
rect 8200 4945 8250 4950
rect 8200 4905 8205 4945
rect 8245 4905 8250 4945
rect 8200 3645 8250 4905
rect 8200 3605 8205 3645
rect 8245 3605 8250 3645
rect 8200 3445 8250 3605
rect 8500 4945 8550 4950
rect 8500 4905 8505 4945
rect 8545 4905 8550 4945
rect 8500 3645 8550 4905
rect 8500 3605 8505 3645
rect 8545 3605 8550 3645
rect 8500 3600 8550 3605
rect 8800 4945 8850 4950
rect 8800 4905 8805 4945
rect 8845 4905 8850 4945
rect 8800 3645 8850 4905
rect 8800 3605 8805 3645
rect 8845 3605 8850 3645
rect 8800 3600 8850 3605
rect 9100 4945 9150 4950
rect 9100 4905 9105 4945
rect 9145 4905 9150 4945
rect 9100 3645 9150 4905
rect 9100 3605 9105 3645
rect 9145 3605 9150 3645
rect 9100 3600 9150 3605
rect 9400 4945 9450 4950
rect 9400 4905 9405 4945
rect 9445 4905 9450 4945
rect 9400 3645 9450 4905
rect 9400 3605 9405 3645
rect 9445 3605 9450 3645
rect 9400 3600 9450 3605
rect 9700 4945 9750 4950
rect 9700 4905 9705 4945
rect 9745 4905 9750 4945
rect 9700 3645 9750 4905
rect 9700 3605 9705 3645
rect 9745 3605 9750 3645
rect 9700 3600 9750 3605
rect 10000 4945 10050 4950
rect 10000 4905 10005 4945
rect 10045 4905 10050 4945
rect 10000 3645 10050 4905
rect 10000 3605 10005 3645
rect 10045 3605 10050 3645
rect 10000 3600 10050 3605
rect 10300 4945 10350 4950
rect 10300 4905 10305 4945
rect 10345 4905 10350 4945
rect 10300 3645 10350 4905
rect 10300 3605 10305 3645
rect 10345 3605 10350 3645
rect 10300 3600 10350 3605
rect 10600 4945 10650 4950
rect 10600 4905 10605 4945
rect 10645 4905 10650 4945
rect 10600 3645 10650 4905
rect 10600 3605 10605 3645
rect 10645 3605 10650 3645
rect 10600 3600 10650 3605
rect 10900 4945 10950 4950
rect 10900 4905 10905 4945
rect 10945 4905 10950 4945
rect 10900 3845 10950 4905
rect 10900 3805 10905 3845
rect 10945 3805 10950 3845
rect 10900 3645 10950 3805
rect 10900 3605 10905 3645
rect 10945 3605 10950 3645
rect 10900 3600 10950 3605
rect 11200 4945 11250 4950
rect 11200 4905 11205 4945
rect 11245 4905 11250 4945
rect 11200 3845 11250 4905
rect 11200 3805 11205 3845
rect 11245 3805 11250 3845
rect 11200 3645 11250 3805
rect 11200 3605 11205 3645
rect 11245 3605 11250 3645
rect 11200 3600 11250 3605
rect 11350 4945 11400 4950
rect 11350 4905 11355 4945
rect 11395 4905 11400 4945
rect 11350 4545 11400 4905
rect 11350 4505 11355 4545
rect 11395 4505 11400 4545
rect 11350 3645 11400 4505
rect 11350 3605 11355 3645
rect 11395 3605 11400 3645
rect 11350 3600 11400 3605
rect 11500 4945 11550 4950
rect 11500 4905 11505 4945
rect 11545 4905 11550 4945
rect 11500 3845 11550 4905
rect 11500 3805 11505 3845
rect 11545 3805 11550 3845
rect 11500 3645 11550 3805
rect 11500 3605 11505 3645
rect 11545 3605 11550 3645
rect 11500 3600 11550 3605
rect 11800 4945 11850 4950
rect 11800 4905 11805 4945
rect 11845 4905 11850 4945
rect 11800 3845 11850 4905
rect 11800 3805 11805 3845
rect 11845 3805 11850 3845
rect 11800 3645 11850 3805
rect 11800 3605 11805 3645
rect 11845 3605 11850 3645
rect 11800 3600 11850 3605
rect 12100 4945 12150 4950
rect 12100 4905 12105 4945
rect 12145 4905 12150 4945
rect 12100 3845 12150 4905
rect 12100 3805 12105 3845
rect 12145 3805 12150 3845
rect 12100 3645 12150 3805
rect 12100 3605 12105 3645
rect 12145 3605 12150 3645
rect 12100 3600 12150 3605
rect 12400 4945 12450 4950
rect 12400 4905 12405 4945
rect 12445 4905 12450 4945
rect 12400 3845 12450 4905
rect 12550 4945 12600 4950
rect 12550 4905 12555 4945
rect 12595 4905 12600 4945
rect 12550 4900 12600 4905
rect 12700 4945 12750 4950
rect 12700 4905 12705 4945
rect 12745 4905 12750 4945
rect 12400 3805 12405 3845
rect 12445 3805 12450 3845
rect 12400 3645 12450 3805
rect 12400 3605 12405 3645
rect 12445 3605 12450 3645
rect 12400 3600 12450 3605
rect 12550 4545 12600 4550
rect 12550 4505 12555 4545
rect 12595 4505 12600 4545
rect 12550 3645 12600 4505
rect 12550 3605 12555 3645
rect 12595 3605 12600 3645
rect 8200 3405 8205 3445
rect 8245 3405 8250 3445
rect 8200 3400 8250 3405
rect 7600 3305 7605 3345
rect 7645 3305 7650 3345
rect 7600 3300 7650 3305
rect 9550 3345 9600 3350
rect 9550 3305 9555 3345
rect 9595 3305 9600 3345
rect 6400 3205 6405 3245
rect 6445 3205 6450 3245
rect 6400 3200 6450 3205
rect -200 3105 -195 3145
rect -155 3105 -150 3145
rect -200 3100 -150 3105
rect -500 1345 -450 1350
rect -500 1305 -495 1345
rect -455 1305 -450 1345
rect -500 845 -450 1305
rect -200 1345 -150 1350
rect -200 1305 -195 1345
rect -155 1305 -150 1345
rect -500 805 -495 845
rect -455 805 -450 845
rect -500 -855 -450 805
rect -500 -895 -495 -855
rect -455 -895 -450 -855
rect -500 -900 -450 -895
rect -350 1045 -300 1050
rect -350 1005 -345 1045
rect -305 1005 -300 1045
rect -350 845 -300 1005
rect -350 805 -345 845
rect -305 805 -300 845
rect -350 -855 -300 805
rect -350 -895 -345 -855
rect -305 -895 -300 -855
rect -350 -950 -300 -895
rect -200 845 -150 1305
rect 3700 1245 3750 1250
rect 3700 1205 3705 1245
rect 3745 1205 3750 1245
rect 1300 1145 1350 1150
rect 1300 1105 1305 1145
rect 1345 1105 1350 1145
rect -200 805 -195 845
rect -155 805 -150 845
rect -200 -855 -150 805
rect -200 -895 -195 -855
rect -155 -895 -150 -855
rect -200 -900 -150 -895
rect 100 1045 150 1050
rect 100 1005 105 1045
rect 145 1005 150 1045
rect 100 845 150 1005
rect 100 805 105 845
rect 145 805 150 845
rect 100 -855 150 805
rect 100 -895 105 -855
rect 145 -895 150 -855
rect 100 -900 150 -895
rect 400 1045 450 1050
rect 400 1005 405 1045
rect 445 1005 450 1045
rect 400 845 450 1005
rect 400 805 405 845
rect 445 805 450 845
rect 400 -855 450 805
rect 400 -895 405 -855
rect 445 -895 450 -855
rect 400 -900 450 -895
rect 700 1045 750 1050
rect 700 1005 705 1045
rect 745 1005 750 1045
rect 700 845 750 1005
rect 700 805 705 845
rect 745 805 750 845
rect 700 -855 750 805
rect 700 -895 705 -855
rect 745 -895 750 -855
rect 700 -900 750 -895
rect 1000 1045 1050 1050
rect 1000 1005 1005 1045
rect 1045 1005 1050 1045
rect 1000 845 1050 1005
rect 1000 805 1005 845
rect 1045 805 1050 845
rect 1000 -855 1050 805
rect 1000 -895 1005 -855
rect 1045 -895 1050 -855
rect 1000 -900 1050 -895
rect 1300 845 1350 1105
rect 1300 805 1305 845
rect 1345 805 1350 845
rect 1300 -855 1350 805
rect 1300 -895 1305 -855
rect 1345 -895 1350 -855
rect 1300 -900 1350 -895
rect 1600 1145 1650 1150
rect 1600 1105 1605 1145
rect 1645 1105 1650 1145
rect 1600 845 1650 1105
rect 1600 805 1605 845
rect 1645 805 1650 845
rect 1600 -855 1650 805
rect 1600 -895 1605 -855
rect 1645 -895 1650 -855
rect 1600 -900 1650 -895
rect 1900 1145 1950 1150
rect 1900 1105 1905 1145
rect 1945 1105 1950 1145
rect 1900 845 1950 1105
rect 1900 805 1905 845
rect 1945 805 1950 845
rect 1900 -855 1950 805
rect 1900 -895 1905 -855
rect 1945 -895 1950 -855
rect 1900 -900 1950 -895
rect 2200 1145 2250 1150
rect 2200 1105 2205 1145
rect 2245 1105 2250 1145
rect 2200 845 2250 1105
rect 2200 805 2205 845
rect 2245 805 2250 845
rect 2200 -855 2250 805
rect 2200 -895 2205 -855
rect 2245 -895 2250 -855
rect 2200 -900 2250 -895
rect 2350 1145 2400 1150
rect 2350 1105 2355 1145
rect 2395 1105 2400 1145
rect 2350 845 2400 1105
rect 2350 805 2355 845
rect 2395 805 2400 845
rect 2350 -855 2400 805
rect 2350 -895 2355 -855
rect 2395 -895 2400 -855
rect 2350 -900 2400 -895
rect 2500 1145 2550 1150
rect 2500 1105 2505 1145
rect 2545 1105 2550 1145
rect 2500 845 2550 1105
rect 2500 805 2505 845
rect 2545 805 2550 845
rect 2500 -855 2550 805
rect 2500 -895 2505 -855
rect 2545 -895 2550 -855
rect 2500 -900 2550 -895
rect 2800 1145 2850 1150
rect 2800 1105 2805 1145
rect 2845 1105 2850 1145
rect 2800 845 2850 1105
rect 2800 805 2805 845
rect 2845 805 2850 845
rect 2800 -855 2850 805
rect 2800 -895 2805 -855
rect 2845 -895 2850 -855
rect 2800 -900 2850 -895
rect 3100 1145 3150 1150
rect 3100 1105 3105 1145
rect 3145 1105 3150 1145
rect 3100 845 3150 1105
rect 3100 805 3105 845
rect 3145 805 3150 845
rect 3100 -855 3150 805
rect 3100 -895 3105 -855
rect 3145 -895 3150 -855
rect 3100 -900 3150 -895
rect 3400 1145 3450 1150
rect 3400 1105 3405 1145
rect 3445 1105 3450 1145
rect 3400 845 3450 1105
rect 3400 805 3405 845
rect 3445 805 3450 845
rect 3400 -855 3450 805
rect 3400 -895 3405 -855
rect 3445 -895 3450 -855
rect 3400 -900 3450 -895
rect 3700 845 3750 1205
rect 4000 1245 4050 1250
rect 4000 1205 4005 1245
rect 4045 1205 4050 1245
rect 3700 805 3705 845
rect 3745 805 3750 845
rect 3700 -855 3750 805
rect 3700 -895 3705 -855
rect 3745 -895 3750 -855
rect 3700 -900 3750 -895
rect 3850 1045 3900 1050
rect 3850 1005 3855 1045
rect 3895 1005 3900 1045
rect 3850 845 3900 1005
rect 3850 805 3855 845
rect 3895 805 3900 845
rect 3850 -855 3900 805
rect 3850 -895 3855 -855
rect 3895 -895 3900 -855
rect 3850 -900 3900 -895
rect 4000 845 4050 1205
rect 4000 805 4005 845
rect 4045 805 4050 845
rect 4000 -855 4050 805
rect 4000 -895 4005 -855
rect 4045 -895 4050 -855
rect 4000 -900 4050 -895
rect 4300 1245 4350 1250
rect 4300 1205 4305 1245
rect 4345 1205 4350 1245
rect 4300 845 4350 1205
rect 4600 1245 4650 1250
rect 4600 1205 4605 1245
rect 4645 1205 4650 1245
rect 4300 805 4305 845
rect 4345 805 4350 845
rect 4300 -855 4350 805
rect 4300 -895 4305 -855
rect 4345 -895 4350 -855
rect 4300 -900 4350 -895
rect 4450 1045 4500 1050
rect 4450 1005 4455 1045
rect 4495 1005 4500 1045
rect 4450 845 4500 1005
rect 4450 805 4455 845
rect 4495 805 4500 845
rect 4450 -855 4500 805
rect 4450 -895 4455 -855
rect 4495 -895 4500 -855
rect 4450 -900 4500 -895
rect 4600 845 4650 1205
rect 4600 805 4605 845
rect 4645 805 4650 845
rect 4600 -855 4650 805
rect 4600 -895 4605 -855
rect 4645 -895 4650 -855
rect 4600 -900 4650 -895
rect 4900 1145 4950 1150
rect 4900 1105 4905 1145
rect 4945 1105 4950 1145
rect 4900 845 4950 1105
rect 4900 805 4905 845
rect 4945 805 4950 845
rect 4900 -855 4950 805
rect 4900 -895 4905 -855
rect 4945 -895 4950 -855
rect 4900 -900 4950 -895
rect 5200 1145 5250 1150
rect 5200 1105 5205 1145
rect 5245 1105 5250 1145
rect 5200 845 5250 1105
rect 5200 805 5205 845
rect 5245 805 5250 845
rect 5200 -855 5250 805
rect 5200 -895 5205 -855
rect 5245 -895 5250 -855
rect 5200 -900 5250 -895
rect 5500 1145 5550 1150
rect 5500 1105 5505 1145
rect 5545 1105 5550 1145
rect 5500 845 5550 1105
rect 5500 805 5505 845
rect 5545 805 5550 845
rect 5500 -855 5550 805
rect 5500 -895 5505 -855
rect 5545 -895 5550 -855
rect 5500 -900 5550 -895
rect 5800 1145 5850 1150
rect 5800 1105 5805 1145
rect 5845 1105 5850 1145
rect 5800 845 5850 1105
rect 5800 805 5805 845
rect 5845 805 5850 845
rect 5800 -855 5850 805
rect 5800 -895 5805 -855
rect 5845 -895 5850 -855
rect 5800 -900 5850 -895
rect 5950 1145 6000 1150
rect 5950 1105 5955 1145
rect 5995 1105 6000 1145
rect 5950 845 6000 1105
rect 5950 805 5955 845
rect 5995 805 6000 845
rect 5950 -855 6000 805
rect 5950 -895 5955 -855
rect 5995 -895 6000 -855
rect 5950 -900 6000 -895
rect 6100 1145 6150 1150
rect 6100 1105 6105 1145
rect 6145 1105 6150 1145
rect 6100 845 6150 1105
rect 6100 805 6105 845
rect 6145 805 6150 845
rect 6100 -855 6150 805
rect 6100 -895 6105 -855
rect 6145 -895 6150 -855
rect 6100 -900 6150 -895
rect 6400 1145 6450 1150
rect 6400 1105 6405 1145
rect 6445 1105 6450 1145
rect 6400 845 6450 1105
rect 6400 805 6405 845
rect 6445 805 6450 845
rect 6400 -855 6450 805
rect 6400 -895 6405 -855
rect 6445 -895 6450 -855
rect 6400 -900 6450 -895
rect 6700 1145 6750 1150
rect 6700 1105 6705 1145
rect 6745 1105 6750 1145
rect 6700 845 6750 1105
rect 6700 805 6705 845
rect 6745 805 6750 845
rect 6700 -855 6750 805
rect 6700 -895 6705 -855
rect 6745 -895 6750 -855
rect 6700 -900 6750 -895
rect 7000 1145 7050 1150
rect 7000 1105 7005 1145
rect 7045 1105 7050 1145
rect 7000 845 7050 1105
rect 7000 805 7005 845
rect 7045 805 7050 845
rect 7000 -855 7050 805
rect 7000 -895 7005 -855
rect 7045 -895 7050 -855
rect 7000 -900 7050 -895
rect 7300 1045 7350 1050
rect 7300 1005 7305 1045
rect 7345 1005 7350 1045
rect 7300 845 7350 1005
rect 7300 805 7305 845
rect 7345 805 7350 845
rect 7300 -855 7350 805
rect 7300 -895 7305 -855
rect 7345 -895 7350 -855
rect 7300 -900 7350 -895
rect 7600 1045 7650 1050
rect 7600 1005 7605 1045
rect 7645 1005 7650 1045
rect 7600 845 7650 1005
rect 7600 805 7605 845
rect 7645 805 7650 845
rect 7600 -855 7650 805
rect 7600 -895 7605 -855
rect 7645 -895 7650 -855
rect 7600 -900 7650 -895
rect 7900 1045 7950 1050
rect 7900 1005 7905 1045
rect 7945 1005 7950 1045
rect 7900 845 7950 1005
rect 7900 805 7905 845
rect 7945 805 7950 845
rect 7900 -855 7950 805
rect 7900 -895 7905 -855
rect 7945 -895 7950 -855
rect 7900 -900 7950 -895
rect 8200 1045 8250 1050
rect 8200 1005 8205 1045
rect 8245 1005 8250 1045
rect 8200 845 8250 1005
rect 8200 805 8205 845
rect 8245 805 8250 845
rect 8200 -855 8250 805
rect 8200 -895 8205 -855
rect 8245 -895 8250 -855
rect 8200 -900 8250 -895
rect 8500 1045 8550 1050
rect 8500 1005 8505 1045
rect 8545 1005 8550 1045
rect 8500 845 8550 1005
rect 8500 805 8505 845
rect 8545 805 8550 845
rect 8500 -855 8550 805
rect 8500 -895 8505 -855
rect 8545 -895 8550 -855
rect 8500 -900 8550 -895
rect 8800 1045 8850 1050
rect 8800 1005 8805 1045
rect 8845 1005 8850 1045
rect 8800 845 8850 1005
rect 8800 805 8805 845
rect 8845 805 8850 845
rect 8800 -855 8850 805
rect 8800 -895 8805 -855
rect 8845 -895 8850 -855
rect 8800 -900 8850 -895
rect 9100 1045 9150 1050
rect 9100 1005 9105 1045
rect 9145 1005 9150 1045
rect 9100 845 9150 1005
rect 9100 805 9105 845
rect 9145 805 9150 845
rect 9100 -855 9150 805
rect 9100 -895 9105 -855
rect 9145 -895 9150 -855
rect 9100 -900 9150 -895
rect 9400 1045 9450 1050
rect 9400 1005 9405 1045
rect 9445 1005 9450 1045
rect 9400 845 9450 1005
rect 9400 805 9405 845
rect 9445 805 9450 845
rect 9400 -855 9450 805
rect 9400 -895 9405 -855
rect 9445 -895 9450 -855
rect 9400 -900 9450 -895
rect 9550 845 9600 3305
rect 12100 2145 12150 2150
rect 12100 2105 12105 2145
rect 12145 2105 12150 2145
rect 9550 805 9555 845
rect 9595 805 9600 845
rect 9550 -855 9600 805
rect 9550 -895 9555 -855
rect 9595 -895 9600 -855
rect 9550 -900 9600 -895
rect 9700 1045 9750 1050
rect 9700 1005 9705 1045
rect 9745 1005 9750 1045
rect 9700 845 9750 1005
rect 9700 805 9705 845
rect 9745 805 9750 845
rect 9700 -855 9750 805
rect 9700 -895 9705 -855
rect 9745 -895 9750 -855
rect 9700 -900 9750 -895
rect 10000 1045 10050 1050
rect 10000 1005 10005 1045
rect 10045 1005 10050 1045
rect 10000 845 10050 1005
rect 10000 805 10005 845
rect 10045 805 10050 845
rect 10000 -855 10050 805
rect 10000 -895 10005 -855
rect 10045 -895 10050 -855
rect 10000 -900 10050 -895
rect 10300 1045 10350 1050
rect 10300 1005 10305 1045
rect 10345 1005 10350 1045
rect 10300 845 10350 1005
rect 10300 805 10305 845
rect 10345 805 10350 845
rect 10300 -855 10350 805
rect 10300 -895 10305 -855
rect 10345 -895 10350 -855
rect 10300 -900 10350 -895
rect 10600 1045 10650 1050
rect 10600 1005 10605 1045
rect 10645 1005 10650 1045
rect 10600 845 10650 1005
rect 10600 805 10605 845
rect 10645 805 10650 845
rect 10600 -855 10650 805
rect 10600 -895 10605 -855
rect 10645 -895 10650 -855
rect 10600 -900 10650 -895
rect 10900 1045 10950 1050
rect 10900 1005 10905 1045
rect 10945 1005 10950 1045
rect 10900 845 10950 1005
rect 10900 805 10905 845
rect 10945 805 10950 845
rect 10900 -855 10950 805
rect 10900 -895 10905 -855
rect 10945 -895 10950 -855
rect 10900 -900 10950 -895
rect 11200 1045 11250 1050
rect 11200 1005 11205 1045
rect 11245 1005 11250 1045
rect 11200 845 11250 1005
rect 11200 805 11205 845
rect 11245 805 11250 845
rect 11200 -855 11250 805
rect 11200 -895 11205 -855
rect 11245 -895 11250 -855
rect 11200 -900 11250 -895
rect 11500 1045 11550 1050
rect 11500 1005 11505 1045
rect 11545 1005 11550 1045
rect 11500 845 11550 1005
rect 11500 805 11505 845
rect 11545 805 11550 845
rect 11500 -855 11550 805
rect 11500 -895 11505 -855
rect 11545 -895 11550 -855
rect 11500 -900 11550 -895
rect 11800 1045 11850 1050
rect 11800 1005 11805 1045
rect 11845 1005 11850 1045
rect 11800 845 11850 1005
rect 11800 805 11805 845
rect 11845 805 11850 845
rect 11800 -855 11850 805
rect 11800 -895 11805 -855
rect 11845 -895 11850 -855
rect 11800 -900 11850 -895
rect 12100 845 12150 2105
rect 12100 805 12105 845
rect 12145 805 12150 845
rect 12100 -855 12150 805
rect 12100 -895 12105 -855
rect 12145 -895 12150 -855
rect 12100 -900 12150 -895
rect 12400 2145 12450 2150
rect 12400 2105 12405 2145
rect 12445 2105 12450 2145
rect 12400 845 12450 2105
rect 12400 805 12405 845
rect 12445 805 12450 845
rect 12400 -855 12450 805
rect 12400 -895 12405 -855
rect 12445 -895 12450 -855
rect 12400 -900 12450 -895
rect 12550 845 12600 3605
rect 12700 3845 12750 4905
rect 12700 3805 12705 3845
rect 12745 3805 12750 3845
rect 12700 3645 12750 3805
rect 12700 3605 12705 3645
rect 12745 3605 12750 3645
rect 12700 3600 12750 3605
rect 13000 4945 13050 4950
rect 13000 4905 13005 4945
rect 13045 4905 13050 4945
rect 13000 3845 13050 4905
rect 13000 3805 13005 3845
rect 13045 3805 13050 3845
rect 13000 3645 13050 3805
rect 13000 3605 13005 3645
rect 13045 3605 13050 3645
rect 13000 3600 13050 3605
rect 13300 4945 13350 4950
rect 13300 4905 13305 4945
rect 13345 4905 13350 4945
rect 13300 3845 13350 4905
rect 13300 3805 13305 3845
rect 13345 3805 13350 3845
rect 13300 3645 13350 3805
rect 13300 3605 13305 3645
rect 13345 3605 13350 3645
rect 13300 3600 13350 3605
rect 13600 4945 13650 4950
rect 13600 4905 13605 4945
rect 13645 4905 13650 4945
rect 13600 3845 13650 4905
rect 13750 4945 13800 4950
rect 13750 4905 13755 4945
rect 13795 4905 13800 4945
rect 13750 4900 13800 4905
rect 13900 4945 13950 4950
rect 13900 4905 13905 4945
rect 13945 4905 13950 4945
rect 13600 3805 13605 3845
rect 13645 3805 13650 3845
rect 13600 3645 13650 3805
rect 13600 3605 13605 3645
rect 13645 3605 13650 3645
rect 13600 3600 13650 3605
rect 13750 4745 13800 4750
rect 13750 4705 13755 4745
rect 13795 4705 13800 4745
rect 13750 3645 13800 4705
rect 13750 3605 13755 3645
rect 13795 3605 13800 3645
rect 13300 2745 13350 2750
rect 13300 2705 13305 2745
rect 13345 2705 13350 2745
rect 12550 805 12555 845
rect 12595 805 12600 845
rect 12550 -855 12600 805
rect 12550 -895 12555 -855
rect 12595 -895 12600 -855
rect 12550 -900 12600 -895
rect 12700 2145 12750 2150
rect 12700 2105 12705 2145
rect 12745 2105 12750 2145
rect 12700 845 12750 2105
rect 12700 805 12705 845
rect 12745 805 12750 845
rect 12700 -855 12750 805
rect 12700 -895 12705 -855
rect 12745 -895 12750 -855
rect 12700 -900 12750 -895
rect 13000 2145 13050 2150
rect 13000 2105 13005 2145
rect 13045 2105 13050 2145
rect 13000 845 13050 2105
rect 13000 805 13005 845
rect 13045 805 13050 845
rect 13000 -855 13050 805
rect 13000 -895 13005 -855
rect 13045 -895 13050 -855
rect 13000 -900 13050 -895
rect 13300 845 13350 2705
rect 13300 805 13305 845
rect 13345 805 13350 845
rect 13300 -855 13350 805
rect 13300 -895 13305 -855
rect 13345 -895 13350 -855
rect 13300 -900 13350 -895
rect 13600 2745 13650 2750
rect 13600 2705 13605 2745
rect 13645 2705 13650 2745
rect 13600 845 13650 2705
rect 13600 805 13605 845
rect 13645 805 13650 845
rect 13600 -855 13650 805
rect 13600 -895 13605 -855
rect 13645 -895 13650 -855
rect 13600 -900 13650 -895
rect 13750 845 13800 3605
rect 13900 3845 13950 4905
rect 13900 3805 13905 3845
rect 13945 3805 13950 3845
rect 13900 3645 13950 3805
rect 13900 3605 13905 3645
rect 13945 3605 13950 3645
rect 13900 3600 13950 3605
rect 14200 4945 14250 4950
rect 14200 4905 14205 4945
rect 14245 4905 14250 4945
rect 14200 3845 14250 4905
rect 14200 3805 14205 3845
rect 14245 3805 14250 3845
rect 14200 3645 14250 3805
rect 14200 3605 14205 3645
rect 14245 3605 14250 3645
rect 14200 3600 14250 3605
rect 14500 4945 14550 4950
rect 14500 4905 14505 4945
rect 14545 4905 14550 4945
rect 14500 3845 14550 4905
rect 14500 3805 14505 3845
rect 14545 3805 14550 3845
rect 14500 3645 14550 3805
rect 14500 3605 14505 3645
rect 14545 3605 14550 3645
rect 14500 3600 14550 3605
rect 14800 4945 14850 4950
rect 14800 4905 14805 4945
rect 14845 4905 14850 4945
rect 14800 3845 14850 4905
rect 14800 3805 14805 3845
rect 14845 3805 14850 3845
rect 14800 3645 14850 3805
rect 14800 3605 14805 3645
rect 14845 3605 14850 3645
rect 14800 3600 14850 3605
rect 14950 4945 15000 4950
rect 14950 4905 14955 4945
rect 14995 4905 15000 4945
rect 14950 4745 15000 4905
rect 14950 4705 14955 4745
rect 14995 4705 15000 4745
rect 14950 3645 15000 4705
rect 15100 4945 15150 4950
rect 15100 4905 15105 4945
rect 15145 4905 15150 4945
rect 15100 4050 15150 4905
rect 15400 4945 15450 4950
rect 15400 4905 15405 4945
rect 15445 4905 15450 4945
rect 15400 4050 15450 4905
rect 15700 4945 15750 4950
rect 15700 4905 15705 4945
rect 15745 4905 15750 4945
rect 14950 3605 14955 3645
rect 14995 3605 15000 3645
rect 14950 3600 15000 3605
rect 15100 3645 15150 4000
rect 15100 3605 15105 3645
rect 15145 3605 15150 3645
rect 15100 3600 15150 3605
rect 15400 3645 15450 4000
rect 15400 3605 15405 3645
rect 15445 3605 15450 3645
rect 15400 3600 15450 3605
rect 15700 3645 15750 4905
rect 15700 3605 15705 3645
rect 15745 3605 15750 3645
rect 15700 3600 15750 3605
rect 16000 4945 16050 4950
rect 16000 4905 16005 4945
rect 16045 4905 16050 4945
rect 16000 3645 16050 4905
rect 16000 3605 16005 3645
rect 16045 3605 16050 3645
rect 16000 3600 16050 3605
rect 16300 4945 16350 5500
rect 16300 4905 16305 4945
rect 16345 4905 16350 4945
rect 16300 3645 16350 4905
rect 16300 3605 16305 3645
rect 16345 3605 16350 3645
rect 13750 805 13755 845
rect 13795 805 13800 845
rect 13750 -855 13800 805
rect 13750 -895 13755 -855
rect 13795 -895 13800 -855
rect 13750 -900 13800 -895
rect 13900 2745 13950 2750
rect 13900 2705 13905 2745
rect 13945 2705 13950 2745
rect 13900 845 13950 2705
rect 13900 805 13905 845
rect 13945 805 13950 845
rect 13900 -855 13950 805
rect 13900 -895 13905 -855
rect 13945 -895 13950 -855
rect 13900 -900 13950 -895
rect 14200 2745 14250 2750
rect 14200 2705 14205 2745
rect 14245 2705 14250 2745
rect 14200 845 14250 2705
rect 16300 2145 16350 3605
rect 16300 2105 16305 2145
rect 16345 2105 16350 2145
rect 16300 2100 16350 2105
rect 16600 4945 16650 5500
rect 16600 4905 16605 4945
rect 16645 4905 16650 4945
rect 16600 3645 16650 4905
rect 16600 3605 16605 3645
rect 16645 3605 16650 3645
rect 16600 2145 16650 3605
rect 16600 2105 16605 2145
rect 16645 2105 16650 2145
rect 16600 2100 16650 2105
rect 16750 4945 16800 4950
rect 16750 4905 16755 4945
rect 16795 4905 16800 4945
rect 16750 3645 16800 4905
rect 16750 3605 16755 3645
rect 16795 3605 16800 3645
rect 14200 805 14205 845
rect 14245 805 14250 845
rect 14200 -855 14250 805
rect 14200 -895 14205 -855
rect 14245 -895 14250 -855
rect 14200 -900 14250 -895
rect 14500 1045 14550 1050
rect 14500 1005 14505 1045
rect 14545 1005 14550 1045
rect 14500 845 14550 1005
rect 14500 805 14505 845
rect 14545 805 14550 845
rect 14500 -855 14550 805
rect 14500 -895 14505 -855
rect 14545 -895 14550 -855
rect 14500 -900 14550 -895
rect 14800 1045 14850 1050
rect 14800 1005 14805 1045
rect 14845 1005 14850 1045
rect 14800 845 14850 1005
rect 14800 805 14805 845
rect 14845 805 14850 845
rect 14800 -855 14850 805
rect 14800 -895 14805 -855
rect 14845 -895 14850 -855
rect 14800 -900 14850 -895
rect 15100 1045 15150 1050
rect 15100 1005 15105 1045
rect 15145 1005 15150 1045
rect 15100 845 15150 1005
rect 15100 805 15105 845
rect 15145 805 15150 845
rect 15100 -855 15150 805
rect 15100 -895 15105 -855
rect 15145 -895 15150 -855
rect 15100 -900 15150 -895
rect 15400 1045 15450 1050
rect 15400 1005 15405 1045
rect 15445 1005 15450 1045
rect 15400 845 15450 1005
rect 15400 805 15405 845
rect 15445 805 15450 845
rect 15400 -855 15450 805
rect 15400 -895 15405 -855
rect 15445 -895 15450 -855
rect 15400 -900 15450 -895
rect 15700 845 15750 850
rect 15700 805 15705 845
rect 15745 805 15750 845
rect 15700 645 15750 805
rect 15700 605 15705 645
rect 15745 605 15750 645
rect 15700 -855 15750 605
rect 15700 -895 15705 -855
rect 15745 -895 15750 -855
rect 15700 -900 15750 -895
rect 16000 845 16050 850
rect 16000 805 16005 845
rect 16045 805 16050 845
rect 16000 645 16050 805
rect 16000 605 16005 645
rect 16045 605 16050 645
rect 16000 -855 16050 605
rect 16000 -895 16005 -855
rect 16045 -895 16050 -855
rect 16000 -900 16050 -895
rect 16300 845 16350 850
rect 16300 805 16305 845
rect 16345 805 16350 845
rect 16300 645 16350 805
rect 16300 605 16305 645
rect 16345 605 16350 645
rect 16300 -855 16350 605
rect 16300 -895 16305 -855
rect 16345 -895 16350 -855
rect 16300 -900 16350 -895
rect 16600 845 16650 850
rect 16600 805 16605 845
rect 16645 805 16650 845
rect 16600 645 16650 805
rect 16600 605 16605 645
rect 16645 605 16650 645
rect 16600 -855 16650 605
rect 16600 -895 16605 -855
rect 16645 -895 16650 -855
rect 16600 -900 16650 -895
rect 16750 845 16800 3605
rect 16900 4945 16950 5500
rect 16900 4905 16905 4945
rect 16945 4905 16950 4945
rect 16900 3645 16950 4905
rect 16900 3605 16905 3645
rect 16945 3605 16950 3645
rect 16900 2145 16950 3605
rect 16900 2105 16905 2145
rect 16945 2105 16950 2145
rect 16900 2100 16950 2105
rect 17200 4945 17250 5500
rect 17200 4905 17205 4945
rect 17245 4905 17250 4945
rect 17200 3645 17250 4905
rect 17200 3605 17205 3645
rect 17245 3605 17250 3645
rect 17200 2145 17250 3605
rect 17500 4945 17550 4950
rect 17500 4905 17505 4945
rect 17545 4905 17550 4945
rect 17500 3645 17550 4905
rect 17500 3605 17505 3645
rect 17545 3605 17550 3645
rect 17500 3600 17550 3605
rect 17800 4945 17850 4950
rect 17800 4905 17805 4945
rect 17845 4905 17850 4945
rect 17800 3645 17850 4905
rect 17800 3605 17805 3645
rect 17845 3605 17850 3645
rect 17800 3600 17850 3605
rect 18100 4945 18150 4950
rect 18100 4905 18105 4945
rect 18145 4905 18150 4945
rect 18100 3645 18150 4905
rect 18100 3605 18105 3645
rect 18145 3605 18150 3645
rect 18100 3445 18150 3605
rect 18100 3405 18105 3445
rect 18145 3405 18150 3445
rect 18100 3400 18150 3405
rect 18400 4945 18450 4950
rect 18400 4905 18405 4945
rect 18445 4905 18450 4945
rect 18400 3645 18450 4905
rect 18400 3605 18405 3645
rect 18445 3605 18450 3645
rect 18400 3445 18450 3605
rect 18400 3405 18405 3445
rect 18445 3405 18450 3445
rect 18400 3400 18450 3405
rect 18700 4945 18750 5500
rect 18700 4905 18705 4945
rect 18745 4905 18750 4945
rect 18700 3645 18750 4905
rect 18700 3605 18705 3645
rect 18745 3605 18750 3645
rect 18700 2745 18750 3605
rect 18700 2705 18705 2745
rect 18745 2705 18750 2745
rect 18700 2700 18750 2705
rect 19000 4945 19050 5500
rect 19000 4905 19005 4945
rect 19045 4905 19050 4945
rect 19000 3645 19050 4905
rect 19000 3605 19005 3645
rect 19045 3605 19050 3645
rect 19000 2745 19050 3605
rect 19000 2705 19005 2745
rect 19045 2705 19050 2745
rect 19000 2700 19050 2705
rect 19150 4945 19200 4950
rect 19150 4905 19155 4945
rect 19195 4905 19200 4945
rect 19150 3645 19200 4905
rect 19150 3605 19155 3645
rect 19195 3605 19200 3645
rect 17200 2105 17205 2145
rect 17245 2105 17250 2145
rect 17200 2100 17250 2105
rect 16750 805 16755 845
rect 16795 805 16800 845
rect 16750 -455 16800 805
rect 16750 -495 16755 -455
rect 16795 -495 16800 -455
rect 16750 -855 16800 -495
rect 16750 -895 16755 -855
rect 16795 -895 16800 -855
rect 16750 -900 16800 -895
rect 16900 845 16950 850
rect 16900 805 16905 845
rect 16945 805 16950 845
rect 16900 645 16950 805
rect 16900 605 16905 645
rect 16945 605 16950 645
rect 16900 -855 16950 605
rect 16900 -895 16905 -855
rect 16945 -895 16950 -855
rect 16900 -900 16950 -895
rect 17200 845 17250 850
rect 17200 805 17205 845
rect 17245 805 17250 845
rect 17200 645 17250 805
rect 17200 605 17205 645
rect 17245 605 17250 645
rect 17200 -855 17250 605
rect 17200 -895 17205 -855
rect 17245 -895 17250 -855
rect 17200 -900 17250 -895
rect 17500 845 17550 850
rect 17500 805 17505 845
rect 17545 805 17550 845
rect 17500 645 17550 805
rect 17500 605 17505 645
rect 17545 605 17550 645
rect 17500 -855 17550 605
rect 17500 -895 17505 -855
rect 17545 -895 17550 -855
rect 17500 -900 17550 -895
rect 17800 845 17850 850
rect 17800 805 17805 845
rect 17845 805 17850 845
rect 17800 645 17850 805
rect 17800 605 17805 645
rect 17845 605 17850 645
rect 17800 -855 17850 605
rect 17800 -895 17805 -855
rect 17845 -895 17850 -855
rect 17800 -900 17850 -895
rect 18100 845 18150 850
rect 18100 805 18105 845
rect 18145 805 18150 845
rect 18100 645 18150 805
rect 18100 605 18105 645
rect 18145 605 18150 645
rect 18100 -855 18150 605
rect 18100 -895 18105 -855
rect 18145 -895 18150 -855
rect 18100 -900 18150 -895
rect 18400 845 18450 850
rect 18400 805 18405 845
rect 18445 805 18450 845
rect 18400 645 18450 805
rect 18400 605 18405 645
rect 18445 605 18450 645
rect 18400 -855 18450 605
rect 18400 -895 18405 -855
rect 18445 -895 18450 -855
rect 18400 -900 18450 -895
rect 18700 845 18750 850
rect 18700 805 18705 845
rect 18745 805 18750 845
rect 18700 645 18750 805
rect 18700 605 18705 645
rect 18745 605 18750 645
rect 18700 -855 18750 605
rect 18700 -895 18705 -855
rect 18745 -895 18750 -855
rect 18700 -900 18750 -895
rect 19000 845 19050 850
rect 19000 805 19005 845
rect 19045 805 19050 845
rect 19000 645 19050 805
rect 19000 605 19005 645
rect 19045 605 19050 645
rect 19000 -855 19050 605
rect 19000 -895 19005 -855
rect 19045 -895 19050 -855
rect 19000 -900 19050 -895
rect 19150 845 19200 3605
rect 19300 4945 19350 5500
rect 19300 4905 19305 4945
rect 19345 4905 19350 4945
rect 19300 3645 19350 4905
rect 19300 3605 19305 3645
rect 19345 3605 19350 3645
rect 19300 2745 19350 3605
rect 19300 2705 19305 2745
rect 19345 2705 19350 2745
rect 19300 2700 19350 2705
rect 19600 4945 19650 5500
rect 19600 4905 19605 4945
rect 19645 4905 19650 4945
rect 19600 3645 19650 4905
rect 19600 3605 19605 3645
rect 19645 3605 19650 3645
rect 19600 2700 19650 3605
rect 19900 4945 19950 4950
rect 19900 4905 19905 4945
rect 19945 4905 19950 4945
rect 19900 3645 19950 4905
rect 19900 3605 19905 3645
rect 19945 3605 19950 3645
rect 19900 3445 19950 3605
rect 19900 3405 19905 3445
rect 19945 3405 19950 3445
rect 19900 3400 19950 3405
rect 20200 4945 20250 4950
rect 20200 4905 20205 4945
rect 20245 4905 20250 4945
rect 20200 3645 20250 4905
rect 20200 3605 20205 3645
rect 20245 3605 20250 3645
rect 20200 3445 20250 3605
rect 20500 4945 20550 4950
rect 20500 4905 20505 4945
rect 20545 4905 20550 4945
rect 20500 3845 20550 4905
rect 20500 3805 20505 3845
rect 20545 3805 20550 3845
rect 20500 3645 20550 3805
rect 20500 3605 20505 3645
rect 20545 3605 20550 3645
rect 20500 3600 20550 3605
rect 20800 4945 20850 4950
rect 20800 4905 20805 4945
rect 20845 4905 20850 4945
rect 20800 3845 20850 4905
rect 20800 3805 20805 3845
rect 20845 3805 20850 3845
rect 20800 3645 20850 3805
rect 20800 3605 20805 3645
rect 20845 3605 20850 3645
rect 20800 3600 20850 3605
rect 20950 4945 21000 4950
rect 20950 4905 20955 4945
rect 20995 4905 21000 4945
rect 20950 4545 21000 4905
rect 20950 4505 20955 4545
rect 20995 4505 21000 4545
rect 20950 3645 21000 4505
rect 20950 3605 20955 3645
rect 20995 3605 21000 3645
rect 20950 3600 21000 3605
rect 21100 4945 21150 4950
rect 21100 4905 21105 4945
rect 21145 4905 21150 4945
rect 21100 3845 21150 4905
rect 21100 3805 21105 3845
rect 21145 3805 21150 3845
rect 21100 3645 21150 3805
rect 21100 3605 21105 3645
rect 21145 3605 21150 3645
rect 21100 3600 21150 3605
rect 21400 3845 21450 4950
rect 21400 3805 21405 3845
rect 21445 3805 21450 3845
rect 21400 3600 21450 3805
rect 21700 4945 21750 4950
rect 21700 4905 21705 4945
rect 21745 4905 21750 4945
rect 21700 3845 21750 4905
rect 21700 3805 21705 3845
rect 21745 3805 21750 3845
rect 21700 3645 21750 3805
rect 21700 3605 21705 3645
rect 21745 3605 21750 3645
rect 21700 3600 21750 3605
rect 21850 4945 21900 4950
rect 21850 4905 21855 4945
rect 21895 4905 21900 4945
rect 21850 4545 21900 4905
rect 21850 4505 21855 4545
rect 21895 4505 21900 4545
rect 21850 3645 21900 4505
rect 21850 3605 21855 3645
rect 21895 3605 21900 3645
rect 21850 3600 21900 3605
rect 22000 4945 22050 4950
rect 22000 4905 22005 4945
rect 22045 4905 22050 4945
rect 22000 3845 22050 4905
rect 22000 3805 22005 3845
rect 22045 3805 22050 3845
rect 22000 3645 22050 3805
rect 22000 3605 22005 3645
rect 22045 3605 22050 3645
rect 22000 3600 22050 3605
rect 22300 4945 22350 4950
rect 22300 4905 22305 4945
rect 22345 4905 22350 4945
rect 22300 3845 22350 4905
rect 22600 4945 22650 4950
rect 22600 4905 22605 4945
rect 22645 4905 22650 4945
rect 22300 3805 22305 3845
rect 22345 3805 22350 3845
rect 22300 3645 22350 3805
rect 22300 3605 22305 3645
rect 22345 3605 22350 3645
rect 22300 3600 22350 3605
rect 22450 3845 22500 3850
rect 22450 3805 22455 3845
rect 22495 3805 22500 3845
rect 20200 3405 20205 3445
rect 20245 3405 20250 3445
rect 20200 3400 20250 3405
rect 21700 1145 21750 1150
rect 21700 1105 21705 1145
rect 21745 1105 21750 1145
rect 20500 1045 20550 1050
rect 20500 1005 20505 1045
rect 20545 1005 20550 1045
rect 19150 805 19155 845
rect 19195 805 19200 845
rect 19150 -855 19200 805
rect 19150 -895 19155 -855
rect 19195 -895 19200 -855
rect 19150 -900 19200 -895
rect 19300 845 19350 850
rect 19300 805 19305 845
rect 19345 805 19350 845
rect 19300 645 19350 805
rect 19300 605 19305 645
rect 19345 605 19350 645
rect 19300 -855 19350 605
rect 19300 -895 19305 -855
rect 19345 -895 19350 -855
rect 19300 -900 19350 -895
rect 19600 845 19650 850
rect 19600 805 19605 845
rect 19645 805 19650 845
rect 19600 645 19650 805
rect 19600 605 19605 645
rect 19645 605 19650 645
rect 19600 -855 19650 605
rect 19600 -895 19605 -855
rect 19645 -895 19650 -855
rect 19600 -900 19650 -895
rect 19900 845 19950 850
rect 19900 805 19905 845
rect 19945 805 19950 845
rect 19900 645 19950 805
rect 19900 605 19905 645
rect 19945 605 19950 645
rect 19900 -855 19950 605
rect 19900 -895 19905 -855
rect 19945 -895 19950 -855
rect 19900 -900 19950 -895
rect 20200 845 20250 850
rect 20200 805 20205 845
rect 20245 805 20250 845
rect 20200 645 20250 805
rect 20200 605 20205 645
rect 20245 605 20250 645
rect 20200 -855 20250 605
rect 20200 -895 20205 -855
rect 20245 -895 20250 -855
rect 20200 -900 20250 -895
rect 20500 845 20550 1005
rect 20500 805 20505 845
rect 20545 805 20550 845
rect 20500 -855 20550 805
rect 20500 -895 20505 -855
rect 20545 -895 20550 -855
rect 20500 -900 20550 -895
rect 20800 1045 20850 1050
rect 20800 1005 20805 1045
rect 20845 1005 20850 1045
rect 20800 845 20850 1005
rect 20800 805 20805 845
rect 20845 805 20850 845
rect 20800 -855 20850 805
rect 20800 -895 20805 -855
rect 20845 -895 20850 -855
rect 20800 -900 20850 -895
rect 21100 1045 21150 1050
rect 21100 1005 21105 1045
rect 21145 1005 21150 1045
rect 21100 845 21150 1005
rect 21100 805 21105 845
rect 21145 805 21150 845
rect 21100 -855 21150 805
rect 21100 -895 21105 -855
rect 21145 -895 21150 -855
rect 21100 -900 21150 -895
rect 21400 1045 21450 1050
rect 21400 1005 21405 1045
rect 21445 1005 21450 1045
rect 21400 845 21450 1005
rect 21400 805 21405 845
rect 21445 805 21450 845
rect 21400 -855 21450 805
rect 21400 -895 21405 -855
rect 21445 -895 21450 -855
rect 21400 -900 21450 -895
rect 21700 845 21750 1105
rect 21700 805 21705 845
rect 21745 805 21750 845
rect 21700 -855 21750 805
rect 21700 -895 21705 -855
rect 21745 -895 21750 -855
rect 21700 -900 21750 -895
rect 22000 1145 22050 1150
rect 22000 1105 22005 1145
rect 22045 1105 22050 1145
rect 22000 845 22050 1105
rect 22000 805 22005 845
rect 22045 805 22050 845
rect 22000 -855 22050 805
rect 22000 -895 22005 -855
rect 22045 -895 22050 -855
rect 22000 -900 22050 -895
rect 22300 1145 22350 1150
rect 22300 1105 22305 1145
rect 22345 1105 22350 1145
rect 22300 845 22350 1105
rect 22300 805 22305 845
rect 22345 805 22350 845
rect 22300 -855 22350 805
rect 22300 -895 22305 -855
rect 22345 -895 22350 -855
rect 22300 -900 22350 -895
rect 22450 845 22500 3805
rect 22600 3845 22650 4905
rect 22600 3805 22605 3845
rect 22645 3805 22650 3845
rect 22600 3645 22650 3805
rect 22600 3605 22605 3645
rect 22645 3605 22650 3645
rect 22600 3600 22650 3605
rect 22900 4945 22950 4950
rect 22900 4905 22905 4945
rect 22945 4905 22950 4945
rect 22900 3845 22950 4905
rect 22900 3805 22905 3845
rect 22945 3805 22950 3845
rect 22900 3645 22950 3805
rect 22900 3605 22905 3645
rect 22945 3605 22950 3645
rect 22900 3600 22950 3605
rect 23050 4945 23100 4950
rect 23050 4905 23055 4945
rect 23095 4905 23100 4945
rect 23050 4545 23100 4905
rect 23050 4505 23055 4545
rect 23095 4505 23100 4545
rect 23050 3645 23100 4505
rect 23050 3605 23055 3645
rect 23095 3605 23100 3645
rect 23050 3600 23100 3605
rect 23200 4945 23250 4950
rect 23200 4905 23205 4945
rect 23245 4905 23250 4945
rect 23200 3845 23250 4905
rect 23350 4945 23400 4950
rect 23350 4905 23355 4945
rect 23395 4905 23400 4945
rect 23350 4900 23400 4905
rect 23200 3805 23205 3845
rect 23245 3805 23250 3845
rect 23200 3645 23250 3805
rect 23500 3845 23550 4950
rect 23650 4945 23700 4950
rect 23650 4905 23655 4945
rect 23695 4905 23700 4945
rect 23650 4900 23700 4905
rect 23800 4945 23850 4950
rect 23800 4905 23805 4945
rect 23845 4905 23850 4945
rect 23500 3805 23505 3845
rect 23545 3805 23550 3845
rect 23200 3605 23205 3645
rect 23245 3605 23250 3645
rect 23200 3600 23250 3605
rect 23350 3645 23400 3650
rect 23350 3605 23355 3645
rect 23395 3605 23400 3645
rect 23350 3600 23400 3605
rect 23500 3600 23550 3805
rect 23800 3845 23850 4905
rect 23800 3805 23805 3845
rect 23845 3805 23850 3845
rect 23650 3645 23700 3650
rect 23650 3605 23655 3645
rect 23695 3605 23700 3645
rect 23650 3600 23700 3605
rect 23800 3645 23850 3805
rect 23800 3605 23805 3645
rect 23845 3605 23850 3645
rect 23800 3600 23850 3605
rect 23950 4945 24000 4950
rect 23950 4905 23955 4945
rect 23995 4905 24000 4945
rect 23950 4545 24000 4905
rect 23950 4505 23955 4545
rect 23995 4505 24000 4545
rect 23950 3645 24000 4505
rect 23950 3605 23955 3645
rect 23995 3605 24000 3645
rect 23950 3600 24000 3605
rect 24100 4945 24150 4950
rect 24100 4905 24105 4945
rect 24145 4905 24150 4945
rect 24100 3845 24150 4905
rect 24100 3805 24105 3845
rect 24145 3805 24150 3845
rect 24100 3645 24150 3805
rect 24100 3605 24105 3645
rect 24145 3605 24150 3645
rect 24100 3600 24150 3605
rect 24400 4945 24450 4950
rect 24400 4905 24405 4945
rect 24445 4905 24450 4945
rect 24400 3845 24450 4905
rect 24400 3805 24405 3845
rect 24445 3805 24450 3845
rect 24400 3645 24450 3805
rect 24400 3605 24405 3645
rect 24445 3605 24450 3645
rect 24400 3600 24450 3605
rect 24700 4945 24750 4950
rect 24700 4905 24705 4945
rect 24745 4905 24750 4945
rect 24700 3645 24750 4905
rect 24700 3605 24705 3645
rect 24745 3605 24750 3645
rect 24700 3445 24750 3605
rect 24700 3405 24705 3445
rect 24745 3405 24750 3445
rect 24700 3400 24750 3405
rect 25000 4945 25050 4950
rect 25000 4905 25005 4945
rect 25045 4905 25050 4945
rect 25000 3645 25050 4905
rect 25000 3605 25005 3645
rect 25045 3605 25050 3645
rect 25000 3445 25050 3605
rect 25000 3405 25005 3445
rect 25045 3405 25050 3445
rect 25000 3400 25050 3405
rect 25450 4945 25500 4950
rect 25450 4905 25455 4945
rect 25495 4905 25500 4945
rect 25450 3645 25500 4905
rect 25450 3605 25455 3645
rect 25495 3605 25500 3645
rect 25450 3345 25500 3605
rect 25450 3305 25455 3345
rect 25495 3305 25500 3345
rect 25450 3300 25500 3305
rect 25600 4945 25650 4950
rect 25600 4905 25605 4945
rect 25645 4905 25650 4945
rect 25600 3645 25650 4905
rect 25600 3605 25605 3645
rect 25645 3605 25650 3645
rect 22450 805 22455 845
rect 22495 805 22500 845
rect 22450 -855 22500 805
rect 22450 -895 22455 -855
rect 22495 -895 22500 -855
rect 22450 -900 22500 -895
rect 22600 1145 22650 1150
rect 22600 1105 22605 1145
rect 22645 1105 22650 1145
rect 22600 845 22650 1105
rect 22600 805 22605 845
rect 22645 805 22650 845
rect 22600 -855 22650 805
rect 22600 -895 22605 -855
rect 22645 -895 22650 -855
rect 22600 -900 22650 -895
rect 22900 1145 22950 1150
rect 22900 1105 22905 1145
rect 22945 1105 22950 1145
rect 22900 845 22950 1105
rect 22900 805 22905 845
rect 22945 805 22950 845
rect 22900 -855 22950 805
rect 22900 -895 22905 -855
rect 22945 -895 22950 -855
rect 22900 -900 22950 -895
rect 23200 1145 23250 1150
rect 23200 1105 23205 1145
rect 23245 1105 23250 1145
rect 23200 845 23250 1105
rect 23200 805 23205 845
rect 23245 805 23250 845
rect 23200 -855 23250 805
rect 23200 -895 23205 -855
rect 23245 -895 23250 -855
rect 23200 -900 23250 -895
rect 23500 1045 23550 1050
rect 23500 1005 23505 1045
rect 23545 1005 23550 1045
rect 23500 845 23550 1005
rect 23500 805 23505 845
rect 23545 805 23550 845
rect 23500 -855 23550 805
rect 23500 -895 23505 -855
rect 23545 -895 23550 -855
rect 23500 -900 23550 -895
rect 23800 1045 23850 1050
rect 23800 1005 23805 1045
rect 23845 1005 23850 1045
rect 23800 845 23850 1005
rect 23800 805 23805 845
rect 23845 805 23850 845
rect 23800 -855 23850 805
rect 23800 -895 23805 -855
rect 23845 -895 23850 -855
rect 23800 -900 23850 -895
rect 24100 1045 24150 1050
rect 24100 1005 24105 1045
rect 24145 1005 24150 1045
rect 24100 845 24150 1005
rect 24100 805 24105 845
rect 24145 805 24150 845
rect 24100 -855 24150 805
rect 24100 -895 24105 -855
rect 24145 -895 24150 -855
rect 24100 -900 24150 -895
rect 24400 1045 24450 1050
rect 24400 1005 24405 1045
rect 24445 1005 24450 1045
rect 24400 845 24450 1005
rect 24400 805 24405 845
rect 24445 805 24450 845
rect 24400 -855 24450 805
rect 24400 -895 24405 -855
rect 24445 -895 24450 -855
rect 24400 -900 24450 -895
rect 24700 845 24750 850
rect 24700 805 24705 845
rect 24745 805 24750 845
rect 24700 645 24750 805
rect 24700 605 24705 645
rect 24745 605 24750 645
rect 24700 -855 24750 605
rect 24700 -895 24705 -855
rect 24745 -895 24750 -855
rect 24700 -900 24750 -895
rect 25000 845 25050 850
rect 25000 805 25005 845
rect 25045 805 25050 845
rect 25000 645 25050 805
rect 25000 605 25005 645
rect 25045 605 25050 645
rect 25000 -855 25050 605
rect 25000 -895 25005 -855
rect 25045 -895 25050 -855
rect 25000 -900 25050 -895
rect 25300 845 25350 850
rect 25300 805 25305 845
rect 25345 805 25350 845
rect 25300 645 25350 805
rect 25300 605 25305 645
rect 25345 605 25350 645
rect 25300 -855 25350 605
rect 25300 -895 25305 -855
rect 25345 -895 25350 -855
rect 25300 -900 25350 -895
rect 25600 845 25650 3605
rect 25750 4945 25800 4950
rect 25750 4905 25755 4945
rect 25795 4905 25800 4945
rect 25750 3645 25800 4905
rect 25750 3605 25755 3645
rect 25795 3605 25800 3645
rect 25750 3345 25800 3605
rect 26200 4945 26250 4950
rect 26200 4905 26205 4945
rect 26245 4905 26250 4945
rect 26200 3645 26250 4905
rect 26200 3605 26205 3645
rect 26245 3605 26250 3645
rect 26200 3445 26250 3605
rect 26200 3405 26205 3445
rect 26245 3405 26250 3445
rect 26200 3400 26250 3405
rect 26500 4945 26550 4950
rect 26500 4905 26505 4945
rect 26545 4905 26550 4945
rect 26500 3645 26550 4905
rect 26500 3605 26505 3645
rect 26545 3605 26550 3645
rect 26500 3445 26550 3605
rect 26500 3405 26505 3445
rect 26545 3405 26550 3445
rect 26500 3400 26550 3405
rect 26800 4945 26850 4950
rect 26800 4905 26805 4945
rect 26845 4905 26850 4945
rect 26800 3645 26850 4905
rect 26800 3605 26805 3645
rect 26845 3605 26850 3645
rect 26800 3445 26850 3605
rect 26800 3405 26805 3445
rect 26845 3405 26850 3445
rect 26800 3400 26850 3405
rect 27100 4945 27150 4950
rect 27100 4905 27105 4945
rect 27145 4905 27150 4945
rect 27100 3645 27150 4905
rect 27100 3605 27105 3645
rect 27145 3605 27150 3645
rect 27100 3445 27150 3605
rect 27100 3405 27105 3445
rect 27145 3405 27150 3445
rect 27100 3400 27150 3405
rect 27550 4945 27600 4950
rect 27550 4905 27555 4945
rect 27595 4905 27600 4945
rect 27550 3645 27600 4905
rect 27550 3605 27555 3645
rect 27595 3605 27600 3645
rect 25750 3305 25755 3345
rect 25795 3305 25800 3345
rect 25750 3300 25800 3305
rect 27550 3345 27600 3605
rect 27550 3305 27555 3345
rect 27595 3305 27600 3345
rect 27550 3300 27600 3305
rect 27700 4945 27750 4950
rect 27700 4905 27705 4945
rect 27745 4905 27750 4945
rect 27700 3645 27750 4905
rect 27700 3605 27705 3645
rect 27745 3605 27750 3645
rect 25600 805 25605 845
rect 25645 805 25650 845
rect 25600 645 25650 805
rect 25600 605 25605 645
rect 25645 605 25650 645
rect 25600 -855 25650 605
rect 25600 -895 25605 -855
rect 25645 -895 25650 -855
rect 25600 -900 25650 -895
rect 25750 845 25800 1600
rect 25750 805 25755 845
rect 25795 805 25800 845
rect 25750 -455 25800 805
rect 25750 -495 25755 -455
rect 25795 -495 25800 -455
rect 25750 -855 25800 -495
rect 25750 -895 25755 -855
rect 25795 -895 25800 -855
rect 25750 -900 25800 -895
rect 25900 845 25950 850
rect 25900 805 25905 845
rect 25945 805 25950 845
rect 25900 645 25950 805
rect 25900 605 25905 645
rect 25945 605 25950 645
rect 25900 -855 25950 605
rect 25900 -895 25905 -855
rect 25945 -895 25950 -855
rect 25900 -900 25950 -895
rect 26200 845 26250 850
rect 26200 805 26205 845
rect 26245 805 26250 845
rect 26200 645 26250 805
rect 26200 605 26205 645
rect 26245 605 26250 645
rect 26200 -855 26250 605
rect 26200 -895 26205 -855
rect 26245 -895 26250 -855
rect 26200 -900 26250 -895
rect 26500 845 26550 850
rect 26500 805 26505 845
rect 26545 805 26550 845
rect 26500 645 26550 805
rect 26500 605 26505 645
rect 26545 605 26550 645
rect 26500 -855 26550 605
rect 26500 -895 26505 -855
rect 26545 -895 26550 -855
rect 26500 -900 26550 -895
rect 26650 845 26700 850
rect 26650 805 26655 845
rect 26695 805 26700 845
rect 26650 645 26700 805
rect 26650 605 26655 645
rect 26695 605 26700 645
rect 26650 -855 26700 605
rect 26650 -895 26655 -855
rect 26695 -895 26700 -855
rect 26650 -900 26700 -895
rect 26800 845 26850 850
rect 26800 805 26805 845
rect 26845 805 26850 845
rect 26800 645 26850 805
rect 26800 605 26805 645
rect 26845 605 26850 645
rect 26800 -855 26850 605
rect 26800 -895 26805 -855
rect 26845 -895 26850 -855
rect 26800 -900 26850 -895
rect 27100 845 27150 850
rect 27100 805 27105 845
rect 27145 805 27150 845
rect 27100 645 27150 805
rect 27100 605 27105 645
rect 27145 605 27150 645
rect 27100 -855 27150 605
rect 27100 -895 27105 -855
rect 27145 -895 27150 -855
rect 27100 -900 27150 -895
rect 27400 845 27450 850
rect 27400 805 27405 845
rect 27445 805 27450 845
rect 27400 645 27450 805
rect 27400 605 27405 645
rect 27445 605 27450 645
rect 27400 -855 27450 605
rect 27400 -895 27405 -855
rect 27445 -895 27450 -855
rect 27400 -900 27450 -895
rect 27550 845 27600 850
rect 27550 805 27555 845
rect 27595 805 27600 845
rect 27550 -455 27600 805
rect 27550 -495 27555 -455
rect 27595 -495 27600 -455
rect 27550 -855 27600 -495
rect 27550 -895 27555 -855
rect 27595 -895 27600 -855
rect 27550 -900 27600 -895
rect 27700 845 27750 3605
rect 27850 4945 27900 4950
rect 27850 4905 27855 4945
rect 27895 4905 27900 4945
rect 27850 3645 27900 4905
rect 27850 3605 27855 3645
rect 27895 3605 27900 3645
rect 27850 3345 27900 3605
rect 28300 4945 28350 4950
rect 28300 4905 28305 4945
rect 28345 4905 28350 4945
rect 28300 3845 28350 4905
rect 28300 3805 28305 3845
rect 28345 3805 28350 3845
rect 28300 3645 28350 3805
rect 28300 3605 28305 3645
rect 28345 3605 28350 3645
rect 28300 3600 28350 3605
rect 28600 4945 28650 4950
rect 28600 4905 28605 4945
rect 28645 4905 28650 4945
rect 28600 3845 28650 4905
rect 28600 3805 28605 3845
rect 28645 3805 28650 3845
rect 28600 3645 28650 3805
rect 28600 3605 28605 3645
rect 28645 3605 28650 3645
rect 28600 3600 28650 3605
rect 28750 4945 28800 4950
rect 28750 4905 28755 4945
rect 28795 4905 28800 4945
rect 28750 4545 28800 4905
rect 28750 4505 28755 4545
rect 28795 4505 28800 4545
rect 28750 3645 28800 4505
rect 28750 3605 28755 3645
rect 28795 3605 28800 3645
rect 28750 3600 28800 3605
rect 28900 4945 28950 4950
rect 28900 4905 28905 4945
rect 28945 4905 28950 4945
rect 28900 3845 28950 4905
rect 28900 3805 28905 3845
rect 28945 3805 28950 3845
rect 28900 3645 28950 3805
rect 28900 3605 28905 3645
rect 28945 3605 28950 3645
rect 28900 3600 28950 3605
rect 29200 4945 29250 4950
rect 29200 4905 29205 4945
rect 29245 4905 29250 4945
rect 29200 3845 29250 4905
rect 29200 3805 29205 3845
rect 29245 3805 29250 3845
rect 29200 3645 29250 3805
rect 29200 3605 29205 3645
rect 29245 3605 29250 3645
rect 29200 3600 29250 3605
rect 29350 4945 29400 4950
rect 29350 4905 29355 4945
rect 29395 4905 29400 4945
rect 29350 4745 29400 4905
rect 29350 4705 29355 4745
rect 29395 4705 29400 4745
rect 29350 3645 29400 4705
rect 29350 3605 29355 3645
rect 29395 3605 29400 3645
rect 29350 3600 29400 3605
rect 29650 4945 29700 4950
rect 29650 4905 29655 4945
rect 29695 4905 29700 4945
rect 29650 3845 29700 4905
rect 29650 3805 29655 3845
rect 29695 3805 29700 3845
rect 29650 3645 29700 3805
rect 29650 3605 29655 3645
rect 29695 3605 29700 3645
rect 29650 3600 29700 3605
rect 29950 4945 30000 4950
rect 29950 4905 29955 4945
rect 29995 4905 30000 4945
rect 29950 3645 30000 4905
rect 29950 3605 29955 3645
rect 29995 3605 30000 3645
rect 27850 3305 27855 3345
rect 27895 3305 27900 3345
rect 27850 3300 27900 3305
rect 29950 3345 30000 3605
rect 29950 3305 29955 3345
rect 29995 3305 30000 3345
rect 29950 3300 30000 3305
rect 30250 4945 30300 4950
rect 30250 4905 30255 4945
rect 30295 4905 30300 4945
rect 30250 3645 30300 4905
rect 30250 3605 30255 3645
rect 30295 3605 30300 3645
rect 30250 3345 30300 3605
rect 30250 3305 30255 3345
rect 30295 3305 30300 3345
rect 30250 3300 30300 3305
rect 30550 4945 30600 4950
rect 30550 4905 30555 4945
rect 30595 4905 30600 4945
rect 30550 3645 30600 4905
rect 30550 3605 30555 3645
rect 30595 3605 30600 3645
rect 30550 3345 30600 3605
rect 30550 3305 30555 3345
rect 30595 3305 30600 3345
rect 30550 3300 30600 3305
rect 30850 4945 30900 4950
rect 30850 4905 30855 4945
rect 30895 4905 30900 4945
rect 30850 3645 30900 4905
rect 30850 3605 30855 3645
rect 30895 3605 30900 3645
rect 30850 3345 30900 3605
rect 31000 4945 31050 4950
rect 31000 4905 31005 4945
rect 31045 4905 31050 4945
rect 31000 4045 31050 4905
rect 31000 4005 31005 4045
rect 31045 4005 31050 4045
rect 31000 3645 31050 4005
rect 31000 3605 31005 3645
rect 31045 3605 31050 3645
rect 31000 3600 31050 3605
rect 31450 4945 31500 4950
rect 31450 4905 31455 4945
rect 31495 4905 31500 4945
rect 31450 4745 31500 4905
rect 31450 4705 31455 4745
rect 31495 4705 31500 4745
rect 31450 3645 31500 4705
rect 31450 3605 31455 3645
rect 31495 3605 31500 3645
rect 31450 3600 31500 3605
rect 31600 4945 31650 4950
rect 31600 4905 31605 4945
rect 31645 4905 31650 4945
rect 31600 3845 31650 4905
rect 31600 3805 31605 3845
rect 31645 3805 31650 3845
rect 31600 3645 31650 3805
rect 31600 3605 31605 3645
rect 31645 3605 31650 3645
rect 31600 3600 31650 3605
rect 31900 4945 31950 4950
rect 31900 4905 31905 4945
rect 31945 4905 31950 4945
rect 31900 3845 31950 4905
rect 31900 3805 31905 3845
rect 31945 3805 31950 3845
rect 31900 3645 31950 3805
rect 31900 3605 31905 3645
rect 31945 3605 31950 3645
rect 31900 3600 31950 3605
rect 32050 4945 32100 4950
rect 32050 4905 32055 4945
rect 32095 4905 32100 4945
rect 32050 4545 32100 4905
rect 32050 4505 32055 4545
rect 32095 4505 32100 4545
rect 32050 3645 32100 4505
rect 32050 3605 32055 3645
rect 32095 3605 32100 3645
rect 32050 3600 32100 3605
rect 30850 3305 30855 3345
rect 30895 3305 30900 3345
rect 30850 3300 30900 3305
rect 27700 805 27705 845
rect 27745 805 27750 845
rect 27700 645 27750 805
rect 27700 605 27705 645
rect 27745 605 27750 645
rect 27700 -855 27750 605
rect 27700 -895 27705 -855
rect 27745 -895 27750 -855
rect 27700 -900 27750 -895
rect 28000 845 28050 850
rect 28000 805 28005 845
rect 28045 805 28050 845
rect 28000 645 28050 805
rect 28000 605 28005 645
rect 28045 605 28050 645
rect 28000 -855 28050 605
rect 28000 -895 28005 -855
rect 28045 -895 28050 -855
rect 28000 -900 28050 -895
rect 28300 845 28350 850
rect 28300 805 28305 845
rect 28345 805 28350 845
rect 28300 645 28350 805
rect 28300 605 28305 645
rect 28345 605 28350 645
rect 28300 -855 28350 605
rect 28300 -895 28305 -855
rect 28345 -895 28350 -855
rect 28300 -900 28350 -895
rect 28600 845 28650 850
rect 28600 805 28605 845
rect 28645 805 28650 845
rect 28600 645 28650 805
rect 28600 605 28605 645
rect 28645 605 28650 645
rect 28600 -855 28650 605
rect 28600 -895 28605 -855
rect 28645 -895 28650 -855
rect 28600 -900 28650 -895
<< end >>
