* num: #num corner: #corner vdd: #vdd temp: #temp

* Include SkyWater sky130 device models
.lib /usr/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice #corner
.temp #temp

.include ../../netlists/lpopamp.cc.spice

* Simulation parameters
.param xavdd  = #vdd
.param xavss  = 0
.param xen    = 1
.param xvin   = {xavdd/2}
.param xvout  = {xavdd/2}

.param xavdd_ac = 0
.param xvin_ac  = 0
.param xvout_ac = 0

.param xibias = 10u

.param xcl    = 30p
.param xrl    = 5k

.param xcl    = 30p
.param xrl    = 5k

.param xamp  = {xavdd-100m}
.param xvlo  = {xavdd/2-xamp/2}
.param xvhi  = {xavdd/2+xamp/2}
.param xper  = {40u}
.param xtdel = {xper/4}
.param xtr   = {xper/1000}
.param xpw   = {xper/2-xtr}

* Design under test
*.subckt lpopamp im o ib vsub avss avdd enb en ip
Xdut out out ibias avss avss avdd enb en in lpopamp
v_avss GND avss xavss
v_avdd avdd avss dc {xavdd} ac {xavdd_ac} 
v_in in avss pulse({xvlo} {xvhi} {xtdel} {xtr} {xtr} {xpw} {xper}) 
v_en en avss {xen*xavdd} 
v_enb enb avss {(1-xen)*xavdd} 
i_ibias avdd ibias {xen*xibias} 
CL out avss 'xcl' m=1 
v_out out_ avss dc {xvout} ac {xvout_ac} 
RL out out_ 'xrl' m=1 

* Simulation control
.option gmin=1e-12
.option rshunt=1e12
.option method=Gear
.param xtstart = 0
.param xtend   = {xper}
.param xtstep  = {xper/100}
.tran {xtstep} {xtend} {xtstart}

.save v(in) v(out)
.control
  run
  plot in out

  let avdd = 3.3
  let vhi  = avdd-50m
  let vlo  = 50m
  let vmax = vlo+0.9*(vhi-vlo)
  let vmin = vlo+0.1*(vhi-vlo)
  let dv   = vmax-vmin

  meas tran slewp trig v(out) rise=1 val=vmin targ v(out) rise=1 val=vmax
  meas tran slewm trig v(out) fall=1 val=vmax targ v(out) fall=1 val=vmin

  let slewrp = abs(dv/slewp)
  let slewrm = abs(dv/slewm)
  let slewr  = (slewrp+slewrm)/2

  print slewrp slewrm slewr

  echo "num,corner,vdd,temp,slewrp,slewrm,slewr"           >  ../meas/tb_lpopamp_buf_tran_step_large_cc.meas#num
  echo "#num,#corner,#vdd,#temp,$&slewrp,$&slewrm,$&slewr" >> ../meas/tb_lpopamp_buf_tran_step_large_cc.meas#num

  wrdata ../data/tb_lpopamp_buf_tran_sine_cc.dat#num v(in) v(out)

.endc

.GLOBAL GND 
.end 
