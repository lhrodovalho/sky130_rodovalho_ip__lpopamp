* expanding   symbol:  lpopampa.sym # of pins=8
* sym_path: /home/rodovalho/git/sky130_rodovalho_ip__lpopamp/xschem/lpopampa.sym
* sch_path: /home/rodovalho/git/sky130_rodovalho_ip__lpopamp/xschem/lpopampa.sch
.subckt lpopampa  im  ip  o  avdd  avss  en  enb  ibias
*.iopin avdd
*.iopin avss
*.iopin ip
*.iopin im
*.iopin o
*.iopin ibias
*.iopin en
*.iopin enb
xslice_1 im ip o avdd avss en enb bpa bpb bnb bna xp ypm ypp zpm zpp xn ynm ynp znm znp avss
+ lpopamp_slice
xslice_0 im ip o avdd avss en enb bpa bpb bnb bna xp ypm ypp zpm zpp xn ynm ynp znm znp avss
+ lpopamp_slice
ralias_ibias ibias bnb 1 m=1
XCp o zpm sky130_fd_pr__cap_mim_m3_1 W=90 L=90 MF=1 m=1
XCn o znm sky130_fd_pr__cap_mim_m3_1 W=90 L=90 MF=1 m=1
.ends
