magic
tech sky130A
timestamp 1714587215
<< locali >>
rect 0 0 50 50
<< metal1 >>
rect 39800 11340 39850 11350
rect 39800 11310 39810 11340
rect 39840 11310 39850 11340
rect 39800 11300 39850 11310
rect 39900 11240 40900 11250
rect 39900 11210 39910 11240
rect 39940 11210 39960 11240
rect 39990 11210 40010 11240
rect 40040 11210 40060 11240
rect 40090 11210 40110 11240
rect 40140 11210 40160 11240
rect 40190 11210 40210 11240
rect 40240 11210 40260 11240
rect 40290 11210 40310 11240
rect 40340 11210 40360 11240
rect 40390 11210 40410 11240
rect 40440 11210 40460 11240
rect 40490 11210 40510 11240
rect 40540 11210 40560 11240
rect 40590 11210 40610 11240
rect 40640 11210 40660 11240
rect 40690 11210 40710 11240
rect 40740 11210 40760 11240
rect 40790 11210 40810 11240
rect 40840 11210 40860 11240
rect 40890 11210 40900 11240
rect 39900 11190 40900 11210
rect 39900 11160 39910 11190
rect 39940 11160 39960 11190
rect 39990 11160 40010 11190
rect 40040 11160 40060 11190
rect 40090 11160 40110 11190
rect 40140 11160 40160 11190
rect 40190 11160 40210 11190
rect 40240 11160 40260 11190
rect 40290 11160 40310 11190
rect 40340 11160 40360 11190
rect 40390 11160 40410 11190
rect 40440 11160 40460 11190
rect 40490 11160 40510 11190
rect 40540 11160 40560 11190
rect 40590 11160 40610 11190
rect 40640 11160 40660 11190
rect 40690 11160 40710 11190
rect 40740 11160 40760 11190
rect 40790 11160 40810 11190
rect 40840 11160 40860 11190
rect 40890 11160 40900 11190
rect 39900 11140 40900 11160
rect 39900 11110 39910 11140
rect 39940 11110 39960 11140
rect 39990 11110 40010 11140
rect 40040 11110 40060 11140
rect 40090 11110 40110 11140
rect 40140 11110 40160 11140
rect 40190 11110 40210 11140
rect 40240 11110 40260 11140
rect 40290 11110 40310 11140
rect 40340 11110 40360 11140
rect 40390 11110 40410 11140
rect 40440 11110 40460 11140
rect 40490 11110 40510 11140
rect 40540 11110 40560 11140
rect 40590 11110 40610 11140
rect 40640 11110 40660 11140
rect 40690 11110 40710 11140
rect 40740 11110 40760 11140
rect 40790 11110 40810 11140
rect 40840 11110 40860 11140
rect 40890 11110 40900 11140
rect 39900 11090 40900 11110
rect 39900 11060 39910 11090
rect 39940 11060 39960 11090
rect 39990 11060 40010 11090
rect 40040 11060 40060 11090
rect 40090 11060 40110 11090
rect 40140 11060 40160 11090
rect 40190 11060 40210 11090
rect 40240 11060 40260 11090
rect 40290 11060 40310 11090
rect 40340 11060 40360 11090
rect 40390 11060 40410 11090
rect 40440 11060 40460 11090
rect 40490 11060 40510 11090
rect 40540 11060 40560 11090
rect 40590 11060 40610 11090
rect 40640 11060 40660 11090
rect 40690 11060 40710 11090
rect 40740 11060 40760 11090
rect 40790 11060 40810 11090
rect 40840 11060 40860 11090
rect 40890 11060 40900 11090
rect 39900 11040 40900 11060
rect 39900 11010 39910 11040
rect 39940 11010 39960 11040
rect 39990 11010 40010 11040
rect 40040 11010 40060 11040
rect 40090 11010 40110 11040
rect 40140 11010 40160 11040
rect 40190 11010 40210 11040
rect 40240 11010 40260 11040
rect 40290 11010 40310 11040
rect 40340 11010 40360 11040
rect 40390 11010 40410 11040
rect 40440 11010 40460 11040
rect 40490 11010 40510 11040
rect 40540 11010 40560 11040
rect 40590 11010 40610 11040
rect 40640 11010 40660 11040
rect 40690 11010 40710 11040
rect 40740 11010 40760 11040
rect 40790 11010 40810 11040
rect 40840 11010 40860 11040
rect 40890 11010 40900 11040
rect 39900 11000 40900 11010
rect 39800 10940 39850 10950
rect 39800 10910 39810 10940
rect 39840 10910 39850 10940
rect 39800 10900 39850 10910
rect 39800 4740 39850 4750
rect 39800 4710 39810 4740
rect 39840 4710 39850 4740
rect 39800 4700 39850 4710
rect 39900 4640 40900 4650
rect 39900 4610 39910 4640
rect 39940 4610 39960 4640
rect 39990 4610 40010 4640
rect 40040 4610 40060 4640
rect 40090 4610 40110 4640
rect 40140 4610 40160 4640
rect 40190 4610 40210 4640
rect 40240 4610 40260 4640
rect 40290 4610 40310 4640
rect 40340 4610 40360 4640
rect 40390 4610 40410 4640
rect 40440 4610 40460 4640
rect 40490 4610 40510 4640
rect 40540 4610 40560 4640
rect 40590 4610 40610 4640
rect 40640 4610 40660 4640
rect 40690 4610 40710 4640
rect 40740 4610 40760 4640
rect 40790 4610 40810 4640
rect 40840 4610 40860 4640
rect 40890 4610 40900 4640
rect 39900 4590 40900 4610
rect 39900 4560 39910 4590
rect 39940 4560 39960 4590
rect 39990 4560 40010 4590
rect 40040 4560 40060 4590
rect 40090 4560 40110 4590
rect 40140 4560 40160 4590
rect 40190 4560 40210 4590
rect 40240 4560 40260 4590
rect 40290 4560 40310 4590
rect 40340 4560 40360 4590
rect 40390 4560 40410 4590
rect 40440 4560 40460 4590
rect 40490 4560 40510 4590
rect 40540 4560 40560 4590
rect 40590 4560 40610 4590
rect 40640 4560 40660 4590
rect 40690 4560 40710 4590
rect 40740 4560 40760 4590
rect 40790 4560 40810 4590
rect 40840 4560 40860 4590
rect 40890 4560 40900 4590
rect 39900 4540 40900 4560
rect 39900 4510 39910 4540
rect 39940 4510 39960 4540
rect 39990 4510 40010 4540
rect 40040 4510 40060 4540
rect 40090 4510 40110 4540
rect 40140 4510 40160 4540
rect 40190 4510 40210 4540
rect 40240 4510 40260 4540
rect 40290 4510 40310 4540
rect 40340 4510 40360 4540
rect 40390 4510 40410 4540
rect 40440 4510 40460 4540
rect 40490 4510 40510 4540
rect 40540 4510 40560 4540
rect 40590 4510 40610 4540
rect 40640 4510 40660 4540
rect 40690 4510 40710 4540
rect 40740 4510 40760 4540
rect 40790 4510 40810 4540
rect 40840 4510 40860 4540
rect 40890 4510 40900 4540
rect 39900 4490 40900 4510
rect 39900 4460 39910 4490
rect 39940 4460 39960 4490
rect 39990 4460 40010 4490
rect 40040 4460 40060 4490
rect 40090 4460 40110 4490
rect 40140 4460 40160 4490
rect 40190 4460 40210 4490
rect 40240 4460 40260 4490
rect 40290 4460 40310 4490
rect 40340 4460 40360 4490
rect 40390 4460 40410 4490
rect 40440 4460 40460 4490
rect 40490 4460 40510 4490
rect 40540 4460 40560 4490
rect 40590 4460 40610 4490
rect 40640 4460 40660 4490
rect 40690 4460 40710 4490
rect 40740 4460 40760 4490
rect 40790 4460 40810 4490
rect 40840 4460 40860 4490
rect 40890 4460 40900 4490
rect 39900 4440 40900 4460
rect 39900 4410 39910 4440
rect 39940 4410 39960 4440
rect 39990 4410 40010 4440
rect 40040 4410 40060 4440
rect 40090 4410 40110 4440
rect 40140 4410 40160 4440
rect 40190 4410 40210 4440
rect 40240 4410 40260 4440
rect 40290 4410 40310 4440
rect 40340 4410 40360 4440
rect 40390 4410 40410 4440
rect 40440 4410 40460 4440
rect 40490 4410 40510 4440
rect 40540 4410 40560 4440
rect 40590 4410 40610 4440
rect 40640 4410 40660 4440
rect 40690 4410 40710 4440
rect 40740 4410 40760 4440
rect 40790 4410 40810 4440
rect 40840 4410 40860 4440
rect 40890 4410 40900 4440
rect 39900 4400 40900 4410
rect 39800 4340 39850 4350
rect 39800 4310 39810 4340
rect 39840 4310 39850 4340
rect 39800 4300 39850 4310
<< via1 >>
rect 39810 11310 39840 11340
rect 39910 11210 39940 11240
rect 39960 11210 39990 11240
rect 40010 11210 40040 11240
rect 40060 11210 40090 11240
rect 40110 11210 40140 11240
rect 40160 11210 40190 11240
rect 40210 11210 40240 11240
rect 40260 11210 40290 11240
rect 40310 11210 40340 11240
rect 40360 11210 40390 11240
rect 40410 11210 40440 11240
rect 40460 11210 40490 11240
rect 40510 11210 40540 11240
rect 40560 11210 40590 11240
rect 40610 11210 40640 11240
rect 40660 11210 40690 11240
rect 40710 11210 40740 11240
rect 40760 11210 40790 11240
rect 40810 11210 40840 11240
rect 40860 11210 40890 11240
rect 39910 11160 39940 11190
rect 39960 11160 39990 11190
rect 40010 11160 40040 11190
rect 40060 11160 40090 11190
rect 40110 11160 40140 11190
rect 40160 11160 40190 11190
rect 40210 11160 40240 11190
rect 40260 11160 40290 11190
rect 40310 11160 40340 11190
rect 40360 11160 40390 11190
rect 40410 11160 40440 11190
rect 40460 11160 40490 11190
rect 40510 11160 40540 11190
rect 40560 11160 40590 11190
rect 40610 11160 40640 11190
rect 40660 11160 40690 11190
rect 40710 11160 40740 11190
rect 40760 11160 40790 11190
rect 40810 11160 40840 11190
rect 40860 11160 40890 11190
rect 39910 11110 39940 11140
rect 39960 11110 39990 11140
rect 40010 11110 40040 11140
rect 40060 11110 40090 11140
rect 40110 11110 40140 11140
rect 40160 11110 40190 11140
rect 40210 11110 40240 11140
rect 40260 11110 40290 11140
rect 40310 11110 40340 11140
rect 40360 11110 40390 11140
rect 40410 11110 40440 11140
rect 40460 11110 40490 11140
rect 40510 11110 40540 11140
rect 40560 11110 40590 11140
rect 40610 11110 40640 11140
rect 40660 11110 40690 11140
rect 40710 11110 40740 11140
rect 40760 11110 40790 11140
rect 40810 11110 40840 11140
rect 40860 11110 40890 11140
rect 39910 11060 39940 11090
rect 39960 11060 39990 11090
rect 40010 11060 40040 11090
rect 40060 11060 40090 11090
rect 40110 11060 40140 11090
rect 40160 11060 40190 11090
rect 40210 11060 40240 11090
rect 40260 11060 40290 11090
rect 40310 11060 40340 11090
rect 40360 11060 40390 11090
rect 40410 11060 40440 11090
rect 40460 11060 40490 11090
rect 40510 11060 40540 11090
rect 40560 11060 40590 11090
rect 40610 11060 40640 11090
rect 40660 11060 40690 11090
rect 40710 11060 40740 11090
rect 40760 11060 40790 11090
rect 40810 11060 40840 11090
rect 40860 11060 40890 11090
rect 39910 11010 39940 11040
rect 39960 11010 39990 11040
rect 40010 11010 40040 11040
rect 40060 11010 40090 11040
rect 40110 11010 40140 11040
rect 40160 11010 40190 11040
rect 40210 11010 40240 11040
rect 40260 11010 40290 11040
rect 40310 11010 40340 11040
rect 40360 11010 40390 11040
rect 40410 11010 40440 11040
rect 40460 11010 40490 11040
rect 40510 11010 40540 11040
rect 40560 11010 40590 11040
rect 40610 11010 40640 11040
rect 40660 11010 40690 11040
rect 40710 11010 40740 11040
rect 40760 11010 40790 11040
rect 40810 11010 40840 11040
rect 40860 11010 40890 11040
rect 39810 10910 39840 10940
rect 39810 4710 39840 4740
rect 39910 4610 39940 4640
rect 39960 4610 39990 4640
rect 40010 4610 40040 4640
rect 40060 4610 40090 4640
rect 40110 4610 40140 4640
rect 40160 4610 40190 4640
rect 40210 4610 40240 4640
rect 40260 4610 40290 4640
rect 40310 4610 40340 4640
rect 40360 4610 40390 4640
rect 40410 4610 40440 4640
rect 40460 4610 40490 4640
rect 40510 4610 40540 4640
rect 40560 4610 40590 4640
rect 40610 4610 40640 4640
rect 40660 4610 40690 4640
rect 40710 4610 40740 4640
rect 40760 4610 40790 4640
rect 40810 4610 40840 4640
rect 40860 4610 40890 4640
rect 39910 4560 39940 4590
rect 39960 4560 39990 4590
rect 40010 4560 40040 4590
rect 40060 4560 40090 4590
rect 40110 4560 40140 4590
rect 40160 4560 40190 4590
rect 40210 4560 40240 4590
rect 40260 4560 40290 4590
rect 40310 4560 40340 4590
rect 40360 4560 40390 4590
rect 40410 4560 40440 4590
rect 40460 4560 40490 4590
rect 40510 4560 40540 4590
rect 40560 4560 40590 4590
rect 40610 4560 40640 4590
rect 40660 4560 40690 4590
rect 40710 4560 40740 4590
rect 40760 4560 40790 4590
rect 40810 4560 40840 4590
rect 40860 4560 40890 4590
rect 39910 4510 39940 4540
rect 39960 4510 39990 4540
rect 40010 4510 40040 4540
rect 40060 4510 40090 4540
rect 40110 4510 40140 4540
rect 40160 4510 40190 4540
rect 40210 4510 40240 4540
rect 40260 4510 40290 4540
rect 40310 4510 40340 4540
rect 40360 4510 40390 4540
rect 40410 4510 40440 4540
rect 40460 4510 40490 4540
rect 40510 4510 40540 4540
rect 40560 4510 40590 4540
rect 40610 4510 40640 4540
rect 40660 4510 40690 4540
rect 40710 4510 40740 4540
rect 40760 4510 40790 4540
rect 40810 4510 40840 4540
rect 40860 4510 40890 4540
rect 39910 4460 39940 4490
rect 39960 4460 39990 4490
rect 40010 4460 40040 4490
rect 40060 4460 40090 4490
rect 40110 4460 40140 4490
rect 40160 4460 40190 4490
rect 40210 4460 40240 4490
rect 40260 4460 40290 4490
rect 40310 4460 40340 4490
rect 40360 4460 40390 4490
rect 40410 4460 40440 4490
rect 40460 4460 40490 4490
rect 40510 4460 40540 4490
rect 40560 4460 40590 4490
rect 40610 4460 40640 4490
rect 40660 4460 40690 4490
rect 40710 4460 40740 4490
rect 40760 4460 40790 4490
rect 40810 4460 40840 4490
rect 40860 4460 40890 4490
rect 39910 4410 39940 4440
rect 39960 4410 39990 4440
rect 40010 4410 40040 4440
rect 40060 4410 40090 4440
rect 40110 4410 40140 4440
rect 40160 4410 40190 4440
rect 40210 4410 40240 4440
rect 40260 4410 40290 4440
rect 40310 4410 40340 4440
rect 40360 4410 40390 4440
rect 40410 4410 40440 4440
rect 40460 4410 40490 4440
rect 40510 4410 40540 4440
rect 40560 4410 40590 4440
rect 40610 4410 40640 4440
rect 40660 4410 40690 4440
rect 40710 4410 40740 4440
rect 40760 4410 40790 4440
rect 40810 4410 40840 4440
rect 40860 4410 40890 4440
rect 39810 4310 39840 4340
<< metal2 >>
rect -3500 17010 -50 17020
rect -3500 16980 -3490 17010
rect -3460 16980 -3290 17010
rect -3260 16980 -3090 17010
rect -3060 16980 -1590 17010
rect -1560 16980 -1190 17010
rect -1160 16980 -1090 17010
rect -1060 16980 -990 17010
rect -960 16980 -890 17010
rect -860 16980 -790 17010
rect -760 16980 -690 17010
rect -660 16980 -590 17010
rect -560 16980 -490 17010
rect -460 16980 -390 17010
rect -360 16980 -290 17010
rect -260 16980 -190 17010
rect -160 16980 -90 17010
rect -60 16980 -50 17010
rect -3500 16970 -50 16980
rect -3500 15740 -50 15750
rect -3500 15710 -3490 15740
rect -3460 15710 -3290 15740
rect -3260 15710 -3090 15740
rect -3060 15710 -1590 15740
rect -1560 15710 -1190 15740
rect -1160 15710 -1090 15740
rect -1060 15710 -990 15740
rect -960 15710 -890 15740
rect -860 15710 -690 15740
rect -660 15710 -590 15740
rect -560 15710 -490 15740
rect -460 15710 -290 15740
rect -260 15710 -190 15740
rect -160 15710 -90 15740
rect -60 15710 -50 15740
rect -3500 15700 -50 15710
rect -3500 15340 0 15350
rect -3500 15310 -3490 15340
rect -3460 15310 -3290 15340
rect -3260 15310 -3090 15340
rect -3060 15310 -1590 15340
rect -1560 15310 -1090 15340
rect -1060 15310 -890 15340
rect -860 15310 -690 15340
rect -660 15310 -490 15340
rect -460 15310 -290 15340
rect -260 15310 -90 15340
rect -60 15310 0 15340
rect -3500 15290 0 15310
rect -3500 15260 -3490 15290
rect -3460 15260 -3290 15290
rect -3260 15260 -3090 15290
rect -3060 15260 -1590 15290
rect -1560 15260 -1090 15290
rect -1060 15260 -890 15290
rect -860 15260 -690 15290
rect -660 15260 -490 15290
rect -460 15260 -290 15290
rect -260 15260 -90 15290
rect -60 15260 0 15290
rect -3500 15240 0 15260
rect -3500 15210 -3490 15240
rect -3460 15210 -3290 15240
rect -3260 15210 -3090 15240
rect -3060 15210 -1590 15240
rect -1560 15210 -1090 15240
rect -1060 15210 -890 15240
rect -860 15210 -690 15240
rect -660 15210 -490 15240
rect -460 15210 -290 15240
rect -260 15210 -90 15240
rect -60 15210 0 15240
rect -3500 15200 0 15210
rect -3500 13640 0 13650
rect -3500 13610 -3490 13640
rect -3460 13610 -3290 13640
rect -3260 13610 -3090 13640
rect -3060 13610 -1590 13640
rect -1560 13610 -1090 13640
rect -1060 13610 -890 13640
rect -860 13610 -690 13640
rect -660 13610 -490 13640
rect -460 13610 -290 13640
rect -260 13610 -90 13640
rect -60 13610 0 13640
rect -3500 13590 0 13610
rect -3500 13560 -3490 13590
rect -3460 13560 -3290 13590
rect -3260 13560 -3090 13590
rect -3060 13560 -1590 13590
rect -1560 13560 -1090 13590
rect -1060 13560 -890 13590
rect -860 13560 -690 13590
rect -660 13560 -490 13590
rect -460 13560 -290 13590
rect -260 13560 -90 13590
rect -60 13560 0 13590
rect -3500 13540 0 13560
rect -3500 13510 -3490 13540
rect -3460 13510 -3290 13540
rect -3260 13510 -3090 13540
rect -3060 13510 -1590 13540
rect -1560 13510 -1090 13540
rect -1060 13510 -890 13540
rect -860 13510 -690 13540
rect -660 13510 -490 13540
rect -460 13510 -290 13540
rect -260 13510 -90 13540
rect -60 13510 0 13540
rect -3500 13500 0 13510
rect -3500 11940 0 11950
rect -3500 11910 -3490 11940
rect -3460 11910 -3290 11940
rect -3260 11910 -3090 11940
rect -3060 11910 -1590 11940
rect -1560 11910 -1090 11940
rect -1060 11910 -890 11940
rect -860 11910 -690 11940
rect -660 11910 -490 11940
rect -460 11910 -290 11940
rect -260 11910 -90 11940
rect -60 11910 0 11940
rect -3500 11890 0 11910
rect -3500 11860 -3490 11890
rect -3460 11860 -3290 11890
rect -3260 11860 -3090 11890
rect -3060 11860 -1590 11890
rect -1560 11860 -1090 11890
rect -1060 11860 -890 11890
rect -860 11860 -690 11890
rect -660 11860 -490 11890
rect -460 11860 -290 11890
rect -260 11860 -90 11890
rect -60 11860 0 11890
rect -3500 11840 0 11860
rect -3500 11810 -3490 11840
rect -3460 11810 -3290 11840
rect -3260 11810 -3090 11840
rect -3060 11810 -1590 11840
rect -1560 11810 -1090 11840
rect -1060 11810 -890 11840
rect -860 11810 -690 11840
rect -660 11810 -490 11840
rect -460 11810 -290 11840
rect -260 11810 -90 11840
rect -60 11810 0 11840
rect -3500 11800 0 11810
rect 39750 11340 39900 11350
rect 39750 11310 39810 11340
rect 39840 11310 39900 11340
rect 39750 11300 39900 11310
rect 39750 11240 40900 11250
rect 39750 11210 39910 11240
rect 39940 11210 39960 11240
rect 39990 11210 40010 11240
rect 40040 11210 40060 11240
rect 40090 11210 40110 11240
rect 40140 11210 40160 11240
rect 40190 11210 40210 11240
rect 40240 11210 40260 11240
rect 40290 11210 40310 11240
rect 40340 11210 40360 11240
rect 40390 11210 40410 11240
rect 40440 11210 40460 11240
rect 40490 11210 40510 11240
rect 40540 11210 40560 11240
rect 40590 11210 40610 11240
rect 40640 11210 40660 11240
rect 40690 11210 40710 11240
rect 40740 11210 40760 11240
rect 40790 11210 40810 11240
rect 40840 11210 40860 11240
rect 40890 11210 40900 11240
rect 39750 11190 40900 11210
rect 39750 11160 39910 11190
rect 39940 11160 39960 11190
rect 39990 11160 40010 11190
rect 40040 11160 40060 11190
rect 40090 11160 40110 11190
rect 40140 11160 40160 11190
rect 40190 11160 40210 11190
rect 40240 11160 40260 11190
rect 40290 11160 40310 11190
rect 40340 11160 40360 11190
rect 40390 11160 40410 11190
rect 40440 11160 40460 11190
rect 40490 11160 40510 11190
rect 40540 11160 40560 11190
rect 40590 11160 40610 11190
rect 40640 11160 40660 11190
rect 40690 11160 40710 11190
rect 40740 11160 40760 11190
rect 40790 11160 40810 11190
rect 40840 11160 40860 11190
rect 40890 11160 40900 11190
rect 39750 11140 40900 11160
rect 39750 11110 39910 11140
rect 39940 11110 39960 11140
rect 39990 11110 40010 11140
rect 40040 11110 40060 11140
rect 40090 11110 40110 11140
rect 40140 11110 40160 11140
rect 40190 11110 40210 11140
rect 40240 11110 40260 11140
rect 40290 11110 40310 11140
rect 40340 11110 40360 11140
rect 40390 11110 40410 11140
rect 40440 11110 40460 11140
rect 40490 11110 40510 11140
rect 40540 11110 40560 11140
rect 40590 11110 40610 11140
rect 40640 11110 40660 11140
rect 40690 11110 40710 11140
rect 40740 11110 40760 11140
rect 40790 11110 40810 11140
rect 40840 11110 40860 11140
rect 40890 11110 40900 11140
rect 39750 11090 40900 11110
rect 39750 11060 39910 11090
rect 39940 11060 39960 11090
rect 39990 11060 40010 11090
rect 40040 11060 40060 11090
rect 40090 11060 40110 11090
rect 40140 11060 40160 11090
rect 40190 11060 40210 11090
rect 40240 11060 40260 11090
rect 40290 11060 40310 11090
rect 40340 11060 40360 11090
rect 40390 11060 40410 11090
rect 40440 11060 40460 11090
rect 40490 11060 40510 11090
rect 40540 11060 40560 11090
rect 40590 11060 40610 11090
rect 40640 11060 40660 11090
rect 40690 11060 40710 11090
rect 40740 11060 40760 11090
rect 40790 11060 40810 11090
rect 40840 11060 40860 11090
rect 40890 11060 40900 11090
rect 39750 11040 40900 11060
rect 39750 11010 39910 11040
rect 39940 11010 39960 11040
rect 39990 11010 40010 11040
rect 40040 11010 40060 11040
rect 40090 11010 40110 11040
rect 40140 11010 40160 11040
rect 40190 11010 40210 11040
rect 40240 11010 40260 11040
rect 40290 11010 40310 11040
rect 40340 11010 40360 11040
rect 40390 11010 40410 11040
rect 40440 11010 40460 11040
rect 40490 11010 40510 11040
rect 40540 11010 40560 11040
rect 40590 11010 40610 11040
rect 40640 11010 40660 11040
rect 40690 11010 40710 11040
rect 40740 11010 40760 11040
rect 40790 11010 40810 11040
rect 40840 11010 40860 11040
rect 40890 11010 40900 11040
rect 39750 11000 40900 11010
rect 39750 10940 39900 10950
rect 39750 10910 39810 10940
rect 39840 10910 39900 10940
rect 39750 10900 39900 10910
rect -3100 10640 0 10650
rect -3100 10610 -2990 10640
rect -2960 10610 -2790 10640
rect -2760 10610 -2590 10640
rect -2560 10610 -2390 10640
rect -2360 10610 -2190 10640
rect -2160 10610 -1990 10640
rect -1960 10610 -1690 10640
rect -1660 10610 0 10640
rect -3100 10590 0 10610
rect -3100 10560 -2990 10590
rect -2960 10560 -2790 10590
rect -2760 10560 -2590 10590
rect -2560 10560 -2390 10590
rect -2360 10560 -2190 10590
rect -2160 10560 -1990 10590
rect -1960 10560 -1690 10590
rect -1660 10560 0 10590
rect -3100 10540 0 10560
rect -3100 10510 -2990 10540
rect -2960 10510 -2790 10540
rect -2760 10510 -2590 10540
rect -2560 10510 -2390 10540
rect -2360 10510 -2190 10540
rect -2160 10510 -1990 10540
rect -1960 10510 -1690 10540
rect -1660 10510 0 10540
rect -3100 10500 0 10510
rect -3100 9340 0 9350
rect -3100 9310 -2990 9340
rect -2960 9310 -2790 9340
rect -2760 9310 -2590 9340
rect -2560 9310 -2390 9340
rect -2360 9310 -2190 9340
rect -2160 9310 -1990 9340
rect -1960 9310 -1690 9340
rect -1660 9310 0 9340
rect -3100 9290 0 9310
rect -3100 9260 -2990 9290
rect -2960 9260 -2790 9290
rect -2760 9260 -2590 9290
rect -2560 9260 -2390 9290
rect -2360 9260 -2190 9290
rect -2160 9260 -1990 9290
rect -1960 9260 -1690 9290
rect -1660 9260 0 9290
rect -3100 9240 0 9260
rect -3100 9210 -2990 9240
rect -2960 9210 -2790 9240
rect -2760 9210 -2590 9240
rect -2560 9210 -2390 9240
rect -2360 9210 -2190 9240
rect -2160 9210 -1990 9240
rect -1960 9210 -1690 9240
rect -1660 9210 0 9240
rect -3100 9200 0 9210
rect -3100 8040 0 8050
rect -3100 8010 -2990 8040
rect -2960 8010 -2790 8040
rect -2760 8010 -2590 8040
rect -2560 8010 -2390 8040
rect -2360 8010 -2190 8040
rect -2160 8010 -1990 8040
rect -1960 8010 -1690 8040
rect -1660 8010 0 8040
rect -3100 7990 0 8010
rect -3100 7960 -2990 7990
rect -2960 7960 -2790 7990
rect -2760 7960 -2590 7990
rect -2560 7960 -2390 7990
rect -2360 7960 -2190 7990
rect -2160 7960 -1990 7990
rect -1960 7960 -1690 7990
rect -1660 7960 0 7990
rect -3100 7940 0 7960
rect -3100 7910 -2990 7940
rect -2960 7910 -2790 7940
rect -2760 7910 -2590 7940
rect -2560 7910 -2390 7940
rect -2360 7910 -2190 7940
rect -2160 7910 -1990 7940
rect -1960 7910 -1690 7940
rect -1660 7910 0 7940
rect -3100 7900 0 7910
rect -3100 7740 0 7750
rect -3100 7710 -2990 7740
rect -2960 7710 -2790 7740
rect -2760 7710 -2590 7740
rect -2560 7710 -2390 7740
rect -2360 7710 -2190 7740
rect -2160 7710 -1990 7740
rect -1960 7710 -1690 7740
rect -1660 7710 0 7740
rect -3100 7690 0 7710
rect -3100 7660 -2990 7690
rect -2960 7660 -2790 7690
rect -2760 7660 -2590 7690
rect -2560 7660 -2390 7690
rect -2360 7660 -2190 7690
rect -2160 7660 -1990 7690
rect -1960 7660 -1690 7690
rect -1660 7660 0 7690
rect -3100 7640 0 7660
rect -3100 7610 -2990 7640
rect -2960 7610 -2790 7640
rect -2760 7610 -2590 7640
rect -2560 7610 -2390 7640
rect -2360 7610 -2190 7640
rect -2160 7610 -1990 7640
rect -1960 7610 -1690 7640
rect -1660 7610 0 7640
rect -3100 7600 0 7610
rect -3100 6440 0 6450
rect -3100 6410 -2990 6440
rect -2960 6410 -2790 6440
rect -2760 6410 -2590 6440
rect -2560 6410 -2390 6440
rect -2360 6410 -2190 6440
rect -2160 6410 -1990 6440
rect -1960 6410 -1690 6440
rect -1660 6410 0 6440
rect -3100 6390 0 6410
rect -3100 6360 -2990 6390
rect -2960 6360 -2790 6390
rect -2760 6360 -2590 6390
rect -2560 6360 -2390 6390
rect -2360 6360 -2190 6390
rect -2160 6360 -1990 6390
rect -1960 6360 -1690 6390
rect -1660 6360 0 6390
rect -3100 6340 0 6360
rect -3100 6310 -2990 6340
rect -2960 6310 -2790 6340
rect -2760 6310 -2590 6340
rect -2560 6310 -2390 6340
rect -2360 6310 -2190 6340
rect -2160 6310 -1990 6340
rect -1960 6310 -1690 6340
rect -1660 6310 0 6340
rect -3100 6300 0 6310
rect -3100 5140 0 5150
rect -3100 5110 -2990 5140
rect -2960 5110 -2790 5140
rect -2760 5110 -2590 5140
rect -2560 5110 -2390 5140
rect -2360 5110 -2190 5140
rect -2160 5110 -1990 5140
rect -1960 5110 -1690 5140
rect -1660 5110 0 5140
rect -3100 5090 0 5110
rect -3100 5060 -2990 5090
rect -2960 5060 -2790 5090
rect -2760 5060 -2590 5090
rect -2560 5060 -2390 5090
rect -2360 5060 -2190 5090
rect -2160 5060 -1990 5090
rect -1960 5060 -1690 5090
rect -1660 5060 0 5090
rect -3100 5040 0 5060
rect -3100 5010 -2990 5040
rect -2960 5010 -2790 5040
rect -2760 5010 -2590 5040
rect -2560 5010 -2390 5040
rect -2360 5010 -2190 5040
rect -2160 5010 -1990 5040
rect -1960 5010 -1690 5040
rect -1660 5010 0 5040
rect -3100 5000 0 5010
rect 39750 4740 39900 4750
rect 39750 4710 39810 4740
rect 39840 4710 39900 4740
rect 39750 4700 39900 4710
rect 39750 4640 40900 4650
rect 39750 4610 39910 4640
rect 39940 4610 39960 4640
rect 39990 4610 40010 4640
rect 40040 4610 40060 4640
rect 40090 4610 40110 4640
rect 40140 4610 40160 4640
rect 40190 4610 40210 4640
rect 40240 4610 40260 4640
rect 40290 4610 40310 4640
rect 40340 4610 40360 4640
rect 40390 4610 40410 4640
rect 40440 4610 40460 4640
rect 40490 4610 40510 4640
rect 40540 4610 40560 4640
rect 40590 4610 40610 4640
rect 40640 4610 40660 4640
rect 40690 4610 40710 4640
rect 40740 4610 40760 4640
rect 40790 4610 40810 4640
rect 40840 4610 40860 4640
rect 40890 4610 40900 4640
rect 39750 4590 40900 4610
rect 39750 4560 39910 4590
rect 39940 4560 39960 4590
rect 39990 4560 40010 4590
rect 40040 4560 40060 4590
rect 40090 4560 40110 4590
rect 40140 4560 40160 4590
rect 40190 4560 40210 4590
rect 40240 4560 40260 4590
rect 40290 4560 40310 4590
rect 40340 4560 40360 4590
rect 40390 4560 40410 4590
rect 40440 4560 40460 4590
rect 40490 4560 40510 4590
rect 40540 4560 40560 4590
rect 40590 4560 40610 4590
rect 40640 4560 40660 4590
rect 40690 4560 40710 4590
rect 40740 4560 40760 4590
rect 40790 4560 40810 4590
rect 40840 4560 40860 4590
rect 40890 4560 40900 4590
rect 39750 4540 40900 4560
rect 39750 4510 39910 4540
rect 39940 4510 39960 4540
rect 39990 4510 40010 4540
rect 40040 4510 40060 4540
rect 40090 4510 40110 4540
rect 40140 4510 40160 4540
rect 40190 4510 40210 4540
rect 40240 4510 40260 4540
rect 40290 4510 40310 4540
rect 40340 4510 40360 4540
rect 40390 4510 40410 4540
rect 40440 4510 40460 4540
rect 40490 4510 40510 4540
rect 40540 4510 40560 4540
rect 40590 4510 40610 4540
rect 40640 4510 40660 4540
rect 40690 4510 40710 4540
rect 40740 4510 40760 4540
rect 40790 4510 40810 4540
rect 40840 4510 40860 4540
rect 40890 4510 40900 4540
rect 39750 4490 40900 4510
rect 39750 4460 39910 4490
rect 39940 4460 39960 4490
rect 39990 4460 40010 4490
rect 40040 4460 40060 4490
rect 40090 4460 40110 4490
rect 40140 4460 40160 4490
rect 40190 4460 40210 4490
rect 40240 4460 40260 4490
rect 40290 4460 40310 4490
rect 40340 4460 40360 4490
rect 40390 4460 40410 4490
rect 40440 4460 40460 4490
rect 40490 4460 40510 4490
rect 40540 4460 40560 4490
rect 40590 4460 40610 4490
rect 40640 4460 40660 4490
rect 40690 4460 40710 4490
rect 40740 4460 40760 4490
rect 40790 4460 40810 4490
rect 40840 4460 40860 4490
rect 40890 4460 40900 4490
rect 39750 4440 40900 4460
rect 39750 4410 39910 4440
rect 39940 4410 39960 4440
rect 39990 4410 40010 4440
rect 40040 4410 40060 4440
rect 40090 4410 40110 4440
rect 40140 4410 40160 4440
rect 40190 4410 40210 4440
rect 40240 4410 40260 4440
rect 40290 4410 40310 4440
rect 40340 4410 40360 4440
rect 40390 4410 40410 4440
rect 40440 4410 40460 4440
rect 40490 4410 40510 4440
rect 40540 4410 40560 4440
rect 40590 4410 40610 4440
rect 40640 4410 40660 4440
rect 40690 4410 40710 4440
rect 40740 4410 40760 4440
rect 40790 4410 40810 4440
rect 40840 4410 40860 4440
rect 40890 4410 40900 4440
rect 39750 4400 40900 4410
rect 39750 4340 39900 4350
rect 39750 4310 39810 4340
rect 39840 4310 39900 4340
rect 39750 4300 39900 4310
rect -3500 3840 0 3850
rect -3500 3810 -3490 3840
rect -3460 3810 -3290 3840
rect -3260 3810 -3090 3840
rect -3060 3810 -1590 3840
rect -1560 3810 -1090 3840
rect -1060 3810 -890 3840
rect -860 3810 -690 3840
rect -660 3810 -490 3840
rect -460 3810 -290 3840
rect -260 3810 -90 3840
rect -60 3810 0 3840
rect -3500 3790 0 3810
rect -3500 3760 -3490 3790
rect -3460 3760 -3290 3790
rect -3260 3760 -3090 3790
rect -3060 3760 -1590 3790
rect -1560 3760 -1090 3790
rect -1060 3760 -890 3790
rect -860 3760 -690 3790
rect -660 3760 -490 3790
rect -460 3760 -290 3790
rect -260 3760 -90 3790
rect -60 3760 0 3790
rect -3500 3740 0 3760
rect -3500 3710 -3490 3740
rect -3460 3710 -3290 3740
rect -3260 3710 -3090 3740
rect -3060 3710 -1590 3740
rect -1560 3710 -1090 3740
rect -1060 3710 -890 3740
rect -860 3710 -690 3740
rect -660 3710 -490 3740
rect -460 3710 -290 3740
rect -260 3710 -90 3740
rect -60 3710 0 3740
rect -3500 3700 0 3710
rect -3500 2140 0 2150
rect -3500 2110 -3490 2140
rect -3460 2110 -3290 2140
rect -3260 2110 -3090 2140
rect -3060 2110 -1590 2140
rect -1560 2110 -1090 2140
rect -1060 2110 -890 2140
rect -860 2110 -690 2140
rect -660 2110 -490 2140
rect -460 2110 -290 2140
rect -260 2110 -90 2140
rect -60 2110 0 2140
rect -3500 2090 0 2110
rect -3500 2060 -3490 2090
rect -3460 2060 -3290 2090
rect -3260 2060 -3090 2090
rect -3060 2060 -1590 2090
rect -1560 2060 -1090 2090
rect -1060 2060 -890 2090
rect -860 2060 -690 2090
rect -660 2060 -490 2090
rect -460 2060 -290 2090
rect -260 2060 -90 2090
rect -60 2060 0 2090
rect -3500 2040 0 2060
rect -3500 2010 -3490 2040
rect -3460 2010 -3290 2040
rect -3260 2010 -3090 2040
rect -3060 2010 -1590 2040
rect -1560 2010 -1090 2040
rect -1060 2010 -890 2040
rect -860 2010 -690 2040
rect -660 2010 -490 2040
rect -460 2010 -290 2040
rect -260 2010 -90 2040
rect -60 2010 0 2040
rect -3500 2000 0 2010
rect -3500 440 0 450
rect -3500 410 -3490 440
rect -3460 410 -3290 440
rect -3260 410 -3090 440
rect -3060 410 -1590 440
rect -1560 410 -1090 440
rect -1060 410 -890 440
rect -860 410 -690 440
rect -660 410 -490 440
rect -460 410 -290 440
rect -260 410 -90 440
rect -60 410 0 440
rect -3500 390 0 410
rect -3500 360 -3490 390
rect -3460 360 -3290 390
rect -3260 360 -3090 390
rect -3060 360 -1590 390
rect -1560 360 -1090 390
rect -1060 360 -890 390
rect -860 360 -690 390
rect -660 360 -490 390
rect -460 360 -290 390
rect -260 360 -90 390
rect -60 360 0 390
rect -3500 340 0 360
rect -3500 310 -3490 340
rect -3460 310 -3290 340
rect -3260 310 -3090 340
rect -3060 310 -1590 340
rect -1560 310 -1090 340
rect -1060 310 -890 340
rect -860 310 -690 340
rect -660 310 -490 340
rect -460 310 -290 340
rect -260 310 -90 340
rect -60 310 0 340
rect -3500 300 0 310
<< via2 >>
rect -3490 16980 -3460 17010
rect -3290 16980 -3260 17010
rect -3090 16980 -3060 17010
rect -1590 16980 -1560 17010
rect -1190 16980 -1160 17010
rect -1090 16980 -1060 17010
rect -990 16980 -960 17010
rect -890 16980 -860 17010
rect -790 16980 -760 17010
rect -690 16980 -660 17010
rect -590 16980 -560 17010
rect -490 16980 -460 17010
rect -390 16980 -360 17010
rect -290 16980 -260 17010
rect -190 16980 -160 17010
rect -90 16980 -60 17010
rect -3490 15710 -3460 15740
rect -3290 15710 -3260 15740
rect -3090 15710 -3060 15740
rect -1590 15710 -1560 15740
rect -1190 15710 -1160 15740
rect -1090 15710 -1060 15740
rect -990 15710 -960 15740
rect -890 15710 -860 15740
rect -690 15710 -660 15740
rect -590 15710 -560 15740
rect -490 15710 -460 15740
rect -290 15710 -260 15740
rect -190 15710 -160 15740
rect -90 15710 -60 15740
rect -3490 15310 -3460 15340
rect -3290 15310 -3260 15340
rect -3090 15310 -3060 15340
rect -1590 15310 -1560 15340
rect -1090 15310 -1060 15340
rect -890 15310 -860 15340
rect -690 15310 -660 15340
rect -490 15310 -460 15340
rect -290 15310 -260 15340
rect -90 15310 -60 15340
rect -3490 15260 -3460 15290
rect -3290 15260 -3260 15290
rect -3090 15260 -3060 15290
rect -1590 15260 -1560 15290
rect -1090 15260 -1060 15290
rect -890 15260 -860 15290
rect -690 15260 -660 15290
rect -490 15260 -460 15290
rect -290 15260 -260 15290
rect -90 15260 -60 15290
rect -3490 15210 -3460 15240
rect -3290 15210 -3260 15240
rect -3090 15210 -3060 15240
rect -1590 15210 -1560 15240
rect -1090 15210 -1060 15240
rect -890 15210 -860 15240
rect -690 15210 -660 15240
rect -490 15210 -460 15240
rect -290 15210 -260 15240
rect -90 15210 -60 15240
rect -3490 13610 -3460 13640
rect -3290 13610 -3260 13640
rect -3090 13610 -3060 13640
rect -1590 13610 -1560 13640
rect -1090 13610 -1060 13640
rect -890 13610 -860 13640
rect -690 13610 -660 13640
rect -490 13610 -460 13640
rect -290 13610 -260 13640
rect -90 13610 -60 13640
rect -3490 13560 -3460 13590
rect -3290 13560 -3260 13590
rect -3090 13560 -3060 13590
rect -1590 13560 -1560 13590
rect -1090 13560 -1060 13590
rect -890 13560 -860 13590
rect -690 13560 -660 13590
rect -490 13560 -460 13590
rect -290 13560 -260 13590
rect -90 13560 -60 13590
rect -3490 13510 -3460 13540
rect -3290 13510 -3260 13540
rect -3090 13510 -3060 13540
rect -1590 13510 -1560 13540
rect -1090 13510 -1060 13540
rect -890 13510 -860 13540
rect -690 13510 -660 13540
rect -490 13510 -460 13540
rect -290 13510 -260 13540
rect -90 13510 -60 13540
rect -3490 11910 -3460 11940
rect -3290 11910 -3260 11940
rect -3090 11910 -3060 11940
rect -1590 11910 -1560 11940
rect -1090 11910 -1060 11940
rect -890 11910 -860 11940
rect -690 11910 -660 11940
rect -490 11910 -460 11940
rect -290 11910 -260 11940
rect -90 11910 -60 11940
rect -3490 11860 -3460 11890
rect -3290 11860 -3260 11890
rect -3090 11860 -3060 11890
rect -1590 11860 -1560 11890
rect -1090 11860 -1060 11890
rect -890 11860 -860 11890
rect -690 11860 -660 11890
rect -490 11860 -460 11890
rect -290 11860 -260 11890
rect -90 11860 -60 11890
rect -3490 11810 -3460 11840
rect -3290 11810 -3260 11840
rect -3090 11810 -3060 11840
rect -1590 11810 -1560 11840
rect -1090 11810 -1060 11840
rect -890 11810 -860 11840
rect -690 11810 -660 11840
rect -490 11810 -460 11840
rect -290 11810 -260 11840
rect -90 11810 -60 11840
rect 39810 11310 39840 11340
rect 39910 11210 39940 11240
rect 39960 11210 39990 11240
rect 40010 11210 40040 11240
rect 40060 11210 40090 11240
rect 40110 11210 40140 11240
rect 40160 11210 40190 11240
rect 40210 11210 40240 11240
rect 40260 11210 40290 11240
rect 40310 11210 40340 11240
rect 40360 11210 40390 11240
rect 40410 11210 40440 11240
rect 40460 11210 40490 11240
rect 40510 11210 40540 11240
rect 40560 11210 40590 11240
rect 40610 11210 40640 11240
rect 40660 11210 40690 11240
rect 40710 11210 40740 11240
rect 40760 11210 40790 11240
rect 40810 11210 40840 11240
rect 40860 11210 40890 11240
rect 39910 11160 39940 11190
rect 39960 11160 39990 11190
rect 40010 11160 40040 11190
rect 40060 11160 40090 11190
rect 40110 11160 40140 11190
rect 40160 11160 40190 11190
rect 40210 11160 40240 11190
rect 40260 11160 40290 11190
rect 40310 11160 40340 11190
rect 40360 11160 40390 11190
rect 40410 11160 40440 11190
rect 40460 11160 40490 11190
rect 40510 11160 40540 11190
rect 40560 11160 40590 11190
rect 40610 11160 40640 11190
rect 40660 11160 40690 11190
rect 40710 11160 40740 11190
rect 40760 11160 40790 11190
rect 40810 11160 40840 11190
rect 40860 11160 40890 11190
rect 39910 11110 39940 11140
rect 39960 11110 39990 11140
rect 40010 11110 40040 11140
rect 40060 11110 40090 11140
rect 40110 11110 40140 11140
rect 40160 11110 40190 11140
rect 40210 11110 40240 11140
rect 40260 11110 40290 11140
rect 40310 11110 40340 11140
rect 40360 11110 40390 11140
rect 40410 11110 40440 11140
rect 40460 11110 40490 11140
rect 40510 11110 40540 11140
rect 40560 11110 40590 11140
rect 40610 11110 40640 11140
rect 40660 11110 40690 11140
rect 40710 11110 40740 11140
rect 40760 11110 40790 11140
rect 40810 11110 40840 11140
rect 40860 11110 40890 11140
rect 39910 11060 39940 11090
rect 39960 11060 39990 11090
rect 40010 11060 40040 11090
rect 40060 11060 40090 11090
rect 40110 11060 40140 11090
rect 40160 11060 40190 11090
rect 40210 11060 40240 11090
rect 40260 11060 40290 11090
rect 40310 11060 40340 11090
rect 40360 11060 40390 11090
rect 40410 11060 40440 11090
rect 40460 11060 40490 11090
rect 40510 11060 40540 11090
rect 40560 11060 40590 11090
rect 40610 11060 40640 11090
rect 40660 11060 40690 11090
rect 40710 11060 40740 11090
rect 40760 11060 40790 11090
rect 40810 11060 40840 11090
rect 40860 11060 40890 11090
rect 39910 11010 39940 11040
rect 39960 11010 39990 11040
rect 40010 11010 40040 11040
rect 40060 11010 40090 11040
rect 40110 11010 40140 11040
rect 40160 11010 40190 11040
rect 40210 11010 40240 11040
rect 40260 11010 40290 11040
rect 40310 11010 40340 11040
rect 40360 11010 40390 11040
rect 40410 11010 40440 11040
rect 40460 11010 40490 11040
rect 40510 11010 40540 11040
rect 40560 11010 40590 11040
rect 40610 11010 40640 11040
rect 40660 11010 40690 11040
rect 40710 11010 40740 11040
rect 40760 11010 40790 11040
rect 40810 11010 40840 11040
rect 40860 11010 40890 11040
rect 39810 10910 39840 10940
rect -2990 10610 -2960 10640
rect -2790 10610 -2760 10640
rect -2590 10610 -2560 10640
rect -2390 10610 -2360 10640
rect -2190 10610 -2160 10640
rect -1990 10610 -1960 10640
rect -1690 10610 -1660 10640
rect -2990 10560 -2960 10590
rect -2790 10560 -2760 10590
rect -2590 10560 -2560 10590
rect -2390 10560 -2360 10590
rect -2190 10560 -2160 10590
rect -1990 10560 -1960 10590
rect -1690 10560 -1660 10590
rect -2990 10510 -2960 10540
rect -2790 10510 -2760 10540
rect -2590 10510 -2560 10540
rect -2390 10510 -2360 10540
rect -2190 10510 -2160 10540
rect -1990 10510 -1960 10540
rect -1690 10510 -1660 10540
rect -2990 9310 -2960 9340
rect -2790 9310 -2760 9340
rect -2590 9310 -2560 9340
rect -2390 9310 -2360 9340
rect -2190 9310 -2160 9340
rect -1990 9310 -1960 9340
rect -1690 9310 -1660 9340
rect -2990 9260 -2960 9290
rect -2790 9260 -2760 9290
rect -2590 9260 -2560 9290
rect -2390 9260 -2360 9290
rect -2190 9260 -2160 9290
rect -1990 9260 -1960 9290
rect -1690 9260 -1660 9290
rect -2990 9210 -2960 9240
rect -2790 9210 -2760 9240
rect -2590 9210 -2560 9240
rect -2390 9210 -2360 9240
rect -2190 9210 -2160 9240
rect -1990 9210 -1960 9240
rect -1690 9210 -1660 9240
rect -2990 8010 -2960 8040
rect -2790 8010 -2760 8040
rect -2590 8010 -2560 8040
rect -2390 8010 -2360 8040
rect -2190 8010 -2160 8040
rect -1990 8010 -1960 8040
rect -1690 8010 -1660 8040
rect -2990 7960 -2960 7990
rect -2790 7960 -2760 7990
rect -2590 7960 -2560 7990
rect -2390 7960 -2360 7990
rect -2190 7960 -2160 7990
rect -1990 7960 -1960 7990
rect -1690 7960 -1660 7990
rect -2990 7910 -2960 7940
rect -2790 7910 -2760 7940
rect -2590 7910 -2560 7940
rect -2390 7910 -2360 7940
rect -2190 7910 -2160 7940
rect -1990 7910 -1960 7940
rect -1690 7910 -1660 7940
rect -2990 7710 -2960 7740
rect -2790 7710 -2760 7740
rect -2590 7710 -2560 7740
rect -2390 7710 -2360 7740
rect -2190 7710 -2160 7740
rect -1990 7710 -1960 7740
rect -1690 7710 -1660 7740
rect -2990 7660 -2960 7690
rect -2790 7660 -2760 7690
rect -2590 7660 -2560 7690
rect -2390 7660 -2360 7690
rect -2190 7660 -2160 7690
rect -1990 7660 -1960 7690
rect -1690 7660 -1660 7690
rect -2990 7610 -2960 7640
rect -2790 7610 -2760 7640
rect -2590 7610 -2560 7640
rect -2390 7610 -2360 7640
rect -2190 7610 -2160 7640
rect -1990 7610 -1960 7640
rect -1690 7610 -1660 7640
rect -2990 6410 -2960 6440
rect -2790 6410 -2760 6440
rect -2590 6410 -2560 6440
rect -2390 6410 -2360 6440
rect -2190 6410 -2160 6440
rect -1990 6410 -1960 6440
rect -1690 6410 -1660 6440
rect -2990 6360 -2960 6390
rect -2790 6360 -2760 6390
rect -2590 6360 -2560 6390
rect -2390 6360 -2360 6390
rect -2190 6360 -2160 6390
rect -1990 6360 -1960 6390
rect -1690 6360 -1660 6390
rect -2990 6310 -2960 6340
rect -2790 6310 -2760 6340
rect -2590 6310 -2560 6340
rect -2390 6310 -2360 6340
rect -2190 6310 -2160 6340
rect -1990 6310 -1960 6340
rect -1690 6310 -1660 6340
rect -2990 5110 -2960 5140
rect -2790 5110 -2760 5140
rect -2590 5110 -2560 5140
rect -2390 5110 -2360 5140
rect -2190 5110 -2160 5140
rect -1990 5110 -1960 5140
rect -1690 5110 -1660 5140
rect -2990 5060 -2960 5090
rect -2790 5060 -2760 5090
rect -2590 5060 -2560 5090
rect -2390 5060 -2360 5090
rect -2190 5060 -2160 5090
rect -1990 5060 -1960 5090
rect -1690 5060 -1660 5090
rect -2990 5010 -2960 5040
rect -2790 5010 -2760 5040
rect -2590 5010 -2560 5040
rect -2390 5010 -2360 5040
rect -2190 5010 -2160 5040
rect -1990 5010 -1960 5040
rect -1690 5010 -1660 5040
rect 39810 4710 39840 4740
rect 39910 4610 39940 4640
rect 39960 4610 39990 4640
rect 40010 4610 40040 4640
rect 40060 4610 40090 4640
rect 40110 4610 40140 4640
rect 40160 4610 40190 4640
rect 40210 4610 40240 4640
rect 40260 4610 40290 4640
rect 40310 4610 40340 4640
rect 40360 4610 40390 4640
rect 40410 4610 40440 4640
rect 40460 4610 40490 4640
rect 40510 4610 40540 4640
rect 40560 4610 40590 4640
rect 40610 4610 40640 4640
rect 40660 4610 40690 4640
rect 40710 4610 40740 4640
rect 40760 4610 40790 4640
rect 40810 4610 40840 4640
rect 40860 4610 40890 4640
rect 39910 4560 39940 4590
rect 39960 4560 39990 4590
rect 40010 4560 40040 4590
rect 40060 4560 40090 4590
rect 40110 4560 40140 4590
rect 40160 4560 40190 4590
rect 40210 4560 40240 4590
rect 40260 4560 40290 4590
rect 40310 4560 40340 4590
rect 40360 4560 40390 4590
rect 40410 4560 40440 4590
rect 40460 4560 40490 4590
rect 40510 4560 40540 4590
rect 40560 4560 40590 4590
rect 40610 4560 40640 4590
rect 40660 4560 40690 4590
rect 40710 4560 40740 4590
rect 40760 4560 40790 4590
rect 40810 4560 40840 4590
rect 40860 4560 40890 4590
rect 39910 4510 39940 4540
rect 39960 4510 39990 4540
rect 40010 4510 40040 4540
rect 40060 4510 40090 4540
rect 40110 4510 40140 4540
rect 40160 4510 40190 4540
rect 40210 4510 40240 4540
rect 40260 4510 40290 4540
rect 40310 4510 40340 4540
rect 40360 4510 40390 4540
rect 40410 4510 40440 4540
rect 40460 4510 40490 4540
rect 40510 4510 40540 4540
rect 40560 4510 40590 4540
rect 40610 4510 40640 4540
rect 40660 4510 40690 4540
rect 40710 4510 40740 4540
rect 40760 4510 40790 4540
rect 40810 4510 40840 4540
rect 40860 4510 40890 4540
rect 39910 4460 39940 4490
rect 39960 4460 39990 4490
rect 40010 4460 40040 4490
rect 40060 4460 40090 4490
rect 40110 4460 40140 4490
rect 40160 4460 40190 4490
rect 40210 4460 40240 4490
rect 40260 4460 40290 4490
rect 40310 4460 40340 4490
rect 40360 4460 40390 4490
rect 40410 4460 40440 4490
rect 40460 4460 40490 4490
rect 40510 4460 40540 4490
rect 40560 4460 40590 4490
rect 40610 4460 40640 4490
rect 40660 4460 40690 4490
rect 40710 4460 40740 4490
rect 40760 4460 40790 4490
rect 40810 4460 40840 4490
rect 40860 4460 40890 4490
rect 39910 4410 39940 4440
rect 39960 4410 39990 4440
rect 40010 4410 40040 4440
rect 40060 4410 40090 4440
rect 40110 4410 40140 4440
rect 40160 4410 40190 4440
rect 40210 4410 40240 4440
rect 40260 4410 40290 4440
rect 40310 4410 40340 4440
rect 40360 4410 40390 4440
rect 40410 4410 40440 4440
rect 40460 4410 40490 4440
rect 40510 4410 40540 4440
rect 40560 4410 40590 4440
rect 40610 4410 40640 4440
rect 40660 4410 40690 4440
rect 40710 4410 40740 4440
rect 40760 4410 40790 4440
rect 40810 4410 40840 4440
rect 40860 4410 40890 4440
rect 39810 4310 39840 4340
rect -3490 3810 -3460 3840
rect -3290 3810 -3260 3840
rect -3090 3810 -3060 3840
rect -1590 3810 -1560 3840
rect -1090 3810 -1060 3840
rect -890 3810 -860 3840
rect -690 3810 -660 3840
rect -490 3810 -460 3840
rect -290 3810 -260 3840
rect -90 3810 -60 3840
rect -3490 3760 -3460 3790
rect -3290 3760 -3260 3790
rect -3090 3760 -3060 3790
rect -1590 3760 -1560 3790
rect -1090 3760 -1060 3790
rect -890 3760 -860 3790
rect -690 3760 -660 3790
rect -490 3760 -460 3790
rect -290 3760 -260 3790
rect -90 3760 -60 3790
rect -3490 3710 -3460 3740
rect -3290 3710 -3260 3740
rect -3090 3710 -3060 3740
rect -1590 3710 -1560 3740
rect -1090 3710 -1060 3740
rect -890 3710 -860 3740
rect -690 3710 -660 3740
rect -490 3710 -460 3740
rect -290 3710 -260 3740
rect -90 3710 -60 3740
rect -3490 2110 -3460 2140
rect -3290 2110 -3260 2140
rect -3090 2110 -3060 2140
rect -1590 2110 -1560 2140
rect -1090 2110 -1060 2140
rect -890 2110 -860 2140
rect -690 2110 -660 2140
rect -490 2110 -460 2140
rect -290 2110 -260 2140
rect -90 2110 -60 2140
rect -3490 2060 -3460 2090
rect -3290 2060 -3260 2090
rect -3090 2060 -3060 2090
rect -1590 2060 -1560 2090
rect -1090 2060 -1060 2090
rect -890 2060 -860 2090
rect -690 2060 -660 2090
rect -490 2060 -460 2090
rect -290 2060 -260 2090
rect -90 2060 -60 2090
rect -3490 2010 -3460 2040
rect -3290 2010 -3260 2040
rect -3090 2010 -3060 2040
rect -1590 2010 -1560 2040
rect -1090 2010 -1060 2040
rect -890 2010 -860 2040
rect -690 2010 -660 2040
rect -490 2010 -460 2040
rect -290 2010 -260 2040
rect -90 2010 -60 2040
rect -3490 410 -3460 440
rect -3290 410 -3260 440
rect -3090 410 -3060 440
rect -1590 410 -1560 440
rect -1090 410 -1060 440
rect -890 410 -860 440
rect -690 410 -660 440
rect -490 410 -460 440
rect -290 410 -260 440
rect -90 410 -60 440
rect -3490 360 -3460 390
rect -3290 360 -3260 390
rect -3090 360 -3060 390
rect -1590 360 -1560 390
rect -1090 360 -1060 390
rect -890 360 -860 390
rect -690 360 -660 390
rect -490 360 -460 390
rect -290 360 -260 390
rect -90 360 -60 390
rect -3490 310 -3460 340
rect -3290 310 -3260 340
rect -3090 310 -3060 340
rect -1590 310 -1560 340
rect -1090 310 -1060 340
rect -890 310 -860 340
rect -690 310 -660 340
rect -490 310 -460 340
rect -290 310 -260 340
rect -90 310 -60 340
<< metal3 >>
rect 0 18285 40900 18290
rect 0 18245 5 18285
rect 45 18245 55 18285
rect 95 18245 105 18285
rect 145 18245 155 18285
rect 195 18245 205 18285
rect 245 18245 255 18285
rect 295 18245 305 18285
rect 345 18245 355 18285
rect 395 18245 405 18285
rect 445 18245 455 18285
rect 495 18245 505 18285
rect 545 18245 555 18285
rect 595 18245 605 18285
rect 645 18245 655 18285
rect 695 18245 705 18285
rect 745 18245 755 18285
rect 795 18245 805 18285
rect 845 18245 855 18285
rect 895 18245 905 18285
rect 945 18245 955 18285
rect 995 18245 1005 18285
rect 1045 18245 1055 18285
rect 1095 18245 1105 18285
rect 1145 18245 1155 18285
rect 1195 18245 1205 18285
rect 1245 18245 1255 18285
rect 1295 18245 1305 18285
rect 1345 18245 1355 18285
rect 1395 18245 1405 18285
rect 1445 18245 1455 18285
rect 1495 18245 1505 18285
rect 1545 18245 1555 18285
rect 1595 18245 1605 18285
rect 1645 18245 1655 18285
rect 1695 18245 1705 18285
rect 1745 18245 1755 18285
rect 1795 18245 1805 18285
rect 1845 18245 1855 18285
rect 1895 18245 1905 18285
rect 1945 18245 1955 18285
rect 1995 18245 2005 18285
rect 2045 18245 2055 18285
rect 2095 18245 2105 18285
rect 2145 18245 2155 18285
rect 2195 18245 2205 18285
rect 2245 18245 2255 18285
rect 2295 18245 2305 18285
rect 2345 18245 2355 18285
rect 2395 18245 2405 18285
rect 2445 18245 2455 18285
rect 2495 18245 2505 18285
rect 2545 18245 2555 18285
rect 2595 18245 2605 18285
rect 2645 18245 2655 18285
rect 2695 18245 2705 18285
rect 2745 18245 2755 18285
rect 2795 18245 2805 18285
rect 2845 18245 2855 18285
rect 2895 18245 2905 18285
rect 2945 18245 2955 18285
rect 2995 18245 3005 18285
rect 3045 18245 3055 18285
rect 3095 18245 3105 18285
rect 3145 18245 3155 18285
rect 3195 18245 3205 18285
rect 3245 18245 3255 18285
rect 3295 18245 3305 18285
rect 3345 18245 3355 18285
rect 3395 18245 3405 18285
rect 3445 18245 3455 18285
rect 3495 18245 3505 18285
rect 3545 18245 3555 18285
rect 3595 18245 3605 18285
rect 3645 18245 3655 18285
rect 3695 18245 3705 18285
rect 3745 18245 3755 18285
rect 3795 18245 3805 18285
rect 3845 18245 3855 18285
rect 3895 18245 3905 18285
rect 3945 18245 3955 18285
rect 3995 18245 4005 18285
rect 4045 18245 4055 18285
rect 4095 18245 4105 18285
rect 4145 18245 4155 18285
rect 4195 18245 4205 18285
rect 4245 18245 4255 18285
rect 4295 18245 4305 18285
rect 4345 18245 4355 18285
rect 4395 18245 4405 18285
rect 4445 18245 4455 18285
rect 4495 18245 4505 18285
rect 4545 18245 4555 18285
rect 4595 18245 4605 18285
rect 4645 18245 4655 18285
rect 4695 18245 4705 18285
rect 4745 18245 4755 18285
rect 4795 18245 4805 18285
rect 4845 18245 4855 18285
rect 4895 18245 4905 18285
rect 4945 18245 4955 18285
rect 4995 18245 5005 18285
rect 5045 18245 5055 18285
rect 5095 18245 5105 18285
rect 5145 18245 5155 18285
rect 5195 18245 5205 18285
rect 5245 18245 5255 18285
rect 5295 18245 5305 18285
rect 5345 18245 5355 18285
rect 5395 18245 5405 18285
rect 5445 18245 5455 18285
rect 5495 18245 5505 18285
rect 5545 18245 5555 18285
rect 5595 18245 5605 18285
rect 5645 18245 5655 18285
rect 5695 18245 5705 18285
rect 5745 18245 5755 18285
rect 5795 18245 5805 18285
rect 5845 18245 5855 18285
rect 5895 18245 5905 18285
rect 5945 18245 5955 18285
rect 5995 18245 6005 18285
rect 6045 18245 6055 18285
rect 6095 18245 6105 18285
rect 6145 18245 6155 18285
rect 6195 18245 6205 18285
rect 6245 18245 6255 18285
rect 6295 18245 6305 18285
rect 6345 18245 6355 18285
rect 6395 18245 6405 18285
rect 6445 18245 6455 18285
rect 6495 18245 6505 18285
rect 6545 18245 6555 18285
rect 6595 18245 6605 18285
rect 6645 18245 6655 18285
rect 6695 18245 6705 18285
rect 6745 18245 6755 18285
rect 6795 18245 6805 18285
rect 6845 18245 6855 18285
rect 6895 18245 6905 18285
rect 6945 18245 6955 18285
rect 6995 18245 7005 18285
rect 7045 18245 7055 18285
rect 7095 18245 7105 18285
rect 7145 18245 7155 18285
rect 7195 18245 7205 18285
rect 7245 18245 7255 18285
rect 7295 18245 7305 18285
rect 7345 18245 7355 18285
rect 7395 18245 7405 18285
rect 7445 18245 7455 18285
rect 7495 18245 7505 18285
rect 7545 18245 7555 18285
rect 7595 18245 7605 18285
rect 7645 18245 7655 18285
rect 7695 18245 7705 18285
rect 7745 18245 7755 18285
rect 7795 18245 7805 18285
rect 7845 18245 7855 18285
rect 7895 18245 7905 18285
rect 7945 18245 7955 18285
rect 7995 18245 8005 18285
rect 8045 18245 8055 18285
rect 8095 18245 8105 18285
rect 8145 18245 8155 18285
rect 8195 18245 8205 18285
rect 8245 18245 8255 18285
rect 8295 18245 8305 18285
rect 8345 18245 8355 18285
rect 8395 18245 8405 18285
rect 8445 18245 8455 18285
rect 8495 18245 8505 18285
rect 8545 18245 8555 18285
rect 8595 18245 8605 18285
rect 8645 18245 8655 18285
rect 8695 18245 8705 18285
rect 8745 18245 8755 18285
rect 8795 18245 8805 18285
rect 8845 18245 8855 18285
rect 8895 18245 8905 18285
rect 8945 18245 8955 18285
rect 8995 18245 9005 18285
rect 9045 18245 9055 18285
rect 9095 18245 9105 18285
rect 9145 18245 9155 18285
rect 9195 18245 9205 18285
rect 9245 18245 9255 18285
rect 9295 18245 9305 18285
rect 9345 18245 9355 18285
rect 9395 18245 9405 18285
rect 9445 18245 9455 18285
rect 9495 18245 9505 18285
rect 9545 18245 9555 18285
rect 9595 18245 9605 18285
rect 9645 18245 9655 18285
rect 9695 18245 9705 18285
rect 9745 18245 9755 18285
rect 9795 18245 9805 18285
rect 9845 18245 9855 18285
rect 9895 18245 9905 18285
rect 9945 18245 9955 18285
rect 9995 18245 10005 18285
rect 10045 18245 10055 18285
rect 10095 18245 10105 18285
rect 10145 18245 10155 18285
rect 10195 18245 10205 18285
rect 10245 18245 10255 18285
rect 10295 18245 10305 18285
rect 10345 18245 10355 18285
rect 10395 18245 10405 18285
rect 10445 18245 10455 18285
rect 10495 18245 10505 18285
rect 10545 18245 10555 18285
rect 10595 18245 10605 18285
rect 10645 18245 10655 18285
rect 10695 18245 10705 18285
rect 10745 18245 10755 18285
rect 10795 18245 10805 18285
rect 10845 18245 10855 18285
rect 10895 18245 10905 18285
rect 10945 18245 10955 18285
rect 10995 18245 11005 18285
rect 11045 18245 11055 18285
rect 11095 18245 11105 18285
rect 11145 18245 11155 18285
rect 11195 18245 11205 18285
rect 11245 18245 11255 18285
rect 11295 18245 11305 18285
rect 11345 18245 11355 18285
rect 11395 18245 11405 18285
rect 11445 18245 11455 18285
rect 11495 18245 11505 18285
rect 11545 18245 11555 18285
rect 11595 18245 11605 18285
rect 11645 18245 11655 18285
rect 11695 18245 11705 18285
rect 11745 18245 11755 18285
rect 11795 18245 11805 18285
rect 11845 18245 11855 18285
rect 11895 18245 11905 18285
rect 11945 18245 11955 18285
rect 11995 18245 12005 18285
rect 12045 18245 12055 18285
rect 12095 18245 12105 18285
rect 12145 18245 12155 18285
rect 12195 18245 12205 18285
rect 12245 18245 12255 18285
rect 12295 18245 12305 18285
rect 12345 18245 12355 18285
rect 12395 18245 12405 18285
rect 12445 18245 12455 18285
rect 12495 18245 12505 18285
rect 12545 18245 12555 18285
rect 12595 18245 12605 18285
rect 12645 18245 12655 18285
rect 12695 18245 12705 18285
rect 12745 18245 12755 18285
rect 12795 18245 12805 18285
rect 12845 18245 12855 18285
rect 12895 18245 12905 18285
rect 12945 18245 12955 18285
rect 12995 18245 13005 18285
rect 13045 18245 13055 18285
rect 13095 18245 13105 18285
rect 13145 18245 13155 18285
rect 13195 18245 13205 18285
rect 13245 18245 13255 18285
rect 13295 18245 13305 18285
rect 13345 18245 13355 18285
rect 13395 18245 13405 18285
rect 13445 18245 13455 18285
rect 13495 18245 13505 18285
rect 13545 18245 13555 18285
rect 13595 18245 13605 18285
rect 13645 18245 13655 18285
rect 13695 18245 13705 18285
rect 13745 18245 13755 18285
rect 13795 18245 13805 18285
rect 13845 18245 13855 18285
rect 13895 18245 13905 18285
rect 13945 18245 13955 18285
rect 13995 18245 14005 18285
rect 14045 18245 14055 18285
rect 14095 18245 14105 18285
rect 14145 18245 14155 18285
rect 14195 18245 14205 18285
rect 14245 18245 14255 18285
rect 14295 18245 14305 18285
rect 14345 18245 14355 18285
rect 14395 18245 14405 18285
rect 14445 18245 14455 18285
rect 14495 18245 14505 18285
rect 14545 18245 14555 18285
rect 14595 18245 14605 18285
rect 14645 18245 14655 18285
rect 14695 18245 14705 18285
rect 14745 18245 14755 18285
rect 14795 18245 14805 18285
rect 14845 18245 14855 18285
rect 14895 18245 14905 18285
rect 14945 18245 14955 18285
rect 14995 18245 15005 18285
rect 15045 18245 15055 18285
rect 15095 18245 15105 18285
rect 15145 18245 15155 18285
rect 15195 18245 15205 18285
rect 15245 18245 15255 18285
rect 15295 18245 15305 18285
rect 15345 18245 15355 18285
rect 15395 18245 15405 18285
rect 15445 18245 15455 18285
rect 15495 18245 15505 18285
rect 15545 18245 15555 18285
rect 15595 18245 15605 18285
rect 15645 18245 15655 18285
rect 15695 18245 15705 18285
rect 15745 18245 15755 18285
rect 15795 18245 15805 18285
rect 15845 18245 15855 18285
rect 15895 18245 15905 18285
rect 15945 18245 15955 18285
rect 15995 18245 16005 18285
rect 16045 18245 16055 18285
rect 16095 18245 16105 18285
rect 16145 18245 16155 18285
rect 16195 18245 16205 18285
rect 16245 18245 16255 18285
rect 16295 18245 16305 18285
rect 16345 18245 16355 18285
rect 16395 18245 16405 18285
rect 16445 18245 16455 18285
rect 16495 18245 16505 18285
rect 16545 18245 16555 18285
rect 16595 18245 16605 18285
rect 16645 18245 16655 18285
rect 16695 18245 16705 18285
rect 16745 18245 16755 18285
rect 16795 18245 16805 18285
rect 16845 18245 16855 18285
rect 16895 18245 16905 18285
rect 16945 18245 16955 18285
rect 16995 18245 17005 18285
rect 17045 18245 17055 18285
rect 17095 18245 17105 18285
rect 17145 18245 17155 18285
rect 17195 18245 17205 18285
rect 17245 18245 17255 18285
rect 17295 18245 17305 18285
rect 17345 18245 17355 18285
rect 17395 18245 17405 18285
rect 17445 18245 17455 18285
rect 17495 18245 17505 18285
rect 17545 18245 17555 18285
rect 17595 18245 17605 18285
rect 17645 18245 17655 18285
rect 17695 18245 17705 18285
rect 17745 18245 17755 18285
rect 17795 18245 17805 18285
rect 17845 18245 17855 18285
rect 17895 18245 17905 18285
rect 17945 18245 17955 18285
rect 17995 18245 18005 18285
rect 18045 18245 18055 18285
rect 18095 18245 18105 18285
rect 18145 18245 18155 18285
rect 18195 18245 18205 18285
rect 18245 18245 18255 18285
rect 18295 18245 18305 18285
rect 18345 18245 18355 18285
rect 18395 18245 18405 18285
rect 18445 18245 18455 18285
rect 18495 18245 18505 18285
rect 18545 18245 18555 18285
rect 18595 18245 18605 18285
rect 18645 18245 18655 18285
rect 18695 18245 18705 18285
rect 18745 18245 18755 18285
rect 18795 18245 18805 18285
rect 18845 18245 18855 18285
rect 18895 18245 18905 18285
rect 18945 18245 18955 18285
rect 18995 18245 19005 18285
rect 19045 18245 19055 18285
rect 19095 18245 19105 18285
rect 19145 18245 19155 18285
rect 19195 18245 19205 18285
rect 19245 18245 19255 18285
rect 19295 18245 19305 18285
rect 19345 18245 19355 18285
rect 19395 18245 19405 18285
rect 19445 18245 19455 18285
rect 19495 18245 19505 18285
rect 19545 18245 19555 18285
rect 19595 18245 19605 18285
rect 19645 18245 19655 18285
rect 19695 18245 19705 18285
rect 19745 18245 19755 18285
rect 19795 18245 19805 18285
rect 19845 18245 19855 18285
rect 19895 18245 19905 18285
rect 19945 18245 19955 18285
rect 19995 18245 20005 18285
rect 20045 18245 20055 18285
rect 20095 18245 20105 18285
rect 20145 18245 20155 18285
rect 20195 18245 20205 18285
rect 20245 18245 20255 18285
rect 20295 18245 20305 18285
rect 20345 18245 20355 18285
rect 20395 18245 20405 18285
rect 20445 18245 20455 18285
rect 20495 18245 20505 18285
rect 20545 18245 20555 18285
rect 20595 18245 20605 18285
rect 20645 18245 20655 18285
rect 20695 18245 20705 18285
rect 20745 18245 20755 18285
rect 20795 18245 20805 18285
rect 20845 18245 20855 18285
rect 20895 18245 20905 18285
rect 20945 18245 20955 18285
rect 20995 18245 21005 18285
rect 21045 18245 21055 18285
rect 21095 18245 21105 18285
rect 21145 18245 21155 18285
rect 21195 18245 21205 18285
rect 21245 18245 21255 18285
rect 21295 18245 21305 18285
rect 21345 18245 21355 18285
rect 21395 18245 21405 18285
rect 21445 18245 21455 18285
rect 21495 18245 21505 18285
rect 21545 18245 21555 18285
rect 21595 18245 21605 18285
rect 21645 18245 21655 18285
rect 21695 18245 21705 18285
rect 21745 18245 21755 18285
rect 21795 18245 21805 18285
rect 21845 18245 21855 18285
rect 21895 18245 21905 18285
rect 21945 18245 21955 18285
rect 21995 18245 22005 18285
rect 22045 18245 22055 18285
rect 22095 18245 22105 18285
rect 22145 18245 22155 18285
rect 22195 18245 22205 18285
rect 22245 18245 22255 18285
rect 22295 18245 22305 18285
rect 22345 18245 22355 18285
rect 22395 18245 22405 18285
rect 22445 18245 22455 18285
rect 22495 18245 22505 18285
rect 22545 18245 22555 18285
rect 22595 18245 22605 18285
rect 22645 18245 22655 18285
rect 22695 18245 22705 18285
rect 22745 18245 22755 18285
rect 22795 18245 22805 18285
rect 22845 18245 22855 18285
rect 22895 18245 22905 18285
rect 22945 18245 22955 18285
rect 22995 18245 23005 18285
rect 23045 18245 23055 18285
rect 23095 18245 23105 18285
rect 23145 18245 23155 18285
rect 23195 18245 23205 18285
rect 23245 18245 23255 18285
rect 23295 18245 23305 18285
rect 23345 18245 23355 18285
rect 23395 18245 23405 18285
rect 23445 18245 23455 18285
rect 23495 18245 23505 18285
rect 23545 18245 23555 18285
rect 23595 18245 23605 18285
rect 23645 18245 23655 18285
rect 23695 18245 23705 18285
rect 23745 18245 23755 18285
rect 23795 18245 23805 18285
rect 23845 18245 23855 18285
rect 23895 18245 23905 18285
rect 23945 18245 23955 18285
rect 23995 18245 24005 18285
rect 24045 18245 24055 18285
rect 24095 18245 24105 18285
rect 24145 18245 24155 18285
rect 24195 18245 24205 18285
rect 24245 18245 24255 18285
rect 24295 18245 24305 18285
rect 24345 18245 24355 18285
rect 24395 18245 24405 18285
rect 24445 18245 24455 18285
rect 24495 18245 24505 18285
rect 24545 18245 24555 18285
rect 24595 18245 24605 18285
rect 24645 18245 24655 18285
rect 24695 18245 24705 18285
rect 24745 18245 24755 18285
rect 24795 18245 24805 18285
rect 24845 18245 24855 18285
rect 24895 18245 24905 18285
rect 24945 18245 24955 18285
rect 24995 18245 25005 18285
rect 25045 18245 25055 18285
rect 25095 18245 25105 18285
rect 25145 18245 25155 18285
rect 25195 18245 25205 18285
rect 25245 18245 25255 18285
rect 25295 18245 25305 18285
rect 25345 18245 25355 18285
rect 25395 18245 25405 18285
rect 25445 18245 25455 18285
rect 25495 18245 25505 18285
rect 25545 18245 25555 18285
rect 25595 18245 25605 18285
rect 25645 18245 25655 18285
rect 25695 18245 25705 18285
rect 25745 18245 25755 18285
rect 25795 18245 25805 18285
rect 25845 18245 25855 18285
rect 25895 18245 25905 18285
rect 25945 18245 25955 18285
rect 25995 18245 26005 18285
rect 26045 18245 26055 18285
rect 26095 18245 26105 18285
rect 26145 18245 26155 18285
rect 26195 18245 26205 18285
rect 26245 18245 26255 18285
rect 26295 18245 26305 18285
rect 26345 18245 26355 18285
rect 26395 18245 26405 18285
rect 26445 18245 26455 18285
rect 26495 18245 26505 18285
rect 26545 18245 26555 18285
rect 26595 18245 26605 18285
rect 26645 18245 26655 18285
rect 26695 18245 26705 18285
rect 26745 18245 26755 18285
rect 26795 18245 26805 18285
rect 26845 18245 26855 18285
rect 26895 18245 26905 18285
rect 26945 18245 26955 18285
rect 26995 18245 27005 18285
rect 27045 18245 27055 18285
rect 27095 18245 27105 18285
rect 27145 18245 27155 18285
rect 27195 18245 27205 18285
rect 27245 18245 27255 18285
rect 27295 18245 27305 18285
rect 27345 18245 27355 18285
rect 27395 18245 27405 18285
rect 27445 18245 27455 18285
rect 27495 18245 27505 18285
rect 27545 18245 27555 18285
rect 27595 18245 27605 18285
rect 27645 18245 27655 18285
rect 27695 18245 27705 18285
rect 27745 18245 27755 18285
rect 27795 18245 27805 18285
rect 27845 18245 27855 18285
rect 27895 18245 27905 18285
rect 27945 18245 27955 18285
rect 27995 18245 28005 18285
rect 28045 18245 28055 18285
rect 28095 18245 28105 18285
rect 28145 18245 28155 18285
rect 28195 18245 28205 18285
rect 28245 18245 28255 18285
rect 28295 18245 28305 18285
rect 28345 18245 28355 18285
rect 28395 18245 28405 18285
rect 28445 18245 28455 18285
rect 28495 18245 28505 18285
rect 28545 18245 28555 18285
rect 28595 18245 28605 18285
rect 28645 18245 28655 18285
rect 28695 18245 28705 18285
rect 28745 18245 28755 18285
rect 28795 18245 28805 18285
rect 28845 18245 28855 18285
rect 28895 18245 28905 18285
rect 28945 18245 28955 18285
rect 28995 18245 29005 18285
rect 29045 18245 29055 18285
rect 29095 18245 29105 18285
rect 29145 18245 29155 18285
rect 29195 18245 29205 18285
rect 29245 18245 29255 18285
rect 29295 18245 29305 18285
rect 29345 18245 29355 18285
rect 29395 18245 29405 18285
rect 29445 18245 29455 18285
rect 29495 18245 29505 18285
rect 29545 18245 29555 18285
rect 29595 18245 29605 18285
rect 29645 18245 29655 18285
rect 29695 18245 29705 18285
rect 29745 18245 29755 18285
rect 29795 18245 29805 18285
rect 29845 18245 29855 18285
rect 29895 18245 29905 18285
rect 29945 18245 29955 18285
rect 29995 18245 30005 18285
rect 30045 18245 30055 18285
rect 30095 18245 30105 18285
rect 30145 18245 30155 18285
rect 30195 18245 30205 18285
rect 30245 18245 30255 18285
rect 30295 18245 30305 18285
rect 30345 18245 30355 18285
rect 30395 18245 30405 18285
rect 30445 18245 30455 18285
rect 30495 18245 30505 18285
rect 30545 18245 30555 18285
rect 30595 18245 30605 18285
rect 30645 18245 30655 18285
rect 30695 18245 30705 18285
rect 30745 18245 30755 18285
rect 30795 18245 30805 18285
rect 30845 18245 30855 18285
rect 30895 18245 30905 18285
rect 30945 18245 30955 18285
rect 30995 18245 31005 18285
rect 31045 18245 31055 18285
rect 31095 18245 31105 18285
rect 31145 18245 31155 18285
rect 31195 18245 31205 18285
rect 31245 18245 31255 18285
rect 31295 18245 31305 18285
rect 31345 18245 31355 18285
rect 31395 18245 31405 18285
rect 31445 18245 31455 18285
rect 31495 18245 31505 18285
rect 31545 18245 31555 18285
rect 31595 18245 31605 18285
rect 31645 18245 31655 18285
rect 31695 18245 31705 18285
rect 31745 18245 31755 18285
rect 31795 18245 31805 18285
rect 31845 18245 31855 18285
rect 31895 18245 31905 18285
rect 31945 18245 31955 18285
rect 31995 18245 32005 18285
rect 32045 18245 32055 18285
rect 32095 18245 32105 18285
rect 32145 18245 32155 18285
rect 32195 18245 32205 18285
rect 32245 18245 32255 18285
rect 32295 18245 32305 18285
rect 32345 18245 32355 18285
rect 32395 18245 32405 18285
rect 32445 18245 32455 18285
rect 32495 18245 32505 18285
rect 32545 18245 32555 18285
rect 32595 18245 32605 18285
rect 32645 18245 32655 18285
rect 32695 18245 32705 18285
rect 32745 18245 32755 18285
rect 32795 18245 32805 18285
rect 32845 18245 32855 18285
rect 32895 18245 32905 18285
rect 32945 18245 32955 18285
rect 32995 18245 33005 18285
rect 33045 18245 33055 18285
rect 33095 18245 33105 18285
rect 33145 18245 33155 18285
rect 33195 18245 33205 18285
rect 33245 18245 33255 18285
rect 33295 18245 33305 18285
rect 33345 18245 33355 18285
rect 33395 18245 33405 18285
rect 33445 18245 33455 18285
rect 33495 18245 33505 18285
rect 33545 18245 33555 18285
rect 33595 18245 33605 18285
rect 33645 18245 33655 18285
rect 33695 18245 33705 18285
rect 33745 18245 33755 18285
rect 33795 18245 33805 18285
rect 33845 18245 33855 18285
rect 33895 18245 33905 18285
rect 33945 18245 33955 18285
rect 33995 18245 34005 18285
rect 34045 18245 34055 18285
rect 34095 18245 34105 18285
rect 34145 18245 34155 18285
rect 34195 18245 34205 18285
rect 34245 18245 34255 18285
rect 34295 18245 34305 18285
rect 34345 18245 34355 18285
rect 34395 18245 34405 18285
rect 34445 18245 34455 18285
rect 34495 18245 34505 18285
rect 34545 18245 34555 18285
rect 34595 18245 34605 18285
rect 34645 18245 34655 18285
rect 34695 18245 34705 18285
rect 34745 18245 34755 18285
rect 34795 18245 34805 18285
rect 34845 18245 34855 18285
rect 34895 18245 34905 18285
rect 34945 18245 34955 18285
rect 34995 18245 35005 18285
rect 35045 18245 35055 18285
rect 35095 18245 35105 18285
rect 35145 18245 35155 18285
rect 35195 18245 35205 18285
rect 35245 18245 35255 18285
rect 35295 18245 35305 18285
rect 35345 18245 35355 18285
rect 35395 18245 35405 18285
rect 35445 18245 35455 18285
rect 35495 18245 35505 18285
rect 35545 18245 35555 18285
rect 35595 18245 35605 18285
rect 35645 18245 35655 18285
rect 35695 18245 35705 18285
rect 35745 18245 35755 18285
rect 35795 18245 35805 18285
rect 35845 18245 35855 18285
rect 35895 18245 35905 18285
rect 35945 18245 35955 18285
rect 35995 18245 36005 18285
rect 36045 18245 36055 18285
rect 36095 18245 36105 18285
rect 36145 18245 36155 18285
rect 36195 18245 36205 18285
rect 36245 18245 36255 18285
rect 36295 18245 36305 18285
rect 36345 18245 36355 18285
rect 36395 18245 36405 18285
rect 36445 18245 36455 18285
rect 36495 18245 36505 18285
rect 36545 18245 36555 18285
rect 36595 18245 36605 18285
rect 36645 18245 36655 18285
rect 36695 18245 36705 18285
rect 36745 18245 36755 18285
rect 36795 18245 36805 18285
rect 36845 18245 36855 18285
rect 36895 18245 36905 18285
rect 36945 18245 36955 18285
rect 36995 18245 37005 18285
rect 37045 18245 37055 18285
rect 37095 18245 37105 18285
rect 37145 18245 37155 18285
rect 37195 18245 37205 18285
rect 37245 18245 37255 18285
rect 37295 18245 37305 18285
rect 37345 18245 37355 18285
rect 37395 18245 37405 18285
rect 37445 18245 37455 18285
rect 37495 18245 37505 18285
rect 37545 18245 37555 18285
rect 37595 18245 37605 18285
rect 37645 18245 37655 18285
rect 37695 18245 37705 18285
rect 37745 18245 37755 18285
rect 37795 18245 37805 18285
rect 37845 18245 37855 18285
rect 37895 18245 37905 18285
rect 37945 18245 37955 18285
rect 37995 18245 38005 18285
rect 38045 18245 38055 18285
rect 38095 18245 38105 18285
rect 38145 18245 38155 18285
rect 38195 18245 38205 18285
rect 38245 18245 38255 18285
rect 38295 18245 38305 18285
rect 38345 18245 38355 18285
rect 38395 18245 38405 18285
rect 38445 18245 38455 18285
rect 38495 18245 38505 18285
rect 38545 18245 38555 18285
rect 38595 18245 38605 18285
rect 38645 18245 38655 18285
rect 38695 18245 38705 18285
rect 38745 18245 38755 18285
rect 38795 18245 38805 18285
rect 38845 18245 38855 18285
rect 38895 18245 38905 18285
rect 38945 18245 38955 18285
rect 38995 18245 39005 18285
rect 39045 18245 39055 18285
rect 39095 18245 39105 18285
rect 39145 18245 39155 18285
rect 39195 18245 39205 18285
rect 39245 18245 39255 18285
rect 39295 18245 39305 18285
rect 39345 18245 39355 18285
rect 39395 18245 39405 18285
rect 39445 18245 39455 18285
rect 39495 18245 39505 18285
rect 39545 18245 39555 18285
rect 39595 18245 39605 18285
rect 39645 18245 39655 18285
rect 39695 18245 39705 18285
rect 39745 18245 39905 18285
rect 39945 18245 39955 18285
rect 39995 18245 40005 18285
rect 40045 18245 40055 18285
rect 40095 18245 40105 18285
rect 40145 18245 40155 18285
rect 40195 18245 40205 18285
rect 40245 18245 40255 18285
rect 40295 18245 40305 18285
rect 40345 18245 40355 18285
rect 40395 18245 40405 18285
rect 40445 18245 40455 18285
rect 40495 18245 40505 18285
rect 40545 18245 40555 18285
rect 40595 18245 40605 18285
rect 40645 18245 40655 18285
rect 40695 18245 40705 18285
rect 40745 18245 40755 18285
rect 40795 18245 40805 18285
rect 40845 18245 40855 18285
rect 40895 18245 40900 18285
rect 0 18240 40900 18245
rect 0 18185 39750 18190
rect 0 18145 5 18185
rect 45 18145 55 18185
rect 95 18145 105 18185
rect 145 18145 155 18185
rect 195 18145 205 18185
rect 245 18145 255 18185
rect 295 18145 305 18185
rect 345 18145 355 18185
rect 395 18145 405 18185
rect 445 18145 455 18185
rect 495 18145 505 18185
rect 545 18145 555 18185
rect 595 18145 605 18185
rect 645 18145 655 18185
rect 695 18145 705 18185
rect 745 18145 755 18185
rect 795 18145 805 18185
rect 845 18145 855 18185
rect 895 18145 905 18185
rect 945 18145 955 18185
rect 995 18145 1005 18185
rect 1045 18145 1055 18185
rect 1095 18145 1105 18185
rect 1145 18145 1155 18185
rect 1195 18145 1205 18185
rect 1245 18145 1255 18185
rect 1295 18145 1305 18185
rect 1345 18145 1355 18185
rect 1395 18145 1405 18185
rect 1445 18145 1455 18185
rect 1495 18145 1505 18185
rect 1545 18145 1555 18185
rect 1595 18145 1605 18185
rect 1645 18145 1655 18185
rect 1695 18145 1705 18185
rect 1745 18145 1755 18185
rect 1795 18145 1805 18185
rect 1845 18145 1855 18185
rect 1895 18145 1905 18185
rect 1945 18145 1955 18185
rect 1995 18145 2005 18185
rect 2045 18145 2055 18185
rect 2095 18145 2105 18185
rect 2145 18145 2155 18185
rect 2195 18145 2205 18185
rect 2245 18145 2255 18185
rect 2295 18145 2305 18185
rect 2345 18145 2355 18185
rect 2395 18145 2405 18185
rect 2445 18145 2455 18185
rect 2495 18145 2505 18185
rect 2545 18145 2555 18185
rect 2595 18145 2605 18185
rect 2645 18145 2655 18185
rect 2695 18145 2705 18185
rect 2745 18145 2755 18185
rect 2795 18145 2805 18185
rect 2845 18145 2855 18185
rect 2895 18145 2905 18185
rect 2945 18145 2955 18185
rect 2995 18145 3005 18185
rect 3045 18145 3055 18185
rect 3095 18145 3105 18185
rect 3145 18145 3155 18185
rect 3195 18145 3205 18185
rect 3245 18145 3255 18185
rect 3295 18145 3305 18185
rect 3345 18145 3355 18185
rect 3395 18145 3405 18185
rect 3445 18145 3455 18185
rect 3495 18145 3505 18185
rect 3545 18145 3555 18185
rect 3595 18145 3605 18185
rect 3645 18145 3655 18185
rect 3695 18145 3705 18185
rect 3745 18145 3755 18185
rect 3795 18145 3805 18185
rect 3845 18145 3855 18185
rect 3895 18145 3905 18185
rect 3945 18145 3955 18185
rect 3995 18145 4005 18185
rect 4045 18145 4055 18185
rect 4095 18145 4105 18185
rect 4145 18145 4155 18185
rect 4195 18145 4205 18185
rect 4245 18145 4255 18185
rect 4295 18145 4305 18185
rect 4345 18145 4355 18185
rect 4395 18145 4405 18185
rect 4445 18145 4455 18185
rect 4495 18145 4505 18185
rect 4545 18145 4555 18185
rect 4595 18145 4605 18185
rect 4645 18145 4655 18185
rect 4695 18145 4705 18185
rect 4745 18145 4755 18185
rect 4795 18145 4805 18185
rect 4845 18145 4855 18185
rect 4895 18145 4905 18185
rect 4945 18145 4955 18185
rect 4995 18145 5005 18185
rect 5045 18145 5055 18185
rect 5095 18145 5105 18185
rect 5145 18145 5155 18185
rect 5195 18145 5205 18185
rect 5245 18145 5255 18185
rect 5295 18145 5305 18185
rect 5345 18145 5355 18185
rect 5395 18145 5405 18185
rect 5445 18145 5455 18185
rect 5495 18145 5505 18185
rect 5545 18145 5555 18185
rect 5595 18145 5605 18185
rect 5645 18145 5655 18185
rect 5695 18145 5705 18185
rect 5745 18145 5755 18185
rect 5795 18145 5805 18185
rect 5845 18145 5855 18185
rect 5895 18145 5905 18185
rect 5945 18145 5955 18185
rect 5995 18145 6005 18185
rect 6045 18145 6055 18185
rect 6095 18145 6105 18185
rect 6145 18145 6155 18185
rect 6195 18145 6205 18185
rect 6245 18145 6255 18185
rect 6295 18145 6305 18185
rect 6345 18145 6355 18185
rect 6395 18145 6405 18185
rect 6445 18145 6455 18185
rect 6495 18145 6505 18185
rect 6545 18145 6555 18185
rect 6595 18145 6605 18185
rect 6645 18145 6655 18185
rect 6695 18145 6705 18185
rect 6745 18145 6755 18185
rect 6795 18145 6805 18185
rect 6845 18145 6855 18185
rect 6895 18145 6905 18185
rect 6945 18145 6955 18185
rect 6995 18145 7005 18185
rect 7045 18145 7055 18185
rect 7095 18145 7105 18185
rect 7145 18145 7155 18185
rect 7195 18145 7205 18185
rect 7245 18145 7255 18185
rect 7295 18145 7305 18185
rect 7345 18145 7355 18185
rect 7395 18145 7405 18185
rect 7445 18145 7455 18185
rect 7495 18145 7505 18185
rect 7545 18145 7555 18185
rect 7595 18145 7605 18185
rect 7645 18145 7655 18185
rect 7695 18145 7705 18185
rect 7745 18145 7755 18185
rect 7795 18145 7805 18185
rect 7845 18145 7855 18185
rect 7895 18145 7905 18185
rect 7945 18145 7955 18185
rect 7995 18145 8005 18185
rect 8045 18145 8055 18185
rect 8095 18145 8105 18185
rect 8145 18145 8155 18185
rect 8195 18145 8205 18185
rect 8245 18145 8255 18185
rect 8295 18145 8305 18185
rect 8345 18145 8355 18185
rect 8395 18145 8405 18185
rect 8445 18145 8455 18185
rect 8495 18145 8505 18185
rect 8545 18145 8555 18185
rect 8595 18145 8605 18185
rect 8645 18145 8655 18185
rect 8695 18145 8705 18185
rect 8745 18145 8755 18185
rect 8795 18145 8805 18185
rect 8845 18145 8855 18185
rect 8895 18145 8905 18185
rect 8945 18145 8955 18185
rect 8995 18145 9005 18185
rect 9045 18145 9055 18185
rect 9095 18145 9105 18185
rect 9145 18145 9155 18185
rect 9195 18145 9205 18185
rect 9245 18145 9255 18185
rect 9295 18145 9305 18185
rect 9345 18145 9355 18185
rect 9395 18145 9405 18185
rect 9445 18145 9455 18185
rect 9495 18145 9505 18185
rect 9545 18145 9555 18185
rect 9595 18145 9605 18185
rect 9645 18145 9655 18185
rect 9695 18145 9705 18185
rect 9745 18145 9755 18185
rect 9795 18145 9805 18185
rect 9845 18145 9855 18185
rect 9895 18145 9905 18185
rect 9945 18145 9955 18185
rect 9995 18145 10005 18185
rect 10045 18145 10055 18185
rect 10095 18145 10105 18185
rect 10145 18145 10155 18185
rect 10195 18145 10205 18185
rect 10245 18145 10255 18185
rect 10295 18145 10305 18185
rect 10345 18145 10355 18185
rect 10395 18145 10405 18185
rect 10445 18145 10455 18185
rect 10495 18145 10505 18185
rect 10545 18145 10555 18185
rect 10595 18145 10605 18185
rect 10645 18145 10655 18185
rect 10695 18145 10705 18185
rect 10745 18145 10755 18185
rect 10795 18145 10805 18185
rect 10845 18145 10855 18185
rect 10895 18145 10905 18185
rect 10945 18145 10955 18185
rect 10995 18145 11005 18185
rect 11045 18145 11055 18185
rect 11095 18145 11105 18185
rect 11145 18145 11155 18185
rect 11195 18145 11205 18185
rect 11245 18145 11255 18185
rect 11295 18145 11305 18185
rect 11345 18145 11355 18185
rect 11395 18145 11405 18185
rect 11445 18145 11455 18185
rect 11495 18145 11505 18185
rect 11545 18145 11555 18185
rect 11595 18145 11605 18185
rect 11645 18145 11655 18185
rect 11695 18145 11705 18185
rect 11745 18145 11755 18185
rect 11795 18145 11805 18185
rect 11845 18145 11855 18185
rect 11895 18145 11905 18185
rect 11945 18145 11955 18185
rect 11995 18145 12005 18185
rect 12045 18145 12055 18185
rect 12095 18145 12105 18185
rect 12145 18145 12155 18185
rect 12195 18145 12205 18185
rect 12245 18145 12255 18185
rect 12295 18145 12305 18185
rect 12345 18145 12355 18185
rect 12395 18145 12405 18185
rect 12445 18145 12455 18185
rect 12495 18145 12505 18185
rect 12545 18145 12555 18185
rect 12595 18145 12605 18185
rect 12645 18145 12655 18185
rect 12695 18145 12705 18185
rect 12745 18145 12755 18185
rect 12795 18145 12805 18185
rect 12845 18145 12855 18185
rect 12895 18145 12905 18185
rect 12945 18145 12955 18185
rect 12995 18145 13005 18185
rect 13045 18145 13055 18185
rect 13095 18145 13105 18185
rect 13145 18145 13155 18185
rect 13195 18145 13205 18185
rect 13245 18145 13255 18185
rect 13295 18145 13305 18185
rect 13345 18145 13355 18185
rect 13395 18145 13405 18185
rect 13445 18145 13455 18185
rect 13495 18145 13505 18185
rect 13545 18145 13555 18185
rect 13595 18145 13605 18185
rect 13645 18145 13655 18185
rect 13695 18145 13705 18185
rect 13745 18145 13755 18185
rect 13795 18145 13805 18185
rect 13845 18145 13855 18185
rect 13895 18145 13905 18185
rect 13945 18145 13955 18185
rect 13995 18145 14005 18185
rect 14045 18145 14055 18185
rect 14095 18145 14105 18185
rect 14145 18145 14155 18185
rect 14195 18145 14205 18185
rect 14245 18145 14255 18185
rect 14295 18145 14305 18185
rect 14345 18145 14355 18185
rect 14395 18145 14405 18185
rect 14445 18145 14455 18185
rect 14495 18145 14505 18185
rect 14545 18145 14555 18185
rect 14595 18145 14605 18185
rect 14645 18145 14655 18185
rect 14695 18145 14705 18185
rect 14745 18145 14755 18185
rect 14795 18145 14805 18185
rect 14845 18145 14855 18185
rect 14895 18145 14905 18185
rect 14945 18145 14955 18185
rect 14995 18145 15005 18185
rect 15045 18145 15055 18185
rect 15095 18145 15105 18185
rect 15145 18145 15155 18185
rect 15195 18145 15205 18185
rect 15245 18145 15255 18185
rect 15295 18145 15305 18185
rect 15345 18145 15355 18185
rect 15395 18145 15405 18185
rect 15445 18145 15455 18185
rect 15495 18145 15505 18185
rect 15545 18145 15555 18185
rect 15595 18145 15605 18185
rect 15645 18145 15655 18185
rect 15695 18145 15705 18185
rect 15745 18145 15755 18185
rect 15795 18145 15805 18185
rect 15845 18145 15855 18185
rect 15895 18145 15905 18185
rect 15945 18145 15955 18185
rect 15995 18145 16005 18185
rect 16045 18145 16055 18185
rect 16095 18145 16105 18185
rect 16145 18145 16155 18185
rect 16195 18145 16205 18185
rect 16245 18145 16255 18185
rect 16295 18145 16305 18185
rect 16345 18145 16355 18185
rect 16395 18145 16405 18185
rect 16445 18145 16455 18185
rect 16495 18145 16505 18185
rect 16545 18145 16555 18185
rect 16595 18145 16605 18185
rect 16645 18145 16655 18185
rect 16695 18145 16705 18185
rect 16745 18145 16755 18185
rect 16795 18145 16805 18185
rect 16845 18145 16855 18185
rect 16895 18145 16905 18185
rect 16945 18145 16955 18185
rect 16995 18145 17005 18185
rect 17045 18145 17055 18185
rect 17095 18145 17105 18185
rect 17145 18145 17155 18185
rect 17195 18145 17205 18185
rect 17245 18145 17255 18185
rect 17295 18145 17305 18185
rect 17345 18145 17355 18185
rect 17395 18145 17405 18185
rect 17445 18145 17455 18185
rect 17495 18145 17505 18185
rect 17545 18145 17555 18185
rect 17595 18145 17605 18185
rect 17645 18145 17655 18185
rect 17695 18145 17705 18185
rect 17745 18145 17755 18185
rect 17795 18145 17805 18185
rect 17845 18145 17855 18185
rect 17895 18145 17905 18185
rect 17945 18145 17955 18185
rect 17995 18145 18005 18185
rect 18045 18145 18055 18185
rect 18095 18145 18105 18185
rect 18145 18145 18155 18185
rect 18195 18145 18205 18185
rect 18245 18145 18255 18185
rect 18295 18145 18305 18185
rect 18345 18145 18355 18185
rect 18395 18145 18405 18185
rect 18445 18145 18455 18185
rect 18495 18145 18505 18185
rect 18545 18145 18555 18185
rect 18595 18145 18605 18185
rect 18645 18145 18655 18185
rect 18695 18145 18705 18185
rect 18745 18145 18755 18185
rect 18795 18145 18805 18185
rect 18845 18145 18855 18185
rect 18895 18145 18905 18185
rect 18945 18145 18955 18185
rect 18995 18145 19005 18185
rect 19045 18145 19055 18185
rect 19095 18145 19105 18185
rect 19145 18145 19155 18185
rect 19195 18145 19205 18185
rect 19245 18145 19255 18185
rect 19295 18145 19305 18185
rect 19345 18145 19355 18185
rect 19395 18145 19405 18185
rect 19445 18145 19455 18185
rect 19495 18145 19505 18185
rect 19545 18145 19555 18185
rect 19595 18145 19605 18185
rect 19645 18145 19655 18185
rect 19695 18145 19705 18185
rect 19745 18145 19755 18185
rect 19795 18145 19805 18185
rect 19845 18145 19855 18185
rect 19895 18145 19905 18185
rect 19945 18145 19955 18185
rect 19995 18145 20005 18185
rect 20045 18145 20055 18185
rect 20095 18145 20105 18185
rect 20145 18145 20155 18185
rect 20195 18145 20205 18185
rect 20245 18145 20255 18185
rect 20295 18145 20305 18185
rect 20345 18145 20355 18185
rect 20395 18145 20405 18185
rect 20445 18145 20455 18185
rect 20495 18145 20505 18185
rect 20545 18145 20555 18185
rect 20595 18145 20605 18185
rect 20645 18145 20655 18185
rect 20695 18145 20705 18185
rect 20745 18145 20755 18185
rect 20795 18145 20805 18185
rect 20845 18145 20855 18185
rect 20895 18145 20905 18185
rect 20945 18145 20955 18185
rect 20995 18145 21005 18185
rect 21045 18145 21055 18185
rect 21095 18145 21105 18185
rect 21145 18145 21155 18185
rect 21195 18145 21205 18185
rect 21245 18145 21255 18185
rect 21295 18145 21305 18185
rect 21345 18145 21355 18185
rect 21395 18145 21405 18185
rect 21445 18145 21455 18185
rect 21495 18145 21505 18185
rect 21545 18145 21555 18185
rect 21595 18145 21605 18185
rect 21645 18145 21655 18185
rect 21695 18145 21705 18185
rect 21745 18145 21755 18185
rect 21795 18145 21805 18185
rect 21845 18145 21855 18185
rect 21895 18145 21905 18185
rect 21945 18145 21955 18185
rect 21995 18145 22005 18185
rect 22045 18145 22055 18185
rect 22095 18145 22105 18185
rect 22145 18145 22155 18185
rect 22195 18145 22205 18185
rect 22245 18145 22255 18185
rect 22295 18145 22305 18185
rect 22345 18145 22355 18185
rect 22395 18145 22405 18185
rect 22445 18145 22455 18185
rect 22495 18145 22505 18185
rect 22545 18145 22555 18185
rect 22595 18145 22605 18185
rect 22645 18145 22655 18185
rect 22695 18145 22705 18185
rect 22745 18145 22755 18185
rect 22795 18145 22805 18185
rect 22845 18145 22855 18185
rect 22895 18145 22905 18185
rect 22945 18145 22955 18185
rect 22995 18145 23005 18185
rect 23045 18145 23055 18185
rect 23095 18145 23105 18185
rect 23145 18145 23155 18185
rect 23195 18145 23205 18185
rect 23245 18145 23255 18185
rect 23295 18145 23305 18185
rect 23345 18145 23355 18185
rect 23395 18145 23405 18185
rect 23445 18145 23455 18185
rect 23495 18145 23505 18185
rect 23545 18145 23555 18185
rect 23595 18145 23605 18185
rect 23645 18145 23655 18185
rect 23695 18145 23705 18185
rect 23745 18145 23755 18185
rect 23795 18145 23805 18185
rect 23845 18145 23855 18185
rect 23895 18145 23905 18185
rect 23945 18145 23955 18185
rect 23995 18145 24005 18185
rect 24045 18145 24055 18185
rect 24095 18145 24105 18185
rect 24145 18145 24155 18185
rect 24195 18145 24205 18185
rect 24245 18145 24255 18185
rect 24295 18145 24305 18185
rect 24345 18145 24355 18185
rect 24395 18145 24405 18185
rect 24445 18145 24455 18185
rect 24495 18145 24505 18185
rect 24545 18145 24555 18185
rect 24595 18145 24605 18185
rect 24645 18145 24655 18185
rect 24695 18145 24705 18185
rect 24745 18145 24755 18185
rect 24795 18145 24805 18185
rect 24845 18145 24855 18185
rect 24895 18145 24905 18185
rect 24945 18145 24955 18185
rect 24995 18145 25005 18185
rect 25045 18145 25055 18185
rect 25095 18145 25105 18185
rect 25145 18145 25155 18185
rect 25195 18145 25205 18185
rect 25245 18145 25255 18185
rect 25295 18145 25305 18185
rect 25345 18145 25355 18185
rect 25395 18145 25405 18185
rect 25445 18145 25455 18185
rect 25495 18145 25505 18185
rect 25545 18145 25555 18185
rect 25595 18145 25605 18185
rect 25645 18145 25655 18185
rect 25695 18145 25705 18185
rect 25745 18145 25755 18185
rect 25795 18145 25805 18185
rect 25845 18145 25855 18185
rect 25895 18145 25905 18185
rect 25945 18145 25955 18185
rect 25995 18145 26005 18185
rect 26045 18145 26055 18185
rect 26095 18145 26105 18185
rect 26145 18145 26155 18185
rect 26195 18145 26205 18185
rect 26245 18145 26255 18185
rect 26295 18145 26305 18185
rect 26345 18145 26355 18185
rect 26395 18145 26405 18185
rect 26445 18145 26455 18185
rect 26495 18145 26505 18185
rect 26545 18145 26555 18185
rect 26595 18145 26605 18185
rect 26645 18145 26655 18185
rect 26695 18145 26705 18185
rect 26745 18145 26755 18185
rect 26795 18145 26805 18185
rect 26845 18145 26855 18185
rect 26895 18145 26905 18185
rect 26945 18145 26955 18185
rect 26995 18145 27005 18185
rect 27045 18145 27055 18185
rect 27095 18145 27105 18185
rect 27145 18145 27155 18185
rect 27195 18145 27205 18185
rect 27245 18145 27255 18185
rect 27295 18145 27305 18185
rect 27345 18145 27355 18185
rect 27395 18145 27405 18185
rect 27445 18145 27455 18185
rect 27495 18145 27505 18185
rect 27545 18145 27555 18185
rect 27595 18145 27605 18185
rect 27645 18145 27655 18185
rect 27695 18145 27705 18185
rect 27745 18145 27755 18185
rect 27795 18145 27805 18185
rect 27845 18145 27855 18185
rect 27895 18145 27905 18185
rect 27945 18145 27955 18185
rect 27995 18145 28005 18185
rect 28045 18145 28055 18185
rect 28095 18145 28105 18185
rect 28145 18145 28155 18185
rect 28195 18145 28205 18185
rect 28245 18145 28255 18185
rect 28295 18145 28305 18185
rect 28345 18145 28355 18185
rect 28395 18145 28405 18185
rect 28445 18145 28455 18185
rect 28495 18145 28505 18185
rect 28545 18145 28555 18185
rect 28595 18145 28605 18185
rect 28645 18145 28655 18185
rect 28695 18145 28705 18185
rect 28745 18145 28755 18185
rect 28795 18145 28805 18185
rect 28845 18145 28855 18185
rect 28895 18145 28905 18185
rect 28945 18145 28955 18185
rect 28995 18145 29005 18185
rect 29045 18145 29055 18185
rect 29095 18145 29105 18185
rect 29145 18145 29155 18185
rect 29195 18145 29205 18185
rect 29245 18145 29255 18185
rect 29295 18145 29305 18185
rect 29345 18145 29355 18185
rect 29395 18145 29405 18185
rect 29445 18145 29455 18185
rect 29495 18145 29505 18185
rect 29545 18145 29555 18185
rect 29595 18145 29605 18185
rect 29645 18145 29655 18185
rect 29695 18145 29705 18185
rect 29745 18145 29755 18185
rect 29795 18145 29805 18185
rect 29845 18145 29855 18185
rect 29895 18145 29905 18185
rect 29945 18145 29955 18185
rect 29995 18145 30005 18185
rect 30045 18145 30055 18185
rect 30095 18145 30105 18185
rect 30145 18145 30155 18185
rect 30195 18145 30205 18185
rect 30245 18145 30255 18185
rect 30295 18145 30305 18185
rect 30345 18145 30355 18185
rect 30395 18145 30405 18185
rect 30445 18145 30455 18185
rect 30495 18145 30505 18185
rect 30545 18145 30555 18185
rect 30595 18145 30605 18185
rect 30645 18145 30655 18185
rect 30695 18145 30705 18185
rect 30745 18145 30755 18185
rect 30795 18145 30805 18185
rect 30845 18145 30855 18185
rect 30895 18145 30905 18185
rect 30945 18145 30955 18185
rect 30995 18145 31005 18185
rect 31045 18145 31055 18185
rect 31095 18145 31105 18185
rect 31145 18145 31155 18185
rect 31195 18145 31205 18185
rect 31245 18145 31255 18185
rect 31295 18145 31305 18185
rect 31345 18145 31355 18185
rect 31395 18145 31405 18185
rect 31445 18145 31455 18185
rect 31495 18145 31505 18185
rect 31545 18145 31555 18185
rect 31595 18145 31605 18185
rect 31645 18145 31655 18185
rect 31695 18145 31705 18185
rect 31745 18145 31755 18185
rect 31795 18145 31805 18185
rect 31845 18145 31855 18185
rect 31895 18145 31905 18185
rect 31945 18145 31955 18185
rect 31995 18145 32005 18185
rect 32045 18145 32055 18185
rect 32095 18145 32105 18185
rect 32145 18145 32155 18185
rect 32195 18145 32205 18185
rect 32245 18145 32255 18185
rect 32295 18145 32305 18185
rect 32345 18145 32355 18185
rect 32395 18145 32405 18185
rect 32445 18145 32455 18185
rect 32495 18145 32505 18185
rect 32545 18145 32555 18185
rect 32595 18145 32605 18185
rect 32645 18145 32655 18185
rect 32695 18145 32705 18185
rect 32745 18145 32755 18185
rect 32795 18145 32805 18185
rect 32845 18145 32855 18185
rect 32895 18145 32905 18185
rect 32945 18145 32955 18185
rect 32995 18145 33005 18185
rect 33045 18145 33055 18185
rect 33095 18145 33105 18185
rect 33145 18145 33155 18185
rect 33195 18145 33205 18185
rect 33245 18145 33255 18185
rect 33295 18145 33305 18185
rect 33345 18145 33355 18185
rect 33395 18145 33405 18185
rect 33445 18145 33455 18185
rect 33495 18145 33505 18185
rect 33545 18145 33555 18185
rect 33595 18145 33605 18185
rect 33645 18145 33655 18185
rect 33695 18145 33705 18185
rect 33745 18145 33755 18185
rect 33795 18145 33805 18185
rect 33845 18145 33855 18185
rect 33895 18145 33905 18185
rect 33945 18145 33955 18185
rect 33995 18145 34005 18185
rect 34045 18145 34055 18185
rect 34095 18145 34105 18185
rect 34145 18145 34155 18185
rect 34195 18145 34205 18185
rect 34245 18145 34255 18185
rect 34295 18145 34305 18185
rect 34345 18145 34355 18185
rect 34395 18145 34405 18185
rect 34445 18145 34455 18185
rect 34495 18145 34505 18185
rect 34545 18145 34555 18185
rect 34595 18145 34605 18185
rect 34645 18145 34655 18185
rect 34695 18145 34705 18185
rect 34745 18145 34755 18185
rect 34795 18145 34805 18185
rect 34845 18145 34855 18185
rect 34895 18145 34905 18185
rect 34945 18145 34955 18185
rect 34995 18145 35005 18185
rect 35045 18145 35055 18185
rect 35095 18145 35105 18185
rect 35145 18145 35155 18185
rect 35195 18145 35205 18185
rect 35245 18145 35255 18185
rect 35295 18145 35305 18185
rect 35345 18145 35355 18185
rect 35395 18145 35405 18185
rect 35445 18145 35455 18185
rect 35495 18145 35505 18185
rect 35545 18145 35555 18185
rect 35595 18145 35605 18185
rect 35645 18145 35655 18185
rect 35695 18145 35705 18185
rect 35745 18145 35755 18185
rect 35795 18145 35805 18185
rect 35845 18145 35855 18185
rect 35895 18145 35905 18185
rect 35945 18145 35955 18185
rect 35995 18145 36005 18185
rect 36045 18145 36055 18185
rect 36095 18145 36105 18185
rect 36145 18145 36155 18185
rect 36195 18145 36205 18185
rect 36245 18145 36255 18185
rect 36295 18145 36305 18185
rect 36345 18145 36355 18185
rect 36395 18145 36405 18185
rect 36445 18145 36455 18185
rect 36495 18145 36505 18185
rect 36545 18145 36555 18185
rect 36595 18145 36605 18185
rect 36645 18145 36655 18185
rect 36695 18145 36705 18185
rect 36745 18145 36755 18185
rect 36795 18145 36805 18185
rect 36845 18145 36855 18185
rect 36895 18145 36905 18185
rect 36945 18145 36955 18185
rect 36995 18145 37005 18185
rect 37045 18145 37055 18185
rect 37095 18145 37105 18185
rect 37145 18145 37155 18185
rect 37195 18145 37205 18185
rect 37245 18145 37255 18185
rect 37295 18145 37305 18185
rect 37345 18145 37355 18185
rect 37395 18145 37405 18185
rect 37445 18145 37455 18185
rect 37495 18145 37505 18185
rect 37545 18145 37555 18185
rect 37595 18145 37605 18185
rect 37645 18145 37655 18185
rect 37695 18145 37705 18185
rect 37745 18145 37755 18185
rect 37795 18145 37805 18185
rect 37845 18145 37855 18185
rect 37895 18145 37905 18185
rect 37945 18145 37955 18185
rect 37995 18145 38005 18185
rect 38045 18145 38055 18185
rect 38095 18145 38105 18185
rect 38145 18145 38155 18185
rect 38195 18145 38205 18185
rect 38245 18145 38255 18185
rect 38295 18145 38305 18185
rect 38345 18145 38355 18185
rect 38395 18145 38405 18185
rect 38445 18145 38455 18185
rect 38495 18145 38505 18185
rect 38545 18145 38555 18185
rect 38595 18145 38605 18185
rect 38645 18145 38655 18185
rect 38695 18145 38705 18185
rect 38745 18145 38755 18185
rect 38795 18145 38805 18185
rect 38845 18145 38855 18185
rect 38895 18145 38905 18185
rect 38945 18145 38955 18185
rect 38995 18145 39005 18185
rect 39045 18145 39055 18185
rect 39095 18145 39105 18185
rect 39145 18145 39155 18185
rect 39195 18145 39205 18185
rect 39245 18145 39255 18185
rect 39295 18145 39305 18185
rect 39345 18145 39355 18185
rect 39395 18145 39405 18185
rect 39445 18145 39455 18185
rect 39495 18145 39505 18185
rect 39545 18145 39555 18185
rect 39595 18145 39605 18185
rect 39645 18145 39655 18185
rect 39695 18145 39705 18185
rect 39745 18145 39750 18185
rect 0 18140 39750 18145
rect 100 17240 3200 18140
rect 3350 17240 6450 18140
rect 6600 17240 9700 18140
rect 9850 17240 12950 18140
rect 13100 17240 16200 18140
rect 16350 17240 19450 18140
rect 19600 17240 22700 18140
rect 22850 17240 25950 18140
rect 26100 17240 29200 18140
rect 29350 17240 32450 18140
rect 32600 17240 35700 18140
rect 35850 17240 38950 18140
rect 39100 17240 39750 18140
rect -2700 17115 39750 17120
rect -2700 17075 -2695 17115
rect -2655 17075 105 17115
rect 145 17075 155 17115
rect 195 17075 205 17115
rect 245 17075 255 17115
rect 295 17075 305 17115
rect 345 17075 355 17115
rect 395 17075 405 17115
rect 445 17075 455 17115
rect 495 17075 505 17115
rect 545 17075 555 17115
rect 595 17075 605 17115
rect 645 17075 655 17115
rect 695 17075 705 17115
rect 745 17075 755 17115
rect 795 17075 805 17115
rect 845 17075 855 17115
rect 895 17075 905 17115
rect 945 17075 955 17115
rect 995 17075 1005 17115
rect 1045 17075 1055 17115
rect 1095 17075 1105 17115
rect 1145 17075 1155 17115
rect 1195 17075 1205 17115
rect 1245 17075 1255 17115
rect 1295 17075 1305 17115
rect 1345 17075 1355 17115
rect 1395 17075 1405 17115
rect 1445 17075 1455 17115
rect 1495 17075 1505 17115
rect 1545 17075 1555 17115
rect 1595 17075 1605 17115
rect 1645 17075 1655 17115
rect 1695 17075 1705 17115
rect 1745 17075 1755 17115
rect 1795 17075 1805 17115
rect 1845 17075 1855 17115
rect 1895 17075 1905 17115
rect 1945 17075 1955 17115
rect 1995 17075 2005 17115
rect 2045 17075 2055 17115
rect 2095 17075 2105 17115
rect 2145 17075 2155 17115
rect 2195 17075 2205 17115
rect 2245 17075 2255 17115
rect 2295 17075 2305 17115
rect 2345 17075 2355 17115
rect 2395 17075 2405 17115
rect 2445 17075 2455 17115
rect 2495 17075 2505 17115
rect 2545 17075 2555 17115
rect 2595 17075 2605 17115
rect 2645 17075 2655 17115
rect 2695 17075 2705 17115
rect 2745 17075 2755 17115
rect 2795 17075 2805 17115
rect 2845 17075 2855 17115
rect 2895 17075 2905 17115
rect 2945 17075 2955 17115
rect 2995 17075 3005 17115
rect 3045 17075 3055 17115
rect 3095 17075 3105 17115
rect 3145 17075 3155 17115
rect 3195 17075 3205 17115
rect 3245 17075 3255 17115
rect 3295 17075 3305 17115
rect 3345 17075 3355 17115
rect 3395 17075 3405 17115
rect 3445 17075 3455 17115
rect 3495 17075 3505 17115
rect 3545 17075 3555 17115
rect 3595 17075 3605 17115
rect 3645 17075 3655 17115
rect 3695 17075 3705 17115
rect 3745 17075 3755 17115
rect 3795 17075 3805 17115
rect 3845 17075 3855 17115
rect 3895 17075 3905 17115
rect 3945 17075 3955 17115
rect 3995 17075 4005 17115
rect 4045 17075 4055 17115
rect 4095 17075 4105 17115
rect 4145 17075 4155 17115
rect 4195 17075 4205 17115
rect 4245 17075 4255 17115
rect 4295 17075 4305 17115
rect 4345 17075 4355 17115
rect 4395 17075 4405 17115
rect 4445 17075 4455 17115
rect 4495 17075 4505 17115
rect 4545 17075 4555 17115
rect 4595 17075 4605 17115
rect 4645 17075 4655 17115
rect 4695 17075 4705 17115
rect 4745 17075 4755 17115
rect 4795 17075 4805 17115
rect 4845 17075 4855 17115
rect 4895 17075 4905 17115
rect 4945 17075 4955 17115
rect 4995 17075 5005 17115
rect 5045 17075 5055 17115
rect 5095 17075 5105 17115
rect 5145 17075 5155 17115
rect 5195 17075 5205 17115
rect 5245 17075 5255 17115
rect 5295 17075 5305 17115
rect 5345 17075 5355 17115
rect 5395 17075 5405 17115
rect 5445 17075 5455 17115
rect 5495 17075 5505 17115
rect 5545 17075 5555 17115
rect 5595 17075 5605 17115
rect 5645 17075 5655 17115
rect 5695 17075 5705 17115
rect 5745 17075 5755 17115
rect 5795 17075 5805 17115
rect 5845 17075 5855 17115
rect 5895 17075 5905 17115
rect 5945 17075 5955 17115
rect 5995 17075 6005 17115
rect 6045 17075 6055 17115
rect 6095 17075 6105 17115
rect 6145 17075 6155 17115
rect 6195 17075 6205 17115
rect 6245 17075 6255 17115
rect 6295 17075 6305 17115
rect 6345 17075 6355 17115
rect 6395 17075 6405 17115
rect 6445 17075 6455 17115
rect 6495 17075 6505 17115
rect 6545 17075 6555 17115
rect 6595 17075 6605 17115
rect 6645 17075 6655 17115
rect 6695 17075 6705 17115
rect 6745 17075 6755 17115
rect 6795 17075 6805 17115
rect 6845 17075 6855 17115
rect 6895 17075 6905 17115
rect 6945 17075 6955 17115
rect 6995 17075 7005 17115
rect 7045 17075 7055 17115
rect 7095 17075 7105 17115
rect 7145 17075 7155 17115
rect 7195 17075 7205 17115
rect 7245 17075 7255 17115
rect 7295 17075 7305 17115
rect 7345 17075 7355 17115
rect 7395 17075 7405 17115
rect 7445 17075 7455 17115
rect 7495 17075 7505 17115
rect 7545 17075 7555 17115
rect 7595 17075 7605 17115
rect 7645 17075 7655 17115
rect 7695 17075 7705 17115
rect 7745 17075 7755 17115
rect 7795 17075 7805 17115
rect 7845 17075 7855 17115
rect 7895 17075 7905 17115
rect 7945 17075 7955 17115
rect 7995 17075 8005 17115
rect 8045 17075 8055 17115
rect 8095 17075 8105 17115
rect 8145 17075 8155 17115
rect 8195 17075 8205 17115
rect 8245 17075 8255 17115
rect 8295 17075 8305 17115
rect 8345 17075 8355 17115
rect 8395 17075 8405 17115
rect 8445 17075 8455 17115
rect 8495 17075 8505 17115
rect 8545 17075 8555 17115
rect 8595 17075 8605 17115
rect 8645 17075 8655 17115
rect 8695 17075 8705 17115
rect 8745 17075 8755 17115
rect 8795 17075 8805 17115
rect 8845 17075 8855 17115
rect 8895 17075 8905 17115
rect 8945 17075 8955 17115
rect 8995 17075 9005 17115
rect 9045 17075 9055 17115
rect 9095 17075 9105 17115
rect 9145 17075 9155 17115
rect 9195 17075 9205 17115
rect 9245 17075 9255 17115
rect 9295 17075 9305 17115
rect 9345 17075 9355 17115
rect 9395 17075 9405 17115
rect 9445 17075 9455 17115
rect 9495 17075 9505 17115
rect 9545 17075 9555 17115
rect 9595 17075 9605 17115
rect 9645 17075 9655 17115
rect 9695 17075 9705 17115
rect 9745 17075 9755 17115
rect 9795 17075 9805 17115
rect 9845 17075 9855 17115
rect 9895 17075 9905 17115
rect 9945 17075 9955 17115
rect 9995 17075 10005 17115
rect 10045 17075 10055 17115
rect 10095 17075 10105 17115
rect 10145 17075 10155 17115
rect 10195 17075 10205 17115
rect 10245 17075 10255 17115
rect 10295 17075 10305 17115
rect 10345 17075 10355 17115
rect 10395 17075 10405 17115
rect 10445 17075 10455 17115
rect 10495 17075 10505 17115
rect 10545 17075 10555 17115
rect 10595 17075 10605 17115
rect 10645 17075 10655 17115
rect 10695 17075 10705 17115
rect 10745 17075 10755 17115
rect 10795 17075 10805 17115
rect 10845 17075 10855 17115
rect 10895 17075 10905 17115
rect 10945 17075 10955 17115
rect 10995 17075 11005 17115
rect 11045 17075 11055 17115
rect 11095 17075 11105 17115
rect 11145 17075 11155 17115
rect 11195 17075 11205 17115
rect 11245 17075 11255 17115
rect 11295 17075 11305 17115
rect 11345 17075 11355 17115
rect 11395 17075 11405 17115
rect 11445 17075 11455 17115
rect 11495 17075 11505 17115
rect 11545 17075 11555 17115
rect 11595 17075 11605 17115
rect 11645 17075 11655 17115
rect 11695 17075 11705 17115
rect 11745 17075 11755 17115
rect 11795 17075 11805 17115
rect 11845 17075 11855 17115
rect 11895 17075 11905 17115
rect 11945 17075 11955 17115
rect 11995 17075 12005 17115
rect 12045 17075 12055 17115
rect 12095 17075 12105 17115
rect 12145 17075 12155 17115
rect 12195 17075 12205 17115
rect 12245 17075 12255 17115
rect 12295 17075 12305 17115
rect 12345 17075 12355 17115
rect 12395 17075 12405 17115
rect 12445 17075 12455 17115
rect 12495 17075 12505 17115
rect 12545 17075 12555 17115
rect 12595 17075 12605 17115
rect 12645 17075 12655 17115
rect 12695 17075 12705 17115
rect 12745 17075 12755 17115
rect 12795 17075 12805 17115
rect 12845 17075 12855 17115
rect 12895 17075 12905 17115
rect 12945 17075 12955 17115
rect 12995 17075 13005 17115
rect 13045 17075 13055 17115
rect 13095 17075 13105 17115
rect 13145 17075 13155 17115
rect 13195 17075 13205 17115
rect 13245 17075 13255 17115
rect 13295 17075 13305 17115
rect 13345 17075 13355 17115
rect 13395 17075 13405 17115
rect 13445 17075 13455 17115
rect 13495 17075 13505 17115
rect 13545 17075 13555 17115
rect 13595 17075 13605 17115
rect 13645 17075 13655 17115
rect 13695 17075 13705 17115
rect 13745 17075 13755 17115
rect 13795 17075 13805 17115
rect 13845 17075 13855 17115
rect 13895 17075 13905 17115
rect 13945 17075 13955 17115
rect 13995 17075 14005 17115
rect 14045 17075 14055 17115
rect 14095 17075 14105 17115
rect 14145 17075 14155 17115
rect 14195 17075 14205 17115
rect 14245 17075 14255 17115
rect 14295 17075 14305 17115
rect 14345 17075 14355 17115
rect 14395 17075 14405 17115
rect 14445 17075 14455 17115
rect 14495 17075 14505 17115
rect 14545 17075 14555 17115
rect 14595 17075 14605 17115
rect 14645 17075 14655 17115
rect 14695 17075 14705 17115
rect 14745 17075 14755 17115
rect 14795 17075 14805 17115
rect 14845 17075 14855 17115
rect 14895 17075 14905 17115
rect 14945 17075 14955 17115
rect 14995 17075 15005 17115
rect 15045 17075 15055 17115
rect 15095 17075 15105 17115
rect 15145 17075 15155 17115
rect 15195 17075 15205 17115
rect 15245 17075 15255 17115
rect 15295 17075 15305 17115
rect 15345 17075 15355 17115
rect 15395 17075 15405 17115
rect 15445 17075 15455 17115
rect 15495 17075 15505 17115
rect 15545 17075 15555 17115
rect 15595 17075 15605 17115
rect 15645 17075 15655 17115
rect 15695 17075 15705 17115
rect 15745 17075 15755 17115
rect 15795 17075 15805 17115
rect 15845 17075 15855 17115
rect 15895 17075 15905 17115
rect 15945 17075 15955 17115
rect 15995 17075 16005 17115
rect 16045 17075 16055 17115
rect 16095 17075 16105 17115
rect 16145 17075 16155 17115
rect 16195 17075 16205 17115
rect 16245 17075 16255 17115
rect 16295 17075 16305 17115
rect 16345 17075 16355 17115
rect 16395 17075 16405 17115
rect 16445 17075 16455 17115
rect 16495 17075 16505 17115
rect 16545 17075 16555 17115
rect 16595 17075 16605 17115
rect 16645 17075 16655 17115
rect 16695 17075 16705 17115
rect 16745 17075 16755 17115
rect 16795 17075 16805 17115
rect 16845 17075 16855 17115
rect 16895 17075 16905 17115
rect 16945 17075 16955 17115
rect 16995 17075 17005 17115
rect 17045 17075 17055 17115
rect 17095 17075 17105 17115
rect 17145 17075 17155 17115
rect 17195 17075 17205 17115
rect 17245 17075 17255 17115
rect 17295 17075 17305 17115
rect 17345 17075 17355 17115
rect 17395 17075 17405 17115
rect 17445 17075 17455 17115
rect 17495 17075 17505 17115
rect 17545 17075 17555 17115
rect 17595 17075 17605 17115
rect 17645 17075 17655 17115
rect 17695 17075 17705 17115
rect 17745 17075 17755 17115
rect 17795 17075 17805 17115
rect 17845 17075 17855 17115
rect 17895 17075 17905 17115
rect 17945 17075 17955 17115
rect 17995 17075 18005 17115
rect 18045 17075 18055 17115
rect 18095 17075 18105 17115
rect 18145 17075 18155 17115
rect 18195 17075 18205 17115
rect 18245 17075 18255 17115
rect 18295 17075 18305 17115
rect 18345 17075 18355 17115
rect 18395 17075 18405 17115
rect 18445 17075 18455 17115
rect 18495 17075 18505 17115
rect 18545 17075 18555 17115
rect 18595 17075 18605 17115
rect 18645 17075 18655 17115
rect 18695 17075 18705 17115
rect 18745 17075 18755 17115
rect 18795 17075 18805 17115
rect 18845 17075 18855 17115
rect 18895 17075 18905 17115
rect 18945 17075 18955 17115
rect 18995 17075 19005 17115
rect 19045 17075 19055 17115
rect 19095 17075 19105 17115
rect 19145 17075 19155 17115
rect 19195 17075 19205 17115
rect 19245 17075 19255 17115
rect 19295 17075 19305 17115
rect 19345 17075 19355 17115
rect 19395 17075 19405 17115
rect 19445 17075 19455 17115
rect 19495 17075 19505 17115
rect 19545 17075 19555 17115
rect 19595 17075 19605 17115
rect 19645 17075 19655 17115
rect 19695 17075 19705 17115
rect 19745 17075 19755 17115
rect 19795 17075 19805 17115
rect 19845 17075 19855 17115
rect 19895 17075 19905 17115
rect 19945 17075 19955 17115
rect 19995 17075 20005 17115
rect 20045 17075 20055 17115
rect 20095 17075 20105 17115
rect 20145 17075 20155 17115
rect 20195 17075 20205 17115
rect 20245 17075 20255 17115
rect 20295 17075 20305 17115
rect 20345 17075 20355 17115
rect 20395 17075 20405 17115
rect 20445 17075 20455 17115
rect 20495 17075 20505 17115
rect 20545 17075 20555 17115
rect 20595 17075 20605 17115
rect 20645 17075 20655 17115
rect 20695 17075 20705 17115
rect 20745 17075 20755 17115
rect 20795 17075 20805 17115
rect 20845 17075 20855 17115
rect 20895 17075 20905 17115
rect 20945 17075 20955 17115
rect 20995 17075 21005 17115
rect 21045 17075 21055 17115
rect 21095 17075 21105 17115
rect 21145 17075 21155 17115
rect 21195 17075 21205 17115
rect 21245 17075 21255 17115
rect 21295 17075 21305 17115
rect 21345 17075 21355 17115
rect 21395 17075 21405 17115
rect 21445 17075 21455 17115
rect 21495 17075 21505 17115
rect 21545 17075 21555 17115
rect 21595 17075 21605 17115
rect 21645 17075 21655 17115
rect 21695 17075 21705 17115
rect 21745 17075 21755 17115
rect 21795 17075 21805 17115
rect 21845 17075 21855 17115
rect 21895 17075 21905 17115
rect 21945 17075 21955 17115
rect 21995 17075 22005 17115
rect 22045 17075 22055 17115
rect 22095 17075 22105 17115
rect 22145 17075 22155 17115
rect 22195 17075 22205 17115
rect 22245 17075 22255 17115
rect 22295 17075 22305 17115
rect 22345 17075 22355 17115
rect 22395 17075 22405 17115
rect 22445 17075 22455 17115
rect 22495 17075 22505 17115
rect 22545 17075 22555 17115
rect 22595 17075 22605 17115
rect 22645 17075 22655 17115
rect 22695 17075 22705 17115
rect 22745 17075 22755 17115
rect 22795 17075 22805 17115
rect 22845 17075 22855 17115
rect 22895 17075 22905 17115
rect 22945 17075 22955 17115
rect 22995 17075 23005 17115
rect 23045 17075 23055 17115
rect 23095 17075 23105 17115
rect 23145 17075 23155 17115
rect 23195 17075 23205 17115
rect 23245 17075 23255 17115
rect 23295 17075 23305 17115
rect 23345 17075 23355 17115
rect 23395 17075 23405 17115
rect 23445 17075 23455 17115
rect 23495 17075 23505 17115
rect 23545 17075 23555 17115
rect 23595 17075 23605 17115
rect 23645 17075 23655 17115
rect 23695 17075 23705 17115
rect 23745 17075 23755 17115
rect 23795 17075 23805 17115
rect 23845 17075 23855 17115
rect 23895 17075 23905 17115
rect 23945 17075 23955 17115
rect 23995 17075 24005 17115
rect 24045 17075 24055 17115
rect 24095 17075 24105 17115
rect 24145 17075 24155 17115
rect 24195 17075 24205 17115
rect 24245 17075 24255 17115
rect 24295 17075 24305 17115
rect 24345 17075 24355 17115
rect 24395 17075 24405 17115
rect 24445 17075 24455 17115
rect 24495 17075 24505 17115
rect 24545 17075 24555 17115
rect 24595 17075 24605 17115
rect 24645 17075 24655 17115
rect 24695 17075 24705 17115
rect 24745 17075 24755 17115
rect 24795 17075 24805 17115
rect 24845 17075 24855 17115
rect 24895 17075 24905 17115
rect 24945 17075 24955 17115
rect 24995 17075 25005 17115
rect 25045 17075 25055 17115
rect 25095 17075 25105 17115
rect 25145 17075 25155 17115
rect 25195 17075 25205 17115
rect 25245 17075 25255 17115
rect 25295 17075 25305 17115
rect 25345 17075 25355 17115
rect 25395 17075 25405 17115
rect 25445 17075 25455 17115
rect 25495 17075 25505 17115
rect 25545 17075 25555 17115
rect 25595 17075 25605 17115
rect 25645 17075 25655 17115
rect 25695 17075 25705 17115
rect 25745 17075 25755 17115
rect 25795 17075 25805 17115
rect 25845 17075 25855 17115
rect 25895 17075 25905 17115
rect 25945 17075 25955 17115
rect 25995 17075 26005 17115
rect 26045 17075 26055 17115
rect 26095 17075 26105 17115
rect 26145 17075 26155 17115
rect 26195 17075 26205 17115
rect 26245 17075 26255 17115
rect 26295 17075 26305 17115
rect 26345 17075 26355 17115
rect 26395 17075 26405 17115
rect 26445 17075 26455 17115
rect 26495 17075 26505 17115
rect 26545 17075 26555 17115
rect 26595 17075 26605 17115
rect 26645 17075 26655 17115
rect 26695 17075 26705 17115
rect 26745 17075 26755 17115
rect 26795 17075 26805 17115
rect 26845 17075 26855 17115
rect 26895 17075 26905 17115
rect 26945 17075 26955 17115
rect 26995 17075 27005 17115
rect 27045 17075 27055 17115
rect 27095 17075 27105 17115
rect 27145 17075 27155 17115
rect 27195 17075 27205 17115
rect 27245 17075 27255 17115
rect 27295 17075 27305 17115
rect 27345 17075 27355 17115
rect 27395 17075 27405 17115
rect 27445 17075 27455 17115
rect 27495 17075 27505 17115
rect 27545 17075 27555 17115
rect 27595 17075 27605 17115
rect 27645 17075 27655 17115
rect 27695 17075 27705 17115
rect 27745 17075 27755 17115
rect 27795 17075 27805 17115
rect 27845 17075 27855 17115
rect 27895 17075 27905 17115
rect 27945 17075 27955 17115
rect 27995 17075 28005 17115
rect 28045 17075 28055 17115
rect 28095 17075 28105 17115
rect 28145 17075 28155 17115
rect 28195 17075 28205 17115
rect 28245 17075 28255 17115
rect 28295 17075 28305 17115
rect 28345 17075 28355 17115
rect 28395 17075 28405 17115
rect 28445 17075 28455 17115
rect 28495 17075 28505 17115
rect 28545 17075 28555 17115
rect 28595 17075 28605 17115
rect 28645 17075 28655 17115
rect 28695 17075 28705 17115
rect 28745 17075 28755 17115
rect 28795 17075 28805 17115
rect 28845 17075 28855 17115
rect 28895 17075 28905 17115
rect 28945 17075 28955 17115
rect 28995 17075 29005 17115
rect 29045 17075 29055 17115
rect 29095 17075 29105 17115
rect 29145 17075 29155 17115
rect 29195 17075 29205 17115
rect 29245 17075 29255 17115
rect 29295 17075 29305 17115
rect 29345 17075 29355 17115
rect 29395 17075 29405 17115
rect 29445 17075 29455 17115
rect 29495 17075 29505 17115
rect 29545 17075 29555 17115
rect 29595 17075 29605 17115
rect 29645 17075 29655 17115
rect 29695 17075 29705 17115
rect 29745 17075 29755 17115
rect 29795 17075 29805 17115
rect 29845 17075 29855 17115
rect 29895 17075 29905 17115
rect 29945 17075 29955 17115
rect 29995 17075 30005 17115
rect 30045 17075 30055 17115
rect 30095 17075 30105 17115
rect 30145 17075 30155 17115
rect 30195 17075 30205 17115
rect 30245 17075 30255 17115
rect 30295 17075 30305 17115
rect 30345 17075 30355 17115
rect 30395 17075 30405 17115
rect 30445 17075 30455 17115
rect 30495 17075 30505 17115
rect 30545 17075 30555 17115
rect 30595 17075 30605 17115
rect 30645 17075 30655 17115
rect 30695 17075 30705 17115
rect 30745 17075 30755 17115
rect 30795 17075 30805 17115
rect 30845 17075 30855 17115
rect 30895 17075 30905 17115
rect 30945 17075 30955 17115
rect 30995 17075 31005 17115
rect 31045 17075 31055 17115
rect 31095 17075 31105 17115
rect 31145 17075 31155 17115
rect 31195 17075 31205 17115
rect 31245 17075 31255 17115
rect 31295 17075 31305 17115
rect 31345 17075 31355 17115
rect 31395 17075 31405 17115
rect 31445 17075 31455 17115
rect 31495 17075 31505 17115
rect 31545 17075 31555 17115
rect 31595 17075 31605 17115
rect 31645 17075 31655 17115
rect 31695 17075 31705 17115
rect 31745 17075 31755 17115
rect 31795 17075 31805 17115
rect 31845 17075 31855 17115
rect 31895 17075 31905 17115
rect 31945 17075 31955 17115
rect 31995 17075 32005 17115
rect 32045 17075 32055 17115
rect 32095 17075 32105 17115
rect 32145 17075 32155 17115
rect 32195 17075 32205 17115
rect 32245 17075 32255 17115
rect 32295 17075 32305 17115
rect 32345 17075 32355 17115
rect 32395 17075 32405 17115
rect 32445 17075 32455 17115
rect 32495 17075 32505 17115
rect 32545 17075 32555 17115
rect 32595 17075 32605 17115
rect 32645 17075 32655 17115
rect 32695 17075 32705 17115
rect 32745 17075 32755 17115
rect 32795 17075 32805 17115
rect 32845 17075 32855 17115
rect 32895 17075 32905 17115
rect 32945 17075 32955 17115
rect 32995 17075 33005 17115
rect 33045 17075 33055 17115
rect 33095 17075 33105 17115
rect 33145 17075 33155 17115
rect 33195 17075 33205 17115
rect 33245 17075 33255 17115
rect 33295 17075 33305 17115
rect 33345 17075 33355 17115
rect 33395 17075 33405 17115
rect 33445 17075 33455 17115
rect 33495 17075 33505 17115
rect 33545 17075 33555 17115
rect 33595 17075 33605 17115
rect 33645 17075 33655 17115
rect 33695 17075 33705 17115
rect 33745 17075 33755 17115
rect 33795 17075 33805 17115
rect 33845 17075 33855 17115
rect 33895 17075 33905 17115
rect 33945 17075 33955 17115
rect 33995 17075 34005 17115
rect 34045 17075 34055 17115
rect 34095 17075 34105 17115
rect 34145 17075 34155 17115
rect 34195 17075 34205 17115
rect 34245 17075 34255 17115
rect 34295 17075 34305 17115
rect 34345 17075 34355 17115
rect 34395 17075 34405 17115
rect 34445 17075 34455 17115
rect 34495 17075 34505 17115
rect 34545 17075 34555 17115
rect 34595 17075 34605 17115
rect 34645 17075 34655 17115
rect 34695 17075 34705 17115
rect 34745 17075 34755 17115
rect 34795 17075 34805 17115
rect 34845 17075 34855 17115
rect 34895 17075 34905 17115
rect 34945 17075 34955 17115
rect 34995 17075 35005 17115
rect 35045 17075 35055 17115
rect 35095 17075 35105 17115
rect 35145 17075 35155 17115
rect 35195 17075 35205 17115
rect 35245 17075 35255 17115
rect 35295 17075 35305 17115
rect 35345 17075 35355 17115
rect 35395 17075 35405 17115
rect 35445 17075 35455 17115
rect 35495 17075 35505 17115
rect 35545 17075 35555 17115
rect 35595 17075 35605 17115
rect 35645 17075 35655 17115
rect 35695 17075 35705 17115
rect 35745 17075 35755 17115
rect 35795 17075 35805 17115
rect 35845 17075 35855 17115
rect 35895 17075 35905 17115
rect 35945 17075 35955 17115
rect 35995 17075 36005 17115
rect 36045 17075 36055 17115
rect 36095 17075 36105 17115
rect 36145 17075 36155 17115
rect 36195 17075 36205 17115
rect 36245 17075 36255 17115
rect 36295 17075 36305 17115
rect 36345 17075 36355 17115
rect 36395 17075 36405 17115
rect 36445 17075 36455 17115
rect 36495 17075 36505 17115
rect 36545 17075 36555 17115
rect 36595 17075 36605 17115
rect 36645 17075 36655 17115
rect 36695 17075 36705 17115
rect 36745 17075 36755 17115
rect 36795 17075 36805 17115
rect 36845 17075 36855 17115
rect 36895 17075 36905 17115
rect 36945 17075 36955 17115
rect 36995 17075 37005 17115
rect 37045 17075 37055 17115
rect 37095 17075 37105 17115
rect 37145 17075 37155 17115
rect 37195 17075 37205 17115
rect 37245 17075 37255 17115
rect 37295 17075 37305 17115
rect 37345 17075 37355 17115
rect 37395 17075 37405 17115
rect 37445 17075 37455 17115
rect 37495 17075 37505 17115
rect 37545 17075 37555 17115
rect 37595 17075 37605 17115
rect 37645 17075 37655 17115
rect 37695 17075 37705 17115
rect 37745 17075 37755 17115
rect 37795 17075 37805 17115
rect 37845 17075 37855 17115
rect 37895 17075 37905 17115
rect 37945 17075 37955 17115
rect 37995 17075 38005 17115
rect 38045 17075 38055 17115
rect 38095 17075 38105 17115
rect 38145 17075 38155 17115
rect 38195 17075 38205 17115
rect 38245 17075 38255 17115
rect 38295 17075 38305 17115
rect 38345 17075 38355 17115
rect 38395 17075 38405 17115
rect 38445 17075 38455 17115
rect 38495 17075 38505 17115
rect 38545 17075 38555 17115
rect 38595 17075 38605 17115
rect 38645 17075 38655 17115
rect 38695 17075 38705 17115
rect 38745 17075 38755 17115
rect 38795 17075 38805 17115
rect 38845 17075 38855 17115
rect 38895 17075 38905 17115
rect 38945 17075 38955 17115
rect 38995 17075 39005 17115
rect 39045 17075 39055 17115
rect 39095 17075 39105 17115
rect 39145 17075 39155 17115
rect 39195 17075 39205 17115
rect 39245 17075 39255 17115
rect 39295 17075 39305 17115
rect 39345 17075 39355 17115
rect 39395 17075 39405 17115
rect 39445 17075 39455 17115
rect 39495 17075 39505 17115
rect 39545 17075 39555 17115
rect 39595 17075 39605 17115
rect 39645 17075 39655 17115
rect 39695 17075 39705 17115
rect 39745 17075 39750 17115
rect -2700 17070 39750 17075
rect -3500 17015 -50 17020
rect -3500 16975 -3495 17015
rect -3455 16975 -3295 17015
rect -3255 16975 -3095 17015
rect -3055 16975 -1595 17015
rect -1555 16975 -1195 17015
rect -1155 16975 -1095 17015
rect -1055 16975 -995 17015
rect -955 16975 -895 17015
rect -855 16975 -795 17015
rect -755 16975 -695 17015
rect -655 16975 -595 17015
rect -555 16975 -495 17015
rect -455 16975 -395 17015
rect -355 16975 -295 17015
rect -255 16975 -195 17015
rect -155 16975 -95 17015
rect -55 16975 -50 17015
rect -3500 16970 -50 16975
rect 0 17015 40900 17020
rect 0 16975 5 17015
rect 45 16975 55 17015
rect 95 16975 105 17015
rect 145 16975 155 17015
rect 195 16975 205 17015
rect 245 16975 255 17015
rect 295 16975 305 17015
rect 345 16975 355 17015
rect 395 16975 405 17015
rect 445 16975 455 17015
rect 495 16975 505 17015
rect 545 16975 555 17015
rect 595 16975 605 17015
rect 645 16975 655 17015
rect 695 16975 705 17015
rect 745 16975 755 17015
rect 795 16975 805 17015
rect 845 16975 855 17015
rect 895 16975 905 17015
rect 945 16975 955 17015
rect 995 16975 1005 17015
rect 1045 16975 1055 17015
rect 1095 16975 1105 17015
rect 1145 16975 1155 17015
rect 1195 16975 1205 17015
rect 1245 16975 1255 17015
rect 1295 16975 1305 17015
rect 1345 16975 1355 17015
rect 1395 16975 1405 17015
rect 1445 16975 1455 17015
rect 1495 16975 1505 17015
rect 1545 16975 1555 17015
rect 1595 16975 1605 17015
rect 1645 16975 1655 17015
rect 1695 16975 1705 17015
rect 1745 16975 1755 17015
rect 1795 16975 1805 17015
rect 1845 16975 1855 17015
rect 1895 16975 1905 17015
rect 1945 16975 1955 17015
rect 1995 16975 2005 17015
rect 2045 16975 2055 17015
rect 2095 16975 2105 17015
rect 2145 16975 2155 17015
rect 2195 16975 2205 17015
rect 2245 16975 2255 17015
rect 2295 16975 2305 17015
rect 2345 16975 2355 17015
rect 2395 16975 2405 17015
rect 2445 16975 2455 17015
rect 2495 16975 2505 17015
rect 2545 16975 2555 17015
rect 2595 16975 2605 17015
rect 2645 16975 2655 17015
rect 2695 16975 2705 17015
rect 2745 16975 2755 17015
rect 2795 16975 2805 17015
rect 2845 16975 2855 17015
rect 2895 16975 2905 17015
rect 2945 16975 2955 17015
rect 2995 16975 3005 17015
rect 3045 16975 3055 17015
rect 3095 16975 3105 17015
rect 3145 16975 3155 17015
rect 3195 16975 3205 17015
rect 3245 16975 3255 17015
rect 3295 16975 3305 17015
rect 3345 16975 3355 17015
rect 3395 16975 3405 17015
rect 3445 16975 3455 17015
rect 3495 16975 3505 17015
rect 3545 16975 3555 17015
rect 3595 16975 3605 17015
rect 3645 16975 3655 17015
rect 3695 16975 3705 17015
rect 3745 16975 3755 17015
rect 3795 16975 3805 17015
rect 3845 16975 3855 17015
rect 3895 16975 3905 17015
rect 3945 16975 3955 17015
rect 3995 16975 4005 17015
rect 4045 16975 4055 17015
rect 4095 16975 4105 17015
rect 4145 16975 4155 17015
rect 4195 16975 4205 17015
rect 4245 16975 4255 17015
rect 4295 16975 4305 17015
rect 4345 16975 4355 17015
rect 4395 16975 4405 17015
rect 4445 16975 4455 17015
rect 4495 16975 4505 17015
rect 4545 16975 4555 17015
rect 4595 16975 4605 17015
rect 4645 16975 4655 17015
rect 4695 16975 4705 17015
rect 4745 16975 4755 17015
rect 4795 16975 4805 17015
rect 4845 16975 4855 17015
rect 4895 16975 4905 17015
rect 4945 16975 4955 17015
rect 4995 16975 5005 17015
rect 5045 16975 5055 17015
rect 5095 16975 5105 17015
rect 5145 16975 5155 17015
rect 5195 16975 5205 17015
rect 5245 16975 5255 17015
rect 5295 16975 5305 17015
rect 5345 16975 5355 17015
rect 5395 16975 5405 17015
rect 5445 16975 5455 17015
rect 5495 16975 5505 17015
rect 5545 16975 5555 17015
rect 5595 16975 5605 17015
rect 5645 16975 5655 17015
rect 5695 16975 5705 17015
rect 5745 16975 5755 17015
rect 5795 16975 5805 17015
rect 5845 16975 5855 17015
rect 5895 16975 5905 17015
rect 5945 16975 5955 17015
rect 5995 16975 6005 17015
rect 6045 16975 6055 17015
rect 6095 16975 6105 17015
rect 6145 16975 6155 17015
rect 6195 16975 6205 17015
rect 6245 16975 6255 17015
rect 6295 16975 6305 17015
rect 6345 16975 6355 17015
rect 6395 16975 6405 17015
rect 6445 16975 6455 17015
rect 6495 16975 6505 17015
rect 6545 16975 6555 17015
rect 6595 16975 6605 17015
rect 6645 16975 6655 17015
rect 6695 16975 6705 17015
rect 6745 16975 6755 17015
rect 6795 16975 6805 17015
rect 6845 16975 6855 17015
rect 6895 16975 6905 17015
rect 6945 16975 6955 17015
rect 6995 16975 7005 17015
rect 7045 16975 7055 17015
rect 7095 16975 7105 17015
rect 7145 16975 7155 17015
rect 7195 16975 7205 17015
rect 7245 16975 7255 17015
rect 7295 16975 7305 17015
rect 7345 16975 7355 17015
rect 7395 16975 7405 17015
rect 7445 16975 7455 17015
rect 7495 16975 7505 17015
rect 7545 16975 7555 17015
rect 7595 16975 7605 17015
rect 7645 16975 7655 17015
rect 7695 16975 7705 17015
rect 7745 16975 7755 17015
rect 7795 16975 7805 17015
rect 7845 16975 7855 17015
rect 7895 16975 7905 17015
rect 7945 16975 7955 17015
rect 7995 16975 8005 17015
rect 8045 16975 8055 17015
rect 8095 16975 8105 17015
rect 8145 16975 8155 17015
rect 8195 16975 8205 17015
rect 8245 16975 8255 17015
rect 8295 16975 8305 17015
rect 8345 16975 8355 17015
rect 8395 16975 8405 17015
rect 8445 16975 8455 17015
rect 8495 16975 8505 17015
rect 8545 16975 8555 17015
rect 8595 16975 8605 17015
rect 8645 16975 8655 17015
rect 8695 16975 8705 17015
rect 8745 16975 8755 17015
rect 8795 16975 8805 17015
rect 8845 16975 8855 17015
rect 8895 16975 8905 17015
rect 8945 16975 8955 17015
rect 8995 16975 9005 17015
rect 9045 16975 9055 17015
rect 9095 16975 9105 17015
rect 9145 16975 9155 17015
rect 9195 16975 9205 17015
rect 9245 16975 9255 17015
rect 9295 16975 9305 17015
rect 9345 16975 9355 17015
rect 9395 16975 9405 17015
rect 9445 16975 9455 17015
rect 9495 16975 9505 17015
rect 9545 16975 9555 17015
rect 9595 16975 9605 17015
rect 9645 16975 9655 17015
rect 9695 16975 9705 17015
rect 9745 16975 9755 17015
rect 9795 16975 9805 17015
rect 9845 16975 9855 17015
rect 9895 16975 9905 17015
rect 9945 16975 9955 17015
rect 9995 16975 10005 17015
rect 10045 16975 10055 17015
rect 10095 16975 10105 17015
rect 10145 16975 10155 17015
rect 10195 16975 10205 17015
rect 10245 16975 10255 17015
rect 10295 16975 10305 17015
rect 10345 16975 10355 17015
rect 10395 16975 10405 17015
rect 10445 16975 10455 17015
rect 10495 16975 10505 17015
rect 10545 16975 10555 17015
rect 10595 16975 10605 17015
rect 10645 16975 10655 17015
rect 10695 16975 10705 17015
rect 10745 16975 10755 17015
rect 10795 16975 10805 17015
rect 10845 16975 10855 17015
rect 10895 16975 10905 17015
rect 10945 16975 10955 17015
rect 10995 16975 11005 17015
rect 11045 16975 11055 17015
rect 11095 16975 11105 17015
rect 11145 16975 11155 17015
rect 11195 16975 11205 17015
rect 11245 16975 11255 17015
rect 11295 16975 11305 17015
rect 11345 16975 11355 17015
rect 11395 16975 11405 17015
rect 11445 16975 11455 17015
rect 11495 16975 11505 17015
rect 11545 16975 11555 17015
rect 11595 16975 11605 17015
rect 11645 16975 11655 17015
rect 11695 16975 11705 17015
rect 11745 16975 11755 17015
rect 11795 16975 11805 17015
rect 11845 16975 11855 17015
rect 11895 16975 11905 17015
rect 11945 16975 11955 17015
rect 11995 16975 12005 17015
rect 12045 16975 12055 17015
rect 12095 16975 12105 17015
rect 12145 16975 12155 17015
rect 12195 16975 12205 17015
rect 12245 16975 12255 17015
rect 12295 16975 12305 17015
rect 12345 16975 12355 17015
rect 12395 16975 12405 17015
rect 12445 16975 12455 17015
rect 12495 16975 12505 17015
rect 12545 16975 12555 17015
rect 12595 16975 12605 17015
rect 12645 16975 12655 17015
rect 12695 16975 12705 17015
rect 12745 16975 12755 17015
rect 12795 16975 12805 17015
rect 12845 16975 12855 17015
rect 12895 16975 12905 17015
rect 12945 16975 12955 17015
rect 12995 16975 13005 17015
rect 13045 16975 13055 17015
rect 13095 16975 13105 17015
rect 13145 16975 13155 17015
rect 13195 16975 13205 17015
rect 13245 16975 13255 17015
rect 13295 16975 13305 17015
rect 13345 16975 13355 17015
rect 13395 16975 13405 17015
rect 13445 16975 13455 17015
rect 13495 16975 13505 17015
rect 13545 16975 13555 17015
rect 13595 16975 13605 17015
rect 13645 16975 13655 17015
rect 13695 16975 13705 17015
rect 13745 16975 13755 17015
rect 13795 16975 13805 17015
rect 13845 16975 13855 17015
rect 13895 16975 13905 17015
rect 13945 16975 13955 17015
rect 13995 16975 14005 17015
rect 14045 16975 14055 17015
rect 14095 16975 14105 17015
rect 14145 16975 14155 17015
rect 14195 16975 14205 17015
rect 14245 16975 14255 17015
rect 14295 16975 14305 17015
rect 14345 16975 14355 17015
rect 14395 16975 14405 17015
rect 14445 16975 14455 17015
rect 14495 16975 14505 17015
rect 14545 16975 14555 17015
rect 14595 16975 14605 17015
rect 14645 16975 14655 17015
rect 14695 16975 14705 17015
rect 14745 16975 14755 17015
rect 14795 16975 14805 17015
rect 14845 16975 14855 17015
rect 14895 16975 14905 17015
rect 14945 16975 14955 17015
rect 14995 16975 15005 17015
rect 15045 16975 15055 17015
rect 15095 16975 15105 17015
rect 15145 16975 15155 17015
rect 15195 16975 15205 17015
rect 15245 16975 15255 17015
rect 15295 16975 15305 17015
rect 15345 16975 15355 17015
rect 15395 16975 15405 17015
rect 15445 16975 15455 17015
rect 15495 16975 15505 17015
rect 15545 16975 15555 17015
rect 15595 16975 15605 17015
rect 15645 16975 15655 17015
rect 15695 16975 15705 17015
rect 15745 16975 15755 17015
rect 15795 16975 15805 17015
rect 15845 16975 15855 17015
rect 15895 16975 15905 17015
rect 15945 16975 15955 17015
rect 15995 16975 16005 17015
rect 16045 16975 16055 17015
rect 16095 16975 16105 17015
rect 16145 16975 16155 17015
rect 16195 16975 16205 17015
rect 16245 16975 16255 17015
rect 16295 16975 16305 17015
rect 16345 16975 16355 17015
rect 16395 16975 16405 17015
rect 16445 16975 16455 17015
rect 16495 16975 16505 17015
rect 16545 16975 16555 17015
rect 16595 16975 16605 17015
rect 16645 16975 16655 17015
rect 16695 16975 16705 17015
rect 16745 16975 16755 17015
rect 16795 16975 16805 17015
rect 16845 16975 16855 17015
rect 16895 16975 16905 17015
rect 16945 16975 16955 17015
rect 16995 16975 17005 17015
rect 17045 16975 17055 17015
rect 17095 16975 17105 17015
rect 17145 16975 17155 17015
rect 17195 16975 17205 17015
rect 17245 16975 17255 17015
rect 17295 16975 17305 17015
rect 17345 16975 17355 17015
rect 17395 16975 17405 17015
rect 17445 16975 17455 17015
rect 17495 16975 17505 17015
rect 17545 16975 17555 17015
rect 17595 16975 17605 17015
rect 17645 16975 17655 17015
rect 17695 16975 17705 17015
rect 17745 16975 17755 17015
rect 17795 16975 17805 17015
rect 17845 16975 17855 17015
rect 17895 16975 17905 17015
rect 17945 16975 17955 17015
rect 17995 16975 18005 17015
rect 18045 16975 18055 17015
rect 18095 16975 18105 17015
rect 18145 16975 18155 17015
rect 18195 16975 18205 17015
rect 18245 16975 18255 17015
rect 18295 16975 18305 17015
rect 18345 16975 18355 17015
rect 18395 16975 18405 17015
rect 18445 16975 18455 17015
rect 18495 16975 18505 17015
rect 18545 16975 18555 17015
rect 18595 16975 18605 17015
rect 18645 16975 18655 17015
rect 18695 16975 18705 17015
rect 18745 16975 18755 17015
rect 18795 16975 18805 17015
rect 18845 16975 18855 17015
rect 18895 16975 18905 17015
rect 18945 16975 18955 17015
rect 18995 16975 19005 17015
rect 19045 16975 19055 17015
rect 19095 16975 19105 17015
rect 19145 16975 19155 17015
rect 19195 16975 19205 17015
rect 19245 16975 19255 17015
rect 19295 16975 19305 17015
rect 19345 16975 19355 17015
rect 19395 16975 19405 17015
rect 19445 16975 19455 17015
rect 19495 16975 19505 17015
rect 19545 16975 19555 17015
rect 19595 16975 19605 17015
rect 19645 16975 19655 17015
rect 19695 16975 19705 17015
rect 19745 16975 19755 17015
rect 19795 16975 19805 17015
rect 19845 16975 19855 17015
rect 19895 16975 19905 17015
rect 19945 16975 19955 17015
rect 19995 16975 20005 17015
rect 20045 16975 20055 17015
rect 20095 16975 20105 17015
rect 20145 16975 20155 17015
rect 20195 16975 20205 17015
rect 20245 16975 20255 17015
rect 20295 16975 20305 17015
rect 20345 16975 20355 17015
rect 20395 16975 20405 17015
rect 20445 16975 20455 17015
rect 20495 16975 20505 17015
rect 20545 16975 20555 17015
rect 20595 16975 20605 17015
rect 20645 16975 20655 17015
rect 20695 16975 20705 17015
rect 20745 16975 20755 17015
rect 20795 16975 20805 17015
rect 20845 16975 20855 17015
rect 20895 16975 20905 17015
rect 20945 16975 20955 17015
rect 20995 16975 21005 17015
rect 21045 16975 21055 17015
rect 21095 16975 21105 17015
rect 21145 16975 21155 17015
rect 21195 16975 21205 17015
rect 21245 16975 21255 17015
rect 21295 16975 21305 17015
rect 21345 16975 21355 17015
rect 21395 16975 21405 17015
rect 21445 16975 21455 17015
rect 21495 16975 21505 17015
rect 21545 16975 21555 17015
rect 21595 16975 21605 17015
rect 21645 16975 21655 17015
rect 21695 16975 21705 17015
rect 21745 16975 21755 17015
rect 21795 16975 21805 17015
rect 21845 16975 21855 17015
rect 21895 16975 21905 17015
rect 21945 16975 21955 17015
rect 21995 16975 22005 17015
rect 22045 16975 22055 17015
rect 22095 16975 22105 17015
rect 22145 16975 22155 17015
rect 22195 16975 22205 17015
rect 22245 16975 22255 17015
rect 22295 16975 22305 17015
rect 22345 16975 22355 17015
rect 22395 16975 22405 17015
rect 22445 16975 22455 17015
rect 22495 16975 22505 17015
rect 22545 16975 22555 17015
rect 22595 16975 22605 17015
rect 22645 16975 22655 17015
rect 22695 16975 22705 17015
rect 22745 16975 22755 17015
rect 22795 16975 22805 17015
rect 22845 16975 22855 17015
rect 22895 16975 22905 17015
rect 22945 16975 22955 17015
rect 22995 16975 23005 17015
rect 23045 16975 23055 17015
rect 23095 16975 23105 17015
rect 23145 16975 23155 17015
rect 23195 16975 23205 17015
rect 23245 16975 23255 17015
rect 23295 16975 23305 17015
rect 23345 16975 23355 17015
rect 23395 16975 23405 17015
rect 23445 16975 23455 17015
rect 23495 16975 23505 17015
rect 23545 16975 23555 17015
rect 23595 16975 23605 17015
rect 23645 16975 23655 17015
rect 23695 16975 23705 17015
rect 23745 16975 23755 17015
rect 23795 16975 23805 17015
rect 23845 16975 23855 17015
rect 23895 16975 23905 17015
rect 23945 16975 23955 17015
rect 23995 16975 24005 17015
rect 24045 16975 24055 17015
rect 24095 16975 24105 17015
rect 24145 16975 24155 17015
rect 24195 16975 24205 17015
rect 24245 16975 24255 17015
rect 24295 16975 24305 17015
rect 24345 16975 24355 17015
rect 24395 16975 24405 17015
rect 24445 16975 24455 17015
rect 24495 16975 24505 17015
rect 24545 16975 24555 17015
rect 24595 16975 24605 17015
rect 24645 16975 24655 17015
rect 24695 16975 24705 17015
rect 24745 16975 24755 17015
rect 24795 16975 24805 17015
rect 24845 16975 24855 17015
rect 24895 16975 24905 17015
rect 24945 16975 24955 17015
rect 24995 16975 25005 17015
rect 25045 16975 25055 17015
rect 25095 16975 25105 17015
rect 25145 16975 25155 17015
rect 25195 16975 25205 17015
rect 25245 16975 25255 17015
rect 25295 16975 25305 17015
rect 25345 16975 25355 17015
rect 25395 16975 25405 17015
rect 25445 16975 25455 17015
rect 25495 16975 25505 17015
rect 25545 16975 25555 17015
rect 25595 16975 25605 17015
rect 25645 16975 25655 17015
rect 25695 16975 25705 17015
rect 25745 16975 25755 17015
rect 25795 16975 25805 17015
rect 25845 16975 25855 17015
rect 25895 16975 25905 17015
rect 25945 16975 25955 17015
rect 25995 16975 26005 17015
rect 26045 16975 26055 17015
rect 26095 16975 26105 17015
rect 26145 16975 26155 17015
rect 26195 16975 26205 17015
rect 26245 16975 26255 17015
rect 26295 16975 26305 17015
rect 26345 16975 26355 17015
rect 26395 16975 26405 17015
rect 26445 16975 26455 17015
rect 26495 16975 26505 17015
rect 26545 16975 26555 17015
rect 26595 16975 26605 17015
rect 26645 16975 26655 17015
rect 26695 16975 26705 17015
rect 26745 16975 26755 17015
rect 26795 16975 26805 17015
rect 26845 16975 26855 17015
rect 26895 16975 26905 17015
rect 26945 16975 26955 17015
rect 26995 16975 27005 17015
rect 27045 16975 27055 17015
rect 27095 16975 27105 17015
rect 27145 16975 27155 17015
rect 27195 16975 27205 17015
rect 27245 16975 27255 17015
rect 27295 16975 27305 17015
rect 27345 16975 27355 17015
rect 27395 16975 27405 17015
rect 27445 16975 27455 17015
rect 27495 16975 27505 17015
rect 27545 16975 27555 17015
rect 27595 16975 27605 17015
rect 27645 16975 27655 17015
rect 27695 16975 27705 17015
rect 27745 16975 27755 17015
rect 27795 16975 27805 17015
rect 27845 16975 27855 17015
rect 27895 16975 27905 17015
rect 27945 16975 27955 17015
rect 27995 16975 28005 17015
rect 28045 16975 28055 17015
rect 28095 16975 28105 17015
rect 28145 16975 28155 17015
rect 28195 16975 28205 17015
rect 28245 16975 28255 17015
rect 28295 16975 28305 17015
rect 28345 16975 28355 17015
rect 28395 16975 28405 17015
rect 28445 16975 28455 17015
rect 28495 16975 28505 17015
rect 28545 16975 28555 17015
rect 28595 16975 28605 17015
rect 28645 16975 28655 17015
rect 28695 16975 28705 17015
rect 28745 16975 28755 17015
rect 28795 16975 28805 17015
rect 28845 16975 28855 17015
rect 28895 16975 28905 17015
rect 28945 16975 28955 17015
rect 28995 16975 29005 17015
rect 29045 16975 29055 17015
rect 29095 16975 29105 17015
rect 29145 16975 29155 17015
rect 29195 16975 29205 17015
rect 29245 16975 29255 17015
rect 29295 16975 29305 17015
rect 29345 16975 29355 17015
rect 29395 16975 29405 17015
rect 29445 16975 29455 17015
rect 29495 16975 29505 17015
rect 29545 16975 29555 17015
rect 29595 16975 29605 17015
rect 29645 16975 29655 17015
rect 29695 16975 29705 17015
rect 29745 16975 29755 17015
rect 29795 16975 29805 17015
rect 29845 16975 29855 17015
rect 29895 16975 29905 17015
rect 29945 16975 29955 17015
rect 29995 16975 30005 17015
rect 30045 16975 30055 17015
rect 30095 16975 30105 17015
rect 30145 16975 30155 17015
rect 30195 16975 30205 17015
rect 30245 16975 30255 17015
rect 30295 16975 30305 17015
rect 30345 16975 30355 17015
rect 30395 16975 30405 17015
rect 30445 16975 30455 17015
rect 30495 16975 30505 17015
rect 30545 16975 30555 17015
rect 30595 16975 30605 17015
rect 30645 16975 30655 17015
rect 30695 16975 30705 17015
rect 30745 16975 30755 17015
rect 30795 16975 30805 17015
rect 30845 16975 30855 17015
rect 30895 16975 30905 17015
rect 30945 16975 30955 17015
rect 30995 16975 31005 17015
rect 31045 16975 31055 17015
rect 31095 16975 31105 17015
rect 31145 16975 31155 17015
rect 31195 16975 31205 17015
rect 31245 16975 31255 17015
rect 31295 16975 31305 17015
rect 31345 16975 31355 17015
rect 31395 16975 31405 17015
rect 31445 16975 31455 17015
rect 31495 16975 31505 17015
rect 31545 16975 31555 17015
rect 31595 16975 31605 17015
rect 31645 16975 31655 17015
rect 31695 16975 31705 17015
rect 31745 16975 31755 17015
rect 31795 16975 31805 17015
rect 31845 16975 31855 17015
rect 31895 16975 31905 17015
rect 31945 16975 31955 17015
rect 31995 16975 32005 17015
rect 32045 16975 32055 17015
rect 32095 16975 32105 17015
rect 32145 16975 32155 17015
rect 32195 16975 32205 17015
rect 32245 16975 32255 17015
rect 32295 16975 32305 17015
rect 32345 16975 32355 17015
rect 32395 16975 32405 17015
rect 32445 16975 32455 17015
rect 32495 16975 32505 17015
rect 32545 16975 32555 17015
rect 32595 16975 32605 17015
rect 32645 16975 32655 17015
rect 32695 16975 32705 17015
rect 32745 16975 32755 17015
rect 32795 16975 32805 17015
rect 32845 16975 32855 17015
rect 32895 16975 32905 17015
rect 32945 16975 32955 17015
rect 32995 16975 33005 17015
rect 33045 16975 33055 17015
rect 33095 16975 33105 17015
rect 33145 16975 33155 17015
rect 33195 16975 33205 17015
rect 33245 16975 33255 17015
rect 33295 16975 33305 17015
rect 33345 16975 33355 17015
rect 33395 16975 33405 17015
rect 33445 16975 33455 17015
rect 33495 16975 33505 17015
rect 33545 16975 33555 17015
rect 33595 16975 33605 17015
rect 33645 16975 33655 17015
rect 33695 16975 33705 17015
rect 33745 16975 33755 17015
rect 33795 16975 33805 17015
rect 33845 16975 33855 17015
rect 33895 16975 33905 17015
rect 33945 16975 33955 17015
rect 33995 16975 34005 17015
rect 34045 16975 34055 17015
rect 34095 16975 34105 17015
rect 34145 16975 34155 17015
rect 34195 16975 34205 17015
rect 34245 16975 34255 17015
rect 34295 16975 34305 17015
rect 34345 16975 34355 17015
rect 34395 16975 34405 17015
rect 34445 16975 34455 17015
rect 34495 16975 34505 17015
rect 34545 16975 34555 17015
rect 34595 16975 34605 17015
rect 34645 16975 34655 17015
rect 34695 16975 34705 17015
rect 34745 16975 34755 17015
rect 34795 16975 34805 17015
rect 34845 16975 34855 17015
rect 34895 16975 34905 17015
rect 34945 16975 34955 17015
rect 34995 16975 35005 17015
rect 35045 16975 35055 17015
rect 35095 16975 35105 17015
rect 35145 16975 35155 17015
rect 35195 16975 35205 17015
rect 35245 16975 35255 17015
rect 35295 16975 35305 17015
rect 35345 16975 35355 17015
rect 35395 16975 35405 17015
rect 35445 16975 35455 17015
rect 35495 16975 35505 17015
rect 35545 16975 35555 17015
rect 35595 16975 35605 17015
rect 35645 16975 35655 17015
rect 35695 16975 35705 17015
rect 35745 16975 35755 17015
rect 35795 16975 35805 17015
rect 35845 16975 35855 17015
rect 35895 16975 35905 17015
rect 35945 16975 35955 17015
rect 35995 16975 36005 17015
rect 36045 16975 36055 17015
rect 36095 16975 36105 17015
rect 36145 16975 36155 17015
rect 36195 16975 36205 17015
rect 36245 16975 36255 17015
rect 36295 16975 36305 17015
rect 36345 16975 36355 17015
rect 36395 16975 36405 17015
rect 36445 16975 36455 17015
rect 36495 16975 36505 17015
rect 36545 16975 36555 17015
rect 36595 16975 36605 17015
rect 36645 16975 36655 17015
rect 36695 16975 36705 17015
rect 36745 16975 36755 17015
rect 36795 16975 36805 17015
rect 36845 16975 36855 17015
rect 36895 16975 36905 17015
rect 36945 16975 36955 17015
rect 36995 16975 37005 17015
rect 37045 16975 37055 17015
rect 37095 16975 37105 17015
rect 37145 16975 37155 17015
rect 37195 16975 37205 17015
rect 37245 16975 37255 17015
rect 37295 16975 37305 17015
rect 37345 16975 37355 17015
rect 37395 16975 37405 17015
rect 37445 16975 37455 17015
rect 37495 16975 37505 17015
rect 37545 16975 37555 17015
rect 37595 16975 37605 17015
rect 37645 16975 37655 17015
rect 37695 16975 37705 17015
rect 37745 16975 37755 17015
rect 37795 16975 37805 17015
rect 37845 16975 37855 17015
rect 37895 16975 37905 17015
rect 37945 16975 37955 17015
rect 37995 16975 38005 17015
rect 38045 16975 38055 17015
rect 38095 16975 38105 17015
rect 38145 16975 38155 17015
rect 38195 16975 38205 17015
rect 38245 16975 38255 17015
rect 38295 16975 38305 17015
rect 38345 16975 38355 17015
rect 38395 16975 38405 17015
rect 38445 16975 38455 17015
rect 38495 16975 38505 17015
rect 38545 16975 38555 17015
rect 38595 16975 38605 17015
rect 38645 16975 38655 17015
rect 38695 16975 38705 17015
rect 38745 16975 38755 17015
rect 38795 16975 38805 17015
rect 38845 16975 38855 17015
rect 38895 16975 38905 17015
rect 38945 16975 38955 17015
rect 38995 16975 39005 17015
rect 39045 16975 39055 17015
rect 39095 16975 39105 17015
rect 39145 16975 39155 17015
rect 39195 16975 39205 17015
rect 39245 16975 39255 17015
rect 39295 16975 39305 17015
rect 39345 16975 39355 17015
rect 39395 16975 39405 17015
rect 39445 16975 39455 17015
rect 39495 16975 39505 17015
rect 39545 16975 39555 17015
rect 39595 16975 39605 17015
rect 39645 16975 39655 17015
rect 39695 16975 39705 17015
rect 39745 16975 39905 17015
rect 39945 16975 39955 17015
rect 39995 16975 40005 17015
rect 40045 16975 40055 17015
rect 40095 16975 40105 17015
rect 40145 16975 40155 17015
rect 40195 16975 40205 17015
rect 40245 16975 40255 17015
rect 40295 16975 40305 17015
rect 40345 16975 40355 17015
rect 40395 16975 40405 17015
rect 40445 16975 40455 17015
rect 40495 16975 40505 17015
rect 40545 16975 40555 17015
rect 40595 16975 40605 17015
rect 40645 16975 40655 17015
rect 40695 16975 40705 17015
rect 40745 16975 40755 17015
rect 40795 16975 40805 17015
rect 40845 16975 40855 17015
rect 40895 16975 40900 17015
rect 0 16970 40900 16975
rect -400 16915 39750 16920
rect -400 16875 -395 16915
rect -355 16875 105 16915
rect 145 16875 155 16915
rect 195 16875 205 16915
rect 245 16875 255 16915
rect 295 16875 305 16915
rect 345 16875 355 16915
rect 395 16875 405 16915
rect 445 16875 455 16915
rect 495 16875 505 16915
rect 545 16875 555 16915
rect 595 16875 605 16915
rect 645 16875 655 16915
rect 695 16875 705 16915
rect 745 16875 755 16915
rect 795 16875 805 16915
rect 845 16875 855 16915
rect 895 16875 905 16915
rect 945 16875 955 16915
rect 995 16875 1005 16915
rect 1045 16875 1055 16915
rect 1095 16875 1105 16915
rect 1145 16875 1155 16915
rect 1195 16875 1205 16915
rect 1245 16875 1255 16915
rect 1295 16875 1305 16915
rect 1345 16875 1355 16915
rect 1395 16875 1405 16915
rect 1445 16875 1455 16915
rect 1495 16875 1505 16915
rect 1545 16875 1555 16915
rect 1595 16875 1605 16915
rect 1645 16875 1655 16915
rect 1695 16875 1705 16915
rect 1745 16875 1755 16915
rect 1795 16875 1805 16915
rect 1845 16875 1855 16915
rect 1895 16875 1905 16915
rect 1945 16875 1955 16915
rect 1995 16875 2005 16915
rect 2045 16875 2055 16915
rect 2095 16875 2105 16915
rect 2145 16875 2155 16915
rect 2195 16875 2205 16915
rect 2245 16875 2255 16915
rect 2295 16875 2305 16915
rect 2345 16875 2355 16915
rect 2395 16875 2405 16915
rect 2445 16875 2455 16915
rect 2495 16875 2505 16915
rect 2545 16875 2555 16915
rect 2595 16875 2605 16915
rect 2645 16875 2655 16915
rect 2695 16875 2705 16915
rect 2745 16875 2755 16915
rect 2795 16875 2805 16915
rect 2845 16875 2855 16915
rect 2895 16875 2905 16915
rect 2945 16875 2955 16915
rect 2995 16875 3005 16915
rect 3045 16875 3055 16915
rect 3095 16875 3105 16915
rect 3145 16875 3155 16915
rect 3195 16875 3205 16915
rect 3245 16875 3255 16915
rect 3295 16875 3305 16915
rect 3345 16875 3355 16915
rect 3395 16875 3405 16915
rect 3445 16875 3455 16915
rect 3495 16875 3505 16915
rect 3545 16875 3555 16915
rect 3595 16875 3605 16915
rect 3645 16875 3655 16915
rect 3695 16875 3705 16915
rect 3745 16875 3755 16915
rect 3795 16875 3805 16915
rect 3845 16875 3855 16915
rect 3895 16875 3905 16915
rect 3945 16875 3955 16915
rect 3995 16875 4005 16915
rect 4045 16875 4055 16915
rect 4095 16875 4105 16915
rect 4145 16875 4155 16915
rect 4195 16875 4205 16915
rect 4245 16875 4255 16915
rect 4295 16875 4305 16915
rect 4345 16875 4355 16915
rect 4395 16875 4405 16915
rect 4445 16875 4455 16915
rect 4495 16875 4505 16915
rect 4545 16875 4555 16915
rect 4595 16875 4605 16915
rect 4645 16875 4655 16915
rect 4695 16875 4705 16915
rect 4745 16875 4755 16915
rect 4795 16875 4805 16915
rect 4845 16875 4855 16915
rect 4895 16875 4905 16915
rect 4945 16875 4955 16915
rect 4995 16875 5005 16915
rect 5045 16875 5055 16915
rect 5095 16875 5105 16915
rect 5145 16875 5155 16915
rect 5195 16875 5205 16915
rect 5245 16875 5255 16915
rect 5295 16875 5305 16915
rect 5345 16875 5355 16915
rect 5395 16875 5405 16915
rect 5445 16875 5455 16915
rect 5495 16875 5505 16915
rect 5545 16875 5555 16915
rect 5595 16875 5605 16915
rect 5645 16875 5655 16915
rect 5695 16875 5705 16915
rect 5745 16875 5755 16915
rect 5795 16875 5805 16915
rect 5845 16875 5855 16915
rect 5895 16875 5905 16915
rect 5945 16875 5955 16915
rect 5995 16875 6005 16915
rect 6045 16875 6055 16915
rect 6095 16875 6105 16915
rect 6145 16875 6155 16915
rect 6195 16875 6205 16915
rect 6245 16875 6255 16915
rect 6295 16875 6305 16915
rect 6345 16875 6355 16915
rect 6395 16875 6405 16915
rect 6445 16875 6455 16915
rect 6495 16875 6505 16915
rect 6545 16875 6555 16915
rect 6595 16875 6605 16915
rect 6645 16875 6655 16915
rect 6695 16875 6705 16915
rect 6745 16875 6755 16915
rect 6795 16875 6805 16915
rect 6845 16875 6855 16915
rect 6895 16875 6905 16915
rect 6945 16875 6955 16915
rect 6995 16875 7005 16915
rect 7045 16875 7055 16915
rect 7095 16875 7105 16915
rect 7145 16875 7155 16915
rect 7195 16875 7205 16915
rect 7245 16875 7255 16915
rect 7295 16875 7305 16915
rect 7345 16875 7355 16915
rect 7395 16875 7405 16915
rect 7445 16875 7455 16915
rect 7495 16875 7505 16915
rect 7545 16875 7555 16915
rect 7595 16875 7605 16915
rect 7645 16875 7655 16915
rect 7695 16875 7705 16915
rect 7745 16875 7755 16915
rect 7795 16875 7805 16915
rect 7845 16875 7855 16915
rect 7895 16875 7905 16915
rect 7945 16875 7955 16915
rect 7995 16875 8005 16915
rect 8045 16875 8055 16915
rect 8095 16875 8105 16915
rect 8145 16875 8155 16915
rect 8195 16875 8205 16915
rect 8245 16875 8255 16915
rect 8295 16875 8305 16915
rect 8345 16875 8355 16915
rect 8395 16875 8405 16915
rect 8445 16875 8455 16915
rect 8495 16875 8505 16915
rect 8545 16875 8555 16915
rect 8595 16875 8605 16915
rect 8645 16875 8655 16915
rect 8695 16875 8705 16915
rect 8745 16875 8755 16915
rect 8795 16875 8805 16915
rect 8845 16875 8855 16915
rect 8895 16875 8905 16915
rect 8945 16875 8955 16915
rect 8995 16875 9005 16915
rect 9045 16875 9055 16915
rect 9095 16875 9105 16915
rect 9145 16875 9155 16915
rect 9195 16875 9205 16915
rect 9245 16875 9255 16915
rect 9295 16875 9305 16915
rect 9345 16875 9355 16915
rect 9395 16875 9405 16915
rect 9445 16875 9455 16915
rect 9495 16875 9505 16915
rect 9545 16875 9555 16915
rect 9595 16875 9605 16915
rect 9645 16875 9655 16915
rect 9695 16875 9705 16915
rect 9745 16875 9755 16915
rect 9795 16875 9805 16915
rect 9845 16875 9855 16915
rect 9895 16875 9905 16915
rect 9945 16875 9955 16915
rect 9995 16875 10005 16915
rect 10045 16875 10055 16915
rect 10095 16875 10105 16915
rect 10145 16875 10155 16915
rect 10195 16875 10205 16915
rect 10245 16875 10255 16915
rect 10295 16875 10305 16915
rect 10345 16875 10355 16915
rect 10395 16875 10405 16915
rect 10445 16875 10455 16915
rect 10495 16875 10505 16915
rect 10545 16875 10555 16915
rect 10595 16875 10605 16915
rect 10645 16875 10655 16915
rect 10695 16875 10705 16915
rect 10745 16875 10755 16915
rect 10795 16875 10805 16915
rect 10845 16875 10855 16915
rect 10895 16875 10905 16915
rect 10945 16875 10955 16915
rect 10995 16875 11005 16915
rect 11045 16875 11055 16915
rect 11095 16875 11105 16915
rect 11145 16875 11155 16915
rect 11195 16875 11205 16915
rect 11245 16875 11255 16915
rect 11295 16875 11305 16915
rect 11345 16875 11355 16915
rect 11395 16875 11405 16915
rect 11445 16875 11455 16915
rect 11495 16875 11505 16915
rect 11545 16875 11555 16915
rect 11595 16875 11605 16915
rect 11645 16875 11655 16915
rect 11695 16875 11705 16915
rect 11745 16875 11755 16915
rect 11795 16875 11805 16915
rect 11845 16875 11855 16915
rect 11895 16875 11905 16915
rect 11945 16875 11955 16915
rect 11995 16875 12005 16915
rect 12045 16875 12055 16915
rect 12095 16875 12105 16915
rect 12145 16875 12155 16915
rect 12195 16875 12205 16915
rect 12245 16875 12255 16915
rect 12295 16875 12305 16915
rect 12345 16875 12355 16915
rect 12395 16875 12405 16915
rect 12445 16875 12455 16915
rect 12495 16875 12505 16915
rect 12545 16875 12555 16915
rect 12595 16875 12605 16915
rect 12645 16875 12655 16915
rect 12695 16875 12705 16915
rect 12745 16875 12755 16915
rect 12795 16875 12805 16915
rect 12845 16875 12855 16915
rect 12895 16875 12905 16915
rect 12945 16875 12955 16915
rect 12995 16875 13005 16915
rect 13045 16875 13055 16915
rect 13095 16875 13105 16915
rect 13145 16875 13155 16915
rect 13195 16875 13205 16915
rect 13245 16875 13255 16915
rect 13295 16875 13305 16915
rect 13345 16875 13355 16915
rect 13395 16875 13405 16915
rect 13445 16875 13455 16915
rect 13495 16875 13505 16915
rect 13545 16875 13555 16915
rect 13595 16875 13605 16915
rect 13645 16875 13655 16915
rect 13695 16875 13705 16915
rect 13745 16875 13755 16915
rect 13795 16875 13805 16915
rect 13845 16875 13855 16915
rect 13895 16875 13905 16915
rect 13945 16875 13955 16915
rect 13995 16875 14005 16915
rect 14045 16875 14055 16915
rect 14095 16875 14105 16915
rect 14145 16875 14155 16915
rect 14195 16875 14205 16915
rect 14245 16875 14255 16915
rect 14295 16875 14305 16915
rect 14345 16875 14355 16915
rect 14395 16875 14405 16915
rect 14445 16875 14455 16915
rect 14495 16875 14505 16915
rect 14545 16875 14555 16915
rect 14595 16875 14605 16915
rect 14645 16875 14655 16915
rect 14695 16875 14705 16915
rect 14745 16875 14755 16915
rect 14795 16875 14805 16915
rect 14845 16875 14855 16915
rect 14895 16875 14905 16915
rect 14945 16875 14955 16915
rect 14995 16875 15005 16915
rect 15045 16875 15055 16915
rect 15095 16875 15105 16915
rect 15145 16875 15155 16915
rect 15195 16875 15205 16915
rect 15245 16875 15255 16915
rect 15295 16875 15305 16915
rect 15345 16875 15355 16915
rect 15395 16875 15405 16915
rect 15445 16875 15455 16915
rect 15495 16875 15505 16915
rect 15545 16875 15555 16915
rect 15595 16875 15605 16915
rect 15645 16875 15655 16915
rect 15695 16875 15705 16915
rect 15745 16875 15755 16915
rect 15795 16875 15805 16915
rect 15845 16875 15855 16915
rect 15895 16875 15905 16915
rect 15945 16875 15955 16915
rect 15995 16875 16005 16915
rect 16045 16875 16055 16915
rect 16095 16875 16105 16915
rect 16145 16875 16155 16915
rect 16195 16875 16205 16915
rect 16245 16875 16255 16915
rect 16295 16875 16305 16915
rect 16345 16875 16355 16915
rect 16395 16875 16405 16915
rect 16445 16875 16455 16915
rect 16495 16875 16505 16915
rect 16545 16875 16555 16915
rect 16595 16875 16605 16915
rect 16645 16875 16655 16915
rect 16695 16875 16705 16915
rect 16745 16875 16755 16915
rect 16795 16875 16805 16915
rect 16845 16875 16855 16915
rect 16895 16875 16905 16915
rect 16945 16875 16955 16915
rect 16995 16875 17005 16915
rect 17045 16875 17055 16915
rect 17095 16875 17105 16915
rect 17145 16875 17155 16915
rect 17195 16875 17205 16915
rect 17245 16875 17255 16915
rect 17295 16875 17305 16915
rect 17345 16875 17355 16915
rect 17395 16875 17405 16915
rect 17445 16875 17455 16915
rect 17495 16875 17505 16915
rect 17545 16875 17555 16915
rect 17595 16875 17605 16915
rect 17645 16875 17655 16915
rect 17695 16875 17705 16915
rect 17745 16875 17755 16915
rect 17795 16875 17805 16915
rect 17845 16875 17855 16915
rect 17895 16875 17905 16915
rect 17945 16875 17955 16915
rect 17995 16875 18005 16915
rect 18045 16875 18055 16915
rect 18095 16875 18105 16915
rect 18145 16875 18155 16915
rect 18195 16875 18205 16915
rect 18245 16875 18255 16915
rect 18295 16875 18305 16915
rect 18345 16875 18355 16915
rect 18395 16875 18405 16915
rect 18445 16875 18455 16915
rect 18495 16875 18505 16915
rect 18545 16875 18555 16915
rect 18595 16875 18605 16915
rect 18645 16875 18655 16915
rect 18695 16875 18705 16915
rect 18745 16875 18755 16915
rect 18795 16875 18805 16915
rect 18845 16875 18855 16915
rect 18895 16875 18905 16915
rect 18945 16875 18955 16915
rect 18995 16875 19005 16915
rect 19045 16875 19055 16915
rect 19095 16875 19105 16915
rect 19145 16875 19155 16915
rect 19195 16875 19205 16915
rect 19245 16875 19255 16915
rect 19295 16875 19305 16915
rect 19345 16875 19355 16915
rect 19395 16875 19405 16915
rect 19445 16875 19455 16915
rect 19495 16875 19505 16915
rect 19545 16875 19555 16915
rect 19595 16875 19605 16915
rect 19645 16875 19655 16915
rect 19695 16875 19705 16915
rect 19745 16875 19755 16915
rect 19795 16875 19805 16915
rect 19845 16875 19855 16915
rect 19895 16875 19905 16915
rect 19945 16875 19955 16915
rect 19995 16875 20005 16915
rect 20045 16875 20055 16915
rect 20095 16875 20105 16915
rect 20145 16875 20155 16915
rect 20195 16875 20205 16915
rect 20245 16875 20255 16915
rect 20295 16875 20305 16915
rect 20345 16875 20355 16915
rect 20395 16875 20405 16915
rect 20445 16875 20455 16915
rect 20495 16875 20505 16915
rect 20545 16875 20555 16915
rect 20595 16875 20605 16915
rect 20645 16875 20655 16915
rect 20695 16875 20705 16915
rect 20745 16875 20755 16915
rect 20795 16875 20805 16915
rect 20845 16875 20855 16915
rect 20895 16875 20905 16915
rect 20945 16875 20955 16915
rect 20995 16875 21005 16915
rect 21045 16875 21055 16915
rect 21095 16875 21105 16915
rect 21145 16875 21155 16915
rect 21195 16875 21205 16915
rect 21245 16875 21255 16915
rect 21295 16875 21305 16915
rect 21345 16875 21355 16915
rect 21395 16875 21405 16915
rect 21445 16875 21455 16915
rect 21495 16875 21505 16915
rect 21545 16875 21555 16915
rect 21595 16875 21605 16915
rect 21645 16875 21655 16915
rect 21695 16875 21705 16915
rect 21745 16875 21755 16915
rect 21795 16875 21805 16915
rect 21845 16875 21855 16915
rect 21895 16875 21905 16915
rect 21945 16875 21955 16915
rect 21995 16875 22005 16915
rect 22045 16875 22055 16915
rect 22095 16875 22105 16915
rect 22145 16875 22155 16915
rect 22195 16875 22205 16915
rect 22245 16875 22255 16915
rect 22295 16875 22305 16915
rect 22345 16875 22355 16915
rect 22395 16875 22405 16915
rect 22445 16875 22455 16915
rect 22495 16875 22505 16915
rect 22545 16875 22555 16915
rect 22595 16875 22605 16915
rect 22645 16875 22655 16915
rect 22695 16875 22705 16915
rect 22745 16875 22755 16915
rect 22795 16875 22805 16915
rect 22845 16875 22855 16915
rect 22895 16875 22905 16915
rect 22945 16875 22955 16915
rect 22995 16875 23005 16915
rect 23045 16875 23055 16915
rect 23095 16875 23105 16915
rect 23145 16875 23155 16915
rect 23195 16875 23205 16915
rect 23245 16875 23255 16915
rect 23295 16875 23305 16915
rect 23345 16875 23355 16915
rect 23395 16875 23405 16915
rect 23445 16875 23455 16915
rect 23495 16875 23505 16915
rect 23545 16875 23555 16915
rect 23595 16875 23605 16915
rect 23645 16875 23655 16915
rect 23695 16875 23705 16915
rect 23745 16875 23755 16915
rect 23795 16875 23805 16915
rect 23845 16875 23855 16915
rect 23895 16875 23905 16915
rect 23945 16875 23955 16915
rect 23995 16875 24005 16915
rect 24045 16875 24055 16915
rect 24095 16875 24105 16915
rect 24145 16875 24155 16915
rect 24195 16875 24205 16915
rect 24245 16875 24255 16915
rect 24295 16875 24305 16915
rect 24345 16875 24355 16915
rect 24395 16875 24405 16915
rect 24445 16875 24455 16915
rect 24495 16875 24505 16915
rect 24545 16875 24555 16915
rect 24595 16875 24605 16915
rect 24645 16875 24655 16915
rect 24695 16875 24705 16915
rect 24745 16875 24755 16915
rect 24795 16875 24805 16915
rect 24845 16875 24855 16915
rect 24895 16875 24905 16915
rect 24945 16875 24955 16915
rect 24995 16875 25005 16915
rect 25045 16875 25055 16915
rect 25095 16875 25105 16915
rect 25145 16875 25155 16915
rect 25195 16875 25205 16915
rect 25245 16875 25255 16915
rect 25295 16875 25305 16915
rect 25345 16875 25355 16915
rect 25395 16875 25405 16915
rect 25445 16875 25455 16915
rect 25495 16875 25505 16915
rect 25545 16875 25555 16915
rect 25595 16875 25605 16915
rect 25645 16875 25655 16915
rect 25695 16875 25705 16915
rect 25745 16875 25755 16915
rect 25795 16875 25805 16915
rect 25845 16875 25855 16915
rect 25895 16875 25905 16915
rect 25945 16875 25955 16915
rect 25995 16875 26005 16915
rect 26045 16875 26055 16915
rect 26095 16875 26105 16915
rect 26145 16875 26155 16915
rect 26195 16875 26205 16915
rect 26245 16875 26255 16915
rect 26295 16875 26305 16915
rect 26345 16875 26355 16915
rect 26395 16875 26405 16915
rect 26445 16875 26455 16915
rect 26495 16875 26505 16915
rect 26545 16875 26555 16915
rect 26595 16875 26605 16915
rect 26645 16875 26655 16915
rect 26695 16875 26705 16915
rect 26745 16875 26755 16915
rect 26795 16875 26805 16915
rect 26845 16875 26855 16915
rect 26895 16875 26905 16915
rect 26945 16875 26955 16915
rect 26995 16875 27005 16915
rect 27045 16875 27055 16915
rect 27095 16875 27105 16915
rect 27145 16875 27155 16915
rect 27195 16875 27205 16915
rect 27245 16875 27255 16915
rect 27295 16875 27305 16915
rect 27345 16875 27355 16915
rect 27395 16875 27405 16915
rect 27445 16875 27455 16915
rect 27495 16875 27505 16915
rect 27545 16875 27555 16915
rect 27595 16875 27605 16915
rect 27645 16875 27655 16915
rect 27695 16875 27705 16915
rect 27745 16875 27755 16915
rect 27795 16875 27805 16915
rect 27845 16875 27855 16915
rect 27895 16875 27905 16915
rect 27945 16875 27955 16915
rect 27995 16875 28005 16915
rect 28045 16875 28055 16915
rect 28095 16875 28105 16915
rect 28145 16875 28155 16915
rect 28195 16875 28205 16915
rect 28245 16875 28255 16915
rect 28295 16875 28305 16915
rect 28345 16875 28355 16915
rect 28395 16875 28405 16915
rect 28445 16875 28455 16915
rect 28495 16875 28505 16915
rect 28545 16875 28555 16915
rect 28595 16875 28605 16915
rect 28645 16875 28655 16915
rect 28695 16875 28705 16915
rect 28745 16875 28755 16915
rect 28795 16875 28805 16915
rect 28845 16875 28855 16915
rect 28895 16875 28905 16915
rect 28945 16875 28955 16915
rect 28995 16875 29005 16915
rect 29045 16875 29055 16915
rect 29095 16875 29105 16915
rect 29145 16875 29155 16915
rect 29195 16875 29205 16915
rect 29245 16875 29255 16915
rect 29295 16875 29305 16915
rect 29345 16875 29355 16915
rect 29395 16875 29405 16915
rect 29445 16875 29455 16915
rect 29495 16875 29505 16915
rect 29545 16875 29555 16915
rect 29595 16875 29605 16915
rect 29645 16875 29655 16915
rect 29695 16875 29705 16915
rect 29745 16875 29755 16915
rect 29795 16875 29805 16915
rect 29845 16875 29855 16915
rect 29895 16875 29905 16915
rect 29945 16875 29955 16915
rect 29995 16875 30005 16915
rect 30045 16875 30055 16915
rect 30095 16875 30105 16915
rect 30145 16875 30155 16915
rect 30195 16875 30205 16915
rect 30245 16875 30255 16915
rect 30295 16875 30305 16915
rect 30345 16875 30355 16915
rect 30395 16875 30405 16915
rect 30445 16875 30455 16915
rect 30495 16875 30505 16915
rect 30545 16875 30555 16915
rect 30595 16875 30605 16915
rect 30645 16875 30655 16915
rect 30695 16875 30705 16915
rect 30745 16875 30755 16915
rect 30795 16875 30805 16915
rect 30845 16875 30855 16915
rect 30895 16875 30905 16915
rect 30945 16875 30955 16915
rect 30995 16875 31005 16915
rect 31045 16875 31055 16915
rect 31095 16875 31105 16915
rect 31145 16875 31155 16915
rect 31195 16875 31205 16915
rect 31245 16875 31255 16915
rect 31295 16875 31305 16915
rect 31345 16875 31355 16915
rect 31395 16875 31405 16915
rect 31445 16875 31455 16915
rect 31495 16875 31505 16915
rect 31545 16875 31555 16915
rect 31595 16875 31605 16915
rect 31645 16875 31655 16915
rect 31695 16875 31705 16915
rect 31745 16875 31755 16915
rect 31795 16875 31805 16915
rect 31845 16875 31855 16915
rect 31895 16875 31905 16915
rect 31945 16875 31955 16915
rect 31995 16875 32005 16915
rect 32045 16875 32055 16915
rect 32095 16875 32105 16915
rect 32145 16875 32155 16915
rect 32195 16875 32205 16915
rect 32245 16875 32255 16915
rect 32295 16875 32305 16915
rect 32345 16875 32355 16915
rect 32395 16875 32405 16915
rect 32445 16875 32455 16915
rect 32495 16875 32505 16915
rect 32545 16875 32555 16915
rect 32595 16875 32605 16915
rect 32645 16875 32655 16915
rect 32695 16875 32705 16915
rect 32745 16875 32755 16915
rect 32795 16875 32805 16915
rect 32845 16875 32855 16915
rect 32895 16875 32905 16915
rect 32945 16875 32955 16915
rect 32995 16875 33005 16915
rect 33045 16875 33055 16915
rect 33095 16875 33105 16915
rect 33145 16875 33155 16915
rect 33195 16875 33205 16915
rect 33245 16875 33255 16915
rect 33295 16875 33305 16915
rect 33345 16875 33355 16915
rect 33395 16875 33405 16915
rect 33445 16875 33455 16915
rect 33495 16875 33505 16915
rect 33545 16875 33555 16915
rect 33595 16875 33605 16915
rect 33645 16875 33655 16915
rect 33695 16875 33705 16915
rect 33745 16875 33755 16915
rect 33795 16875 33805 16915
rect 33845 16875 33855 16915
rect 33895 16875 33905 16915
rect 33945 16875 33955 16915
rect 33995 16875 34005 16915
rect 34045 16875 34055 16915
rect 34095 16875 34105 16915
rect 34145 16875 34155 16915
rect 34195 16875 34205 16915
rect 34245 16875 34255 16915
rect 34295 16875 34305 16915
rect 34345 16875 34355 16915
rect 34395 16875 34405 16915
rect 34445 16875 34455 16915
rect 34495 16875 34505 16915
rect 34545 16875 34555 16915
rect 34595 16875 34605 16915
rect 34645 16875 34655 16915
rect 34695 16875 34705 16915
rect 34745 16875 34755 16915
rect 34795 16875 34805 16915
rect 34845 16875 34855 16915
rect 34895 16875 34905 16915
rect 34945 16875 34955 16915
rect 34995 16875 35005 16915
rect 35045 16875 35055 16915
rect 35095 16875 35105 16915
rect 35145 16875 35155 16915
rect 35195 16875 35205 16915
rect 35245 16875 35255 16915
rect 35295 16875 35305 16915
rect 35345 16875 35355 16915
rect 35395 16875 35405 16915
rect 35445 16875 35455 16915
rect 35495 16875 35505 16915
rect 35545 16875 35555 16915
rect 35595 16875 35605 16915
rect 35645 16875 35655 16915
rect 35695 16875 35705 16915
rect 35745 16875 35755 16915
rect 35795 16875 35805 16915
rect 35845 16875 35855 16915
rect 35895 16875 35905 16915
rect 35945 16875 35955 16915
rect 35995 16875 36005 16915
rect 36045 16875 36055 16915
rect 36095 16875 36105 16915
rect 36145 16875 36155 16915
rect 36195 16875 36205 16915
rect 36245 16875 36255 16915
rect 36295 16875 36305 16915
rect 36345 16875 36355 16915
rect 36395 16875 36405 16915
rect 36445 16875 36455 16915
rect 36495 16875 36505 16915
rect 36545 16875 36555 16915
rect 36595 16875 36605 16915
rect 36645 16875 36655 16915
rect 36695 16875 36705 16915
rect 36745 16875 36755 16915
rect 36795 16875 36805 16915
rect 36845 16875 36855 16915
rect 36895 16875 36905 16915
rect 36945 16875 36955 16915
rect 36995 16875 37005 16915
rect 37045 16875 37055 16915
rect 37095 16875 37105 16915
rect 37145 16875 37155 16915
rect 37195 16875 37205 16915
rect 37245 16875 37255 16915
rect 37295 16875 37305 16915
rect 37345 16875 37355 16915
rect 37395 16875 37405 16915
rect 37445 16875 37455 16915
rect 37495 16875 37505 16915
rect 37545 16875 37555 16915
rect 37595 16875 37605 16915
rect 37645 16875 37655 16915
rect 37695 16875 37705 16915
rect 37745 16875 37755 16915
rect 37795 16875 37805 16915
rect 37845 16875 37855 16915
rect 37895 16875 37905 16915
rect 37945 16875 37955 16915
rect 37995 16875 38005 16915
rect 38045 16875 38055 16915
rect 38095 16875 38105 16915
rect 38145 16875 38155 16915
rect 38195 16875 38205 16915
rect 38245 16875 38255 16915
rect 38295 16875 38305 16915
rect 38345 16875 38355 16915
rect 38395 16875 38405 16915
rect 38445 16875 38455 16915
rect 38495 16875 38505 16915
rect 38545 16875 38555 16915
rect 38595 16875 38605 16915
rect 38645 16875 38655 16915
rect 38695 16875 38705 16915
rect 38745 16875 38755 16915
rect 38795 16875 38805 16915
rect 38845 16875 38855 16915
rect 38895 16875 38905 16915
rect 38945 16875 38955 16915
rect 38995 16875 39005 16915
rect 39045 16875 39055 16915
rect 39095 16875 39105 16915
rect 39145 16875 39155 16915
rect 39195 16875 39205 16915
rect 39245 16875 39255 16915
rect 39295 16875 39305 16915
rect 39345 16875 39355 16915
rect 39395 16875 39405 16915
rect 39445 16875 39455 16915
rect 39495 16875 39505 16915
rect 39545 16875 39555 16915
rect 39595 16875 39605 16915
rect 39645 16875 39655 16915
rect 39695 16875 39705 16915
rect 39745 16875 39750 16915
rect -400 16870 39750 16875
rect 100 15850 3200 16750
rect 3350 15850 6450 16750
rect 6600 15850 9700 16750
rect 9850 15850 12950 16750
rect 13100 15850 16200 16750
rect 16350 15850 19450 16750
rect 19600 15850 22700 16750
rect 22850 15850 25950 16750
rect 26100 15850 29200 16750
rect 29350 15850 32450 16750
rect 32600 15850 35700 16750
rect 35850 15850 38950 16750
rect 39100 15850 39750 16750
rect 0 15845 39750 15850
rect 0 15805 5 15845
rect 45 15805 55 15845
rect 95 15805 105 15845
rect 145 15805 155 15845
rect 195 15805 205 15845
rect 245 15805 255 15845
rect 295 15805 305 15845
rect 345 15805 355 15845
rect 395 15805 405 15845
rect 445 15805 455 15845
rect 495 15805 505 15845
rect 545 15805 555 15845
rect 595 15805 605 15845
rect 645 15805 655 15845
rect 695 15805 705 15845
rect 745 15805 755 15845
rect 795 15805 805 15845
rect 845 15805 855 15845
rect 895 15805 905 15845
rect 945 15805 955 15845
rect 995 15805 1005 15845
rect 1045 15805 1055 15845
rect 1095 15805 1105 15845
rect 1145 15805 1155 15845
rect 1195 15805 1205 15845
rect 1245 15805 1255 15845
rect 1295 15805 1305 15845
rect 1345 15805 1355 15845
rect 1395 15805 1405 15845
rect 1445 15805 1455 15845
rect 1495 15805 1505 15845
rect 1545 15805 1555 15845
rect 1595 15805 1605 15845
rect 1645 15805 1655 15845
rect 1695 15805 1705 15845
rect 1745 15805 1755 15845
rect 1795 15805 1805 15845
rect 1845 15805 1855 15845
rect 1895 15805 1905 15845
rect 1945 15805 1955 15845
rect 1995 15805 2005 15845
rect 2045 15805 2055 15845
rect 2095 15805 2105 15845
rect 2145 15805 2155 15845
rect 2195 15805 2205 15845
rect 2245 15805 2255 15845
rect 2295 15805 2305 15845
rect 2345 15805 2355 15845
rect 2395 15805 2405 15845
rect 2445 15805 2455 15845
rect 2495 15805 2505 15845
rect 2545 15805 2555 15845
rect 2595 15805 2605 15845
rect 2645 15805 2655 15845
rect 2695 15805 2705 15845
rect 2745 15805 2755 15845
rect 2795 15805 2805 15845
rect 2845 15805 2855 15845
rect 2895 15805 2905 15845
rect 2945 15805 2955 15845
rect 2995 15805 3005 15845
rect 3045 15805 3055 15845
rect 3095 15805 3105 15845
rect 3145 15805 3155 15845
rect 3195 15805 3205 15845
rect 3245 15805 3255 15845
rect 3295 15805 3305 15845
rect 3345 15805 3355 15845
rect 3395 15805 3405 15845
rect 3445 15805 3455 15845
rect 3495 15805 3505 15845
rect 3545 15805 3555 15845
rect 3595 15805 3605 15845
rect 3645 15805 3655 15845
rect 3695 15805 3705 15845
rect 3745 15805 3755 15845
rect 3795 15805 3805 15845
rect 3845 15805 3855 15845
rect 3895 15805 3905 15845
rect 3945 15805 3955 15845
rect 3995 15805 4005 15845
rect 4045 15805 4055 15845
rect 4095 15805 4105 15845
rect 4145 15805 4155 15845
rect 4195 15805 4205 15845
rect 4245 15805 4255 15845
rect 4295 15805 4305 15845
rect 4345 15805 4355 15845
rect 4395 15805 4405 15845
rect 4445 15805 4455 15845
rect 4495 15805 4505 15845
rect 4545 15805 4555 15845
rect 4595 15805 4605 15845
rect 4645 15805 4655 15845
rect 4695 15805 4705 15845
rect 4745 15805 4755 15845
rect 4795 15805 4805 15845
rect 4845 15805 4855 15845
rect 4895 15805 4905 15845
rect 4945 15805 4955 15845
rect 4995 15805 5005 15845
rect 5045 15805 5055 15845
rect 5095 15805 5105 15845
rect 5145 15805 5155 15845
rect 5195 15805 5205 15845
rect 5245 15805 5255 15845
rect 5295 15805 5305 15845
rect 5345 15805 5355 15845
rect 5395 15805 5405 15845
rect 5445 15805 5455 15845
rect 5495 15805 5505 15845
rect 5545 15805 5555 15845
rect 5595 15805 5605 15845
rect 5645 15805 5655 15845
rect 5695 15805 5705 15845
rect 5745 15805 5755 15845
rect 5795 15805 5805 15845
rect 5845 15805 5855 15845
rect 5895 15805 5905 15845
rect 5945 15805 5955 15845
rect 5995 15805 6005 15845
rect 6045 15805 6055 15845
rect 6095 15805 6105 15845
rect 6145 15805 6155 15845
rect 6195 15805 6205 15845
rect 6245 15805 6255 15845
rect 6295 15805 6305 15845
rect 6345 15805 6355 15845
rect 6395 15805 6405 15845
rect 6445 15805 6455 15845
rect 6495 15805 6505 15845
rect 6545 15805 6555 15845
rect 6595 15805 6605 15845
rect 6645 15805 6655 15845
rect 6695 15805 6705 15845
rect 6745 15805 6755 15845
rect 6795 15805 6805 15845
rect 6845 15805 6855 15845
rect 6895 15805 6905 15845
rect 6945 15805 6955 15845
rect 6995 15805 7005 15845
rect 7045 15805 7055 15845
rect 7095 15805 7105 15845
rect 7145 15805 7155 15845
rect 7195 15805 7205 15845
rect 7245 15805 7255 15845
rect 7295 15805 7305 15845
rect 7345 15805 7355 15845
rect 7395 15805 7405 15845
rect 7445 15805 7455 15845
rect 7495 15805 7505 15845
rect 7545 15805 7555 15845
rect 7595 15805 7605 15845
rect 7645 15805 7655 15845
rect 7695 15805 7705 15845
rect 7745 15805 7755 15845
rect 7795 15805 7805 15845
rect 7845 15805 7855 15845
rect 7895 15805 7905 15845
rect 7945 15805 7955 15845
rect 7995 15805 8005 15845
rect 8045 15805 8055 15845
rect 8095 15805 8105 15845
rect 8145 15805 8155 15845
rect 8195 15805 8205 15845
rect 8245 15805 8255 15845
rect 8295 15805 8305 15845
rect 8345 15805 8355 15845
rect 8395 15805 8405 15845
rect 8445 15805 8455 15845
rect 8495 15805 8505 15845
rect 8545 15805 8555 15845
rect 8595 15805 8605 15845
rect 8645 15805 8655 15845
rect 8695 15805 8705 15845
rect 8745 15805 8755 15845
rect 8795 15805 8805 15845
rect 8845 15805 8855 15845
rect 8895 15805 8905 15845
rect 8945 15805 8955 15845
rect 8995 15805 9005 15845
rect 9045 15805 9055 15845
rect 9095 15805 9105 15845
rect 9145 15805 9155 15845
rect 9195 15805 9205 15845
rect 9245 15805 9255 15845
rect 9295 15805 9305 15845
rect 9345 15805 9355 15845
rect 9395 15805 9405 15845
rect 9445 15805 9455 15845
rect 9495 15805 9505 15845
rect 9545 15805 9555 15845
rect 9595 15805 9605 15845
rect 9645 15805 9655 15845
rect 9695 15805 9705 15845
rect 9745 15805 9755 15845
rect 9795 15805 9805 15845
rect 9845 15805 9855 15845
rect 9895 15805 9905 15845
rect 9945 15805 9955 15845
rect 9995 15805 10005 15845
rect 10045 15805 10055 15845
rect 10095 15805 10105 15845
rect 10145 15805 10155 15845
rect 10195 15805 10205 15845
rect 10245 15805 10255 15845
rect 10295 15805 10305 15845
rect 10345 15805 10355 15845
rect 10395 15805 10405 15845
rect 10445 15805 10455 15845
rect 10495 15805 10505 15845
rect 10545 15805 10555 15845
rect 10595 15805 10605 15845
rect 10645 15805 10655 15845
rect 10695 15805 10705 15845
rect 10745 15805 10755 15845
rect 10795 15805 10805 15845
rect 10845 15805 10855 15845
rect 10895 15805 10905 15845
rect 10945 15805 10955 15845
rect 10995 15805 11005 15845
rect 11045 15805 11055 15845
rect 11095 15805 11105 15845
rect 11145 15805 11155 15845
rect 11195 15805 11205 15845
rect 11245 15805 11255 15845
rect 11295 15805 11305 15845
rect 11345 15805 11355 15845
rect 11395 15805 11405 15845
rect 11445 15805 11455 15845
rect 11495 15805 11505 15845
rect 11545 15805 11555 15845
rect 11595 15805 11605 15845
rect 11645 15805 11655 15845
rect 11695 15805 11705 15845
rect 11745 15805 11755 15845
rect 11795 15805 11805 15845
rect 11845 15805 11855 15845
rect 11895 15805 11905 15845
rect 11945 15805 11955 15845
rect 11995 15805 12005 15845
rect 12045 15805 12055 15845
rect 12095 15805 12105 15845
rect 12145 15805 12155 15845
rect 12195 15805 12205 15845
rect 12245 15805 12255 15845
rect 12295 15805 12305 15845
rect 12345 15805 12355 15845
rect 12395 15805 12405 15845
rect 12445 15805 12455 15845
rect 12495 15805 12505 15845
rect 12545 15805 12555 15845
rect 12595 15805 12605 15845
rect 12645 15805 12655 15845
rect 12695 15805 12705 15845
rect 12745 15805 12755 15845
rect 12795 15805 12805 15845
rect 12845 15805 12855 15845
rect 12895 15805 12905 15845
rect 12945 15805 12955 15845
rect 12995 15805 13005 15845
rect 13045 15805 13055 15845
rect 13095 15805 13105 15845
rect 13145 15805 13155 15845
rect 13195 15805 13205 15845
rect 13245 15805 13255 15845
rect 13295 15805 13305 15845
rect 13345 15805 13355 15845
rect 13395 15805 13405 15845
rect 13445 15805 13455 15845
rect 13495 15805 13505 15845
rect 13545 15805 13555 15845
rect 13595 15805 13605 15845
rect 13645 15805 13655 15845
rect 13695 15805 13705 15845
rect 13745 15805 13755 15845
rect 13795 15805 13805 15845
rect 13845 15805 13855 15845
rect 13895 15805 13905 15845
rect 13945 15805 13955 15845
rect 13995 15805 14005 15845
rect 14045 15805 14055 15845
rect 14095 15805 14105 15845
rect 14145 15805 14155 15845
rect 14195 15805 14205 15845
rect 14245 15805 14255 15845
rect 14295 15805 14305 15845
rect 14345 15805 14355 15845
rect 14395 15805 14405 15845
rect 14445 15805 14455 15845
rect 14495 15805 14505 15845
rect 14545 15805 14555 15845
rect 14595 15805 14605 15845
rect 14645 15805 14655 15845
rect 14695 15805 14705 15845
rect 14745 15805 14755 15845
rect 14795 15805 14805 15845
rect 14845 15805 14855 15845
rect 14895 15805 14905 15845
rect 14945 15805 14955 15845
rect 14995 15805 15005 15845
rect 15045 15805 15055 15845
rect 15095 15805 15105 15845
rect 15145 15805 15155 15845
rect 15195 15805 15205 15845
rect 15245 15805 15255 15845
rect 15295 15805 15305 15845
rect 15345 15805 15355 15845
rect 15395 15805 15405 15845
rect 15445 15805 15455 15845
rect 15495 15805 15505 15845
rect 15545 15805 15555 15845
rect 15595 15805 15605 15845
rect 15645 15805 15655 15845
rect 15695 15805 15705 15845
rect 15745 15805 15755 15845
rect 15795 15805 15805 15845
rect 15845 15805 15855 15845
rect 15895 15805 15905 15845
rect 15945 15805 15955 15845
rect 15995 15805 16005 15845
rect 16045 15805 16055 15845
rect 16095 15805 16105 15845
rect 16145 15805 16155 15845
rect 16195 15805 16205 15845
rect 16245 15805 16255 15845
rect 16295 15805 16305 15845
rect 16345 15805 16355 15845
rect 16395 15805 16405 15845
rect 16445 15805 16455 15845
rect 16495 15805 16505 15845
rect 16545 15805 16555 15845
rect 16595 15805 16605 15845
rect 16645 15805 16655 15845
rect 16695 15805 16705 15845
rect 16745 15805 16755 15845
rect 16795 15805 16805 15845
rect 16845 15805 16855 15845
rect 16895 15805 16905 15845
rect 16945 15805 16955 15845
rect 16995 15805 17005 15845
rect 17045 15805 17055 15845
rect 17095 15805 17105 15845
rect 17145 15805 17155 15845
rect 17195 15805 17205 15845
rect 17245 15805 17255 15845
rect 17295 15805 17305 15845
rect 17345 15805 17355 15845
rect 17395 15805 17405 15845
rect 17445 15805 17455 15845
rect 17495 15805 17505 15845
rect 17545 15805 17555 15845
rect 17595 15805 17605 15845
rect 17645 15805 17655 15845
rect 17695 15805 17705 15845
rect 17745 15805 17755 15845
rect 17795 15805 17805 15845
rect 17845 15805 17855 15845
rect 17895 15805 17905 15845
rect 17945 15805 17955 15845
rect 17995 15805 18005 15845
rect 18045 15805 18055 15845
rect 18095 15805 18105 15845
rect 18145 15805 18155 15845
rect 18195 15805 18205 15845
rect 18245 15805 18255 15845
rect 18295 15805 18305 15845
rect 18345 15805 18355 15845
rect 18395 15805 18405 15845
rect 18445 15805 18455 15845
rect 18495 15805 18505 15845
rect 18545 15805 18555 15845
rect 18595 15805 18605 15845
rect 18645 15805 18655 15845
rect 18695 15805 18705 15845
rect 18745 15805 18755 15845
rect 18795 15805 18805 15845
rect 18845 15805 18855 15845
rect 18895 15805 18905 15845
rect 18945 15805 18955 15845
rect 18995 15805 19005 15845
rect 19045 15805 19055 15845
rect 19095 15805 19105 15845
rect 19145 15805 19155 15845
rect 19195 15805 19205 15845
rect 19245 15805 19255 15845
rect 19295 15805 19305 15845
rect 19345 15805 19355 15845
rect 19395 15805 19405 15845
rect 19445 15805 19455 15845
rect 19495 15805 19505 15845
rect 19545 15805 19555 15845
rect 19595 15805 19605 15845
rect 19645 15805 19655 15845
rect 19695 15805 19705 15845
rect 19745 15805 19755 15845
rect 19795 15805 19805 15845
rect 19845 15805 19855 15845
rect 19895 15805 19905 15845
rect 19945 15805 19955 15845
rect 19995 15805 20005 15845
rect 20045 15805 20055 15845
rect 20095 15805 20105 15845
rect 20145 15805 20155 15845
rect 20195 15805 20205 15845
rect 20245 15805 20255 15845
rect 20295 15805 20305 15845
rect 20345 15805 20355 15845
rect 20395 15805 20405 15845
rect 20445 15805 20455 15845
rect 20495 15805 20505 15845
rect 20545 15805 20555 15845
rect 20595 15805 20605 15845
rect 20645 15805 20655 15845
rect 20695 15805 20705 15845
rect 20745 15805 20755 15845
rect 20795 15805 20805 15845
rect 20845 15805 20855 15845
rect 20895 15805 20905 15845
rect 20945 15805 20955 15845
rect 20995 15805 21005 15845
rect 21045 15805 21055 15845
rect 21095 15805 21105 15845
rect 21145 15805 21155 15845
rect 21195 15805 21205 15845
rect 21245 15805 21255 15845
rect 21295 15805 21305 15845
rect 21345 15805 21355 15845
rect 21395 15805 21405 15845
rect 21445 15805 21455 15845
rect 21495 15805 21505 15845
rect 21545 15805 21555 15845
rect 21595 15805 21605 15845
rect 21645 15805 21655 15845
rect 21695 15805 21705 15845
rect 21745 15805 21755 15845
rect 21795 15805 21805 15845
rect 21845 15805 21855 15845
rect 21895 15805 21905 15845
rect 21945 15805 21955 15845
rect 21995 15805 22005 15845
rect 22045 15805 22055 15845
rect 22095 15805 22105 15845
rect 22145 15805 22155 15845
rect 22195 15805 22205 15845
rect 22245 15805 22255 15845
rect 22295 15805 22305 15845
rect 22345 15805 22355 15845
rect 22395 15805 22405 15845
rect 22445 15805 22455 15845
rect 22495 15805 22505 15845
rect 22545 15805 22555 15845
rect 22595 15805 22605 15845
rect 22645 15805 22655 15845
rect 22695 15805 22705 15845
rect 22745 15805 22755 15845
rect 22795 15805 22805 15845
rect 22845 15805 22855 15845
rect 22895 15805 22905 15845
rect 22945 15805 22955 15845
rect 22995 15805 23005 15845
rect 23045 15805 23055 15845
rect 23095 15805 23105 15845
rect 23145 15805 23155 15845
rect 23195 15805 23205 15845
rect 23245 15805 23255 15845
rect 23295 15805 23305 15845
rect 23345 15805 23355 15845
rect 23395 15805 23405 15845
rect 23445 15805 23455 15845
rect 23495 15805 23505 15845
rect 23545 15805 23555 15845
rect 23595 15805 23605 15845
rect 23645 15805 23655 15845
rect 23695 15805 23705 15845
rect 23745 15805 23755 15845
rect 23795 15805 23805 15845
rect 23845 15805 23855 15845
rect 23895 15805 23905 15845
rect 23945 15805 23955 15845
rect 23995 15805 24005 15845
rect 24045 15805 24055 15845
rect 24095 15805 24105 15845
rect 24145 15805 24155 15845
rect 24195 15805 24205 15845
rect 24245 15805 24255 15845
rect 24295 15805 24305 15845
rect 24345 15805 24355 15845
rect 24395 15805 24405 15845
rect 24445 15805 24455 15845
rect 24495 15805 24505 15845
rect 24545 15805 24555 15845
rect 24595 15805 24605 15845
rect 24645 15805 24655 15845
rect 24695 15805 24705 15845
rect 24745 15805 24755 15845
rect 24795 15805 24805 15845
rect 24845 15805 24855 15845
rect 24895 15805 24905 15845
rect 24945 15805 24955 15845
rect 24995 15805 25005 15845
rect 25045 15805 25055 15845
rect 25095 15805 25105 15845
rect 25145 15805 25155 15845
rect 25195 15805 25205 15845
rect 25245 15805 25255 15845
rect 25295 15805 25305 15845
rect 25345 15805 25355 15845
rect 25395 15805 25405 15845
rect 25445 15805 25455 15845
rect 25495 15805 25505 15845
rect 25545 15805 25555 15845
rect 25595 15805 25605 15845
rect 25645 15805 25655 15845
rect 25695 15805 25705 15845
rect 25745 15805 25755 15845
rect 25795 15805 25805 15845
rect 25845 15805 25855 15845
rect 25895 15805 25905 15845
rect 25945 15805 25955 15845
rect 25995 15805 26005 15845
rect 26045 15805 26055 15845
rect 26095 15805 26105 15845
rect 26145 15805 26155 15845
rect 26195 15805 26205 15845
rect 26245 15805 26255 15845
rect 26295 15805 26305 15845
rect 26345 15805 26355 15845
rect 26395 15805 26405 15845
rect 26445 15805 26455 15845
rect 26495 15805 26505 15845
rect 26545 15805 26555 15845
rect 26595 15805 26605 15845
rect 26645 15805 26655 15845
rect 26695 15805 26705 15845
rect 26745 15805 26755 15845
rect 26795 15805 26805 15845
rect 26845 15805 26855 15845
rect 26895 15805 26905 15845
rect 26945 15805 26955 15845
rect 26995 15805 27005 15845
rect 27045 15805 27055 15845
rect 27095 15805 27105 15845
rect 27145 15805 27155 15845
rect 27195 15805 27205 15845
rect 27245 15805 27255 15845
rect 27295 15805 27305 15845
rect 27345 15805 27355 15845
rect 27395 15805 27405 15845
rect 27445 15805 27455 15845
rect 27495 15805 27505 15845
rect 27545 15805 27555 15845
rect 27595 15805 27605 15845
rect 27645 15805 27655 15845
rect 27695 15805 27705 15845
rect 27745 15805 27755 15845
rect 27795 15805 27805 15845
rect 27845 15805 27855 15845
rect 27895 15805 27905 15845
rect 27945 15805 27955 15845
rect 27995 15805 28005 15845
rect 28045 15805 28055 15845
rect 28095 15805 28105 15845
rect 28145 15805 28155 15845
rect 28195 15805 28205 15845
rect 28245 15805 28255 15845
rect 28295 15805 28305 15845
rect 28345 15805 28355 15845
rect 28395 15805 28405 15845
rect 28445 15805 28455 15845
rect 28495 15805 28505 15845
rect 28545 15805 28555 15845
rect 28595 15805 28605 15845
rect 28645 15805 28655 15845
rect 28695 15805 28705 15845
rect 28745 15805 28755 15845
rect 28795 15805 28805 15845
rect 28845 15805 28855 15845
rect 28895 15805 28905 15845
rect 28945 15805 28955 15845
rect 28995 15805 29005 15845
rect 29045 15805 29055 15845
rect 29095 15805 29105 15845
rect 29145 15805 29155 15845
rect 29195 15805 29205 15845
rect 29245 15805 29255 15845
rect 29295 15805 29305 15845
rect 29345 15805 29355 15845
rect 29395 15805 29405 15845
rect 29445 15805 29455 15845
rect 29495 15805 29505 15845
rect 29545 15805 29555 15845
rect 29595 15805 29605 15845
rect 29645 15805 29655 15845
rect 29695 15805 29705 15845
rect 29745 15805 29755 15845
rect 29795 15805 29805 15845
rect 29845 15805 29855 15845
rect 29895 15805 29905 15845
rect 29945 15805 29955 15845
rect 29995 15805 30005 15845
rect 30045 15805 30055 15845
rect 30095 15805 30105 15845
rect 30145 15805 30155 15845
rect 30195 15805 30205 15845
rect 30245 15805 30255 15845
rect 30295 15805 30305 15845
rect 30345 15805 30355 15845
rect 30395 15805 30405 15845
rect 30445 15805 30455 15845
rect 30495 15805 30505 15845
rect 30545 15805 30555 15845
rect 30595 15805 30605 15845
rect 30645 15805 30655 15845
rect 30695 15805 30705 15845
rect 30745 15805 30755 15845
rect 30795 15805 30805 15845
rect 30845 15805 30855 15845
rect 30895 15805 30905 15845
rect 30945 15805 30955 15845
rect 30995 15805 31005 15845
rect 31045 15805 31055 15845
rect 31095 15805 31105 15845
rect 31145 15805 31155 15845
rect 31195 15805 31205 15845
rect 31245 15805 31255 15845
rect 31295 15805 31305 15845
rect 31345 15805 31355 15845
rect 31395 15805 31405 15845
rect 31445 15805 31455 15845
rect 31495 15805 31505 15845
rect 31545 15805 31555 15845
rect 31595 15805 31605 15845
rect 31645 15805 31655 15845
rect 31695 15805 31705 15845
rect 31745 15805 31755 15845
rect 31795 15805 31805 15845
rect 31845 15805 31855 15845
rect 31895 15805 31905 15845
rect 31945 15805 31955 15845
rect 31995 15805 32005 15845
rect 32045 15805 32055 15845
rect 32095 15805 32105 15845
rect 32145 15805 32155 15845
rect 32195 15805 32205 15845
rect 32245 15805 32255 15845
rect 32295 15805 32305 15845
rect 32345 15805 32355 15845
rect 32395 15805 32405 15845
rect 32445 15805 32455 15845
rect 32495 15805 32505 15845
rect 32545 15805 32555 15845
rect 32595 15805 32605 15845
rect 32645 15805 32655 15845
rect 32695 15805 32705 15845
rect 32745 15805 32755 15845
rect 32795 15805 32805 15845
rect 32845 15805 32855 15845
rect 32895 15805 32905 15845
rect 32945 15805 32955 15845
rect 32995 15805 33005 15845
rect 33045 15805 33055 15845
rect 33095 15805 33105 15845
rect 33145 15805 33155 15845
rect 33195 15805 33205 15845
rect 33245 15805 33255 15845
rect 33295 15805 33305 15845
rect 33345 15805 33355 15845
rect 33395 15805 33405 15845
rect 33445 15805 33455 15845
rect 33495 15805 33505 15845
rect 33545 15805 33555 15845
rect 33595 15805 33605 15845
rect 33645 15805 33655 15845
rect 33695 15805 33705 15845
rect 33745 15805 33755 15845
rect 33795 15805 33805 15845
rect 33845 15805 33855 15845
rect 33895 15805 33905 15845
rect 33945 15805 33955 15845
rect 33995 15805 34005 15845
rect 34045 15805 34055 15845
rect 34095 15805 34105 15845
rect 34145 15805 34155 15845
rect 34195 15805 34205 15845
rect 34245 15805 34255 15845
rect 34295 15805 34305 15845
rect 34345 15805 34355 15845
rect 34395 15805 34405 15845
rect 34445 15805 34455 15845
rect 34495 15805 34505 15845
rect 34545 15805 34555 15845
rect 34595 15805 34605 15845
rect 34645 15805 34655 15845
rect 34695 15805 34705 15845
rect 34745 15805 34755 15845
rect 34795 15805 34805 15845
rect 34845 15805 34855 15845
rect 34895 15805 34905 15845
rect 34945 15805 34955 15845
rect 34995 15805 35005 15845
rect 35045 15805 35055 15845
rect 35095 15805 35105 15845
rect 35145 15805 35155 15845
rect 35195 15805 35205 15845
rect 35245 15805 35255 15845
rect 35295 15805 35305 15845
rect 35345 15805 35355 15845
rect 35395 15805 35405 15845
rect 35445 15805 35455 15845
rect 35495 15805 35505 15845
rect 35545 15805 35555 15845
rect 35595 15805 35605 15845
rect 35645 15805 35655 15845
rect 35695 15805 35705 15845
rect 35745 15805 35755 15845
rect 35795 15805 35805 15845
rect 35845 15805 35855 15845
rect 35895 15805 35905 15845
rect 35945 15805 35955 15845
rect 35995 15805 36005 15845
rect 36045 15805 36055 15845
rect 36095 15805 36105 15845
rect 36145 15805 36155 15845
rect 36195 15805 36205 15845
rect 36245 15805 36255 15845
rect 36295 15805 36305 15845
rect 36345 15805 36355 15845
rect 36395 15805 36405 15845
rect 36445 15805 36455 15845
rect 36495 15805 36505 15845
rect 36545 15805 36555 15845
rect 36595 15805 36605 15845
rect 36645 15805 36655 15845
rect 36695 15805 36705 15845
rect 36745 15805 36755 15845
rect 36795 15805 36805 15845
rect 36845 15805 36855 15845
rect 36895 15805 36905 15845
rect 36945 15805 36955 15845
rect 36995 15805 37005 15845
rect 37045 15805 37055 15845
rect 37095 15805 37105 15845
rect 37145 15805 37155 15845
rect 37195 15805 37205 15845
rect 37245 15805 37255 15845
rect 37295 15805 37305 15845
rect 37345 15805 37355 15845
rect 37395 15805 37405 15845
rect 37445 15805 37455 15845
rect 37495 15805 37505 15845
rect 37545 15805 37555 15845
rect 37595 15805 37605 15845
rect 37645 15805 37655 15845
rect 37695 15805 37705 15845
rect 37745 15805 37755 15845
rect 37795 15805 37805 15845
rect 37845 15805 37855 15845
rect 37895 15805 37905 15845
rect 37945 15805 37955 15845
rect 37995 15805 38005 15845
rect 38045 15805 38055 15845
rect 38095 15805 38105 15845
rect 38145 15805 38155 15845
rect 38195 15805 38205 15845
rect 38245 15805 38255 15845
rect 38295 15805 38305 15845
rect 38345 15805 38355 15845
rect 38395 15805 38405 15845
rect 38445 15805 38455 15845
rect 38495 15805 38505 15845
rect 38545 15805 38555 15845
rect 38595 15805 38605 15845
rect 38645 15805 38655 15845
rect 38695 15805 38705 15845
rect 38745 15805 38755 15845
rect 38795 15805 38805 15845
rect 38845 15805 38855 15845
rect 38895 15805 38905 15845
rect 38945 15805 38955 15845
rect 38995 15805 39005 15845
rect 39045 15805 39055 15845
rect 39095 15805 39105 15845
rect 39145 15805 39155 15845
rect 39195 15805 39205 15845
rect 39245 15805 39255 15845
rect 39295 15805 39305 15845
rect 39345 15805 39355 15845
rect 39395 15805 39405 15845
rect 39445 15805 39455 15845
rect 39495 15805 39505 15845
rect 39545 15805 39555 15845
rect 39595 15805 39605 15845
rect 39645 15805 39655 15845
rect 39695 15805 39705 15845
rect 39745 15805 39750 15845
rect 0 15800 39750 15805
rect -3500 15745 -50 15750
rect -3500 15705 -3495 15745
rect -3455 15705 -3295 15745
rect -3255 15705 -3095 15745
rect -3055 15705 -1595 15745
rect -1555 15705 -1195 15745
rect -1155 15705 -1095 15745
rect -1055 15705 -995 15745
rect -955 15705 -895 15745
rect -855 15705 -695 15745
rect -655 15705 -595 15745
rect -555 15705 -495 15745
rect -455 15705 -295 15745
rect -255 15705 -195 15745
rect -155 15705 -95 15745
rect -55 15705 -50 15745
rect -3500 15700 -50 15705
rect 0 15745 40900 15750
rect 0 15705 5 15745
rect 45 15705 55 15745
rect 95 15705 105 15745
rect 145 15705 155 15745
rect 195 15705 205 15745
rect 245 15705 255 15745
rect 295 15705 305 15745
rect 345 15705 355 15745
rect 395 15705 405 15745
rect 445 15705 455 15745
rect 495 15705 505 15745
rect 545 15705 555 15745
rect 595 15705 605 15745
rect 645 15705 655 15745
rect 695 15705 705 15745
rect 745 15705 755 15745
rect 795 15705 805 15745
rect 845 15705 855 15745
rect 895 15705 905 15745
rect 945 15705 955 15745
rect 995 15705 1005 15745
rect 1045 15705 1055 15745
rect 1095 15705 1105 15745
rect 1145 15705 1155 15745
rect 1195 15705 1205 15745
rect 1245 15705 1255 15745
rect 1295 15705 1305 15745
rect 1345 15705 1355 15745
rect 1395 15705 1405 15745
rect 1445 15705 1455 15745
rect 1495 15705 1505 15745
rect 1545 15705 1555 15745
rect 1595 15705 1605 15745
rect 1645 15705 1655 15745
rect 1695 15705 1705 15745
rect 1745 15705 1755 15745
rect 1795 15705 1805 15745
rect 1845 15705 1855 15745
rect 1895 15705 1905 15745
rect 1945 15705 1955 15745
rect 1995 15705 2005 15745
rect 2045 15705 2055 15745
rect 2095 15705 2105 15745
rect 2145 15705 2155 15745
rect 2195 15705 2205 15745
rect 2245 15705 2255 15745
rect 2295 15705 2305 15745
rect 2345 15705 2355 15745
rect 2395 15705 2405 15745
rect 2445 15705 2455 15745
rect 2495 15705 2505 15745
rect 2545 15705 2555 15745
rect 2595 15705 2605 15745
rect 2645 15705 2655 15745
rect 2695 15705 2705 15745
rect 2745 15705 2755 15745
rect 2795 15705 2805 15745
rect 2845 15705 2855 15745
rect 2895 15705 2905 15745
rect 2945 15705 2955 15745
rect 2995 15705 3005 15745
rect 3045 15705 3055 15745
rect 3095 15705 3105 15745
rect 3145 15705 3155 15745
rect 3195 15705 3205 15745
rect 3245 15705 3255 15745
rect 3295 15705 3305 15745
rect 3345 15705 3355 15745
rect 3395 15705 3405 15745
rect 3445 15705 3455 15745
rect 3495 15705 3505 15745
rect 3545 15705 3555 15745
rect 3595 15705 3605 15745
rect 3645 15705 3655 15745
rect 3695 15705 3705 15745
rect 3745 15705 3755 15745
rect 3795 15705 3805 15745
rect 3845 15705 3855 15745
rect 3895 15705 3905 15745
rect 3945 15705 3955 15745
rect 3995 15705 4005 15745
rect 4045 15705 4055 15745
rect 4095 15705 4105 15745
rect 4145 15705 4155 15745
rect 4195 15705 4205 15745
rect 4245 15705 4255 15745
rect 4295 15705 4305 15745
rect 4345 15705 4355 15745
rect 4395 15705 4405 15745
rect 4445 15705 4455 15745
rect 4495 15705 4505 15745
rect 4545 15705 4555 15745
rect 4595 15705 4605 15745
rect 4645 15705 4655 15745
rect 4695 15705 4705 15745
rect 4745 15705 4755 15745
rect 4795 15705 4805 15745
rect 4845 15705 4855 15745
rect 4895 15705 4905 15745
rect 4945 15705 4955 15745
rect 4995 15705 5005 15745
rect 5045 15705 5055 15745
rect 5095 15705 5105 15745
rect 5145 15705 5155 15745
rect 5195 15705 5205 15745
rect 5245 15705 5255 15745
rect 5295 15705 5305 15745
rect 5345 15705 5355 15745
rect 5395 15705 5405 15745
rect 5445 15705 5455 15745
rect 5495 15705 5505 15745
rect 5545 15705 5555 15745
rect 5595 15705 5605 15745
rect 5645 15705 5655 15745
rect 5695 15705 5705 15745
rect 5745 15705 5755 15745
rect 5795 15705 5805 15745
rect 5845 15705 5855 15745
rect 5895 15705 5905 15745
rect 5945 15705 5955 15745
rect 5995 15705 6005 15745
rect 6045 15705 6055 15745
rect 6095 15705 6105 15745
rect 6145 15705 6155 15745
rect 6195 15705 6205 15745
rect 6245 15705 6255 15745
rect 6295 15705 6305 15745
rect 6345 15705 6355 15745
rect 6395 15705 6405 15745
rect 6445 15705 6455 15745
rect 6495 15705 6505 15745
rect 6545 15705 6555 15745
rect 6595 15705 6605 15745
rect 6645 15705 6655 15745
rect 6695 15705 6705 15745
rect 6745 15705 6755 15745
rect 6795 15705 6805 15745
rect 6845 15705 6855 15745
rect 6895 15705 6905 15745
rect 6945 15705 6955 15745
rect 6995 15705 7005 15745
rect 7045 15705 7055 15745
rect 7095 15705 7105 15745
rect 7145 15705 7155 15745
rect 7195 15705 7205 15745
rect 7245 15705 7255 15745
rect 7295 15705 7305 15745
rect 7345 15705 7355 15745
rect 7395 15705 7405 15745
rect 7445 15705 7455 15745
rect 7495 15705 7505 15745
rect 7545 15705 7555 15745
rect 7595 15705 7605 15745
rect 7645 15705 7655 15745
rect 7695 15705 7705 15745
rect 7745 15705 7755 15745
rect 7795 15705 7805 15745
rect 7845 15705 7855 15745
rect 7895 15705 7905 15745
rect 7945 15705 7955 15745
rect 7995 15705 8005 15745
rect 8045 15705 8055 15745
rect 8095 15705 8105 15745
rect 8145 15705 8155 15745
rect 8195 15705 8205 15745
rect 8245 15705 8255 15745
rect 8295 15705 8305 15745
rect 8345 15705 8355 15745
rect 8395 15705 8405 15745
rect 8445 15705 8455 15745
rect 8495 15705 8505 15745
rect 8545 15705 8555 15745
rect 8595 15705 8605 15745
rect 8645 15705 8655 15745
rect 8695 15705 8705 15745
rect 8745 15705 8755 15745
rect 8795 15705 8805 15745
rect 8845 15705 8855 15745
rect 8895 15705 8905 15745
rect 8945 15705 8955 15745
rect 8995 15705 9005 15745
rect 9045 15705 9055 15745
rect 9095 15705 9105 15745
rect 9145 15705 9155 15745
rect 9195 15705 9205 15745
rect 9245 15705 9255 15745
rect 9295 15705 9305 15745
rect 9345 15705 9355 15745
rect 9395 15705 9405 15745
rect 9445 15705 9455 15745
rect 9495 15705 9505 15745
rect 9545 15705 9555 15745
rect 9595 15705 9605 15745
rect 9645 15705 9655 15745
rect 9695 15705 9705 15745
rect 9745 15705 9755 15745
rect 9795 15705 9805 15745
rect 9845 15705 9855 15745
rect 9895 15705 9905 15745
rect 9945 15705 9955 15745
rect 9995 15705 10005 15745
rect 10045 15705 10055 15745
rect 10095 15705 10105 15745
rect 10145 15705 10155 15745
rect 10195 15705 10205 15745
rect 10245 15705 10255 15745
rect 10295 15705 10305 15745
rect 10345 15705 10355 15745
rect 10395 15705 10405 15745
rect 10445 15705 10455 15745
rect 10495 15705 10505 15745
rect 10545 15705 10555 15745
rect 10595 15705 10605 15745
rect 10645 15705 10655 15745
rect 10695 15705 10705 15745
rect 10745 15705 10755 15745
rect 10795 15705 10805 15745
rect 10845 15705 10855 15745
rect 10895 15705 10905 15745
rect 10945 15705 10955 15745
rect 10995 15705 11005 15745
rect 11045 15705 11055 15745
rect 11095 15705 11105 15745
rect 11145 15705 11155 15745
rect 11195 15705 11205 15745
rect 11245 15705 11255 15745
rect 11295 15705 11305 15745
rect 11345 15705 11355 15745
rect 11395 15705 11405 15745
rect 11445 15705 11455 15745
rect 11495 15705 11505 15745
rect 11545 15705 11555 15745
rect 11595 15705 11605 15745
rect 11645 15705 11655 15745
rect 11695 15705 11705 15745
rect 11745 15705 11755 15745
rect 11795 15705 11805 15745
rect 11845 15705 11855 15745
rect 11895 15705 11905 15745
rect 11945 15705 11955 15745
rect 11995 15705 12005 15745
rect 12045 15705 12055 15745
rect 12095 15705 12105 15745
rect 12145 15705 12155 15745
rect 12195 15705 12205 15745
rect 12245 15705 12255 15745
rect 12295 15705 12305 15745
rect 12345 15705 12355 15745
rect 12395 15705 12405 15745
rect 12445 15705 12455 15745
rect 12495 15705 12505 15745
rect 12545 15705 12555 15745
rect 12595 15705 12605 15745
rect 12645 15705 12655 15745
rect 12695 15705 12705 15745
rect 12745 15705 12755 15745
rect 12795 15705 12805 15745
rect 12845 15705 12855 15745
rect 12895 15705 12905 15745
rect 12945 15705 12955 15745
rect 12995 15705 13005 15745
rect 13045 15705 13055 15745
rect 13095 15705 13105 15745
rect 13145 15705 13155 15745
rect 13195 15705 13205 15745
rect 13245 15705 13255 15745
rect 13295 15705 13305 15745
rect 13345 15705 13355 15745
rect 13395 15705 13405 15745
rect 13445 15705 13455 15745
rect 13495 15705 13505 15745
rect 13545 15705 13555 15745
rect 13595 15705 13605 15745
rect 13645 15705 13655 15745
rect 13695 15705 13705 15745
rect 13745 15705 13755 15745
rect 13795 15705 13805 15745
rect 13845 15705 13855 15745
rect 13895 15705 13905 15745
rect 13945 15705 13955 15745
rect 13995 15705 14005 15745
rect 14045 15705 14055 15745
rect 14095 15705 14105 15745
rect 14145 15705 14155 15745
rect 14195 15705 14205 15745
rect 14245 15705 14255 15745
rect 14295 15705 14305 15745
rect 14345 15705 14355 15745
rect 14395 15705 14405 15745
rect 14445 15705 14455 15745
rect 14495 15705 14505 15745
rect 14545 15705 14555 15745
rect 14595 15705 14605 15745
rect 14645 15705 14655 15745
rect 14695 15705 14705 15745
rect 14745 15705 14755 15745
rect 14795 15705 14805 15745
rect 14845 15705 14855 15745
rect 14895 15705 14905 15745
rect 14945 15705 14955 15745
rect 14995 15705 15005 15745
rect 15045 15705 15055 15745
rect 15095 15705 15105 15745
rect 15145 15705 15155 15745
rect 15195 15705 15205 15745
rect 15245 15705 15255 15745
rect 15295 15705 15305 15745
rect 15345 15705 15355 15745
rect 15395 15705 15405 15745
rect 15445 15705 15455 15745
rect 15495 15705 15505 15745
rect 15545 15705 15555 15745
rect 15595 15705 15605 15745
rect 15645 15705 15655 15745
rect 15695 15705 15705 15745
rect 15745 15705 15755 15745
rect 15795 15705 15805 15745
rect 15845 15705 15855 15745
rect 15895 15705 15905 15745
rect 15945 15705 15955 15745
rect 15995 15705 16005 15745
rect 16045 15705 16055 15745
rect 16095 15705 16105 15745
rect 16145 15705 16155 15745
rect 16195 15705 16205 15745
rect 16245 15705 16255 15745
rect 16295 15705 16305 15745
rect 16345 15705 16355 15745
rect 16395 15705 16405 15745
rect 16445 15705 16455 15745
rect 16495 15705 16505 15745
rect 16545 15705 16555 15745
rect 16595 15705 16605 15745
rect 16645 15705 16655 15745
rect 16695 15705 16705 15745
rect 16745 15705 16755 15745
rect 16795 15705 16805 15745
rect 16845 15705 16855 15745
rect 16895 15705 16905 15745
rect 16945 15705 16955 15745
rect 16995 15705 17005 15745
rect 17045 15705 17055 15745
rect 17095 15705 17105 15745
rect 17145 15705 17155 15745
rect 17195 15705 17205 15745
rect 17245 15705 17255 15745
rect 17295 15705 17305 15745
rect 17345 15705 17355 15745
rect 17395 15705 17405 15745
rect 17445 15705 17455 15745
rect 17495 15705 17505 15745
rect 17545 15705 17555 15745
rect 17595 15705 17605 15745
rect 17645 15705 17655 15745
rect 17695 15705 17705 15745
rect 17745 15705 17755 15745
rect 17795 15705 17805 15745
rect 17845 15705 17855 15745
rect 17895 15705 17905 15745
rect 17945 15705 17955 15745
rect 17995 15705 18005 15745
rect 18045 15705 18055 15745
rect 18095 15705 18105 15745
rect 18145 15705 18155 15745
rect 18195 15705 18205 15745
rect 18245 15705 18255 15745
rect 18295 15705 18305 15745
rect 18345 15705 18355 15745
rect 18395 15705 18405 15745
rect 18445 15705 18455 15745
rect 18495 15705 18505 15745
rect 18545 15705 18555 15745
rect 18595 15705 18605 15745
rect 18645 15705 18655 15745
rect 18695 15705 18705 15745
rect 18745 15705 18755 15745
rect 18795 15705 18805 15745
rect 18845 15705 18855 15745
rect 18895 15705 18905 15745
rect 18945 15705 18955 15745
rect 18995 15705 19005 15745
rect 19045 15705 19055 15745
rect 19095 15705 19105 15745
rect 19145 15705 19155 15745
rect 19195 15705 19205 15745
rect 19245 15705 19255 15745
rect 19295 15705 19305 15745
rect 19345 15705 19355 15745
rect 19395 15705 19405 15745
rect 19445 15705 19455 15745
rect 19495 15705 19505 15745
rect 19545 15705 19555 15745
rect 19595 15705 19605 15745
rect 19645 15705 19655 15745
rect 19695 15705 19705 15745
rect 19745 15705 19755 15745
rect 19795 15705 19805 15745
rect 19845 15705 19855 15745
rect 19895 15705 19905 15745
rect 19945 15705 19955 15745
rect 19995 15705 20005 15745
rect 20045 15705 20055 15745
rect 20095 15705 20105 15745
rect 20145 15705 20155 15745
rect 20195 15705 20205 15745
rect 20245 15705 20255 15745
rect 20295 15705 20305 15745
rect 20345 15705 20355 15745
rect 20395 15705 20405 15745
rect 20445 15705 20455 15745
rect 20495 15705 20505 15745
rect 20545 15705 20555 15745
rect 20595 15705 20605 15745
rect 20645 15705 20655 15745
rect 20695 15705 20705 15745
rect 20745 15705 20755 15745
rect 20795 15705 20805 15745
rect 20845 15705 20855 15745
rect 20895 15705 20905 15745
rect 20945 15705 20955 15745
rect 20995 15705 21005 15745
rect 21045 15705 21055 15745
rect 21095 15705 21105 15745
rect 21145 15705 21155 15745
rect 21195 15705 21205 15745
rect 21245 15705 21255 15745
rect 21295 15705 21305 15745
rect 21345 15705 21355 15745
rect 21395 15705 21405 15745
rect 21445 15705 21455 15745
rect 21495 15705 21505 15745
rect 21545 15705 21555 15745
rect 21595 15705 21605 15745
rect 21645 15705 21655 15745
rect 21695 15705 21705 15745
rect 21745 15705 21755 15745
rect 21795 15705 21805 15745
rect 21845 15705 21855 15745
rect 21895 15705 21905 15745
rect 21945 15705 21955 15745
rect 21995 15705 22005 15745
rect 22045 15705 22055 15745
rect 22095 15705 22105 15745
rect 22145 15705 22155 15745
rect 22195 15705 22205 15745
rect 22245 15705 22255 15745
rect 22295 15705 22305 15745
rect 22345 15705 22355 15745
rect 22395 15705 22405 15745
rect 22445 15705 22455 15745
rect 22495 15705 22505 15745
rect 22545 15705 22555 15745
rect 22595 15705 22605 15745
rect 22645 15705 22655 15745
rect 22695 15705 22705 15745
rect 22745 15705 22755 15745
rect 22795 15705 22805 15745
rect 22845 15705 22855 15745
rect 22895 15705 22905 15745
rect 22945 15705 22955 15745
rect 22995 15705 23005 15745
rect 23045 15705 23055 15745
rect 23095 15705 23105 15745
rect 23145 15705 23155 15745
rect 23195 15705 23205 15745
rect 23245 15705 23255 15745
rect 23295 15705 23305 15745
rect 23345 15705 23355 15745
rect 23395 15705 23405 15745
rect 23445 15705 23455 15745
rect 23495 15705 23505 15745
rect 23545 15705 23555 15745
rect 23595 15705 23605 15745
rect 23645 15705 23655 15745
rect 23695 15705 23705 15745
rect 23745 15705 23755 15745
rect 23795 15705 23805 15745
rect 23845 15705 23855 15745
rect 23895 15705 23905 15745
rect 23945 15705 23955 15745
rect 23995 15705 24005 15745
rect 24045 15705 24055 15745
rect 24095 15705 24105 15745
rect 24145 15705 24155 15745
rect 24195 15705 24205 15745
rect 24245 15705 24255 15745
rect 24295 15705 24305 15745
rect 24345 15705 24355 15745
rect 24395 15705 24405 15745
rect 24445 15705 24455 15745
rect 24495 15705 24505 15745
rect 24545 15705 24555 15745
rect 24595 15705 24605 15745
rect 24645 15705 24655 15745
rect 24695 15705 24705 15745
rect 24745 15705 24755 15745
rect 24795 15705 24805 15745
rect 24845 15705 24855 15745
rect 24895 15705 24905 15745
rect 24945 15705 24955 15745
rect 24995 15705 25005 15745
rect 25045 15705 25055 15745
rect 25095 15705 25105 15745
rect 25145 15705 25155 15745
rect 25195 15705 25205 15745
rect 25245 15705 25255 15745
rect 25295 15705 25305 15745
rect 25345 15705 25355 15745
rect 25395 15705 25405 15745
rect 25445 15705 25455 15745
rect 25495 15705 25505 15745
rect 25545 15705 25555 15745
rect 25595 15705 25605 15745
rect 25645 15705 25655 15745
rect 25695 15705 25705 15745
rect 25745 15705 25755 15745
rect 25795 15705 25805 15745
rect 25845 15705 25855 15745
rect 25895 15705 25905 15745
rect 25945 15705 25955 15745
rect 25995 15705 26005 15745
rect 26045 15705 26055 15745
rect 26095 15705 26105 15745
rect 26145 15705 26155 15745
rect 26195 15705 26205 15745
rect 26245 15705 26255 15745
rect 26295 15705 26305 15745
rect 26345 15705 26355 15745
rect 26395 15705 26405 15745
rect 26445 15705 26455 15745
rect 26495 15705 26505 15745
rect 26545 15705 26555 15745
rect 26595 15705 26605 15745
rect 26645 15705 26655 15745
rect 26695 15705 26705 15745
rect 26745 15705 26755 15745
rect 26795 15705 26805 15745
rect 26845 15705 26855 15745
rect 26895 15705 26905 15745
rect 26945 15705 26955 15745
rect 26995 15705 27005 15745
rect 27045 15705 27055 15745
rect 27095 15705 27105 15745
rect 27145 15705 27155 15745
rect 27195 15705 27205 15745
rect 27245 15705 27255 15745
rect 27295 15705 27305 15745
rect 27345 15705 27355 15745
rect 27395 15705 27405 15745
rect 27445 15705 27455 15745
rect 27495 15705 27505 15745
rect 27545 15705 27555 15745
rect 27595 15705 27605 15745
rect 27645 15705 27655 15745
rect 27695 15705 27705 15745
rect 27745 15705 27755 15745
rect 27795 15705 27805 15745
rect 27845 15705 27855 15745
rect 27895 15705 27905 15745
rect 27945 15705 27955 15745
rect 27995 15705 28005 15745
rect 28045 15705 28055 15745
rect 28095 15705 28105 15745
rect 28145 15705 28155 15745
rect 28195 15705 28205 15745
rect 28245 15705 28255 15745
rect 28295 15705 28305 15745
rect 28345 15705 28355 15745
rect 28395 15705 28405 15745
rect 28445 15705 28455 15745
rect 28495 15705 28505 15745
rect 28545 15705 28555 15745
rect 28595 15705 28605 15745
rect 28645 15705 28655 15745
rect 28695 15705 28705 15745
rect 28745 15705 28755 15745
rect 28795 15705 28805 15745
rect 28845 15705 28855 15745
rect 28895 15705 28905 15745
rect 28945 15705 28955 15745
rect 28995 15705 29005 15745
rect 29045 15705 29055 15745
rect 29095 15705 29105 15745
rect 29145 15705 29155 15745
rect 29195 15705 29205 15745
rect 29245 15705 29255 15745
rect 29295 15705 29305 15745
rect 29345 15705 29355 15745
rect 29395 15705 29405 15745
rect 29445 15705 29455 15745
rect 29495 15705 29505 15745
rect 29545 15705 29555 15745
rect 29595 15705 29605 15745
rect 29645 15705 29655 15745
rect 29695 15705 29705 15745
rect 29745 15705 29755 15745
rect 29795 15705 29805 15745
rect 29845 15705 29855 15745
rect 29895 15705 29905 15745
rect 29945 15705 29955 15745
rect 29995 15705 30005 15745
rect 30045 15705 30055 15745
rect 30095 15705 30105 15745
rect 30145 15705 30155 15745
rect 30195 15705 30205 15745
rect 30245 15705 30255 15745
rect 30295 15705 30305 15745
rect 30345 15705 30355 15745
rect 30395 15705 30405 15745
rect 30445 15705 30455 15745
rect 30495 15705 30505 15745
rect 30545 15705 30555 15745
rect 30595 15705 30605 15745
rect 30645 15705 30655 15745
rect 30695 15705 30705 15745
rect 30745 15705 30755 15745
rect 30795 15705 30805 15745
rect 30845 15705 30855 15745
rect 30895 15705 30905 15745
rect 30945 15705 30955 15745
rect 30995 15705 31005 15745
rect 31045 15705 31055 15745
rect 31095 15705 31105 15745
rect 31145 15705 31155 15745
rect 31195 15705 31205 15745
rect 31245 15705 31255 15745
rect 31295 15705 31305 15745
rect 31345 15705 31355 15745
rect 31395 15705 31405 15745
rect 31445 15705 31455 15745
rect 31495 15705 31505 15745
rect 31545 15705 31555 15745
rect 31595 15705 31605 15745
rect 31645 15705 31655 15745
rect 31695 15705 31705 15745
rect 31745 15705 31755 15745
rect 31795 15705 31805 15745
rect 31845 15705 31855 15745
rect 31895 15705 31905 15745
rect 31945 15705 31955 15745
rect 31995 15705 32005 15745
rect 32045 15705 32055 15745
rect 32095 15705 32105 15745
rect 32145 15705 32155 15745
rect 32195 15705 32205 15745
rect 32245 15705 32255 15745
rect 32295 15705 32305 15745
rect 32345 15705 32355 15745
rect 32395 15705 32405 15745
rect 32445 15705 32455 15745
rect 32495 15705 32505 15745
rect 32545 15705 32555 15745
rect 32595 15705 32605 15745
rect 32645 15705 32655 15745
rect 32695 15705 32705 15745
rect 32745 15705 32755 15745
rect 32795 15705 32805 15745
rect 32845 15705 32855 15745
rect 32895 15705 32905 15745
rect 32945 15705 32955 15745
rect 32995 15705 33005 15745
rect 33045 15705 33055 15745
rect 33095 15705 33105 15745
rect 33145 15705 33155 15745
rect 33195 15705 33205 15745
rect 33245 15705 33255 15745
rect 33295 15705 33305 15745
rect 33345 15705 33355 15745
rect 33395 15705 33405 15745
rect 33445 15705 33455 15745
rect 33495 15705 33505 15745
rect 33545 15705 33555 15745
rect 33595 15705 33605 15745
rect 33645 15705 33655 15745
rect 33695 15705 33705 15745
rect 33745 15705 33755 15745
rect 33795 15705 33805 15745
rect 33845 15705 33855 15745
rect 33895 15705 33905 15745
rect 33945 15705 33955 15745
rect 33995 15705 34005 15745
rect 34045 15705 34055 15745
rect 34095 15705 34105 15745
rect 34145 15705 34155 15745
rect 34195 15705 34205 15745
rect 34245 15705 34255 15745
rect 34295 15705 34305 15745
rect 34345 15705 34355 15745
rect 34395 15705 34405 15745
rect 34445 15705 34455 15745
rect 34495 15705 34505 15745
rect 34545 15705 34555 15745
rect 34595 15705 34605 15745
rect 34645 15705 34655 15745
rect 34695 15705 34705 15745
rect 34745 15705 34755 15745
rect 34795 15705 34805 15745
rect 34845 15705 34855 15745
rect 34895 15705 34905 15745
rect 34945 15705 34955 15745
rect 34995 15705 35005 15745
rect 35045 15705 35055 15745
rect 35095 15705 35105 15745
rect 35145 15705 35155 15745
rect 35195 15705 35205 15745
rect 35245 15705 35255 15745
rect 35295 15705 35305 15745
rect 35345 15705 35355 15745
rect 35395 15705 35405 15745
rect 35445 15705 35455 15745
rect 35495 15705 35505 15745
rect 35545 15705 35555 15745
rect 35595 15705 35605 15745
rect 35645 15705 35655 15745
rect 35695 15705 35705 15745
rect 35745 15705 35755 15745
rect 35795 15705 35805 15745
rect 35845 15705 35855 15745
rect 35895 15705 35905 15745
rect 35945 15705 35955 15745
rect 35995 15705 36005 15745
rect 36045 15705 36055 15745
rect 36095 15705 36105 15745
rect 36145 15705 36155 15745
rect 36195 15705 36205 15745
rect 36245 15705 36255 15745
rect 36295 15705 36305 15745
rect 36345 15705 36355 15745
rect 36395 15705 36405 15745
rect 36445 15705 36455 15745
rect 36495 15705 36505 15745
rect 36545 15705 36555 15745
rect 36595 15705 36605 15745
rect 36645 15705 36655 15745
rect 36695 15705 36705 15745
rect 36745 15705 36755 15745
rect 36795 15705 36805 15745
rect 36845 15705 36855 15745
rect 36895 15705 36905 15745
rect 36945 15705 36955 15745
rect 36995 15705 37005 15745
rect 37045 15705 37055 15745
rect 37095 15705 37105 15745
rect 37145 15705 37155 15745
rect 37195 15705 37205 15745
rect 37245 15705 37255 15745
rect 37295 15705 37305 15745
rect 37345 15705 37355 15745
rect 37395 15705 37405 15745
rect 37445 15705 37455 15745
rect 37495 15705 37505 15745
rect 37545 15705 37555 15745
rect 37595 15705 37605 15745
rect 37645 15705 37655 15745
rect 37695 15705 37705 15745
rect 37745 15705 37755 15745
rect 37795 15705 37805 15745
rect 37845 15705 37855 15745
rect 37895 15705 37905 15745
rect 37945 15705 37955 15745
rect 37995 15705 38005 15745
rect 38045 15705 38055 15745
rect 38095 15705 38105 15745
rect 38145 15705 38155 15745
rect 38195 15705 38205 15745
rect 38245 15705 38255 15745
rect 38295 15705 38305 15745
rect 38345 15705 38355 15745
rect 38395 15705 38405 15745
rect 38445 15705 38455 15745
rect 38495 15705 38505 15745
rect 38545 15705 38555 15745
rect 38595 15705 38605 15745
rect 38645 15705 38655 15745
rect 38695 15705 38705 15745
rect 38745 15705 38755 15745
rect 38795 15705 38805 15745
rect 38845 15705 38855 15745
rect 38895 15705 38905 15745
rect 38945 15705 38955 15745
rect 38995 15705 39005 15745
rect 39045 15705 39055 15745
rect 39095 15705 39105 15745
rect 39145 15705 39155 15745
rect 39195 15705 39205 15745
rect 39245 15705 39255 15745
rect 39295 15705 39305 15745
rect 39345 15705 39355 15745
rect 39395 15705 39405 15745
rect 39445 15705 39455 15745
rect 39495 15705 39505 15745
rect 39545 15705 39555 15745
rect 39595 15705 39605 15745
rect 39645 15705 39655 15745
rect 39695 15705 39705 15745
rect 39745 15705 39905 15745
rect 39945 15705 39955 15745
rect 39995 15705 40005 15745
rect 40045 15705 40055 15745
rect 40095 15705 40105 15745
rect 40145 15705 40155 15745
rect 40195 15705 40205 15745
rect 40245 15705 40255 15745
rect 40295 15705 40305 15745
rect 40345 15705 40355 15745
rect 40395 15705 40405 15745
rect 40445 15705 40455 15745
rect 40495 15705 40505 15745
rect 40545 15705 40555 15745
rect 40595 15705 40605 15745
rect 40645 15705 40655 15745
rect 40695 15705 40705 15745
rect 40745 15705 40755 15745
rect 40795 15705 40805 15745
rect 40845 15705 40855 15745
rect 40895 15705 40900 15745
rect 0 15700 40900 15705
rect -3500 15345 0 15350
rect -3500 15305 -3495 15345
rect -3455 15305 -3295 15345
rect -3255 15305 -3095 15345
rect -3055 15305 -1595 15345
rect -1555 15305 -1095 15345
rect -1055 15305 -895 15345
rect -855 15305 -695 15345
rect -655 15305 -495 15345
rect -455 15305 -295 15345
rect -255 15305 -95 15345
rect -55 15305 0 15345
rect -3500 15295 0 15305
rect -3500 15255 -3495 15295
rect -3455 15255 -3295 15295
rect -3255 15255 -3095 15295
rect -3055 15255 -1595 15295
rect -1555 15255 -1095 15295
rect -1055 15255 -895 15295
rect -855 15255 -695 15295
rect -655 15255 -495 15295
rect -455 15255 -295 15295
rect -255 15255 -95 15295
rect -55 15255 0 15295
rect -3500 15245 0 15255
rect -3500 15205 -3495 15245
rect -3455 15205 -3295 15245
rect -3255 15205 -3095 15245
rect -3055 15205 -1595 15245
rect -1555 15205 -1095 15245
rect -1055 15205 -895 15245
rect -855 15205 -695 15245
rect -655 15205 -495 15245
rect -455 15205 -295 15245
rect -255 15205 -95 15245
rect -55 15205 0 15245
rect -3500 15200 0 15205
rect -200 14645 0 14650
rect -200 14605 -195 14645
rect -155 14605 0 14645
rect -200 14600 0 14605
rect -400 14245 0 14250
rect -400 14205 -395 14245
rect -355 14205 0 14245
rect -400 14200 0 14205
rect -600 14045 0 14050
rect -600 14005 -595 14045
rect -555 14005 0 14045
rect -600 14000 0 14005
rect -3500 13645 0 13650
rect -3500 13605 -3495 13645
rect -3455 13605 -3295 13645
rect -3255 13605 -3095 13645
rect -3055 13605 -1595 13645
rect -1555 13605 -1095 13645
rect -1055 13605 -895 13645
rect -855 13605 -695 13645
rect -655 13605 -495 13645
rect -455 13605 -295 13645
rect -255 13605 -95 13645
rect -55 13605 0 13645
rect -3500 13595 0 13605
rect -3500 13555 -3495 13595
rect -3455 13555 -3295 13595
rect -3255 13555 -3095 13595
rect -3055 13555 -1595 13595
rect -1555 13555 -1095 13595
rect -1055 13555 -895 13595
rect -855 13555 -695 13595
rect -655 13555 -495 13595
rect -455 13555 -295 13595
rect -255 13555 -95 13595
rect -55 13555 0 13595
rect -3500 13545 0 13555
rect -3500 13505 -3495 13545
rect -3455 13505 -3295 13545
rect -3255 13505 -3095 13545
rect -3055 13505 -1595 13545
rect -1555 13505 -1095 13545
rect -1055 13505 -895 13545
rect -855 13505 -695 13545
rect -655 13505 -495 13545
rect -455 13505 -295 13545
rect -255 13505 -95 13545
rect -55 13505 0 13545
rect -3500 13500 0 13505
rect -800 13145 0 13150
rect -800 13105 -795 13145
rect -755 13105 0 13145
rect -800 13100 0 13105
rect -1000 12945 0 12950
rect -1000 12905 -995 12945
rect -955 12905 0 12945
rect -1000 12900 0 12905
rect -1200 12545 0 12550
rect -1200 12505 -1195 12545
rect -1155 12505 0 12545
rect -1200 12500 0 12505
rect -1300 12445 0 12450
rect -1300 12405 -1295 12445
rect -1255 12405 0 12445
rect -1300 12400 0 12405
rect -1400 12345 0 12350
rect -1400 12305 -1395 12345
rect -1355 12305 0 12345
rect -1400 12300 0 12305
rect -1500 12245 0 12250
rect -1500 12205 -1495 12245
rect -1455 12205 0 12245
rect -1500 12200 0 12205
rect -3500 11945 0 11950
rect -3500 11905 -3495 11945
rect -3455 11905 -3295 11945
rect -3255 11905 -3095 11945
rect -3055 11905 -1595 11945
rect -1555 11905 -1095 11945
rect -1055 11905 -895 11945
rect -855 11905 -695 11945
rect -655 11905 -495 11945
rect -455 11905 -295 11945
rect -255 11905 -95 11945
rect -55 11905 0 11945
rect -3500 11895 0 11905
rect -3500 11855 -3495 11895
rect -3455 11855 -3295 11895
rect -3255 11855 -3095 11895
rect -3055 11855 -1595 11895
rect -1555 11855 -1095 11895
rect -1055 11855 -895 11895
rect -855 11855 -695 11895
rect -655 11855 -495 11895
rect -455 11855 -295 11895
rect -255 11855 -95 11895
rect -55 11855 0 11895
rect -3500 11845 0 11855
rect -3500 11805 -3495 11845
rect -3455 11805 -3295 11845
rect -3255 11805 -3095 11845
rect -3055 11805 -1595 11845
rect -1555 11805 -1095 11845
rect -1055 11805 -895 11845
rect -855 11805 -695 11845
rect -655 11805 -495 11845
rect -455 11805 -295 11845
rect -255 11805 -95 11845
rect -55 11805 0 11845
rect -3500 11800 0 11805
rect -3200 11445 0 11450
rect -3200 11405 -3195 11445
rect -3155 11405 0 11445
rect -3200 11400 0 11405
rect 39750 11345 39900 11350
rect 39750 11305 39805 11345
rect 39845 11305 39900 11345
rect 39750 11300 39900 11305
rect 39750 11245 40900 11250
rect 39750 11205 39905 11245
rect 39945 11205 39955 11245
rect 39995 11205 40005 11245
rect 40045 11205 40055 11245
rect 40095 11205 40105 11245
rect 40145 11205 40155 11245
rect 40195 11205 40205 11245
rect 40245 11205 40255 11245
rect 40295 11205 40305 11245
rect 40345 11205 40355 11245
rect 40395 11205 40405 11245
rect 40445 11205 40455 11245
rect 40495 11205 40505 11245
rect 40545 11205 40555 11245
rect 40595 11205 40605 11245
rect 40645 11205 40655 11245
rect 40695 11205 40705 11245
rect 40745 11205 40755 11245
rect 40795 11205 40805 11245
rect 40845 11205 40855 11245
rect 40895 11205 40900 11245
rect 39750 11195 40900 11205
rect 39750 11155 39905 11195
rect 39945 11155 39955 11195
rect 39995 11155 40005 11195
rect 40045 11155 40055 11195
rect 40095 11155 40105 11195
rect 40145 11155 40155 11195
rect 40195 11155 40205 11195
rect 40245 11155 40255 11195
rect 40295 11155 40305 11195
rect 40345 11155 40355 11195
rect 40395 11155 40405 11195
rect 40445 11155 40455 11195
rect 40495 11155 40505 11195
rect 40545 11155 40555 11195
rect 40595 11155 40605 11195
rect 40645 11155 40655 11195
rect 40695 11155 40705 11195
rect 40745 11155 40755 11195
rect 40795 11155 40805 11195
rect 40845 11155 40855 11195
rect 40895 11155 40900 11195
rect 39750 11145 40900 11155
rect 39750 11105 39905 11145
rect 39945 11105 39955 11145
rect 39995 11105 40005 11145
rect 40045 11105 40055 11145
rect 40095 11105 40105 11145
rect 40145 11105 40155 11145
rect 40195 11105 40205 11145
rect 40245 11105 40255 11145
rect 40295 11105 40305 11145
rect 40345 11105 40355 11145
rect 40395 11105 40405 11145
rect 40445 11105 40455 11145
rect 40495 11105 40505 11145
rect 40545 11105 40555 11145
rect 40595 11105 40605 11145
rect 40645 11105 40655 11145
rect 40695 11105 40705 11145
rect 40745 11105 40755 11145
rect 40795 11105 40805 11145
rect 40845 11105 40855 11145
rect 40895 11105 40900 11145
rect 39750 11095 40900 11105
rect 39750 11055 39905 11095
rect 39945 11055 39955 11095
rect 39995 11055 40005 11095
rect 40045 11055 40055 11095
rect 40095 11055 40105 11095
rect 40145 11055 40155 11095
rect 40195 11055 40205 11095
rect 40245 11055 40255 11095
rect 40295 11055 40305 11095
rect 40345 11055 40355 11095
rect 40395 11055 40405 11095
rect 40445 11055 40455 11095
rect 40495 11055 40505 11095
rect 40545 11055 40555 11095
rect 40595 11055 40605 11095
rect 40645 11055 40655 11095
rect 40695 11055 40705 11095
rect 40745 11055 40755 11095
rect 40795 11055 40805 11095
rect 40845 11055 40855 11095
rect 40895 11055 40900 11095
rect 39750 11045 40900 11055
rect 39750 11005 39905 11045
rect 39945 11005 39955 11045
rect 39995 11005 40005 11045
rect 40045 11005 40055 11045
rect 40095 11005 40105 11045
rect 40145 11005 40155 11045
rect 40195 11005 40205 11045
rect 40245 11005 40255 11045
rect 40295 11005 40305 11045
rect 40345 11005 40355 11045
rect 40395 11005 40405 11045
rect 40445 11005 40455 11045
rect 40495 11005 40505 11045
rect 40545 11005 40555 11045
rect 40595 11005 40605 11045
rect 40645 11005 40655 11045
rect 40695 11005 40705 11045
rect 40745 11005 40755 11045
rect 40795 11005 40805 11045
rect 40845 11005 40855 11045
rect 40895 11005 40900 11045
rect 39750 11000 40900 11005
rect 39750 10945 39900 10950
rect 39750 10905 39805 10945
rect 39845 10905 39900 10945
rect 39750 10900 39900 10905
rect -3400 10845 0 10850
rect -3400 10805 -3395 10845
rect -3355 10805 0 10845
rect -3400 10800 0 10805
rect -3100 10645 0 10650
rect -3100 10605 -2995 10645
rect -2955 10605 -2795 10645
rect -2755 10605 -2595 10645
rect -2555 10605 -2395 10645
rect -2355 10605 -2195 10645
rect -2155 10605 -1995 10645
rect -1955 10605 -1695 10645
rect -1655 10605 0 10645
rect -3100 10595 0 10605
rect -3100 10555 -2995 10595
rect -2955 10555 -2795 10595
rect -2755 10555 -2595 10595
rect -2555 10555 -2395 10595
rect -2355 10555 -2195 10595
rect -2155 10555 -1995 10595
rect -1955 10555 -1695 10595
rect -1655 10555 0 10595
rect -3100 10545 0 10555
rect -3100 10505 -2995 10545
rect -2955 10505 -2795 10545
rect -2755 10505 -2595 10545
rect -2555 10505 -2395 10545
rect -2355 10505 -2195 10545
rect -2155 10505 -1995 10545
rect -1955 10505 -1695 10545
rect -1655 10505 0 10545
rect -3100 10500 0 10505
rect -1800 10245 0 10250
rect -1800 10205 -1795 10245
rect -1755 10205 0 10245
rect -1800 10200 0 10205
rect -1900 10145 0 10150
rect -1900 10105 -1895 10145
rect -1855 10105 0 10145
rect -1900 10100 0 10105
rect -2100 9745 0 9750
rect -2100 9705 -2095 9745
rect -2055 9705 0 9745
rect -2100 9700 0 9705
rect -2300 9545 0 9550
rect -2300 9505 -2295 9545
rect -2255 9505 0 9545
rect -2300 9500 0 9505
rect -3100 9345 0 9350
rect -3100 9305 -2995 9345
rect -2955 9305 -2795 9345
rect -2755 9305 -2595 9345
rect -2555 9305 -2395 9345
rect -2355 9305 -2195 9345
rect -2155 9305 -1995 9345
rect -1955 9305 -1695 9345
rect -1655 9305 0 9345
rect -3100 9295 0 9305
rect -3100 9255 -2995 9295
rect -2955 9255 -2795 9295
rect -2755 9255 -2595 9295
rect -2555 9255 -2395 9295
rect -2355 9255 -2195 9295
rect -2155 9255 -1995 9295
rect -1955 9255 -1695 9295
rect -1655 9255 0 9295
rect -3100 9245 0 9255
rect -3100 9205 -2995 9245
rect -2955 9205 -2795 9245
rect -2755 9205 -2595 9245
rect -2555 9205 -2395 9245
rect -2355 9205 -2195 9245
rect -2155 9205 -1995 9245
rect -1955 9205 -1695 9245
rect -1655 9205 0 9245
rect -3100 9200 0 9205
rect -2500 9045 0 9050
rect -2500 9005 -2495 9045
rect -2455 9005 0 9045
rect -2500 9000 0 9005
rect -2700 8845 0 8850
rect -2700 8805 -2695 8845
rect -2655 8805 0 8845
rect -2700 8800 0 8805
rect -2900 8445 0 8450
rect -2900 8405 -2895 8445
rect -2855 8405 0 8445
rect -2900 8400 0 8405
rect -3100 8045 0 8050
rect -3100 8005 -2995 8045
rect -2955 8005 -2795 8045
rect -2755 8005 -2595 8045
rect -2555 8005 -2395 8045
rect -2355 8005 -2195 8045
rect -2155 8005 -1995 8045
rect -1955 8005 -1695 8045
rect -1655 8005 0 8045
rect -3100 7995 0 8005
rect -3100 7955 -2995 7995
rect -2955 7955 -2795 7995
rect -2755 7955 -2595 7995
rect -2555 7955 -2395 7995
rect -2355 7955 -2195 7995
rect -2155 7955 -1995 7995
rect -1955 7955 -1695 7995
rect -1655 7955 0 7995
rect -3100 7945 0 7955
rect -3100 7905 -2995 7945
rect -2955 7905 -2795 7945
rect -2755 7905 -2595 7945
rect -2555 7905 -2395 7945
rect -2355 7905 -2195 7945
rect -2155 7905 -1995 7945
rect -1955 7905 -1695 7945
rect -1655 7905 0 7945
rect -3100 7900 0 7905
rect -3100 7745 0 7750
rect -3100 7705 -2995 7745
rect -2955 7705 -2795 7745
rect -2755 7705 -2595 7745
rect -2555 7705 -2395 7745
rect -2355 7705 -2195 7745
rect -2155 7705 -1995 7745
rect -1955 7705 -1695 7745
rect -1655 7705 0 7745
rect -3100 7695 0 7705
rect -3100 7655 -2995 7695
rect -2955 7655 -2795 7695
rect -2755 7655 -2595 7695
rect -2555 7655 -2395 7695
rect -2355 7655 -2195 7695
rect -2155 7655 -1995 7695
rect -1955 7655 -1695 7695
rect -1655 7655 0 7695
rect -3100 7645 0 7655
rect -3100 7605 -2995 7645
rect -2955 7605 -2795 7645
rect -2755 7605 -2595 7645
rect -2555 7605 -2395 7645
rect -2355 7605 -2195 7645
rect -2155 7605 -1995 7645
rect -1955 7605 -1695 7645
rect -1655 7605 0 7645
rect -3100 7600 0 7605
rect -2900 7245 0 7250
rect -2900 7205 -2895 7245
rect -2855 7205 0 7245
rect -2900 7200 0 7205
rect -2700 6845 0 6850
rect -2700 6805 -2695 6845
rect -2655 6805 0 6845
rect -2700 6800 0 6805
rect -2500 6645 0 6650
rect -2500 6605 -2495 6645
rect -2455 6605 0 6645
rect -2500 6600 0 6605
rect -3100 6445 0 6450
rect -3100 6405 -2995 6445
rect -2955 6405 -2795 6445
rect -2755 6405 -2595 6445
rect -2555 6405 -2395 6445
rect -2355 6405 -2195 6445
rect -2155 6405 -1995 6445
rect -1955 6405 -1695 6445
rect -1655 6405 0 6445
rect -3100 6395 0 6405
rect -3100 6355 -2995 6395
rect -2955 6355 -2795 6395
rect -2755 6355 -2595 6395
rect -2555 6355 -2395 6395
rect -2355 6355 -2195 6395
rect -2155 6355 -1995 6395
rect -1955 6355 -1695 6395
rect -1655 6355 0 6395
rect -3100 6345 0 6355
rect -3100 6305 -2995 6345
rect -2955 6305 -2795 6345
rect -2755 6305 -2595 6345
rect -2555 6305 -2395 6345
rect -2355 6305 -2195 6345
rect -2155 6305 -1995 6345
rect -1955 6305 -1695 6345
rect -1655 6305 0 6345
rect -3100 6300 0 6305
rect -2300 6145 0 6150
rect -2300 6105 -2295 6145
rect -2255 6105 0 6145
rect -2300 6100 0 6105
rect -2100 5945 0 5950
rect -2100 5905 -2095 5945
rect -2055 5905 0 5945
rect -2100 5900 0 5905
rect -1900 5545 0 5550
rect -1900 5505 -1895 5545
rect -1855 5505 0 5545
rect -1900 5500 0 5505
rect -1800 5445 0 5450
rect -1800 5405 -1795 5445
rect -1755 5405 0 5445
rect -1800 5400 0 5405
rect -3100 5145 0 5150
rect -3100 5105 -2995 5145
rect -2955 5105 -2795 5145
rect -2755 5105 -2595 5145
rect -2555 5105 -2395 5145
rect -2355 5105 -2195 5145
rect -2155 5105 -1995 5145
rect -1955 5105 -1695 5145
rect -1655 5105 0 5145
rect -3100 5095 0 5105
rect -3100 5055 -2995 5095
rect -2955 5055 -2795 5095
rect -2755 5055 -2595 5095
rect -2555 5055 -2395 5095
rect -2355 5055 -2195 5095
rect -2155 5055 -1995 5095
rect -1955 5055 -1695 5095
rect -1655 5055 0 5095
rect -3100 5045 0 5055
rect -3100 5005 -2995 5045
rect -2955 5005 -2795 5045
rect -2755 5005 -2595 5045
rect -2555 5005 -2395 5045
rect -2355 5005 -2195 5045
rect -2155 5005 -1995 5045
rect -1955 5005 -1695 5045
rect -1655 5005 0 5045
rect -3100 5000 0 5005
rect -3400 4845 0 4850
rect -3400 4805 -3395 4845
rect -3355 4805 0 4845
rect -3400 4800 0 4805
rect 39750 4745 39900 4750
rect 39750 4705 39805 4745
rect 39845 4705 39900 4745
rect 39750 4700 39900 4705
rect 39750 4645 40900 4650
rect 39750 4605 39905 4645
rect 39945 4605 39955 4645
rect 39995 4605 40005 4645
rect 40045 4605 40055 4645
rect 40095 4605 40105 4645
rect 40145 4605 40155 4645
rect 40195 4605 40205 4645
rect 40245 4605 40255 4645
rect 40295 4605 40305 4645
rect 40345 4605 40355 4645
rect 40395 4605 40405 4645
rect 40445 4605 40455 4645
rect 40495 4605 40505 4645
rect 40545 4605 40555 4645
rect 40595 4605 40605 4645
rect 40645 4605 40655 4645
rect 40695 4605 40705 4645
rect 40745 4605 40755 4645
rect 40795 4605 40805 4645
rect 40845 4605 40855 4645
rect 40895 4605 40900 4645
rect 39750 4595 40900 4605
rect 39750 4555 39905 4595
rect 39945 4555 39955 4595
rect 39995 4555 40005 4595
rect 40045 4555 40055 4595
rect 40095 4555 40105 4595
rect 40145 4555 40155 4595
rect 40195 4555 40205 4595
rect 40245 4555 40255 4595
rect 40295 4555 40305 4595
rect 40345 4555 40355 4595
rect 40395 4555 40405 4595
rect 40445 4555 40455 4595
rect 40495 4555 40505 4595
rect 40545 4555 40555 4595
rect 40595 4555 40605 4595
rect 40645 4555 40655 4595
rect 40695 4555 40705 4595
rect 40745 4555 40755 4595
rect 40795 4555 40805 4595
rect 40845 4555 40855 4595
rect 40895 4555 40900 4595
rect 39750 4545 40900 4555
rect 39750 4505 39905 4545
rect 39945 4505 39955 4545
rect 39995 4505 40005 4545
rect 40045 4505 40055 4545
rect 40095 4505 40105 4545
rect 40145 4505 40155 4545
rect 40195 4505 40205 4545
rect 40245 4505 40255 4545
rect 40295 4505 40305 4545
rect 40345 4505 40355 4545
rect 40395 4505 40405 4545
rect 40445 4505 40455 4545
rect 40495 4505 40505 4545
rect 40545 4505 40555 4545
rect 40595 4505 40605 4545
rect 40645 4505 40655 4545
rect 40695 4505 40705 4545
rect 40745 4505 40755 4545
rect 40795 4505 40805 4545
rect 40845 4505 40855 4545
rect 40895 4505 40900 4545
rect 39750 4495 40900 4505
rect 39750 4455 39905 4495
rect 39945 4455 39955 4495
rect 39995 4455 40005 4495
rect 40045 4455 40055 4495
rect 40095 4455 40105 4495
rect 40145 4455 40155 4495
rect 40195 4455 40205 4495
rect 40245 4455 40255 4495
rect 40295 4455 40305 4495
rect 40345 4455 40355 4495
rect 40395 4455 40405 4495
rect 40445 4455 40455 4495
rect 40495 4455 40505 4495
rect 40545 4455 40555 4495
rect 40595 4455 40605 4495
rect 40645 4455 40655 4495
rect 40695 4455 40705 4495
rect 40745 4455 40755 4495
rect 40795 4455 40805 4495
rect 40845 4455 40855 4495
rect 40895 4455 40900 4495
rect 39750 4445 40900 4455
rect 39750 4405 39905 4445
rect 39945 4405 39955 4445
rect 39995 4405 40005 4445
rect 40045 4405 40055 4445
rect 40095 4405 40105 4445
rect 40145 4405 40155 4445
rect 40195 4405 40205 4445
rect 40245 4405 40255 4445
rect 40295 4405 40305 4445
rect 40345 4405 40355 4445
rect 40395 4405 40405 4445
rect 40445 4405 40455 4445
rect 40495 4405 40505 4445
rect 40545 4405 40555 4445
rect 40595 4405 40605 4445
rect 40645 4405 40655 4445
rect 40695 4405 40705 4445
rect 40745 4405 40755 4445
rect 40795 4405 40805 4445
rect 40845 4405 40855 4445
rect 40895 4405 40900 4445
rect 39750 4400 40900 4405
rect 39750 4345 39900 4350
rect 39750 4305 39805 4345
rect 39845 4305 39900 4345
rect 39750 4300 39900 4305
rect -3200 4245 0 4250
rect -3200 4205 -3195 4245
rect -3155 4205 0 4245
rect -3200 4200 0 4205
rect -3500 3845 0 3850
rect -3500 3805 -3495 3845
rect -3455 3805 -3295 3845
rect -3255 3805 -3095 3845
rect -3055 3805 -1595 3845
rect -1555 3805 -1095 3845
rect -1055 3805 -895 3845
rect -855 3805 -695 3845
rect -655 3805 -495 3845
rect -455 3805 -295 3845
rect -255 3805 -95 3845
rect -55 3805 0 3845
rect -3500 3795 0 3805
rect -3500 3755 -3495 3795
rect -3455 3755 -3295 3795
rect -3255 3755 -3095 3795
rect -3055 3755 -1595 3795
rect -1555 3755 -1095 3795
rect -1055 3755 -895 3795
rect -855 3755 -695 3795
rect -655 3755 -495 3795
rect -455 3755 -295 3795
rect -255 3755 -95 3795
rect -55 3755 0 3795
rect -3500 3745 0 3755
rect -3500 3705 -3495 3745
rect -3455 3705 -3295 3745
rect -3255 3705 -3095 3745
rect -3055 3705 -1595 3745
rect -1555 3705 -1095 3745
rect -1055 3705 -895 3745
rect -855 3705 -695 3745
rect -655 3705 -495 3745
rect -455 3705 -295 3745
rect -255 3705 -95 3745
rect -55 3705 0 3745
rect -3500 3700 0 3705
rect -1500 3445 0 3450
rect -1500 3405 -1495 3445
rect -1455 3405 0 3445
rect -1500 3400 0 3405
rect -1400 3345 0 3350
rect -1400 3305 -1395 3345
rect -1355 3305 0 3345
rect -1400 3300 0 3305
rect -1300 3245 0 3250
rect -1300 3205 -1295 3245
rect -1255 3205 0 3245
rect -1300 3200 0 3205
rect -1200 3145 0 3150
rect -1200 3105 -1195 3145
rect -1155 3105 0 3145
rect -1200 3100 0 3105
rect -1000 2745 0 2750
rect -1000 2705 -995 2745
rect -955 2705 0 2745
rect -1000 2700 0 2705
rect -800 2545 0 2550
rect -800 2505 -795 2545
rect -755 2505 0 2545
rect -800 2500 0 2505
rect -3500 2145 0 2150
rect -3500 2105 -3495 2145
rect -3455 2105 -3295 2145
rect -3255 2105 -3095 2145
rect -3055 2105 -1595 2145
rect -1555 2105 -1095 2145
rect -1055 2105 -895 2145
rect -855 2105 -695 2145
rect -655 2105 -495 2145
rect -455 2105 -295 2145
rect -255 2105 -95 2145
rect -55 2105 0 2145
rect -3500 2095 0 2105
rect -3500 2055 -3495 2095
rect -3455 2055 -3295 2095
rect -3255 2055 -3095 2095
rect -3055 2055 -1595 2095
rect -1555 2055 -1095 2095
rect -1055 2055 -895 2095
rect -855 2055 -695 2095
rect -655 2055 -495 2095
rect -455 2055 -295 2095
rect -255 2055 -95 2095
rect -55 2055 0 2095
rect -3500 2045 0 2055
rect -3500 2005 -3495 2045
rect -3455 2005 -3295 2045
rect -3255 2005 -3095 2045
rect -3055 2005 -1595 2045
rect -1555 2005 -1095 2045
rect -1055 2005 -895 2045
rect -855 2005 -695 2045
rect -655 2005 -495 2045
rect -455 2005 -295 2045
rect -255 2005 -95 2045
rect -55 2005 0 2045
rect -3500 2000 0 2005
rect -600 1645 0 1650
rect -600 1605 -595 1645
rect -555 1605 0 1645
rect -600 1600 0 1605
rect -400 1445 0 1450
rect -400 1405 -395 1445
rect -355 1405 0 1445
rect -400 1400 0 1405
rect -200 1045 0 1050
rect -200 1005 -195 1045
rect -155 1005 0 1045
rect -200 1000 0 1005
rect -3500 445 0 450
rect -3500 405 -3495 445
rect -3455 405 -3295 445
rect -3255 405 -3095 445
rect -3055 405 -1595 445
rect -1555 405 -1095 445
rect -1055 405 -895 445
rect -855 405 -695 445
rect -655 405 -495 445
rect -455 405 -295 445
rect -255 405 -95 445
rect -55 405 0 445
rect -3500 395 0 405
rect -3500 355 -3495 395
rect -3455 355 -3295 395
rect -3255 355 -3095 395
rect -3055 355 -1595 395
rect -1555 355 -1095 395
rect -1055 355 -895 395
rect -855 355 -695 395
rect -655 355 -495 395
rect -455 355 -295 395
rect -255 355 -95 395
rect -55 355 0 395
rect -3500 345 0 355
rect -3500 305 -3495 345
rect -3455 305 -3295 345
rect -3255 305 -3095 345
rect -3055 305 -1595 345
rect -1555 305 -1095 345
rect -1055 305 -895 345
rect -855 305 -695 345
rect -655 305 -495 345
rect -455 305 -295 345
rect -255 305 -95 345
rect -55 305 0 345
rect -3500 300 0 305
<< via3 >>
rect 5 18245 45 18285
rect 55 18245 95 18285
rect 105 18245 145 18285
rect 155 18245 195 18285
rect 205 18245 245 18285
rect 255 18245 295 18285
rect 305 18245 345 18285
rect 355 18245 395 18285
rect 405 18245 445 18285
rect 455 18245 495 18285
rect 505 18245 545 18285
rect 555 18245 595 18285
rect 605 18245 645 18285
rect 655 18245 695 18285
rect 705 18245 745 18285
rect 755 18245 795 18285
rect 805 18245 845 18285
rect 855 18245 895 18285
rect 905 18245 945 18285
rect 955 18245 995 18285
rect 1005 18245 1045 18285
rect 1055 18245 1095 18285
rect 1105 18245 1145 18285
rect 1155 18245 1195 18285
rect 1205 18245 1245 18285
rect 1255 18245 1295 18285
rect 1305 18245 1345 18285
rect 1355 18245 1395 18285
rect 1405 18245 1445 18285
rect 1455 18245 1495 18285
rect 1505 18245 1545 18285
rect 1555 18245 1595 18285
rect 1605 18245 1645 18285
rect 1655 18245 1695 18285
rect 1705 18245 1745 18285
rect 1755 18245 1795 18285
rect 1805 18245 1845 18285
rect 1855 18245 1895 18285
rect 1905 18245 1945 18285
rect 1955 18245 1995 18285
rect 2005 18245 2045 18285
rect 2055 18245 2095 18285
rect 2105 18245 2145 18285
rect 2155 18245 2195 18285
rect 2205 18245 2245 18285
rect 2255 18245 2295 18285
rect 2305 18245 2345 18285
rect 2355 18245 2395 18285
rect 2405 18245 2445 18285
rect 2455 18245 2495 18285
rect 2505 18245 2545 18285
rect 2555 18245 2595 18285
rect 2605 18245 2645 18285
rect 2655 18245 2695 18285
rect 2705 18245 2745 18285
rect 2755 18245 2795 18285
rect 2805 18245 2845 18285
rect 2855 18245 2895 18285
rect 2905 18245 2945 18285
rect 2955 18245 2995 18285
rect 3005 18245 3045 18285
rect 3055 18245 3095 18285
rect 3105 18245 3145 18285
rect 3155 18245 3195 18285
rect 3205 18245 3245 18285
rect 3255 18245 3295 18285
rect 3305 18245 3345 18285
rect 3355 18245 3395 18285
rect 3405 18245 3445 18285
rect 3455 18245 3495 18285
rect 3505 18245 3545 18285
rect 3555 18245 3595 18285
rect 3605 18245 3645 18285
rect 3655 18245 3695 18285
rect 3705 18245 3745 18285
rect 3755 18245 3795 18285
rect 3805 18245 3845 18285
rect 3855 18245 3895 18285
rect 3905 18245 3945 18285
rect 3955 18245 3995 18285
rect 4005 18245 4045 18285
rect 4055 18245 4095 18285
rect 4105 18245 4145 18285
rect 4155 18245 4195 18285
rect 4205 18245 4245 18285
rect 4255 18245 4295 18285
rect 4305 18245 4345 18285
rect 4355 18245 4395 18285
rect 4405 18245 4445 18285
rect 4455 18245 4495 18285
rect 4505 18245 4545 18285
rect 4555 18245 4595 18285
rect 4605 18245 4645 18285
rect 4655 18245 4695 18285
rect 4705 18245 4745 18285
rect 4755 18245 4795 18285
rect 4805 18245 4845 18285
rect 4855 18245 4895 18285
rect 4905 18245 4945 18285
rect 4955 18245 4995 18285
rect 5005 18245 5045 18285
rect 5055 18245 5095 18285
rect 5105 18245 5145 18285
rect 5155 18245 5195 18285
rect 5205 18245 5245 18285
rect 5255 18245 5295 18285
rect 5305 18245 5345 18285
rect 5355 18245 5395 18285
rect 5405 18245 5445 18285
rect 5455 18245 5495 18285
rect 5505 18245 5545 18285
rect 5555 18245 5595 18285
rect 5605 18245 5645 18285
rect 5655 18245 5695 18285
rect 5705 18245 5745 18285
rect 5755 18245 5795 18285
rect 5805 18245 5845 18285
rect 5855 18245 5895 18285
rect 5905 18245 5945 18285
rect 5955 18245 5995 18285
rect 6005 18245 6045 18285
rect 6055 18245 6095 18285
rect 6105 18245 6145 18285
rect 6155 18245 6195 18285
rect 6205 18245 6245 18285
rect 6255 18245 6295 18285
rect 6305 18245 6345 18285
rect 6355 18245 6395 18285
rect 6405 18245 6445 18285
rect 6455 18245 6495 18285
rect 6505 18245 6545 18285
rect 6555 18245 6595 18285
rect 6605 18245 6645 18285
rect 6655 18245 6695 18285
rect 6705 18245 6745 18285
rect 6755 18245 6795 18285
rect 6805 18245 6845 18285
rect 6855 18245 6895 18285
rect 6905 18245 6945 18285
rect 6955 18245 6995 18285
rect 7005 18245 7045 18285
rect 7055 18245 7095 18285
rect 7105 18245 7145 18285
rect 7155 18245 7195 18285
rect 7205 18245 7245 18285
rect 7255 18245 7295 18285
rect 7305 18245 7345 18285
rect 7355 18245 7395 18285
rect 7405 18245 7445 18285
rect 7455 18245 7495 18285
rect 7505 18245 7545 18285
rect 7555 18245 7595 18285
rect 7605 18245 7645 18285
rect 7655 18245 7695 18285
rect 7705 18245 7745 18285
rect 7755 18245 7795 18285
rect 7805 18245 7845 18285
rect 7855 18245 7895 18285
rect 7905 18245 7945 18285
rect 7955 18245 7995 18285
rect 8005 18245 8045 18285
rect 8055 18245 8095 18285
rect 8105 18245 8145 18285
rect 8155 18245 8195 18285
rect 8205 18245 8245 18285
rect 8255 18245 8295 18285
rect 8305 18245 8345 18285
rect 8355 18245 8395 18285
rect 8405 18245 8445 18285
rect 8455 18245 8495 18285
rect 8505 18245 8545 18285
rect 8555 18245 8595 18285
rect 8605 18245 8645 18285
rect 8655 18245 8695 18285
rect 8705 18245 8745 18285
rect 8755 18245 8795 18285
rect 8805 18245 8845 18285
rect 8855 18245 8895 18285
rect 8905 18245 8945 18285
rect 8955 18245 8995 18285
rect 9005 18245 9045 18285
rect 9055 18245 9095 18285
rect 9105 18245 9145 18285
rect 9155 18245 9195 18285
rect 9205 18245 9245 18285
rect 9255 18245 9295 18285
rect 9305 18245 9345 18285
rect 9355 18245 9395 18285
rect 9405 18245 9445 18285
rect 9455 18245 9495 18285
rect 9505 18245 9545 18285
rect 9555 18245 9595 18285
rect 9605 18245 9645 18285
rect 9655 18245 9695 18285
rect 9705 18245 9745 18285
rect 9755 18245 9795 18285
rect 9805 18245 9845 18285
rect 9855 18245 9895 18285
rect 9905 18245 9945 18285
rect 9955 18245 9995 18285
rect 10005 18245 10045 18285
rect 10055 18245 10095 18285
rect 10105 18245 10145 18285
rect 10155 18245 10195 18285
rect 10205 18245 10245 18285
rect 10255 18245 10295 18285
rect 10305 18245 10345 18285
rect 10355 18245 10395 18285
rect 10405 18245 10445 18285
rect 10455 18245 10495 18285
rect 10505 18245 10545 18285
rect 10555 18245 10595 18285
rect 10605 18245 10645 18285
rect 10655 18245 10695 18285
rect 10705 18245 10745 18285
rect 10755 18245 10795 18285
rect 10805 18245 10845 18285
rect 10855 18245 10895 18285
rect 10905 18245 10945 18285
rect 10955 18245 10995 18285
rect 11005 18245 11045 18285
rect 11055 18245 11095 18285
rect 11105 18245 11145 18285
rect 11155 18245 11195 18285
rect 11205 18245 11245 18285
rect 11255 18245 11295 18285
rect 11305 18245 11345 18285
rect 11355 18245 11395 18285
rect 11405 18245 11445 18285
rect 11455 18245 11495 18285
rect 11505 18245 11545 18285
rect 11555 18245 11595 18285
rect 11605 18245 11645 18285
rect 11655 18245 11695 18285
rect 11705 18245 11745 18285
rect 11755 18245 11795 18285
rect 11805 18245 11845 18285
rect 11855 18245 11895 18285
rect 11905 18245 11945 18285
rect 11955 18245 11995 18285
rect 12005 18245 12045 18285
rect 12055 18245 12095 18285
rect 12105 18245 12145 18285
rect 12155 18245 12195 18285
rect 12205 18245 12245 18285
rect 12255 18245 12295 18285
rect 12305 18245 12345 18285
rect 12355 18245 12395 18285
rect 12405 18245 12445 18285
rect 12455 18245 12495 18285
rect 12505 18245 12545 18285
rect 12555 18245 12595 18285
rect 12605 18245 12645 18285
rect 12655 18245 12695 18285
rect 12705 18245 12745 18285
rect 12755 18245 12795 18285
rect 12805 18245 12845 18285
rect 12855 18245 12895 18285
rect 12905 18245 12945 18285
rect 12955 18245 12995 18285
rect 13005 18245 13045 18285
rect 13055 18245 13095 18285
rect 13105 18245 13145 18285
rect 13155 18245 13195 18285
rect 13205 18245 13245 18285
rect 13255 18245 13295 18285
rect 13305 18245 13345 18285
rect 13355 18245 13395 18285
rect 13405 18245 13445 18285
rect 13455 18245 13495 18285
rect 13505 18245 13545 18285
rect 13555 18245 13595 18285
rect 13605 18245 13645 18285
rect 13655 18245 13695 18285
rect 13705 18245 13745 18285
rect 13755 18245 13795 18285
rect 13805 18245 13845 18285
rect 13855 18245 13895 18285
rect 13905 18245 13945 18285
rect 13955 18245 13995 18285
rect 14005 18245 14045 18285
rect 14055 18245 14095 18285
rect 14105 18245 14145 18285
rect 14155 18245 14195 18285
rect 14205 18245 14245 18285
rect 14255 18245 14295 18285
rect 14305 18245 14345 18285
rect 14355 18245 14395 18285
rect 14405 18245 14445 18285
rect 14455 18245 14495 18285
rect 14505 18245 14545 18285
rect 14555 18245 14595 18285
rect 14605 18245 14645 18285
rect 14655 18245 14695 18285
rect 14705 18245 14745 18285
rect 14755 18245 14795 18285
rect 14805 18245 14845 18285
rect 14855 18245 14895 18285
rect 14905 18245 14945 18285
rect 14955 18245 14995 18285
rect 15005 18245 15045 18285
rect 15055 18245 15095 18285
rect 15105 18245 15145 18285
rect 15155 18245 15195 18285
rect 15205 18245 15245 18285
rect 15255 18245 15295 18285
rect 15305 18245 15345 18285
rect 15355 18245 15395 18285
rect 15405 18245 15445 18285
rect 15455 18245 15495 18285
rect 15505 18245 15545 18285
rect 15555 18245 15595 18285
rect 15605 18245 15645 18285
rect 15655 18245 15695 18285
rect 15705 18245 15745 18285
rect 15755 18245 15795 18285
rect 15805 18245 15845 18285
rect 15855 18245 15895 18285
rect 15905 18245 15945 18285
rect 15955 18245 15995 18285
rect 16005 18245 16045 18285
rect 16055 18245 16095 18285
rect 16105 18245 16145 18285
rect 16155 18245 16195 18285
rect 16205 18245 16245 18285
rect 16255 18245 16295 18285
rect 16305 18245 16345 18285
rect 16355 18245 16395 18285
rect 16405 18245 16445 18285
rect 16455 18245 16495 18285
rect 16505 18245 16545 18285
rect 16555 18245 16595 18285
rect 16605 18245 16645 18285
rect 16655 18245 16695 18285
rect 16705 18245 16745 18285
rect 16755 18245 16795 18285
rect 16805 18245 16845 18285
rect 16855 18245 16895 18285
rect 16905 18245 16945 18285
rect 16955 18245 16995 18285
rect 17005 18245 17045 18285
rect 17055 18245 17095 18285
rect 17105 18245 17145 18285
rect 17155 18245 17195 18285
rect 17205 18245 17245 18285
rect 17255 18245 17295 18285
rect 17305 18245 17345 18285
rect 17355 18245 17395 18285
rect 17405 18245 17445 18285
rect 17455 18245 17495 18285
rect 17505 18245 17545 18285
rect 17555 18245 17595 18285
rect 17605 18245 17645 18285
rect 17655 18245 17695 18285
rect 17705 18245 17745 18285
rect 17755 18245 17795 18285
rect 17805 18245 17845 18285
rect 17855 18245 17895 18285
rect 17905 18245 17945 18285
rect 17955 18245 17995 18285
rect 18005 18245 18045 18285
rect 18055 18245 18095 18285
rect 18105 18245 18145 18285
rect 18155 18245 18195 18285
rect 18205 18245 18245 18285
rect 18255 18245 18295 18285
rect 18305 18245 18345 18285
rect 18355 18245 18395 18285
rect 18405 18245 18445 18285
rect 18455 18245 18495 18285
rect 18505 18245 18545 18285
rect 18555 18245 18595 18285
rect 18605 18245 18645 18285
rect 18655 18245 18695 18285
rect 18705 18245 18745 18285
rect 18755 18245 18795 18285
rect 18805 18245 18845 18285
rect 18855 18245 18895 18285
rect 18905 18245 18945 18285
rect 18955 18245 18995 18285
rect 19005 18245 19045 18285
rect 19055 18245 19095 18285
rect 19105 18245 19145 18285
rect 19155 18245 19195 18285
rect 19205 18245 19245 18285
rect 19255 18245 19295 18285
rect 19305 18245 19345 18285
rect 19355 18245 19395 18285
rect 19405 18245 19445 18285
rect 19455 18245 19495 18285
rect 19505 18245 19545 18285
rect 19555 18245 19595 18285
rect 19605 18245 19645 18285
rect 19655 18245 19695 18285
rect 19705 18245 19745 18285
rect 19755 18245 19795 18285
rect 19805 18245 19845 18285
rect 19855 18245 19895 18285
rect 19905 18245 19945 18285
rect 19955 18245 19995 18285
rect 20005 18245 20045 18285
rect 20055 18245 20095 18285
rect 20105 18245 20145 18285
rect 20155 18245 20195 18285
rect 20205 18245 20245 18285
rect 20255 18245 20295 18285
rect 20305 18245 20345 18285
rect 20355 18245 20395 18285
rect 20405 18245 20445 18285
rect 20455 18245 20495 18285
rect 20505 18245 20545 18285
rect 20555 18245 20595 18285
rect 20605 18245 20645 18285
rect 20655 18245 20695 18285
rect 20705 18245 20745 18285
rect 20755 18245 20795 18285
rect 20805 18245 20845 18285
rect 20855 18245 20895 18285
rect 20905 18245 20945 18285
rect 20955 18245 20995 18285
rect 21005 18245 21045 18285
rect 21055 18245 21095 18285
rect 21105 18245 21145 18285
rect 21155 18245 21195 18285
rect 21205 18245 21245 18285
rect 21255 18245 21295 18285
rect 21305 18245 21345 18285
rect 21355 18245 21395 18285
rect 21405 18245 21445 18285
rect 21455 18245 21495 18285
rect 21505 18245 21545 18285
rect 21555 18245 21595 18285
rect 21605 18245 21645 18285
rect 21655 18245 21695 18285
rect 21705 18245 21745 18285
rect 21755 18245 21795 18285
rect 21805 18245 21845 18285
rect 21855 18245 21895 18285
rect 21905 18245 21945 18285
rect 21955 18245 21995 18285
rect 22005 18245 22045 18285
rect 22055 18245 22095 18285
rect 22105 18245 22145 18285
rect 22155 18245 22195 18285
rect 22205 18245 22245 18285
rect 22255 18245 22295 18285
rect 22305 18245 22345 18285
rect 22355 18245 22395 18285
rect 22405 18245 22445 18285
rect 22455 18245 22495 18285
rect 22505 18245 22545 18285
rect 22555 18245 22595 18285
rect 22605 18245 22645 18285
rect 22655 18245 22695 18285
rect 22705 18245 22745 18285
rect 22755 18245 22795 18285
rect 22805 18245 22845 18285
rect 22855 18245 22895 18285
rect 22905 18245 22945 18285
rect 22955 18245 22995 18285
rect 23005 18245 23045 18285
rect 23055 18245 23095 18285
rect 23105 18245 23145 18285
rect 23155 18245 23195 18285
rect 23205 18245 23245 18285
rect 23255 18245 23295 18285
rect 23305 18245 23345 18285
rect 23355 18245 23395 18285
rect 23405 18245 23445 18285
rect 23455 18245 23495 18285
rect 23505 18245 23545 18285
rect 23555 18245 23595 18285
rect 23605 18245 23645 18285
rect 23655 18245 23695 18285
rect 23705 18245 23745 18285
rect 23755 18245 23795 18285
rect 23805 18245 23845 18285
rect 23855 18245 23895 18285
rect 23905 18245 23945 18285
rect 23955 18245 23995 18285
rect 24005 18245 24045 18285
rect 24055 18245 24095 18285
rect 24105 18245 24145 18285
rect 24155 18245 24195 18285
rect 24205 18245 24245 18285
rect 24255 18245 24295 18285
rect 24305 18245 24345 18285
rect 24355 18245 24395 18285
rect 24405 18245 24445 18285
rect 24455 18245 24495 18285
rect 24505 18245 24545 18285
rect 24555 18245 24595 18285
rect 24605 18245 24645 18285
rect 24655 18245 24695 18285
rect 24705 18245 24745 18285
rect 24755 18245 24795 18285
rect 24805 18245 24845 18285
rect 24855 18245 24895 18285
rect 24905 18245 24945 18285
rect 24955 18245 24995 18285
rect 25005 18245 25045 18285
rect 25055 18245 25095 18285
rect 25105 18245 25145 18285
rect 25155 18245 25195 18285
rect 25205 18245 25245 18285
rect 25255 18245 25295 18285
rect 25305 18245 25345 18285
rect 25355 18245 25395 18285
rect 25405 18245 25445 18285
rect 25455 18245 25495 18285
rect 25505 18245 25545 18285
rect 25555 18245 25595 18285
rect 25605 18245 25645 18285
rect 25655 18245 25695 18285
rect 25705 18245 25745 18285
rect 25755 18245 25795 18285
rect 25805 18245 25845 18285
rect 25855 18245 25895 18285
rect 25905 18245 25945 18285
rect 25955 18245 25995 18285
rect 26005 18245 26045 18285
rect 26055 18245 26095 18285
rect 26105 18245 26145 18285
rect 26155 18245 26195 18285
rect 26205 18245 26245 18285
rect 26255 18245 26295 18285
rect 26305 18245 26345 18285
rect 26355 18245 26395 18285
rect 26405 18245 26445 18285
rect 26455 18245 26495 18285
rect 26505 18245 26545 18285
rect 26555 18245 26595 18285
rect 26605 18245 26645 18285
rect 26655 18245 26695 18285
rect 26705 18245 26745 18285
rect 26755 18245 26795 18285
rect 26805 18245 26845 18285
rect 26855 18245 26895 18285
rect 26905 18245 26945 18285
rect 26955 18245 26995 18285
rect 27005 18245 27045 18285
rect 27055 18245 27095 18285
rect 27105 18245 27145 18285
rect 27155 18245 27195 18285
rect 27205 18245 27245 18285
rect 27255 18245 27295 18285
rect 27305 18245 27345 18285
rect 27355 18245 27395 18285
rect 27405 18245 27445 18285
rect 27455 18245 27495 18285
rect 27505 18245 27545 18285
rect 27555 18245 27595 18285
rect 27605 18245 27645 18285
rect 27655 18245 27695 18285
rect 27705 18245 27745 18285
rect 27755 18245 27795 18285
rect 27805 18245 27845 18285
rect 27855 18245 27895 18285
rect 27905 18245 27945 18285
rect 27955 18245 27995 18285
rect 28005 18245 28045 18285
rect 28055 18245 28095 18285
rect 28105 18245 28145 18285
rect 28155 18245 28195 18285
rect 28205 18245 28245 18285
rect 28255 18245 28295 18285
rect 28305 18245 28345 18285
rect 28355 18245 28395 18285
rect 28405 18245 28445 18285
rect 28455 18245 28495 18285
rect 28505 18245 28545 18285
rect 28555 18245 28595 18285
rect 28605 18245 28645 18285
rect 28655 18245 28695 18285
rect 28705 18245 28745 18285
rect 28755 18245 28795 18285
rect 28805 18245 28845 18285
rect 28855 18245 28895 18285
rect 28905 18245 28945 18285
rect 28955 18245 28995 18285
rect 29005 18245 29045 18285
rect 29055 18245 29095 18285
rect 29105 18245 29145 18285
rect 29155 18245 29195 18285
rect 29205 18245 29245 18285
rect 29255 18245 29295 18285
rect 29305 18245 29345 18285
rect 29355 18245 29395 18285
rect 29405 18245 29445 18285
rect 29455 18245 29495 18285
rect 29505 18245 29545 18285
rect 29555 18245 29595 18285
rect 29605 18245 29645 18285
rect 29655 18245 29695 18285
rect 29705 18245 29745 18285
rect 29755 18245 29795 18285
rect 29805 18245 29845 18285
rect 29855 18245 29895 18285
rect 29905 18245 29945 18285
rect 29955 18245 29995 18285
rect 30005 18245 30045 18285
rect 30055 18245 30095 18285
rect 30105 18245 30145 18285
rect 30155 18245 30195 18285
rect 30205 18245 30245 18285
rect 30255 18245 30295 18285
rect 30305 18245 30345 18285
rect 30355 18245 30395 18285
rect 30405 18245 30445 18285
rect 30455 18245 30495 18285
rect 30505 18245 30545 18285
rect 30555 18245 30595 18285
rect 30605 18245 30645 18285
rect 30655 18245 30695 18285
rect 30705 18245 30745 18285
rect 30755 18245 30795 18285
rect 30805 18245 30845 18285
rect 30855 18245 30895 18285
rect 30905 18245 30945 18285
rect 30955 18245 30995 18285
rect 31005 18245 31045 18285
rect 31055 18245 31095 18285
rect 31105 18245 31145 18285
rect 31155 18245 31195 18285
rect 31205 18245 31245 18285
rect 31255 18245 31295 18285
rect 31305 18245 31345 18285
rect 31355 18245 31395 18285
rect 31405 18245 31445 18285
rect 31455 18245 31495 18285
rect 31505 18245 31545 18285
rect 31555 18245 31595 18285
rect 31605 18245 31645 18285
rect 31655 18245 31695 18285
rect 31705 18245 31745 18285
rect 31755 18245 31795 18285
rect 31805 18245 31845 18285
rect 31855 18245 31895 18285
rect 31905 18245 31945 18285
rect 31955 18245 31995 18285
rect 32005 18245 32045 18285
rect 32055 18245 32095 18285
rect 32105 18245 32145 18285
rect 32155 18245 32195 18285
rect 32205 18245 32245 18285
rect 32255 18245 32295 18285
rect 32305 18245 32345 18285
rect 32355 18245 32395 18285
rect 32405 18245 32445 18285
rect 32455 18245 32495 18285
rect 32505 18245 32545 18285
rect 32555 18245 32595 18285
rect 32605 18245 32645 18285
rect 32655 18245 32695 18285
rect 32705 18245 32745 18285
rect 32755 18245 32795 18285
rect 32805 18245 32845 18285
rect 32855 18245 32895 18285
rect 32905 18245 32945 18285
rect 32955 18245 32995 18285
rect 33005 18245 33045 18285
rect 33055 18245 33095 18285
rect 33105 18245 33145 18285
rect 33155 18245 33195 18285
rect 33205 18245 33245 18285
rect 33255 18245 33295 18285
rect 33305 18245 33345 18285
rect 33355 18245 33395 18285
rect 33405 18245 33445 18285
rect 33455 18245 33495 18285
rect 33505 18245 33545 18285
rect 33555 18245 33595 18285
rect 33605 18245 33645 18285
rect 33655 18245 33695 18285
rect 33705 18245 33745 18285
rect 33755 18245 33795 18285
rect 33805 18245 33845 18285
rect 33855 18245 33895 18285
rect 33905 18245 33945 18285
rect 33955 18245 33995 18285
rect 34005 18245 34045 18285
rect 34055 18245 34095 18285
rect 34105 18245 34145 18285
rect 34155 18245 34195 18285
rect 34205 18245 34245 18285
rect 34255 18245 34295 18285
rect 34305 18245 34345 18285
rect 34355 18245 34395 18285
rect 34405 18245 34445 18285
rect 34455 18245 34495 18285
rect 34505 18245 34545 18285
rect 34555 18245 34595 18285
rect 34605 18245 34645 18285
rect 34655 18245 34695 18285
rect 34705 18245 34745 18285
rect 34755 18245 34795 18285
rect 34805 18245 34845 18285
rect 34855 18245 34895 18285
rect 34905 18245 34945 18285
rect 34955 18245 34995 18285
rect 35005 18245 35045 18285
rect 35055 18245 35095 18285
rect 35105 18245 35145 18285
rect 35155 18245 35195 18285
rect 35205 18245 35245 18285
rect 35255 18245 35295 18285
rect 35305 18245 35345 18285
rect 35355 18245 35395 18285
rect 35405 18245 35445 18285
rect 35455 18245 35495 18285
rect 35505 18245 35545 18285
rect 35555 18245 35595 18285
rect 35605 18245 35645 18285
rect 35655 18245 35695 18285
rect 35705 18245 35745 18285
rect 35755 18245 35795 18285
rect 35805 18245 35845 18285
rect 35855 18245 35895 18285
rect 35905 18245 35945 18285
rect 35955 18245 35995 18285
rect 36005 18245 36045 18285
rect 36055 18245 36095 18285
rect 36105 18245 36145 18285
rect 36155 18245 36195 18285
rect 36205 18245 36245 18285
rect 36255 18245 36295 18285
rect 36305 18245 36345 18285
rect 36355 18245 36395 18285
rect 36405 18245 36445 18285
rect 36455 18245 36495 18285
rect 36505 18245 36545 18285
rect 36555 18245 36595 18285
rect 36605 18245 36645 18285
rect 36655 18245 36695 18285
rect 36705 18245 36745 18285
rect 36755 18245 36795 18285
rect 36805 18245 36845 18285
rect 36855 18245 36895 18285
rect 36905 18245 36945 18285
rect 36955 18245 36995 18285
rect 37005 18245 37045 18285
rect 37055 18245 37095 18285
rect 37105 18245 37145 18285
rect 37155 18245 37195 18285
rect 37205 18245 37245 18285
rect 37255 18245 37295 18285
rect 37305 18245 37345 18285
rect 37355 18245 37395 18285
rect 37405 18245 37445 18285
rect 37455 18245 37495 18285
rect 37505 18245 37545 18285
rect 37555 18245 37595 18285
rect 37605 18245 37645 18285
rect 37655 18245 37695 18285
rect 37705 18245 37745 18285
rect 37755 18245 37795 18285
rect 37805 18245 37845 18285
rect 37855 18245 37895 18285
rect 37905 18245 37945 18285
rect 37955 18245 37995 18285
rect 38005 18245 38045 18285
rect 38055 18245 38095 18285
rect 38105 18245 38145 18285
rect 38155 18245 38195 18285
rect 38205 18245 38245 18285
rect 38255 18245 38295 18285
rect 38305 18245 38345 18285
rect 38355 18245 38395 18285
rect 38405 18245 38445 18285
rect 38455 18245 38495 18285
rect 38505 18245 38545 18285
rect 38555 18245 38595 18285
rect 38605 18245 38645 18285
rect 38655 18245 38695 18285
rect 38705 18245 38745 18285
rect 38755 18245 38795 18285
rect 38805 18245 38845 18285
rect 38855 18245 38895 18285
rect 38905 18245 38945 18285
rect 38955 18245 38995 18285
rect 39005 18245 39045 18285
rect 39055 18245 39095 18285
rect 39105 18245 39145 18285
rect 39155 18245 39195 18285
rect 39205 18245 39245 18285
rect 39255 18245 39295 18285
rect 39305 18245 39345 18285
rect 39355 18245 39395 18285
rect 39405 18245 39445 18285
rect 39455 18245 39495 18285
rect 39505 18245 39545 18285
rect 39555 18245 39595 18285
rect 39605 18245 39645 18285
rect 39655 18245 39695 18285
rect 39705 18245 39745 18285
rect 39905 18245 39945 18285
rect 39955 18245 39995 18285
rect 40005 18245 40045 18285
rect 40055 18245 40095 18285
rect 40105 18245 40145 18285
rect 40155 18245 40195 18285
rect 40205 18245 40245 18285
rect 40255 18245 40295 18285
rect 40305 18245 40345 18285
rect 40355 18245 40395 18285
rect 40405 18245 40445 18285
rect 40455 18245 40495 18285
rect 40505 18245 40545 18285
rect 40555 18245 40595 18285
rect 40605 18245 40645 18285
rect 40655 18245 40695 18285
rect 40705 18245 40745 18285
rect 40755 18245 40795 18285
rect 40805 18245 40845 18285
rect 40855 18245 40895 18285
rect 5 18145 45 18185
rect 55 18145 95 18185
rect 105 18145 145 18185
rect 155 18145 195 18185
rect 205 18145 245 18185
rect 255 18145 295 18185
rect 305 18145 345 18185
rect 355 18145 395 18185
rect 405 18145 445 18185
rect 455 18145 495 18185
rect 505 18145 545 18185
rect 555 18145 595 18185
rect 605 18145 645 18185
rect 655 18145 695 18185
rect 705 18145 745 18185
rect 755 18145 795 18185
rect 805 18145 845 18185
rect 855 18145 895 18185
rect 905 18145 945 18185
rect 955 18145 995 18185
rect 1005 18145 1045 18185
rect 1055 18145 1095 18185
rect 1105 18145 1145 18185
rect 1155 18145 1195 18185
rect 1205 18145 1245 18185
rect 1255 18145 1295 18185
rect 1305 18145 1345 18185
rect 1355 18145 1395 18185
rect 1405 18145 1445 18185
rect 1455 18145 1495 18185
rect 1505 18145 1545 18185
rect 1555 18145 1595 18185
rect 1605 18145 1645 18185
rect 1655 18145 1695 18185
rect 1705 18145 1745 18185
rect 1755 18145 1795 18185
rect 1805 18145 1845 18185
rect 1855 18145 1895 18185
rect 1905 18145 1945 18185
rect 1955 18145 1995 18185
rect 2005 18145 2045 18185
rect 2055 18145 2095 18185
rect 2105 18145 2145 18185
rect 2155 18145 2195 18185
rect 2205 18145 2245 18185
rect 2255 18145 2295 18185
rect 2305 18145 2345 18185
rect 2355 18145 2395 18185
rect 2405 18145 2445 18185
rect 2455 18145 2495 18185
rect 2505 18145 2545 18185
rect 2555 18145 2595 18185
rect 2605 18145 2645 18185
rect 2655 18145 2695 18185
rect 2705 18145 2745 18185
rect 2755 18145 2795 18185
rect 2805 18145 2845 18185
rect 2855 18145 2895 18185
rect 2905 18145 2945 18185
rect 2955 18145 2995 18185
rect 3005 18145 3045 18185
rect 3055 18145 3095 18185
rect 3105 18145 3145 18185
rect 3155 18145 3195 18185
rect 3205 18145 3245 18185
rect 3255 18145 3295 18185
rect 3305 18145 3345 18185
rect 3355 18145 3395 18185
rect 3405 18145 3445 18185
rect 3455 18145 3495 18185
rect 3505 18145 3545 18185
rect 3555 18145 3595 18185
rect 3605 18145 3645 18185
rect 3655 18145 3695 18185
rect 3705 18145 3745 18185
rect 3755 18145 3795 18185
rect 3805 18145 3845 18185
rect 3855 18145 3895 18185
rect 3905 18145 3945 18185
rect 3955 18145 3995 18185
rect 4005 18145 4045 18185
rect 4055 18145 4095 18185
rect 4105 18145 4145 18185
rect 4155 18145 4195 18185
rect 4205 18145 4245 18185
rect 4255 18145 4295 18185
rect 4305 18145 4345 18185
rect 4355 18145 4395 18185
rect 4405 18145 4445 18185
rect 4455 18145 4495 18185
rect 4505 18145 4545 18185
rect 4555 18145 4595 18185
rect 4605 18145 4645 18185
rect 4655 18145 4695 18185
rect 4705 18145 4745 18185
rect 4755 18145 4795 18185
rect 4805 18145 4845 18185
rect 4855 18145 4895 18185
rect 4905 18145 4945 18185
rect 4955 18145 4995 18185
rect 5005 18145 5045 18185
rect 5055 18145 5095 18185
rect 5105 18145 5145 18185
rect 5155 18145 5195 18185
rect 5205 18145 5245 18185
rect 5255 18145 5295 18185
rect 5305 18145 5345 18185
rect 5355 18145 5395 18185
rect 5405 18145 5445 18185
rect 5455 18145 5495 18185
rect 5505 18145 5545 18185
rect 5555 18145 5595 18185
rect 5605 18145 5645 18185
rect 5655 18145 5695 18185
rect 5705 18145 5745 18185
rect 5755 18145 5795 18185
rect 5805 18145 5845 18185
rect 5855 18145 5895 18185
rect 5905 18145 5945 18185
rect 5955 18145 5995 18185
rect 6005 18145 6045 18185
rect 6055 18145 6095 18185
rect 6105 18145 6145 18185
rect 6155 18145 6195 18185
rect 6205 18145 6245 18185
rect 6255 18145 6295 18185
rect 6305 18145 6345 18185
rect 6355 18145 6395 18185
rect 6405 18145 6445 18185
rect 6455 18145 6495 18185
rect 6505 18145 6545 18185
rect 6555 18145 6595 18185
rect 6605 18145 6645 18185
rect 6655 18145 6695 18185
rect 6705 18145 6745 18185
rect 6755 18145 6795 18185
rect 6805 18145 6845 18185
rect 6855 18145 6895 18185
rect 6905 18145 6945 18185
rect 6955 18145 6995 18185
rect 7005 18145 7045 18185
rect 7055 18145 7095 18185
rect 7105 18145 7145 18185
rect 7155 18145 7195 18185
rect 7205 18145 7245 18185
rect 7255 18145 7295 18185
rect 7305 18145 7345 18185
rect 7355 18145 7395 18185
rect 7405 18145 7445 18185
rect 7455 18145 7495 18185
rect 7505 18145 7545 18185
rect 7555 18145 7595 18185
rect 7605 18145 7645 18185
rect 7655 18145 7695 18185
rect 7705 18145 7745 18185
rect 7755 18145 7795 18185
rect 7805 18145 7845 18185
rect 7855 18145 7895 18185
rect 7905 18145 7945 18185
rect 7955 18145 7995 18185
rect 8005 18145 8045 18185
rect 8055 18145 8095 18185
rect 8105 18145 8145 18185
rect 8155 18145 8195 18185
rect 8205 18145 8245 18185
rect 8255 18145 8295 18185
rect 8305 18145 8345 18185
rect 8355 18145 8395 18185
rect 8405 18145 8445 18185
rect 8455 18145 8495 18185
rect 8505 18145 8545 18185
rect 8555 18145 8595 18185
rect 8605 18145 8645 18185
rect 8655 18145 8695 18185
rect 8705 18145 8745 18185
rect 8755 18145 8795 18185
rect 8805 18145 8845 18185
rect 8855 18145 8895 18185
rect 8905 18145 8945 18185
rect 8955 18145 8995 18185
rect 9005 18145 9045 18185
rect 9055 18145 9095 18185
rect 9105 18145 9145 18185
rect 9155 18145 9195 18185
rect 9205 18145 9245 18185
rect 9255 18145 9295 18185
rect 9305 18145 9345 18185
rect 9355 18145 9395 18185
rect 9405 18145 9445 18185
rect 9455 18145 9495 18185
rect 9505 18145 9545 18185
rect 9555 18145 9595 18185
rect 9605 18145 9645 18185
rect 9655 18145 9695 18185
rect 9705 18145 9745 18185
rect 9755 18145 9795 18185
rect 9805 18145 9845 18185
rect 9855 18145 9895 18185
rect 9905 18145 9945 18185
rect 9955 18145 9995 18185
rect 10005 18145 10045 18185
rect 10055 18145 10095 18185
rect 10105 18145 10145 18185
rect 10155 18145 10195 18185
rect 10205 18145 10245 18185
rect 10255 18145 10295 18185
rect 10305 18145 10345 18185
rect 10355 18145 10395 18185
rect 10405 18145 10445 18185
rect 10455 18145 10495 18185
rect 10505 18145 10545 18185
rect 10555 18145 10595 18185
rect 10605 18145 10645 18185
rect 10655 18145 10695 18185
rect 10705 18145 10745 18185
rect 10755 18145 10795 18185
rect 10805 18145 10845 18185
rect 10855 18145 10895 18185
rect 10905 18145 10945 18185
rect 10955 18145 10995 18185
rect 11005 18145 11045 18185
rect 11055 18145 11095 18185
rect 11105 18145 11145 18185
rect 11155 18145 11195 18185
rect 11205 18145 11245 18185
rect 11255 18145 11295 18185
rect 11305 18145 11345 18185
rect 11355 18145 11395 18185
rect 11405 18145 11445 18185
rect 11455 18145 11495 18185
rect 11505 18145 11545 18185
rect 11555 18145 11595 18185
rect 11605 18145 11645 18185
rect 11655 18145 11695 18185
rect 11705 18145 11745 18185
rect 11755 18145 11795 18185
rect 11805 18145 11845 18185
rect 11855 18145 11895 18185
rect 11905 18145 11945 18185
rect 11955 18145 11995 18185
rect 12005 18145 12045 18185
rect 12055 18145 12095 18185
rect 12105 18145 12145 18185
rect 12155 18145 12195 18185
rect 12205 18145 12245 18185
rect 12255 18145 12295 18185
rect 12305 18145 12345 18185
rect 12355 18145 12395 18185
rect 12405 18145 12445 18185
rect 12455 18145 12495 18185
rect 12505 18145 12545 18185
rect 12555 18145 12595 18185
rect 12605 18145 12645 18185
rect 12655 18145 12695 18185
rect 12705 18145 12745 18185
rect 12755 18145 12795 18185
rect 12805 18145 12845 18185
rect 12855 18145 12895 18185
rect 12905 18145 12945 18185
rect 12955 18145 12995 18185
rect 13005 18145 13045 18185
rect 13055 18145 13095 18185
rect 13105 18145 13145 18185
rect 13155 18145 13195 18185
rect 13205 18145 13245 18185
rect 13255 18145 13295 18185
rect 13305 18145 13345 18185
rect 13355 18145 13395 18185
rect 13405 18145 13445 18185
rect 13455 18145 13495 18185
rect 13505 18145 13545 18185
rect 13555 18145 13595 18185
rect 13605 18145 13645 18185
rect 13655 18145 13695 18185
rect 13705 18145 13745 18185
rect 13755 18145 13795 18185
rect 13805 18145 13845 18185
rect 13855 18145 13895 18185
rect 13905 18145 13945 18185
rect 13955 18145 13995 18185
rect 14005 18145 14045 18185
rect 14055 18145 14095 18185
rect 14105 18145 14145 18185
rect 14155 18145 14195 18185
rect 14205 18145 14245 18185
rect 14255 18145 14295 18185
rect 14305 18145 14345 18185
rect 14355 18145 14395 18185
rect 14405 18145 14445 18185
rect 14455 18145 14495 18185
rect 14505 18145 14545 18185
rect 14555 18145 14595 18185
rect 14605 18145 14645 18185
rect 14655 18145 14695 18185
rect 14705 18145 14745 18185
rect 14755 18145 14795 18185
rect 14805 18145 14845 18185
rect 14855 18145 14895 18185
rect 14905 18145 14945 18185
rect 14955 18145 14995 18185
rect 15005 18145 15045 18185
rect 15055 18145 15095 18185
rect 15105 18145 15145 18185
rect 15155 18145 15195 18185
rect 15205 18145 15245 18185
rect 15255 18145 15295 18185
rect 15305 18145 15345 18185
rect 15355 18145 15395 18185
rect 15405 18145 15445 18185
rect 15455 18145 15495 18185
rect 15505 18145 15545 18185
rect 15555 18145 15595 18185
rect 15605 18145 15645 18185
rect 15655 18145 15695 18185
rect 15705 18145 15745 18185
rect 15755 18145 15795 18185
rect 15805 18145 15845 18185
rect 15855 18145 15895 18185
rect 15905 18145 15945 18185
rect 15955 18145 15995 18185
rect 16005 18145 16045 18185
rect 16055 18145 16095 18185
rect 16105 18145 16145 18185
rect 16155 18145 16195 18185
rect 16205 18145 16245 18185
rect 16255 18145 16295 18185
rect 16305 18145 16345 18185
rect 16355 18145 16395 18185
rect 16405 18145 16445 18185
rect 16455 18145 16495 18185
rect 16505 18145 16545 18185
rect 16555 18145 16595 18185
rect 16605 18145 16645 18185
rect 16655 18145 16695 18185
rect 16705 18145 16745 18185
rect 16755 18145 16795 18185
rect 16805 18145 16845 18185
rect 16855 18145 16895 18185
rect 16905 18145 16945 18185
rect 16955 18145 16995 18185
rect 17005 18145 17045 18185
rect 17055 18145 17095 18185
rect 17105 18145 17145 18185
rect 17155 18145 17195 18185
rect 17205 18145 17245 18185
rect 17255 18145 17295 18185
rect 17305 18145 17345 18185
rect 17355 18145 17395 18185
rect 17405 18145 17445 18185
rect 17455 18145 17495 18185
rect 17505 18145 17545 18185
rect 17555 18145 17595 18185
rect 17605 18145 17645 18185
rect 17655 18145 17695 18185
rect 17705 18145 17745 18185
rect 17755 18145 17795 18185
rect 17805 18145 17845 18185
rect 17855 18145 17895 18185
rect 17905 18145 17945 18185
rect 17955 18145 17995 18185
rect 18005 18145 18045 18185
rect 18055 18145 18095 18185
rect 18105 18145 18145 18185
rect 18155 18145 18195 18185
rect 18205 18145 18245 18185
rect 18255 18145 18295 18185
rect 18305 18145 18345 18185
rect 18355 18145 18395 18185
rect 18405 18145 18445 18185
rect 18455 18145 18495 18185
rect 18505 18145 18545 18185
rect 18555 18145 18595 18185
rect 18605 18145 18645 18185
rect 18655 18145 18695 18185
rect 18705 18145 18745 18185
rect 18755 18145 18795 18185
rect 18805 18145 18845 18185
rect 18855 18145 18895 18185
rect 18905 18145 18945 18185
rect 18955 18145 18995 18185
rect 19005 18145 19045 18185
rect 19055 18145 19095 18185
rect 19105 18145 19145 18185
rect 19155 18145 19195 18185
rect 19205 18145 19245 18185
rect 19255 18145 19295 18185
rect 19305 18145 19345 18185
rect 19355 18145 19395 18185
rect 19405 18145 19445 18185
rect 19455 18145 19495 18185
rect 19505 18145 19545 18185
rect 19555 18145 19595 18185
rect 19605 18145 19645 18185
rect 19655 18145 19695 18185
rect 19705 18145 19745 18185
rect 19755 18145 19795 18185
rect 19805 18145 19845 18185
rect 19855 18145 19895 18185
rect 19905 18145 19945 18185
rect 19955 18145 19995 18185
rect 20005 18145 20045 18185
rect 20055 18145 20095 18185
rect 20105 18145 20145 18185
rect 20155 18145 20195 18185
rect 20205 18145 20245 18185
rect 20255 18145 20295 18185
rect 20305 18145 20345 18185
rect 20355 18145 20395 18185
rect 20405 18145 20445 18185
rect 20455 18145 20495 18185
rect 20505 18145 20545 18185
rect 20555 18145 20595 18185
rect 20605 18145 20645 18185
rect 20655 18145 20695 18185
rect 20705 18145 20745 18185
rect 20755 18145 20795 18185
rect 20805 18145 20845 18185
rect 20855 18145 20895 18185
rect 20905 18145 20945 18185
rect 20955 18145 20995 18185
rect 21005 18145 21045 18185
rect 21055 18145 21095 18185
rect 21105 18145 21145 18185
rect 21155 18145 21195 18185
rect 21205 18145 21245 18185
rect 21255 18145 21295 18185
rect 21305 18145 21345 18185
rect 21355 18145 21395 18185
rect 21405 18145 21445 18185
rect 21455 18145 21495 18185
rect 21505 18145 21545 18185
rect 21555 18145 21595 18185
rect 21605 18145 21645 18185
rect 21655 18145 21695 18185
rect 21705 18145 21745 18185
rect 21755 18145 21795 18185
rect 21805 18145 21845 18185
rect 21855 18145 21895 18185
rect 21905 18145 21945 18185
rect 21955 18145 21995 18185
rect 22005 18145 22045 18185
rect 22055 18145 22095 18185
rect 22105 18145 22145 18185
rect 22155 18145 22195 18185
rect 22205 18145 22245 18185
rect 22255 18145 22295 18185
rect 22305 18145 22345 18185
rect 22355 18145 22395 18185
rect 22405 18145 22445 18185
rect 22455 18145 22495 18185
rect 22505 18145 22545 18185
rect 22555 18145 22595 18185
rect 22605 18145 22645 18185
rect 22655 18145 22695 18185
rect 22705 18145 22745 18185
rect 22755 18145 22795 18185
rect 22805 18145 22845 18185
rect 22855 18145 22895 18185
rect 22905 18145 22945 18185
rect 22955 18145 22995 18185
rect 23005 18145 23045 18185
rect 23055 18145 23095 18185
rect 23105 18145 23145 18185
rect 23155 18145 23195 18185
rect 23205 18145 23245 18185
rect 23255 18145 23295 18185
rect 23305 18145 23345 18185
rect 23355 18145 23395 18185
rect 23405 18145 23445 18185
rect 23455 18145 23495 18185
rect 23505 18145 23545 18185
rect 23555 18145 23595 18185
rect 23605 18145 23645 18185
rect 23655 18145 23695 18185
rect 23705 18145 23745 18185
rect 23755 18145 23795 18185
rect 23805 18145 23845 18185
rect 23855 18145 23895 18185
rect 23905 18145 23945 18185
rect 23955 18145 23995 18185
rect 24005 18145 24045 18185
rect 24055 18145 24095 18185
rect 24105 18145 24145 18185
rect 24155 18145 24195 18185
rect 24205 18145 24245 18185
rect 24255 18145 24295 18185
rect 24305 18145 24345 18185
rect 24355 18145 24395 18185
rect 24405 18145 24445 18185
rect 24455 18145 24495 18185
rect 24505 18145 24545 18185
rect 24555 18145 24595 18185
rect 24605 18145 24645 18185
rect 24655 18145 24695 18185
rect 24705 18145 24745 18185
rect 24755 18145 24795 18185
rect 24805 18145 24845 18185
rect 24855 18145 24895 18185
rect 24905 18145 24945 18185
rect 24955 18145 24995 18185
rect 25005 18145 25045 18185
rect 25055 18145 25095 18185
rect 25105 18145 25145 18185
rect 25155 18145 25195 18185
rect 25205 18145 25245 18185
rect 25255 18145 25295 18185
rect 25305 18145 25345 18185
rect 25355 18145 25395 18185
rect 25405 18145 25445 18185
rect 25455 18145 25495 18185
rect 25505 18145 25545 18185
rect 25555 18145 25595 18185
rect 25605 18145 25645 18185
rect 25655 18145 25695 18185
rect 25705 18145 25745 18185
rect 25755 18145 25795 18185
rect 25805 18145 25845 18185
rect 25855 18145 25895 18185
rect 25905 18145 25945 18185
rect 25955 18145 25995 18185
rect 26005 18145 26045 18185
rect 26055 18145 26095 18185
rect 26105 18145 26145 18185
rect 26155 18145 26195 18185
rect 26205 18145 26245 18185
rect 26255 18145 26295 18185
rect 26305 18145 26345 18185
rect 26355 18145 26395 18185
rect 26405 18145 26445 18185
rect 26455 18145 26495 18185
rect 26505 18145 26545 18185
rect 26555 18145 26595 18185
rect 26605 18145 26645 18185
rect 26655 18145 26695 18185
rect 26705 18145 26745 18185
rect 26755 18145 26795 18185
rect 26805 18145 26845 18185
rect 26855 18145 26895 18185
rect 26905 18145 26945 18185
rect 26955 18145 26995 18185
rect 27005 18145 27045 18185
rect 27055 18145 27095 18185
rect 27105 18145 27145 18185
rect 27155 18145 27195 18185
rect 27205 18145 27245 18185
rect 27255 18145 27295 18185
rect 27305 18145 27345 18185
rect 27355 18145 27395 18185
rect 27405 18145 27445 18185
rect 27455 18145 27495 18185
rect 27505 18145 27545 18185
rect 27555 18145 27595 18185
rect 27605 18145 27645 18185
rect 27655 18145 27695 18185
rect 27705 18145 27745 18185
rect 27755 18145 27795 18185
rect 27805 18145 27845 18185
rect 27855 18145 27895 18185
rect 27905 18145 27945 18185
rect 27955 18145 27995 18185
rect 28005 18145 28045 18185
rect 28055 18145 28095 18185
rect 28105 18145 28145 18185
rect 28155 18145 28195 18185
rect 28205 18145 28245 18185
rect 28255 18145 28295 18185
rect 28305 18145 28345 18185
rect 28355 18145 28395 18185
rect 28405 18145 28445 18185
rect 28455 18145 28495 18185
rect 28505 18145 28545 18185
rect 28555 18145 28595 18185
rect 28605 18145 28645 18185
rect 28655 18145 28695 18185
rect 28705 18145 28745 18185
rect 28755 18145 28795 18185
rect 28805 18145 28845 18185
rect 28855 18145 28895 18185
rect 28905 18145 28945 18185
rect 28955 18145 28995 18185
rect 29005 18145 29045 18185
rect 29055 18145 29095 18185
rect 29105 18145 29145 18185
rect 29155 18145 29195 18185
rect 29205 18145 29245 18185
rect 29255 18145 29295 18185
rect 29305 18145 29345 18185
rect 29355 18145 29395 18185
rect 29405 18145 29445 18185
rect 29455 18145 29495 18185
rect 29505 18145 29545 18185
rect 29555 18145 29595 18185
rect 29605 18145 29645 18185
rect 29655 18145 29695 18185
rect 29705 18145 29745 18185
rect 29755 18145 29795 18185
rect 29805 18145 29845 18185
rect 29855 18145 29895 18185
rect 29905 18145 29945 18185
rect 29955 18145 29995 18185
rect 30005 18145 30045 18185
rect 30055 18145 30095 18185
rect 30105 18145 30145 18185
rect 30155 18145 30195 18185
rect 30205 18145 30245 18185
rect 30255 18145 30295 18185
rect 30305 18145 30345 18185
rect 30355 18145 30395 18185
rect 30405 18145 30445 18185
rect 30455 18145 30495 18185
rect 30505 18145 30545 18185
rect 30555 18145 30595 18185
rect 30605 18145 30645 18185
rect 30655 18145 30695 18185
rect 30705 18145 30745 18185
rect 30755 18145 30795 18185
rect 30805 18145 30845 18185
rect 30855 18145 30895 18185
rect 30905 18145 30945 18185
rect 30955 18145 30995 18185
rect 31005 18145 31045 18185
rect 31055 18145 31095 18185
rect 31105 18145 31145 18185
rect 31155 18145 31195 18185
rect 31205 18145 31245 18185
rect 31255 18145 31295 18185
rect 31305 18145 31345 18185
rect 31355 18145 31395 18185
rect 31405 18145 31445 18185
rect 31455 18145 31495 18185
rect 31505 18145 31545 18185
rect 31555 18145 31595 18185
rect 31605 18145 31645 18185
rect 31655 18145 31695 18185
rect 31705 18145 31745 18185
rect 31755 18145 31795 18185
rect 31805 18145 31845 18185
rect 31855 18145 31895 18185
rect 31905 18145 31945 18185
rect 31955 18145 31995 18185
rect 32005 18145 32045 18185
rect 32055 18145 32095 18185
rect 32105 18145 32145 18185
rect 32155 18145 32195 18185
rect 32205 18145 32245 18185
rect 32255 18145 32295 18185
rect 32305 18145 32345 18185
rect 32355 18145 32395 18185
rect 32405 18145 32445 18185
rect 32455 18145 32495 18185
rect 32505 18145 32545 18185
rect 32555 18145 32595 18185
rect 32605 18145 32645 18185
rect 32655 18145 32695 18185
rect 32705 18145 32745 18185
rect 32755 18145 32795 18185
rect 32805 18145 32845 18185
rect 32855 18145 32895 18185
rect 32905 18145 32945 18185
rect 32955 18145 32995 18185
rect 33005 18145 33045 18185
rect 33055 18145 33095 18185
rect 33105 18145 33145 18185
rect 33155 18145 33195 18185
rect 33205 18145 33245 18185
rect 33255 18145 33295 18185
rect 33305 18145 33345 18185
rect 33355 18145 33395 18185
rect 33405 18145 33445 18185
rect 33455 18145 33495 18185
rect 33505 18145 33545 18185
rect 33555 18145 33595 18185
rect 33605 18145 33645 18185
rect 33655 18145 33695 18185
rect 33705 18145 33745 18185
rect 33755 18145 33795 18185
rect 33805 18145 33845 18185
rect 33855 18145 33895 18185
rect 33905 18145 33945 18185
rect 33955 18145 33995 18185
rect 34005 18145 34045 18185
rect 34055 18145 34095 18185
rect 34105 18145 34145 18185
rect 34155 18145 34195 18185
rect 34205 18145 34245 18185
rect 34255 18145 34295 18185
rect 34305 18145 34345 18185
rect 34355 18145 34395 18185
rect 34405 18145 34445 18185
rect 34455 18145 34495 18185
rect 34505 18145 34545 18185
rect 34555 18145 34595 18185
rect 34605 18145 34645 18185
rect 34655 18145 34695 18185
rect 34705 18145 34745 18185
rect 34755 18145 34795 18185
rect 34805 18145 34845 18185
rect 34855 18145 34895 18185
rect 34905 18145 34945 18185
rect 34955 18145 34995 18185
rect 35005 18145 35045 18185
rect 35055 18145 35095 18185
rect 35105 18145 35145 18185
rect 35155 18145 35195 18185
rect 35205 18145 35245 18185
rect 35255 18145 35295 18185
rect 35305 18145 35345 18185
rect 35355 18145 35395 18185
rect 35405 18145 35445 18185
rect 35455 18145 35495 18185
rect 35505 18145 35545 18185
rect 35555 18145 35595 18185
rect 35605 18145 35645 18185
rect 35655 18145 35695 18185
rect 35705 18145 35745 18185
rect 35755 18145 35795 18185
rect 35805 18145 35845 18185
rect 35855 18145 35895 18185
rect 35905 18145 35945 18185
rect 35955 18145 35995 18185
rect 36005 18145 36045 18185
rect 36055 18145 36095 18185
rect 36105 18145 36145 18185
rect 36155 18145 36195 18185
rect 36205 18145 36245 18185
rect 36255 18145 36295 18185
rect 36305 18145 36345 18185
rect 36355 18145 36395 18185
rect 36405 18145 36445 18185
rect 36455 18145 36495 18185
rect 36505 18145 36545 18185
rect 36555 18145 36595 18185
rect 36605 18145 36645 18185
rect 36655 18145 36695 18185
rect 36705 18145 36745 18185
rect 36755 18145 36795 18185
rect 36805 18145 36845 18185
rect 36855 18145 36895 18185
rect 36905 18145 36945 18185
rect 36955 18145 36995 18185
rect 37005 18145 37045 18185
rect 37055 18145 37095 18185
rect 37105 18145 37145 18185
rect 37155 18145 37195 18185
rect 37205 18145 37245 18185
rect 37255 18145 37295 18185
rect 37305 18145 37345 18185
rect 37355 18145 37395 18185
rect 37405 18145 37445 18185
rect 37455 18145 37495 18185
rect 37505 18145 37545 18185
rect 37555 18145 37595 18185
rect 37605 18145 37645 18185
rect 37655 18145 37695 18185
rect 37705 18145 37745 18185
rect 37755 18145 37795 18185
rect 37805 18145 37845 18185
rect 37855 18145 37895 18185
rect 37905 18145 37945 18185
rect 37955 18145 37995 18185
rect 38005 18145 38045 18185
rect 38055 18145 38095 18185
rect 38105 18145 38145 18185
rect 38155 18145 38195 18185
rect 38205 18145 38245 18185
rect 38255 18145 38295 18185
rect 38305 18145 38345 18185
rect 38355 18145 38395 18185
rect 38405 18145 38445 18185
rect 38455 18145 38495 18185
rect 38505 18145 38545 18185
rect 38555 18145 38595 18185
rect 38605 18145 38645 18185
rect 38655 18145 38695 18185
rect 38705 18145 38745 18185
rect 38755 18145 38795 18185
rect 38805 18145 38845 18185
rect 38855 18145 38895 18185
rect 38905 18145 38945 18185
rect 38955 18145 38995 18185
rect 39005 18145 39045 18185
rect 39055 18145 39095 18185
rect 39105 18145 39145 18185
rect 39155 18145 39195 18185
rect 39205 18145 39245 18185
rect 39255 18145 39295 18185
rect 39305 18145 39345 18185
rect 39355 18145 39395 18185
rect 39405 18145 39445 18185
rect 39455 18145 39495 18185
rect 39505 18145 39545 18185
rect 39555 18145 39595 18185
rect 39605 18145 39645 18185
rect 39655 18145 39695 18185
rect 39705 18145 39745 18185
rect -2695 17075 -2655 17115
rect 105 17075 145 17115
rect 155 17075 195 17115
rect 205 17075 245 17115
rect 255 17075 295 17115
rect 305 17075 345 17115
rect 355 17075 395 17115
rect 405 17075 445 17115
rect 455 17075 495 17115
rect 505 17075 545 17115
rect 555 17075 595 17115
rect 605 17075 645 17115
rect 655 17075 695 17115
rect 705 17075 745 17115
rect 755 17075 795 17115
rect 805 17075 845 17115
rect 855 17075 895 17115
rect 905 17075 945 17115
rect 955 17075 995 17115
rect 1005 17075 1045 17115
rect 1055 17075 1095 17115
rect 1105 17075 1145 17115
rect 1155 17075 1195 17115
rect 1205 17075 1245 17115
rect 1255 17075 1295 17115
rect 1305 17075 1345 17115
rect 1355 17075 1395 17115
rect 1405 17075 1445 17115
rect 1455 17075 1495 17115
rect 1505 17075 1545 17115
rect 1555 17075 1595 17115
rect 1605 17075 1645 17115
rect 1655 17075 1695 17115
rect 1705 17075 1745 17115
rect 1755 17075 1795 17115
rect 1805 17075 1845 17115
rect 1855 17075 1895 17115
rect 1905 17075 1945 17115
rect 1955 17075 1995 17115
rect 2005 17075 2045 17115
rect 2055 17075 2095 17115
rect 2105 17075 2145 17115
rect 2155 17075 2195 17115
rect 2205 17075 2245 17115
rect 2255 17075 2295 17115
rect 2305 17075 2345 17115
rect 2355 17075 2395 17115
rect 2405 17075 2445 17115
rect 2455 17075 2495 17115
rect 2505 17075 2545 17115
rect 2555 17075 2595 17115
rect 2605 17075 2645 17115
rect 2655 17075 2695 17115
rect 2705 17075 2745 17115
rect 2755 17075 2795 17115
rect 2805 17075 2845 17115
rect 2855 17075 2895 17115
rect 2905 17075 2945 17115
rect 2955 17075 2995 17115
rect 3005 17075 3045 17115
rect 3055 17075 3095 17115
rect 3105 17075 3145 17115
rect 3155 17075 3195 17115
rect 3205 17075 3245 17115
rect 3255 17075 3295 17115
rect 3305 17075 3345 17115
rect 3355 17075 3395 17115
rect 3405 17075 3445 17115
rect 3455 17075 3495 17115
rect 3505 17075 3545 17115
rect 3555 17075 3595 17115
rect 3605 17075 3645 17115
rect 3655 17075 3695 17115
rect 3705 17075 3745 17115
rect 3755 17075 3795 17115
rect 3805 17075 3845 17115
rect 3855 17075 3895 17115
rect 3905 17075 3945 17115
rect 3955 17075 3995 17115
rect 4005 17075 4045 17115
rect 4055 17075 4095 17115
rect 4105 17075 4145 17115
rect 4155 17075 4195 17115
rect 4205 17075 4245 17115
rect 4255 17075 4295 17115
rect 4305 17075 4345 17115
rect 4355 17075 4395 17115
rect 4405 17075 4445 17115
rect 4455 17075 4495 17115
rect 4505 17075 4545 17115
rect 4555 17075 4595 17115
rect 4605 17075 4645 17115
rect 4655 17075 4695 17115
rect 4705 17075 4745 17115
rect 4755 17075 4795 17115
rect 4805 17075 4845 17115
rect 4855 17075 4895 17115
rect 4905 17075 4945 17115
rect 4955 17075 4995 17115
rect 5005 17075 5045 17115
rect 5055 17075 5095 17115
rect 5105 17075 5145 17115
rect 5155 17075 5195 17115
rect 5205 17075 5245 17115
rect 5255 17075 5295 17115
rect 5305 17075 5345 17115
rect 5355 17075 5395 17115
rect 5405 17075 5445 17115
rect 5455 17075 5495 17115
rect 5505 17075 5545 17115
rect 5555 17075 5595 17115
rect 5605 17075 5645 17115
rect 5655 17075 5695 17115
rect 5705 17075 5745 17115
rect 5755 17075 5795 17115
rect 5805 17075 5845 17115
rect 5855 17075 5895 17115
rect 5905 17075 5945 17115
rect 5955 17075 5995 17115
rect 6005 17075 6045 17115
rect 6055 17075 6095 17115
rect 6105 17075 6145 17115
rect 6155 17075 6195 17115
rect 6205 17075 6245 17115
rect 6255 17075 6295 17115
rect 6305 17075 6345 17115
rect 6355 17075 6395 17115
rect 6405 17075 6445 17115
rect 6455 17075 6495 17115
rect 6505 17075 6545 17115
rect 6555 17075 6595 17115
rect 6605 17075 6645 17115
rect 6655 17075 6695 17115
rect 6705 17075 6745 17115
rect 6755 17075 6795 17115
rect 6805 17075 6845 17115
rect 6855 17075 6895 17115
rect 6905 17075 6945 17115
rect 6955 17075 6995 17115
rect 7005 17075 7045 17115
rect 7055 17075 7095 17115
rect 7105 17075 7145 17115
rect 7155 17075 7195 17115
rect 7205 17075 7245 17115
rect 7255 17075 7295 17115
rect 7305 17075 7345 17115
rect 7355 17075 7395 17115
rect 7405 17075 7445 17115
rect 7455 17075 7495 17115
rect 7505 17075 7545 17115
rect 7555 17075 7595 17115
rect 7605 17075 7645 17115
rect 7655 17075 7695 17115
rect 7705 17075 7745 17115
rect 7755 17075 7795 17115
rect 7805 17075 7845 17115
rect 7855 17075 7895 17115
rect 7905 17075 7945 17115
rect 7955 17075 7995 17115
rect 8005 17075 8045 17115
rect 8055 17075 8095 17115
rect 8105 17075 8145 17115
rect 8155 17075 8195 17115
rect 8205 17075 8245 17115
rect 8255 17075 8295 17115
rect 8305 17075 8345 17115
rect 8355 17075 8395 17115
rect 8405 17075 8445 17115
rect 8455 17075 8495 17115
rect 8505 17075 8545 17115
rect 8555 17075 8595 17115
rect 8605 17075 8645 17115
rect 8655 17075 8695 17115
rect 8705 17075 8745 17115
rect 8755 17075 8795 17115
rect 8805 17075 8845 17115
rect 8855 17075 8895 17115
rect 8905 17075 8945 17115
rect 8955 17075 8995 17115
rect 9005 17075 9045 17115
rect 9055 17075 9095 17115
rect 9105 17075 9145 17115
rect 9155 17075 9195 17115
rect 9205 17075 9245 17115
rect 9255 17075 9295 17115
rect 9305 17075 9345 17115
rect 9355 17075 9395 17115
rect 9405 17075 9445 17115
rect 9455 17075 9495 17115
rect 9505 17075 9545 17115
rect 9555 17075 9595 17115
rect 9605 17075 9645 17115
rect 9655 17075 9695 17115
rect 9705 17075 9745 17115
rect 9755 17075 9795 17115
rect 9805 17075 9845 17115
rect 9855 17075 9895 17115
rect 9905 17075 9945 17115
rect 9955 17075 9995 17115
rect 10005 17075 10045 17115
rect 10055 17075 10095 17115
rect 10105 17075 10145 17115
rect 10155 17075 10195 17115
rect 10205 17075 10245 17115
rect 10255 17075 10295 17115
rect 10305 17075 10345 17115
rect 10355 17075 10395 17115
rect 10405 17075 10445 17115
rect 10455 17075 10495 17115
rect 10505 17075 10545 17115
rect 10555 17075 10595 17115
rect 10605 17075 10645 17115
rect 10655 17075 10695 17115
rect 10705 17075 10745 17115
rect 10755 17075 10795 17115
rect 10805 17075 10845 17115
rect 10855 17075 10895 17115
rect 10905 17075 10945 17115
rect 10955 17075 10995 17115
rect 11005 17075 11045 17115
rect 11055 17075 11095 17115
rect 11105 17075 11145 17115
rect 11155 17075 11195 17115
rect 11205 17075 11245 17115
rect 11255 17075 11295 17115
rect 11305 17075 11345 17115
rect 11355 17075 11395 17115
rect 11405 17075 11445 17115
rect 11455 17075 11495 17115
rect 11505 17075 11545 17115
rect 11555 17075 11595 17115
rect 11605 17075 11645 17115
rect 11655 17075 11695 17115
rect 11705 17075 11745 17115
rect 11755 17075 11795 17115
rect 11805 17075 11845 17115
rect 11855 17075 11895 17115
rect 11905 17075 11945 17115
rect 11955 17075 11995 17115
rect 12005 17075 12045 17115
rect 12055 17075 12095 17115
rect 12105 17075 12145 17115
rect 12155 17075 12195 17115
rect 12205 17075 12245 17115
rect 12255 17075 12295 17115
rect 12305 17075 12345 17115
rect 12355 17075 12395 17115
rect 12405 17075 12445 17115
rect 12455 17075 12495 17115
rect 12505 17075 12545 17115
rect 12555 17075 12595 17115
rect 12605 17075 12645 17115
rect 12655 17075 12695 17115
rect 12705 17075 12745 17115
rect 12755 17075 12795 17115
rect 12805 17075 12845 17115
rect 12855 17075 12895 17115
rect 12905 17075 12945 17115
rect 12955 17075 12995 17115
rect 13005 17075 13045 17115
rect 13055 17075 13095 17115
rect 13105 17075 13145 17115
rect 13155 17075 13195 17115
rect 13205 17075 13245 17115
rect 13255 17075 13295 17115
rect 13305 17075 13345 17115
rect 13355 17075 13395 17115
rect 13405 17075 13445 17115
rect 13455 17075 13495 17115
rect 13505 17075 13545 17115
rect 13555 17075 13595 17115
rect 13605 17075 13645 17115
rect 13655 17075 13695 17115
rect 13705 17075 13745 17115
rect 13755 17075 13795 17115
rect 13805 17075 13845 17115
rect 13855 17075 13895 17115
rect 13905 17075 13945 17115
rect 13955 17075 13995 17115
rect 14005 17075 14045 17115
rect 14055 17075 14095 17115
rect 14105 17075 14145 17115
rect 14155 17075 14195 17115
rect 14205 17075 14245 17115
rect 14255 17075 14295 17115
rect 14305 17075 14345 17115
rect 14355 17075 14395 17115
rect 14405 17075 14445 17115
rect 14455 17075 14495 17115
rect 14505 17075 14545 17115
rect 14555 17075 14595 17115
rect 14605 17075 14645 17115
rect 14655 17075 14695 17115
rect 14705 17075 14745 17115
rect 14755 17075 14795 17115
rect 14805 17075 14845 17115
rect 14855 17075 14895 17115
rect 14905 17075 14945 17115
rect 14955 17075 14995 17115
rect 15005 17075 15045 17115
rect 15055 17075 15095 17115
rect 15105 17075 15145 17115
rect 15155 17075 15195 17115
rect 15205 17075 15245 17115
rect 15255 17075 15295 17115
rect 15305 17075 15345 17115
rect 15355 17075 15395 17115
rect 15405 17075 15445 17115
rect 15455 17075 15495 17115
rect 15505 17075 15545 17115
rect 15555 17075 15595 17115
rect 15605 17075 15645 17115
rect 15655 17075 15695 17115
rect 15705 17075 15745 17115
rect 15755 17075 15795 17115
rect 15805 17075 15845 17115
rect 15855 17075 15895 17115
rect 15905 17075 15945 17115
rect 15955 17075 15995 17115
rect 16005 17075 16045 17115
rect 16055 17075 16095 17115
rect 16105 17075 16145 17115
rect 16155 17075 16195 17115
rect 16205 17075 16245 17115
rect 16255 17075 16295 17115
rect 16305 17075 16345 17115
rect 16355 17075 16395 17115
rect 16405 17075 16445 17115
rect 16455 17075 16495 17115
rect 16505 17075 16545 17115
rect 16555 17075 16595 17115
rect 16605 17075 16645 17115
rect 16655 17075 16695 17115
rect 16705 17075 16745 17115
rect 16755 17075 16795 17115
rect 16805 17075 16845 17115
rect 16855 17075 16895 17115
rect 16905 17075 16945 17115
rect 16955 17075 16995 17115
rect 17005 17075 17045 17115
rect 17055 17075 17095 17115
rect 17105 17075 17145 17115
rect 17155 17075 17195 17115
rect 17205 17075 17245 17115
rect 17255 17075 17295 17115
rect 17305 17075 17345 17115
rect 17355 17075 17395 17115
rect 17405 17075 17445 17115
rect 17455 17075 17495 17115
rect 17505 17075 17545 17115
rect 17555 17075 17595 17115
rect 17605 17075 17645 17115
rect 17655 17075 17695 17115
rect 17705 17075 17745 17115
rect 17755 17075 17795 17115
rect 17805 17075 17845 17115
rect 17855 17075 17895 17115
rect 17905 17075 17945 17115
rect 17955 17075 17995 17115
rect 18005 17075 18045 17115
rect 18055 17075 18095 17115
rect 18105 17075 18145 17115
rect 18155 17075 18195 17115
rect 18205 17075 18245 17115
rect 18255 17075 18295 17115
rect 18305 17075 18345 17115
rect 18355 17075 18395 17115
rect 18405 17075 18445 17115
rect 18455 17075 18495 17115
rect 18505 17075 18545 17115
rect 18555 17075 18595 17115
rect 18605 17075 18645 17115
rect 18655 17075 18695 17115
rect 18705 17075 18745 17115
rect 18755 17075 18795 17115
rect 18805 17075 18845 17115
rect 18855 17075 18895 17115
rect 18905 17075 18945 17115
rect 18955 17075 18995 17115
rect 19005 17075 19045 17115
rect 19055 17075 19095 17115
rect 19105 17075 19145 17115
rect 19155 17075 19195 17115
rect 19205 17075 19245 17115
rect 19255 17075 19295 17115
rect 19305 17075 19345 17115
rect 19355 17075 19395 17115
rect 19405 17075 19445 17115
rect 19455 17075 19495 17115
rect 19505 17075 19545 17115
rect 19555 17075 19595 17115
rect 19605 17075 19645 17115
rect 19655 17075 19695 17115
rect 19705 17075 19745 17115
rect 19755 17075 19795 17115
rect 19805 17075 19845 17115
rect 19855 17075 19895 17115
rect 19905 17075 19945 17115
rect 19955 17075 19995 17115
rect 20005 17075 20045 17115
rect 20055 17075 20095 17115
rect 20105 17075 20145 17115
rect 20155 17075 20195 17115
rect 20205 17075 20245 17115
rect 20255 17075 20295 17115
rect 20305 17075 20345 17115
rect 20355 17075 20395 17115
rect 20405 17075 20445 17115
rect 20455 17075 20495 17115
rect 20505 17075 20545 17115
rect 20555 17075 20595 17115
rect 20605 17075 20645 17115
rect 20655 17075 20695 17115
rect 20705 17075 20745 17115
rect 20755 17075 20795 17115
rect 20805 17075 20845 17115
rect 20855 17075 20895 17115
rect 20905 17075 20945 17115
rect 20955 17075 20995 17115
rect 21005 17075 21045 17115
rect 21055 17075 21095 17115
rect 21105 17075 21145 17115
rect 21155 17075 21195 17115
rect 21205 17075 21245 17115
rect 21255 17075 21295 17115
rect 21305 17075 21345 17115
rect 21355 17075 21395 17115
rect 21405 17075 21445 17115
rect 21455 17075 21495 17115
rect 21505 17075 21545 17115
rect 21555 17075 21595 17115
rect 21605 17075 21645 17115
rect 21655 17075 21695 17115
rect 21705 17075 21745 17115
rect 21755 17075 21795 17115
rect 21805 17075 21845 17115
rect 21855 17075 21895 17115
rect 21905 17075 21945 17115
rect 21955 17075 21995 17115
rect 22005 17075 22045 17115
rect 22055 17075 22095 17115
rect 22105 17075 22145 17115
rect 22155 17075 22195 17115
rect 22205 17075 22245 17115
rect 22255 17075 22295 17115
rect 22305 17075 22345 17115
rect 22355 17075 22395 17115
rect 22405 17075 22445 17115
rect 22455 17075 22495 17115
rect 22505 17075 22545 17115
rect 22555 17075 22595 17115
rect 22605 17075 22645 17115
rect 22655 17075 22695 17115
rect 22705 17075 22745 17115
rect 22755 17075 22795 17115
rect 22805 17075 22845 17115
rect 22855 17075 22895 17115
rect 22905 17075 22945 17115
rect 22955 17075 22995 17115
rect 23005 17075 23045 17115
rect 23055 17075 23095 17115
rect 23105 17075 23145 17115
rect 23155 17075 23195 17115
rect 23205 17075 23245 17115
rect 23255 17075 23295 17115
rect 23305 17075 23345 17115
rect 23355 17075 23395 17115
rect 23405 17075 23445 17115
rect 23455 17075 23495 17115
rect 23505 17075 23545 17115
rect 23555 17075 23595 17115
rect 23605 17075 23645 17115
rect 23655 17075 23695 17115
rect 23705 17075 23745 17115
rect 23755 17075 23795 17115
rect 23805 17075 23845 17115
rect 23855 17075 23895 17115
rect 23905 17075 23945 17115
rect 23955 17075 23995 17115
rect 24005 17075 24045 17115
rect 24055 17075 24095 17115
rect 24105 17075 24145 17115
rect 24155 17075 24195 17115
rect 24205 17075 24245 17115
rect 24255 17075 24295 17115
rect 24305 17075 24345 17115
rect 24355 17075 24395 17115
rect 24405 17075 24445 17115
rect 24455 17075 24495 17115
rect 24505 17075 24545 17115
rect 24555 17075 24595 17115
rect 24605 17075 24645 17115
rect 24655 17075 24695 17115
rect 24705 17075 24745 17115
rect 24755 17075 24795 17115
rect 24805 17075 24845 17115
rect 24855 17075 24895 17115
rect 24905 17075 24945 17115
rect 24955 17075 24995 17115
rect 25005 17075 25045 17115
rect 25055 17075 25095 17115
rect 25105 17075 25145 17115
rect 25155 17075 25195 17115
rect 25205 17075 25245 17115
rect 25255 17075 25295 17115
rect 25305 17075 25345 17115
rect 25355 17075 25395 17115
rect 25405 17075 25445 17115
rect 25455 17075 25495 17115
rect 25505 17075 25545 17115
rect 25555 17075 25595 17115
rect 25605 17075 25645 17115
rect 25655 17075 25695 17115
rect 25705 17075 25745 17115
rect 25755 17075 25795 17115
rect 25805 17075 25845 17115
rect 25855 17075 25895 17115
rect 25905 17075 25945 17115
rect 25955 17075 25995 17115
rect 26005 17075 26045 17115
rect 26055 17075 26095 17115
rect 26105 17075 26145 17115
rect 26155 17075 26195 17115
rect 26205 17075 26245 17115
rect 26255 17075 26295 17115
rect 26305 17075 26345 17115
rect 26355 17075 26395 17115
rect 26405 17075 26445 17115
rect 26455 17075 26495 17115
rect 26505 17075 26545 17115
rect 26555 17075 26595 17115
rect 26605 17075 26645 17115
rect 26655 17075 26695 17115
rect 26705 17075 26745 17115
rect 26755 17075 26795 17115
rect 26805 17075 26845 17115
rect 26855 17075 26895 17115
rect 26905 17075 26945 17115
rect 26955 17075 26995 17115
rect 27005 17075 27045 17115
rect 27055 17075 27095 17115
rect 27105 17075 27145 17115
rect 27155 17075 27195 17115
rect 27205 17075 27245 17115
rect 27255 17075 27295 17115
rect 27305 17075 27345 17115
rect 27355 17075 27395 17115
rect 27405 17075 27445 17115
rect 27455 17075 27495 17115
rect 27505 17075 27545 17115
rect 27555 17075 27595 17115
rect 27605 17075 27645 17115
rect 27655 17075 27695 17115
rect 27705 17075 27745 17115
rect 27755 17075 27795 17115
rect 27805 17075 27845 17115
rect 27855 17075 27895 17115
rect 27905 17075 27945 17115
rect 27955 17075 27995 17115
rect 28005 17075 28045 17115
rect 28055 17075 28095 17115
rect 28105 17075 28145 17115
rect 28155 17075 28195 17115
rect 28205 17075 28245 17115
rect 28255 17075 28295 17115
rect 28305 17075 28345 17115
rect 28355 17075 28395 17115
rect 28405 17075 28445 17115
rect 28455 17075 28495 17115
rect 28505 17075 28545 17115
rect 28555 17075 28595 17115
rect 28605 17075 28645 17115
rect 28655 17075 28695 17115
rect 28705 17075 28745 17115
rect 28755 17075 28795 17115
rect 28805 17075 28845 17115
rect 28855 17075 28895 17115
rect 28905 17075 28945 17115
rect 28955 17075 28995 17115
rect 29005 17075 29045 17115
rect 29055 17075 29095 17115
rect 29105 17075 29145 17115
rect 29155 17075 29195 17115
rect 29205 17075 29245 17115
rect 29255 17075 29295 17115
rect 29305 17075 29345 17115
rect 29355 17075 29395 17115
rect 29405 17075 29445 17115
rect 29455 17075 29495 17115
rect 29505 17075 29545 17115
rect 29555 17075 29595 17115
rect 29605 17075 29645 17115
rect 29655 17075 29695 17115
rect 29705 17075 29745 17115
rect 29755 17075 29795 17115
rect 29805 17075 29845 17115
rect 29855 17075 29895 17115
rect 29905 17075 29945 17115
rect 29955 17075 29995 17115
rect 30005 17075 30045 17115
rect 30055 17075 30095 17115
rect 30105 17075 30145 17115
rect 30155 17075 30195 17115
rect 30205 17075 30245 17115
rect 30255 17075 30295 17115
rect 30305 17075 30345 17115
rect 30355 17075 30395 17115
rect 30405 17075 30445 17115
rect 30455 17075 30495 17115
rect 30505 17075 30545 17115
rect 30555 17075 30595 17115
rect 30605 17075 30645 17115
rect 30655 17075 30695 17115
rect 30705 17075 30745 17115
rect 30755 17075 30795 17115
rect 30805 17075 30845 17115
rect 30855 17075 30895 17115
rect 30905 17075 30945 17115
rect 30955 17075 30995 17115
rect 31005 17075 31045 17115
rect 31055 17075 31095 17115
rect 31105 17075 31145 17115
rect 31155 17075 31195 17115
rect 31205 17075 31245 17115
rect 31255 17075 31295 17115
rect 31305 17075 31345 17115
rect 31355 17075 31395 17115
rect 31405 17075 31445 17115
rect 31455 17075 31495 17115
rect 31505 17075 31545 17115
rect 31555 17075 31595 17115
rect 31605 17075 31645 17115
rect 31655 17075 31695 17115
rect 31705 17075 31745 17115
rect 31755 17075 31795 17115
rect 31805 17075 31845 17115
rect 31855 17075 31895 17115
rect 31905 17075 31945 17115
rect 31955 17075 31995 17115
rect 32005 17075 32045 17115
rect 32055 17075 32095 17115
rect 32105 17075 32145 17115
rect 32155 17075 32195 17115
rect 32205 17075 32245 17115
rect 32255 17075 32295 17115
rect 32305 17075 32345 17115
rect 32355 17075 32395 17115
rect 32405 17075 32445 17115
rect 32455 17075 32495 17115
rect 32505 17075 32545 17115
rect 32555 17075 32595 17115
rect 32605 17075 32645 17115
rect 32655 17075 32695 17115
rect 32705 17075 32745 17115
rect 32755 17075 32795 17115
rect 32805 17075 32845 17115
rect 32855 17075 32895 17115
rect 32905 17075 32945 17115
rect 32955 17075 32995 17115
rect 33005 17075 33045 17115
rect 33055 17075 33095 17115
rect 33105 17075 33145 17115
rect 33155 17075 33195 17115
rect 33205 17075 33245 17115
rect 33255 17075 33295 17115
rect 33305 17075 33345 17115
rect 33355 17075 33395 17115
rect 33405 17075 33445 17115
rect 33455 17075 33495 17115
rect 33505 17075 33545 17115
rect 33555 17075 33595 17115
rect 33605 17075 33645 17115
rect 33655 17075 33695 17115
rect 33705 17075 33745 17115
rect 33755 17075 33795 17115
rect 33805 17075 33845 17115
rect 33855 17075 33895 17115
rect 33905 17075 33945 17115
rect 33955 17075 33995 17115
rect 34005 17075 34045 17115
rect 34055 17075 34095 17115
rect 34105 17075 34145 17115
rect 34155 17075 34195 17115
rect 34205 17075 34245 17115
rect 34255 17075 34295 17115
rect 34305 17075 34345 17115
rect 34355 17075 34395 17115
rect 34405 17075 34445 17115
rect 34455 17075 34495 17115
rect 34505 17075 34545 17115
rect 34555 17075 34595 17115
rect 34605 17075 34645 17115
rect 34655 17075 34695 17115
rect 34705 17075 34745 17115
rect 34755 17075 34795 17115
rect 34805 17075 34845 17115
rect 34855 17075 34895 17115
rect 34905 17075 34945 17115
rect 34955 17075 34995 17115
rect 35005 17075 35045 17115
rect 35055 17075 35095 17115
rect 35105 17075 35145 17115
rect 35155 17075 35195 17115
rect 35205 17075 35245 17115
rect 35255 17075 35295 17115
rect 35305 17075 35345 17115
rect 35355 17075 35395 17115
rect 35405 17075 35445 17115
rect 35455 17075 35495 17115
rect 35505 17075 35545 17115
rect 35555 17075 35595 17115
rect 35605 17075 35645 17115
rect 35655 17075 35695 17115
rect 35705 17075 35745 17115
rect 35755 17075 35795 17115
rect 35805 17075 35845 17115
rect 35855 17075 35895 17115
rect 35905 17075 35945 17115
rect 35955 17075 35995 17115
rect 36005 17075 36045 17115
rect 36055 17075 36095 17115
rect 36105 17075 36145 17115
rect 36155 17075 36195 17115
rect 36205 17075 36245 17115
rect 36255 17075 36295 17115
rect 36305 17075 36345 17115
rect 36355 17075 36395 17115
rect 36405 17075 36445 17115
rect 36455 17075 36495 17115
rect 36505 17075 36545 17115
rect 36555 17075 36595 17115
rect 36605 17075 36645 17115
rect 36655 17075 36695 17115
rect 36705 17075 36745 17115
rect 36755 17075 36795 17115
rect 36805 17075 36845 17115
rect 36855 17075 36895 17115
rect 36905 17075 36945 17115
rect 36955 17075 36995 17115
rect 37005 17075 37045 17115
rect 37055 17075 37095 17115
rect 37105 17075 37145 17115
rect 37155 17075 37195 17115
rect 37205 17075 37245 17115
rect 37255 17075 37295 17115
rect 37305 17075 37345 17115
rect 37355 17075 37395 17115
rect 37405 17075 37445 17115
rect 37455 17075 37495 17115
rect 37505 17075 37545 17115
rect 37555 17075 37595 17115
rect 37605 17075 37645 17115
rect 37655 17075 37695 17115
rect 37705 17075 37745 17115
rect 37755 17075 37795 17115
rect 37805 17075 37845 17115
rect 37855 17075 37895 17115
rect 37905 17075 37945 17115
rect 37955 17075 37995 17115
rect 38005 17075 38045 17115
rect 38055 17075 38095 17115
rect 38105 17075 38145 17115
rect 38155 17075 38195 17115
rect 38205 17075 38245 17115
rect 38255 17075 38295 17115
rect 38305 17075 38345 17115
rect 38355 17075 38395 17115
rect 38405 17075 38445 17115
rect 38455 17075 38495 17115
rect 38505 17075 38545 17115
rect 38555 17075 38595 17115
rect 38605 17075 38645 17115
rect 38655 17075 38695 17115
rect 38705 17075 38745 17115
rect 38755 17075 38795 17115
rect 38805 17075 38845 17115
rect 38855 17075 38895 17115
rect 38905 17075 38945 17115
rect 38955 17075 38995 17115
rect 39005 17075 39045 17115
rect 39055 17075 39095 17115
rect 39105 17075 39145 17115
rect 39155 17075 39195 17115
rect 39205 17075 39245 17115
rect 39255 17075 39295 17115
rect 39305 17075 39345 17115
rect 39355 17075 39395 17115
rect 39405 17075 39445 17115
rect 39455 17075 39495 17115
rect 39505 17075 39545 17115
rect 39555 17075 39595 17115
rect 39605 17075 39645 17115
rect 39655 17075 39695 17115
rect 39705 17075 39745 17115
rect -3495 17010 -3455 17015
rect -3495 16980 -3490 17010
rect -3490 16980 -3460 17010
rect -3460 16980 -3455 17010
rect -3495 16975 -3455 16980
rect -3295 17010 -3255 17015
rect -3295 16980 -3290 17010
rect -3290 16980 -3260 17010
rect -3260 16980 -3255 17010
rect -3295 16975 -3255 16980
rect -3095 17010 -3055 17015
rect -3095 16980 -3090 17010
rect -3090 16980 -3060 17010
rect -3060 16980 -3055 17010
rect -3095 16975 -3055 16980
rect -1595 17010 -1555 17015
rect -1595 16980 -1590 17010
rect -1590 16980 -1560 17010
rect -1560 16980 -1555 17010
rect -1595 16975 -1555 16980
rect -1195 17010 -1155 17015
rect -1195 16980 -1190 17010
rect -1190 16980 -1160 17010
rect -1160 16980 -1155 17010
rect -1195 16975 -1155 16980
rect -1095 17010 -1055 17015
rect -1095 16980 -1090 17010
rect -1090 16980 -1060 17010
rect -1060 16980 -1055 17010
rect -1095 16975 -1055 16980
rect -995 17010 -955 17015
rect -995 16980 -990 17010
rect -990 16980 -960 17010
rect -960 16980 -955 17010
rect -995 16975 -955 16980
rect -895 17010 -855 17015
rect -895 16980 -890 17010
rect -890 16980 -860 17010
rect -860 16980 -855 17010
rect -895 16975 -855 16980
rect -795 17010 -755 17015
rect -795 16980 -790 17010
rect -790 16980 -760 17010
rect -760 16980 -755 17010
rect -795 16975 -755 16980
rect -695 17010 -655 17015
rect -695 16980 -690 17010
rect -690 16980 -660 17010
rect -660 16980 -655 17010
rect -695 16975 -655 16980
rect -595 17010 -555 17015
rect -595 16980 -590 17010
rect -590 16980 -560 17010
rect -560 16980 -555 17010
rect -595 16975 -555 16980
rect -495 17010 -455 17015
rect -495 16980 -490 17010
rect -490 16980 -460 17010
rect -460 16980 -455 17010
rect -495 16975 -455 16980
rect -395 17010 -355 17015
rect -395 16980 -390 17010
rect -390 16980 -360 17010
rect -360 16980 -355 17010
rect -395 16975 -355 16980
rect -295 17010 -255 17015
rect -295 16980 -290 17010
rect -290 16980 -260 17010
rect -260 16980 -255 17010
rect -295 16975 -255 16980
rect -195 17010 -155 17015
rect -195 16980 -190 17010
rect -190 16980 -160 17010
rect -160 16980 -155 17010
rect -195 16975 -155 16980
rect -95 17010 -55 17015
rect -95 16980 -90 17010
rect -90 16980 -60 17010
rect -60 16980 -55 17010
rect -95 16975 -55 16980
rect 5 16975 45 17015
rect 55 16975 95 17015
rect 105 16975 145 17015
rect 155 16975 195 17015
rect 205 16975 245 17015
rect 255 16975 295 17015
rect 305 16975 345 17015
rect 355 16975 395 17015
rect 405 16975 445 17015
rect 455 16975 495 17015
rect 505 16975 545 17015
rect 555 16975 595 17015
rect 605 16975 645 17015
rect 655 16975 695 17015
rect 705 16975 745 17015
rect 755 16975 795 17015
rect 805 16975 845 17015
rect 855 16975 895 17015
rect 905 16975 945 17015
rect 955 16975 995 17015
rect 1005 16975 1045 17015
rect 1055 16975 1095 17015
rect 1105 16975 1145 17015
rect 1155 16975 1195 17015
rect 1205 16975 1245 17015
rect 1255 16975 1295 17015
rect 1305 16975 1345 17015
rect 1355 16975 1395 17015
rect 1405 16975 1445 17015
rect 1455 16975 1495 17015
rect 1505 16975 1545 17015
rect 1555 16975 1595 17015
rect 1605 16975 1645 17015
rect 1655 16975 1695 17015
rect 1705 16975 1745 17015
rect 1755 16975 1795 17015
rect 1805 16975 1845 17015
rect 1855 16975 1895 17015
rect 1905 16975 1945 17015
rect 1955 16975 1995 17015
rect 2005 16975 2045 17015
rect 2055 16975 2095 17015
rect 2105 16975 2145 17015
rect 2155 16975 2195 17015
rect 2205 16975 2245 17015
rect 2255 16975 2295 17015
rect 2305 16975 2345 17015
rect 2355 16975 2395 17015
rect 2405 16975 2445 17015
rect 2455 16975 2495 17015
rect 2505 16975 2545 17015
rect 2555 16975 2595 17015
rect 2605 16975 2645 17015
rect 2655 16975 2695 17015
rect 2705 16975 2745 17015
rect 2755 16975 2795 17015
rect 2805 16975 2845 17015
rect 2855 16975 2895 17015
rect 2905 16975 2945 17015
rect 2955 16975 2995 17015
rect 3005 16975 3045 17015
rect 3055 16975 3095 17015
rect 3105 16975 3145 17015
rect 3155 16975 3195 17015
rect 3205 16975 3245 17015
rect 3255 16975 3295 17015
rect 3305 16975 3345 17015
rect 3355 16975 3395 17015
rect 3405 16975 3445 17015
rect 3455 16975 3495 17015
rect 3505 16975 3545 17015
rect 3555 16975 3595 17015
rect 3605 16975 3645 17015
rect 3655 16975 3695 17015
rect 3705 16975 3745 17015
rect 3755 16975 3795 17015
rect 3805 16975 3845 17015
rect 3855 16975 3895 17015
rect 3905 16975 3945 17015
rect 3955 16975 3995 17015
rect 4005 16975 4045 17015
rect 4055 16975 4095 17015
rect 4105 16975 4145 17015
rect 4155 16975 4195 17015
rect 4205 16975 4245 17015
rect 4255 16975 4295 17015
rect 4305 16975 4345 17015
rect 4355 16975 4395 17015
rect 4405 16975 4445 17015
rect 4455 16975 4495 17015
rect 4505 16975 4545 17015
rect 4555 16975 4595 17015
rect 4605 16975 4645 17015
rect 4655 16975 4695 17015
rect 4705 16975 4745 17015
rect 4755 16975 4795 17015
rect 4805 16975 4845 17015
rect 4855 16975 4895 17015
rect 4905 16975 4945 17015
rect 4955 16975 4995 17015
rect 5005 16975 5045 17015
rect 5055 16975 5095 17015
rect 5105 16975 5145 17015
rect 5155 16975 5195 17015
rect 5205 16975 5245 17015
rect 5255 16975 5295 17015
rect 5305 16975 5345 17015
rect 5355 16975 5395 17015
rect 5405 16975 5445 17015
rect 5455 16975 5495 17015
rect 5505 16975 5545 17015
rect 5555 16975 5595 17015
rect 5605 16975 5645 17015
rect 5655 16975 5695 17015
rect 5705 16975 5745 17015
rect 5755 16975 5795 17015
rect 5805 16975 5845 17015
rect 5855 16975 5895 17015
rect 5905 16975 5945 17015
rect 5955 16975 5995 17015
rect 6005 16975 6045 17015
rect 6055 16975 6095 17015
rect 6105 16975 6145 17015
rect 6155 16975 6195 17015
rect 6205 16975 6245 17015
rect 6255 16975 6295 17015
rect 6305 16975 6345 17015
rect 6355 16975 6395 17015
rect 6405 16975 6445 17015
rect 6455 16975 6495 17015
rect 6505 16975 6545 17015
rect 6555 16975 6595 17015
rect 6605 16975 6645 17015
rect 6655 16975 6695 17015
rect 6705 16975 6745 17015
rect 6755 16975 6795 17015
rect 6805 16975 6845 17015
rect 6855 16975 6895 17015
rect 6905 16975 6945 17015
rect 6955 16975 6995 17015
rect 7005 16975 7045 17015
rect 7055 16975 7095 17015
rect 7105 16975 7145 17015
rect 7155 16975 7195 17015
rect 7205 16975 7245 17015
rect 7255 16975 7295 17015
rect 7305 16975 7345 17015
rect 7355 16975 7395 17015
rect 7405 16975 7445 17015
rect 7455 16975 7495 17015
rect 7505 16975 7545 17015
rect 7555 16975 7595 17015
rect 7605 16975 7645 17015
rect 7655 16975 7695 17015
rect 7705 16975 7745 17015
rect 7755 16975 7795 17015
rect 7805 16975 7845 17015
rect 7855 16975 7895 17015
rect 7905 16975 7945 17015
rect 7955 16975 7995 17015
rect 8005 16975 8045 17015
rect 8055 16975 8095 17015
rect 8105 16975 8145 17015
rect 8155 16975 8195 17015
rect 8205 16975 8245 17015
rect 8255 16975 8295 17015
rect 8305 16975 8345 17015
rect 8355 16975 8395 17015
rect 8405 16975 8445 17015
rect 8455 16975 8495 17015
rect 8505 16975 8545 17015
rect 8555 16975 8595 17015
rect 8605 16975 8645 17015
rect 8655 16975 8695 17015
rect 8705 16975 8745 17015
rect 8755 16975 8795 17015
rect 8805 16975 8845 17015
rect 8855 16975 8895 17015
rect 8905 16975 8945 17015
rect 8955 16975 8995 17015
rect 9005 16975 9045 17015
rect 9055 16975 9095 17015
rect 9105 16975 9145 17015
rect 9155 16975 9195 17015
rect 9205 16975 9245 17015
rect 9255 16975 9295 17015
rect 9305 16975 9345 17015
rect 9355 16975 9395 17015
rect 9405 16975 9445 17015
rect 9455 16975 9495 17015
rect 9505 16975 9545 17015
rect 9555 16975 9595 17015
rect 9605 16975 9645 17015
rect 9655 16975 9695 17015
rect 9705 16975 9745 17015
rect 9755 16975 9795 17015
rect 9805 16975 9845 17015
rect 9855 16975 9895 17015
rect 9905 16975 9945 17015
rect 9955 16975 9995 17015
rect 10005 16975 10045 17015
rect 10055 16975 10095 17015
rect 10105 16975 10145 17015
rect 10155 16975 10195 17015
rect 10205 16975 10245 17015
rect 10255 16975 10295 17015
rect 10305 16975 10345 17015
rect 10355 16975 10395 17015
rect 10405 16975 10445 17015
rect 10455 16975 10495 17015
rect 10505 16975 10545 17015
rect 10555 16975 10595 17015
rect 10605 16975 10645 17015
rect 10655 16975 10695 17015
rect 10705 16975 10745 17015
rect 10755 16975 10795 17015
rect 10805 16975 10845 17015
rect 10855 16975 10895 17015
rect 10905 16975 10945 17015
rect 10955 16975 10995 17015
rect 11005 16975 11045 17015
rect 11055 16975 11095 17015
rect 11105 16975 11145 17015
rect 11155 16975 11195 17015
rect 11205 16975 11245 17015
rect 11255 16975 11295 17015
rect 11305 16975 11345 17015
rect 11355 16975 11395 17015
rect 11405 16975 11445 17015
rect 11455 16975 11495 17015
rect 11505 16975 11545 17015
rect 11555 16975 11595 17015
rect 11605 16975 11645 17015
rect 11655 16975 11695 17015
rect 11705 16975 11745 17015
rect 11755 16975 11795 17015
rect 11805 16975 11845 17015
rect 11855 16975 11895 17015
rect 11905 16975 11945 17015
rect 11955 16975 11995 17015
rect 12005 16975 12045 17015
rect 12055 16975 12095 17015
rect 12105 16975 12145 17015
rect 12155 16975 12195 17015
rect 12205 16975 12245 17015
rect 12255 16975 12295 17015
rect 12305 16975 12345 17015
rect 12355 16975 12395 17015
rect 12405 16975 12445 17015
rect 12455 16975 12495 17015
rect 12505 16975 12545 17015
rect 12555 16975 12595 17015
rect 12605 16975 12645 17015
rect 12655 16975 12695 17015
rect 12705 16975 12745 17015
rect 12755 16975 12795 17015
rect 12805 16975 12845 17015
rect 12855 16975 12895 17015
rect 12905 16975 12945 17015
rect 12955 16975 12995 17015
rect 13005 16975 13045 17015
rect 13055 16975 13095 17015
rect 13105 16975 13145 17015
rect 13155 16975 13195 17015
rect 13205 16975 13245 17015
rect 13255 16975 13295 17015
rect 13305 16975 13345 17015
rect 13355 16975 13395 17015
rect 13405 16975 13445 17015
rect 13455 16975 13495 17015
rect 13505 16975 13545 17015
rect 13555 16975 13595 17015
rect 13605 16975 13645 17015
rect 13655 16975 13695 17015
rect 13705 16975 13745 17015
rect 13755 16975 13795 17015
rect 13805 16975 13845 17015
rect 13855 16975 13895 17015
rect 13905 16975 13945 17015
rect 13955 16975 13995 17015
rect 14005 16975 14045 17015
rect 14055 16975 14095 17015
rect 14105 16975 14145 17015
rect 14155 16975 14195 17015
rect 14205 16975 14245 17015
rect 14255 16975 14295 17015
rect 14305 16975 14345 17015
rect 14355 16975 14395 17015
rect 14405 16975 14445 17015
rect 14455 16975 14495 17015
rect 14505 16975 14545 17015
rect 14555 16975 14595 17015
rect 14605 16975 14645 17015
rect 14655 16975 14695 17015
rect 14705 16975 14745 17015
rect 14755 16975 14795 17015
rect 14805 16975 14845 17015
rect 14855 16975 14895 17015
rect 14905 16975 14945 17015
rect 14955 16975 14995 17015
rect 15005 16975 15045 17015
rect 15055 16975 15095 17015
rect 15105 16975 15145 17015
rect 15155 16975 15195 17015
rect 15205 16975 15245 17015
rect 15255 16975 15295 17015
rect 15305 16975 15345 17015
rect 15355 16975 15395 17015
rect 15405 16975 15445 17015
rect 15455 16975 15495 17015
rect 15505 16975 15545 17015
rect 15555 16975 15595 17015
rect 15605 16975 15645 17015
rect 15655 16975 15695 17015
rect 15705 16975 15745 17015
rect 15755 16975 15795 17015
rect 15805 16975 15845 17015
rect 15855 16975 15895 17015
rect 15905 16975 15945 17015
rect 15955 16975 15995 17015
rect 16005 16975 16045 17015
rect 16055 16975 16095 17015
rect 16105 16975 16145 17015
rect 16155 16975 16195 17015
rect 16205 16975 16245 17015
rect 16255 16975 16295 17015
rect 16305 16975 16345 17015
rect 16355 16975 16395 17015
rect 16405 16975 16445 17015
rect 16455 16975 16495 17015
rect 16505 16975 16545 17015
rect 16555 16975 16595 17015
rect 16605 16975 16645 17015
rect 16655 16975 16695 17015
rect 16705 16975 16745 17015
rect 16755 16975 16795 17015
rect 16805 16975 16845 17015
rect 16855 16975 16895 17015
rect 16905 16975 16945 17015
rect 16955 16975 16995 17015
rect 17005 16975 17045 17015
rect 17055 16975 17095 17015
rect 17105 16975 17145 17015
rect 17155 16975 17195 17015
rect 17205 16975 17245 17015
rect 17255 16975 17295 17015
rect 17305 16975 17345 17015
rect 17355 16975 17395 17015
rect 17405 16975 17445 17015
rect 17455 16975 17495 17015
rect 17505 16975 17545 17015
rect 17555 16975 17595 17015
rect 17605 16975 17645 17015
rect 17655 16975 17695 17015
rect 17705 16975 17745 17015
rect 17755 16975 17795 17015
rect 17805 16975 17845 17015
rect 17855 16975 17895 17015
rect 17905 16975 17945 17015
rect 17955 16975 17995 17015
rect 18005 16975 18045 17015
rect 18055 16975 18095 17015
rect 18105 16975 18145 17015
rect 18155 16975 18195 17015
rect 18205 16975 18245 17015
rect 18255 16975 18295 17015
rect 18305 16975 18345 17015
rect 18355 16975 18395 17015
rect 18405 16975 18445 17015
rect 18455 16975 18495 17015
rect 18505 16975 18545 17015
rect 18555 16975 18595 17015
rect 18605 16975 18645 17015
rect 18655 16975 18695 17015
rect 18705 16975 18745 17015
rect 18755 16975 18795 17015
rect 18805 16975 18845 17015
rect 18855 16975 18895 17015
rect 18905 16975 18945 17015
rect 18955 16975 18995 17015
rect 19005 16975 19045 17015
rect 19055 16975 19095 17015
rect 19105 16975 19145 17015
rect 19155 16975 19195 17015
rect 19205 16975 19245 17015
rect 19255 16975 19295 17015
rect 19305 16975 19345 17015
rect 19355 16975 19395 17015
rect 19405 16975 19445 17015
rect 19455 16975 19495 17015
rect 19505 16975 19545 17015
rect 19555 16975 19595 17015
rect 19605 16975 19645 17015
rect 19655 16975 19695 17015
rect 19705 16975 19745 17015
rect 19755 16975 19795 17015
rect 19805 16975 19845 17015
rect 19855 16975 19895 17015
rect 19905 16975 19945 17015
rect 19955 16975 19995 17015
rect 20005 16975 20045 17015
rect 20055 16975 20095 17015
rect 20105 16975 20145 17015
rect 20155 16975 20195 17015
rect 20205 16975 20245 17015
rect 20255 16975 20295 17015
rect 20305 16975 20345 17015
rect 20355 16975 20395 17015
rect 20405 16975 20445 17015
rect 20455 16975 20495 17015
rect 20505 16975 20545 17015
rect 20555 16975 20595 17015
rect 20605 16975 20645 17015
rect 20655 16975 20695 17015
rect 20705 16975 20745 17015
rect 20755 16975 20795 17015
rect 20805 16975 20845 17015
rect 20855 16975 20895 17015
rect 20905 16975 20945 17015
rect 20955 16975 20995 17015
rect 21005 16975 21045 17015
rect 21055 16975 21095 17015
rect 21105 16975 21145 17015
rect 21155 16975 21195 17015
rect 21205 16975 21245 17015
rect 21255 16975 21295 17015
rect 21305 16975 21345 17015
rect 21355 16975 21395 17015
rect 21405 16975 21445 17015
rect 21455 16975 21495 17015
rect 21505 16975 21545 17015
rect 21555 16975 21595 17015
rect 21605 16975 21645 17015
rect 21655 16975 21695 17015
rect 21705 16975 21745 17015
rect 21755 16975 21795 17015
rect 21805 16975 21845 17015
rect 21855 16975 21895 17015
rect 21905 16975 21945 17015
rect 21955 16975 21995 17015
rect 22005 16975 22045 17015
rect 22055 16975 22095 17015
rect 22105 16975 22145 17015
rect 22155 16975 22195 17015
rect 22205 16975 22245 17015
rect 22255 16975 22295 17015
rect 22305 16975 22345 17015
rect 22355 16975 22395 17015
rect 22405 16975 22445 17015
rect 22455 16975 22495 17015
rect 22505 16975 22545 17015
rect 22555 16975 22595 17015
rect 22605 16975 22645 17015
rect 22655 16975 22695 17015
rect 22705 16975 22745 17015
rect 22755 16975 22795 17015
rect 22805 16975 22845 17015
rect 22855 16975 22895 17015
rect 22905 16975 22945 17015
rect 22955 16975 22995 17015
rect 23005 16975 23045 17015
rect 23055 16975 23095 17015
rect 23105 16975 23145 17015
rect 23155 16975 23195 17015
rect 23205 16975 23245 17015
rect 23255 16975 23295 17015
rect 23305 16975 23345 17015
rect 23355 16975 23395 17015
rect 23405 16975 23445 17015
rect 23455 16975 23495 17015
rect 23505 16975 23545 17015
rect 23555 16975 23595 17015
rect 23605 16975 23645 17015
rect 23655 16975 23695 17015
rect 23705 16975 23745 17015
rect 23755 16975 23795 17015
rect 23805 16975 23845 17015
rect 23855 16975 23895 17015
rect 23905 16975 23945 17015
rect 23955 16975 23995 17015
rect 24005 16975 24045 17015
rect 24055 16975 24095 17015
rect 24105 16975 24145 17015
rect 24155 16975 24195 17015
rect 24205 16975 24245 17015
rect 24255 16975 24295 17015
rect 24305 16975 24345 17015
rect 24355 16975 24395 17015
rect 24405 16975 24445 17015
rect 24455 16975 24495 17015
rect 24505 16975 24545 17015
rect 24555 16975 24595 17015
rect 24605 16975 24645 17015
rect 24655 16975 24695 17015
rect 24705 16975 24745 17015
rect 24755 16975 24795 17015
rect 24805 16975 24845 17015
rect 24855 16975 24895 17015
rect 24905 16975 24945 17015
rect 24955 16975 24995 17015
rect 25005 16975 25045 17015
rect 25055 16975 25095 17015
rect 25105 16975 25145 17015
rect 25155 16975 25195 17015
rect 25205 16975 25245 17015
rect 25255 16975 25295 17015
rect 25305 16975 25345 17015
rect 25355 16975 25395 17015
rect 25405 16975 25445 17015
rect 25455 16975 25495 17015
rect 25505 16975 25545 17015
rect 25555 16975 25595 17015
rect 25605 16975 25645 17015
rect 25655 16975 25695 17015
rect 25705 16975 25745 17015
rect 25755 16975 25795 17015
rect 25805 16975 25845 17015
rect 25855 16975 25895 17015
rect 25905 16975 25945 17015
rect 25955 16975 25995 17015
rect 26005 16975 26045 17015
rect 26055 16975 26095 17015
rect 26105 16975 26145 17015
rect 26155 16975 26195 17015
rect 26205 16975 26245 17015
rect 26255 16975 26295 17015
rect 26305 16975 26345 17015
rect 26355 16975 26395 17015
rect 26405 16975 26445 17015
rect 26455 16975 26495 17015
rect 26505 16975 26545 17015
rect 26555 16975 26595 17015
rect 26605 16975 26645 17015
rect 26655 16975 26695 17015
rect 26705 16975 26745 17015
rect 26755 16975 26795 17015
rect 26805 16975 26845 17015
rect 26855 16975 26895 17015
rect 26905 16975 26945 17015
rect 26955 16975 26995 17015
rect 27005 16975 27045 17015
rect 27055 16975 27095 17015
rect 27105 16975 27145 17015
rect 27155 16975 27195 17015
rect 27205 16975 27245 17015
rect 27255 16975 27295 17015
rect 27305 16975 27345 17015
rect 27355 16975 27395 17015
rect 27405 16975 27445 17015
rect 27455 16975 27495 17015
rect 27505 16975 27545 17015
rect 27555 16975 27595 17015
rect 27605 16975 27645 17015
rect 27655 16975 27695 17015
rect 27705 16975 27745 17015
rect 27755 16975 27795 17015
rect 27805 16975 27845 17015
rect 27855 16975 27895 17015
rect 27905 16975 27945 17015
rect 27955 16975 27995 17015
rect 28005 16975 28045 17015
rect 28055 16975 28095 17015
rect 28105 16975 28145 17015
rect 28155 16975 28195 17015
rect 28205 16975 28245 17015
rect 28255 16975 28295 17015
rect 28305 16975 28345 17015
rect 28355 16975 28395 17015
rect 28405 16975 28445 17015
rect 28455 16975 28495 17015
rect 28505 16975 28545 17015
rect 28555 16975 28595 17015
rect 28605 16975 28645 17015
rect 28655 16975 28695 17015
rect 28705 16975 28745 17015
rect 28755 16975 28795 17015
rect 28805 16975 28845 17015
rect 28855 16975 28895 17015
rect 28905 16975 28945 17015
rect 28955 16975 28995 17015
rect 29005 16975 29045 17015
rect 29055 16975 29095 17015
rect 29105 16975 29145 17015
rect 29155 16975 29195 17015
rect 29205 16975 29245 17015
rect 29255 16975 29295 17015
rect 29305 16975 29345 17015
rect 29355 16975 29395 17015
rect 29405 16975 29445 17015
rect 29455 16975 29495 17015
rect 29505 16975 29545 17015
rect 29555 16975 29595 17015
rect 29605 16975 29645 17015
rect 29655 16975 29695 17015
rect 29705 16975 29745 17015
rect 29755 16975 29795 17015
rect 29805 16975 29845 17015
rect 29855 16975 29895 17015
rect 29905 16975 29945 17015
rect 29955 16975 29995 17015
rect 30005 16975 30045 17015
rect 30055 16975 30095 17015
rect 30105 16975 30145 17015
rect 30155 16975 30195 17015
rect 30205 16975 30245 17015
rect 30255 16975 30295 17015
rect 30305 16975 30345 17015
rect 30355 16975 30395 17015
rect 30405 16975 30445 17015
rect 30455 16975 30495 17015
rect 30505 16975 30545 17015
rect 30555 16975 30595 17015
rect 30605 16975 30645 17015
rect 30655 16975 30695 17015
rect 30705 16975 30745 17015
rect 30755 16975 30795 17015
rect 30805 16975 30845 17015
rect 30855 16975 30895 17015
rect 30905 16975 30945 17015
rect 30955 16975 30995 17015
rect 31005 16975 31045 17015
rect 31055 16975 31095 17015
rect 31105 16975 31145 17015
rect 31155 16975 31195 17015
rect 31205 16975 31245 17015
rect 31255 16975 31295 17015
rect 31305 16975 31345 17015
rect 31355 16975 31395 17015
rect 31405 16975 31445 17015
rect 31455 16975 31495 17015
rect 31505 16975 31545 17015
rect 31555 16975 31595 17015
rect 31605 16975 31645 17015
rect 31655 16975 31695 17015
rect 31705 16975 31745 17015
rect 31755 16975 31795 17015
rect 31805 16975 31845 17015
rect 31855 16975 31895 17015
rect 31905 16975 31945 17015
rect 31955 16975 31995 17015
rect 32005 16975 32045 17015
rect 32055 16975 32095 17015
rect 32105 16975 32145 17015
rect 32155 16975 32195 17015
rect 32205 16975 32245 17015
rect 32255 16975 32295 17015
rect 32305 16975 32345 17015
rect 32355 16975 32395 17015
rect 32405 16975 32445 17015
rect 32455 16975 32495 17015
rect 32505 16975 32545 17015
rect 32555 16975 32595 17015
rect 32605 16975 32645 17015
rect 32655 16975 32695 17015
rect 32705 16975 32745 17015
rect 32755 16975 32795 17015
rect 32805 16975 32845 17015
rect 32855 16975 32895 17015
rect 32905 16975 32945 17015
rect 32955 16975 32995 17015
rect 33005 16975 33045 17015
rect 33055 16975 33095 17015
rect 33105 16975 33145 17015
rect 33155 16975 33195 17015
rect 33205 16975 33245 17015
rect 33255 16975 33295 17015
rect 33305 16975 33345 17015
rect 33355 16975 33395 17015
rect 33405 16975 33445 17015
rect 33455 16975 33495 17015
rect 33505 16975 33545 17015
rect 33555 16975 33595 17015
rect 33605 16975 33645 17015
rect 33655 16975 33695 17015
rect 33705 16975 33745 17015
rect 33755 16975 33795 17015
rect 33805 16975 33845 17015
rect 33855 16975 33895 17015
rect 33905 16975 33945 17015
rect 33955 16975 33995 17015
rect 34005 16975 34045 17015
rect 34055 16975 34095 17015
rect 34105 16975 34145 17015
rect 34155 16975 34195 17015
rect 34205 16975 34245 17015
rect 34255 16975 34295 17015
rect 34305 16975 34345 17015
rect 34355 16975 34395 17015
rect 34405 16975 34445 17015
rect 34455 16975 34495 17015
rect 34505 16975 34545 17015
rect 34555 16975 34595 17015
rect 34605 16975 34645 17015
rect 34655 16975 34695 17015
rect 34705 16975 34745 17015
rect 34755 16975 34795 17015
rect 34805 16975 34845 17015
rect 34855 16975 34895 17015
rect 34905 16975 34945 17015
rect 34955 16975 34995 17015
rect 35005 16975 35045 17015
rect 35055 16975 35095 17015
rect 35105 16975 35145 17015
rect 35155 16975 35195 17015
rect 35205 16975 35245 17015
rect 35255 16975 35295 17015
rect 35305 16975 35345 17015
rect 35355 16975 35395 17015
rect 35405 16975 35445 17015
rect 35455 16975 35495 17015
rect 35505 16975 35545 17015
rect 35555 16975 35595 17015
rect 35605 16975 35645 17015
rect 35655 16975 35695 17015
rect 35705 16975 35745 17015
rect 35755 16975 35795 17015
rect 35805 16975 35845 17015
rect 35855 16975 35895 17015
rect 35905 16975 35945 17015
rect 35955 16975 35995 17015
rect 36005 16975 36045 17015
rect 36055 16975 36095 17015
rect 36105 16975 36145 17015
rect 36155 16975 36195 17015
rect 36205 16975 36245 17015
rect 36255 16975 36295 17015
rect 36305 16975 36345 17015
rect 36355 16975 36395 17015
rect 36405 16975 36445 17015
rect 36455 16975 36495 17015
rect 36505 16975 36545 17015
rect 36555 16975 36595 17015
rect 36605 16975 36645 17015
rect 36655 16975 36695 17015
rect 36705 16975 36745 17015
rect 36755 16975 36795 17015
rect 36805 16975 36845 17015
rect 36855 16975 36895 17015
rect 36905 16975 36945 17015
rect 36955 16975 36995 17015
rect 37005 16975 37045 17015
rect 37055 16975 37095 17015
rect 37105 16975 37145 17015
rect 37155 16975 37195 17015
rect 37205 16975 37245 17015
rect 37255 16975 37295 17015
rect 37305 16975 37345 17015
rect 37355 16975 37395 17015
rect 37405 16975 37445 17015
rect 37455 16975 37495 17015
rect 37505 16975 37545 17015
rect 37555 16975 37595 17015
rect 37605 16975 37645 17015
rect 37655 16975 37695 17015
rect 37705 16975 37745 17015
rect 37755 16975 37795 17015
rect 37805 16975 37845 17015
rect 37855 16975 37895 17015
rect 37905 16975 37945 17015
rect 37955 16975 37995 17015
rect 38005 16975 38045 17015
rect 38055 16975 38095 17015
rect 38105 16975 38145 17015
rect 38155 16975 38195 17015
rect 38205 16975 38245 17015
rect 38255 16975 38295 17015
rect 38305 16975 38345 17015
rect 38355 16975 38395 17015
rect 38405 16975 38445 17015
rect 38455 16975 38495 17015
rect 38505 16975 38545 17015
rect 38555 16975 38595 17015
rect 38605 16975 38645 17015
rect 38655 16975 38695 17015
rect 38705 16975 38745 17015
rect 38755 16975 38795 17015
rect 38805 16975 38845 17015
rect 38855 16975 38895 17015
rect 38905 16975 38945 17015
rect 38955 16975 38995 17015
rect 39005 16975 39045 17015
rect 39055 16975 39095 17015
rect 39105 16975 39145 17015
rect 39155 16975 39195 17015
rect 39205 16975 39245 17015
rect 39255 16975 39295 17015
rect 39305 16975 39345 17015
rect 39355 16975 39395 17015
rect 39405 16975 39445 17015
rect 39455 16975 39495 17015
rect 39505 16975 39545 17015
rect 39555 16975 39595 17015
rect 39605 16975 39645 17015
rect 39655 16975 39695 17015
rect 39705 16975 39745 17015
rect 39905 16975 39945 17015
rect 39955 16975 39995 17015
rect 40005 16975 40045 17015
rect 40055 16975 40095 17015
rect 40105 16975 40145 17015
rect 40155 16975 40195 17015
rect 40205 16975 40245 17015
rect 40255 16975 40295 17015
rect 40305 16975 40345 17015
rect 40355 16975 40395 17015
rect 40405 16975 40445 17015
rect 40455 16975 40495 17015
rect 40505 16975 40545 17015
rect 40555 16975 40595 17015
rect 40605 16975 40645 17015
rect 40655 16975 40695 17015
rect 40705 16975 40745 17015
rect 40755 16975 40795 17015
rect 40805 16975 40845 17015
rect 40855 16975 40895 17015
rect -395 16875 -355 16915
rect 105 16875 145 16915
rect 155 16875 195 16915
rect 205 16875 245 16915
rect 255 16875 295 16915
rect 305 16875 345 16915
rect 355 16875 395 16915
rect 405 16875 445 16915
rect 455 16875 495 16915
rect 505 16875 545 16915
rect 555 16875 595 16915
rect 605 16875 645 16915
rect 655 16875 695 16915
rect 705 16875 745 16915
rect 755 16875 795 16915
rect 805 16875 845 16915
rect 855 16875 895 16915
rect 905 16875 945 16915
rect 955 16875 995 16915
rect 1005 16875 1045 16915
rect 1055 16875 1095 16915
rect 1105 16875 1145 16915
rect 1155 16875 1195 16915
rect 1205 16875 1245 16915
rect 1255 16875 1295 16915
rect 1305 16875 1345 16915
rect 1355 16875 1395 16915
rect 1405 16875 1445 16915
rect 1455 16875 1495 16915
rect 1505 16875 1545 16915
rect 1555 16875 1595 16915
rect 1605 16875 1645 16915
rect 1655 16875 1695 16915
rect 1705 16875 1745 16915
rect 1755 16875 1795 16915
rect 1805 16875 1845 16915
rect 1855 16875 1895 16915
rect 1905 16875 1945 16915
rect 1955 16875 1995 16915
rect 2005 16875 2045 16915
rect 2055 16875 2095 16915
rect 2105 16875 2145 16915
rect 2155 16875 2195 16915
rect 2205 16875 2245 16915
rect 2255 16875 2295 16915
rect 2305 16875 2345 16915
rect 2355 16875 2395 16915
rect 2405 16875 2445 16915
rect 2455 16875 2495 16915
rect 2505 16875 2545 16915
rect 2555 16875 2595 16915
rect 2605 16875 2645 16915
rect 2655 16875 2695 16915
rect 2705 16875 2745 16915
rect 2755 16875 2795 16915
rect 2805 16875 2845 16915
rect 2855 16875 2895 16915
rect 2905 16875 2945 16915
rect 2955 16875 2995 16915
rect 3005 16875 3045 16915
rect 3055 16875 3095 16915
rect 3105 16875 3145 16915
rect 3155 16875 3195 16915
rect 3205 16875 3245 16915
rect 3255 16875 3295 16915
rect 3305 16875 3345 16915
rect 3355 16875 3395 16915
rect 3405 16875 3445 16915
rect 3455 16875 3495 16915
rect 3505 16875 3545 16915
rect 3555 16875 3595 16915
rect 3605 16875 3645 16915
rect 3655 16875 3695 16915
rect 3705 16875 3745 16915
rect 3755 16875 3795 16915
rect 3805 16875 3845 16915
rect 3855 16875 3895 16915
rect 3905 16875 3945 16915
rect 3955 16875 3995 16915
rect 4005 16875 4045 16915
rect 4055 16875 4095 16915
rect 4105 16875 4145 16915
rect 4155 16875 4195 16915
rect 4205 16875 4245 16915
rect 4255 16875 4295 16915
rect 4305 16875 4345 16915
rect 4355 16875 4395 16915
rect 4405 16875 4445 16915
rect 4455 16875 4495 16915
rect 4505 16875 4545 16915
rect 4555 16875 4595 16915
rect 4605 16875 4645 16915
rect 4655 16875 4695 16915
rect 4705 16875 4745 16915
rect 4755 16875 4795 16915
rect 4805 16875 4845 16915
rect 4855 16875 4895 16915
rect 4905 16875 4945 16915
rect 4955 16875 4995 16915
rect 5005 16875 5045 16915
rect 5055 16875 5095 16915
rect 5105 16875 5145 16915
rect 5155 16875 5195 16915
rect 5205 16875 5245 16915
rect 5255 16875 5295 16915
rect 5305 16875 5345 16915
rect 5355 16875 5395 16915
rect 5405 16875 5445 16915
rect 5455 16875 5495 16915
rect 5505 16875 5545 16915
rect 5555 16875 5595 16915
rect 5605 16875 5645 16915
rect 5655 16875 5695 16915
rect 5705 16875 5745 16915
rect 5755 16875 5795 16915
rect 5805 16875 5845 16915
rect 5855 16875 5895 16915
rect 5905 16875 5945 16915
rect 5955 16875 5995 16915
rect 6005 16875 6045 16915
rect 6055 16875 6095 16915
rect 6105 16875 6145 16915
rect 6155 16875 6195 16915
rect 6205 16875 6245 16915
rect 6255 16875 6295 16915
rect 6305 16875 6345 16915
rect 6355 16875 6395 16915
rect 6405 16875 6445 16915
rect 6455 16875 6495 16915
rect 6505 16875 6545 16915
rect 6555 16875 6595 16915
rect 6605 16875 6645 16915
rect 6655 16875 6695 16915
rect 6705 16875 6745 16915
rect 6755 16875 6795 16915
rect 6805 16875 6845 16915
rect 6855 16875 6895 16915
rect 6905 16875 6945 16915
rect 6955 16875 6995 16915
rect 7005 16875 7045 16915
rect 7055 16875 7095 16915
rect 7105 16875 7145 16915
rect 7155 16875 7195 16915
rect 7205 16875 7245 16915
rect 7255 16875 7295 16915
rect 7305 16875 7345 16915
rect 7355 16875 7395 16915
rect 7405 16875 7445 16915
rect 7455 16875 7495 16915
rect 7505 16875 7545 16915
rect 7555 16875 7595 16915
rect 7605 16875 7645 16915
rect 7655 16875 7695 16915
rect 7705 16875 7745 16915
rect 7755 16875 7795 16915
rect 7805 16875 7845 16915
rect 7855 16875 7895 16915
rect 7905 16875 7945 16915
rect 7955 16875 7995 16915
rect 8005 16875 8045 16915
rect 8055 16875 8095 16915
rect 8105 16875 8145 16915
rect 8155 16875 8195 16915
rect 8205 16875 8245 16915
rect 8255 16875 8295 16915
rect 8305 16875 8345 16915
rect 8355 16875 8395 16915
rect 8405 16875 8445 16915
rect 8455 16875 8495 16915
rect 8505 16875 8545 16915
rect 8555 16875 8595 16915
rect 8605 16875 8645 16915
rect 8655 16875 8695 16915
rect 8705 16875 8745 16915
rect 8755 16875 8795 16915
rect 8805 16875 8845 16915
rect 8855 16875 8895 16915
rect 8905 16875 8945 16915
rect 8955 16875 8995 16915
rect 9005 16875 9045 16915
rect 9055 16875 9095 16915
rect 9105 16875 9145 16915
rect 9155 16875 9195 16915
rect 9205 16875 9245 16915
rect 9255 16875 9295 16915
rect 9305 16875 9345 16915
rect 9355 16875 9395 16915
rect 9405 16875 9445 16915
rect 9455 16875 9495 16915
rect 9505 16875 9545 16915
rect 9555 16875 9595 16915
rect 9605 16875 9645 16915
rect 9655 16875 9695 16915
rect 9705 16875 9745 16915
rect 9755 16875 9795 16915
rect 9805 16875 9845 16915
rect 9855 16875 9895 16915
rect 9905 16875 9945 16915
rect 9955 16875 9995 16915
rect 10005 16875 10045 16915
rect 10055 16875 10095 16915
rect 10105 16875 10145 16915
rect 10155 16875 10195 16915
rect 10205 16875 10245 16915
rect 10255 16875 10295 16915
rect 10305 16875 10345 16915
rect 10355 16875 10395 16915
rect 10405 16875 10445 16915
rect 10455 16875 10495 16915
rect 10505 16875 10545 16915
rect 10555 16875 10595 16915
rect 10605 16875 10645 16915
rect 10655 16875 10695 16915
rect 10705 16875 10745 16915
rect 10755 16875 10795 16915
rect 10805 16875 10845 16915
rect 10855 16875 10895 16915
rect 10905 16875 10945 16915
rect 10955 16875 10995 16915
rect 11005 16875 11045 16915
rect 11055 16875 11095 16915
rect 11105 16875 11145 16915
rect 11155 16875 11195 16915
rect 11205 16875 11245 16915
rect 11255 16875 11295 16915
rect 11305 16875 11345 16915
rect 11355 16875 11395 16915
rect 11405 16875 11445 16915
rect 11455 16875 11495 16915
rect 11505 16875 11545 16915
rect 11555 16875 11595 16915
rect 11605 16875 11645 16915
rect 11655 16875 11695 16915
rect 11705 16875 11745 16915
rect 11755 16875 11795 16915
rect 11805 16875 11845 16915
rect 11855 16875 11895 16915
rect 11905 16875 11945 16915
rect 11955 16875 11995 16915
rect 12005 16875 12045 16915
rect 12055 16875 12095 16915
rect 12105 16875 12145 16915
rect 12155 16875 12195 16915
rect 12205 16875 12245 16915
rect 12255 16875 12295 16915
rect 12305 16875 12345 16915
rect 12355 16875 12395 16915
rect 12405 16875 12445 16915
rect 12455 16875 12495 16915
rect 12505 16875 12545 16915
rect 12555 16875 12595 16915
rect 12605 16875 12645 16915
rect 12655 16875 12695 16915
rect 12705 16875 12745 16915
rect 12755 16875 12795 16915
rect 12805 16875 12845 16915
rect 12855 16875 12895 16915
rect 12905 16875 12945 16915
rect 12955 16875 12995 16915
rect 13005 16875 13045 16915
rect 13055 16875 13095 16915
rect 13105 16875 13145 16915
rect 13155 16875 13195 16915
rect 13205 16875 13245 16915
rect 13255 16875 13295 16915
rect 13305 16875 13345 16915
rect 13355 16875 13395 16915
rect 13405 16875 13445 16915
rect 13455 16875 13495 16915
rect 13505 16875 13545 16915
rect 13555 16875 13595 16915
rect 13605 16875 13645 16915
rect 13655 16875 13695 16915
rect 13705 16875 13745 16915
rect 13755 16875 13795 16915
rect 13805 16875 13845 16915
rect 13855 16875 13895 16915
rect 13905 16875 13945 16915
rect 13955 16875 13995 16915
rect 14005 16875 14045 16915
rect 14055 16875 14095 16915
rect 14105 16875 14145 16915
rect 14155 16875 14195 16915
rect 14205 16875 14245 16915
rect 14255 16875 14295 16915
rect 14305 16875 14345 16915
rect 14355 16875 14395 16915
rect 14405 16875 14445 16915
rect 14455 16875 14495 16915
rect 14505 16875 14545 16915
rect 14555 16875 14595 16915
rect 14605 16875 14645 16915
rect 14655 16875 14695 16915
rect 14705 16875 14745 16915
rect 14755 16875 14795 16915
rect 14805 16875 14845 16915
rect 14855 16875 14895 16915
rect 14905 16875 14945 16915
rect 14955 16875 14995 16915
rect 15005 16875 15045 16915
rect 15055 16875 15095 16915
rect 15105 16875 15145 16915
rect 15155 16875 15195 16915
rect 15205 16875 15245 16915
rect 15255 16875 15295 16915
rect 15305 16875 15345 16915
rect 15355 16875 15395 16915
rect 15405 16875 15445 16915
rect 15455 16875 15495 16915
rect 15505 16875 15545 16915
rect 15555 16875 15595 16915
rect 15605 16875 15645 16915
rect 15655 16875 15695 16915
rect 15705 16875 15745 16915
rect 15755 16875 15795 16915
rect 15805 16875 15845 16915
rect 15855 16875 15895 16915
rect 15905 16875 15945 16915
rect 15955 16875 15995 16915
rect 16005 16875 16045 16915
rect 16055 16875 16095 16915
rect 16105 16875 16145 16915
rect 16155 16875 16195 16915
rect 16205 16875 16245 16915
rect 16255 16875 16295 16915
rect 16305 16875 16345 16915
rect 16355 16875 16395 16915
rect 16405 16875 16445 16915
rect 16455 16875 16495 16915
rect 16505 16875 16545 16915
rect 16555 16875 16595 16915
rect 16605 16875 16645 16915
rect 16655 16875 16695 16915
rect 16705 16875 16745 16915
rect 16755 16875 16795 16915
rect 16805 16875 16845 16915
rect 16855 16875 16895 16915
rect 16905 16875 16945 16915
rect 16955 16875 16995 16915
rect 17005 16875 17045 16915
rect 17055 16875 17095 16915
rect 17105 16875 17145 16915
rect 17155 16875 17195 16915
rect 17205 16875 17245 16915
rect 17255 16875 17295 16915
rect 17305 16875 17345 16915
rect 17355 16875 17395 16915
rect 17405 16875 17445 16915
rect 17455 16875 17495 16915
rect 17505 16875 17545 16915
rect 17555 16875 17595 16915
rect 17605 16875 17645 16915
rect 17655 16875 17695 16915
rect 17705 16875 17745 16915
rect 17755 16875 17795 16915
rect 17805 16875 17845 16915
rect 17855 16875 17895 16915
rect 17905 16875 17945 16915
rect 17955 16875 17995 16915
rect 18005 16875 18045 16915
rect 18055 16875 18095 16915
rect 18105 16875 18145 16915
rect 18155 16875 18195 16915
rect 18205 16875 18245 16915
rect 18255 16875 18295 16915
rect 18305 16875 18345 16915
rect 18355 16875 18395 16915
rect 18405 16875 18445 16915
rect 18455 16875 18495 16915
rect 18505 16875 18545 16915
rect 18555 16875 18595 16915
rect 18605 16875 18645 16915
rect 18655 16875 18695 16915
rect 18705 16875 18745 16915
rect 18755 16875 18795 16915
rect 18805 16875 18845 16915
rect 18855 16875 18895 16915
rect 18905 16875 18945 16915
rect 18955 16875 18995 16915
rect 19005 16875 19045 16915
rect 19055 16875 19095 16915
rect 19105 16875 19145 16915
rect 19155 16875 19195 16915
rect 19205 16875 19245 16915
rect 19255 16875 19295 16915
rect 19305 16875 19345 16915
rect 19355 16875 19395 16915
rect 19405 16875 19445 16915
rect 19455 16875 19495 16915
rect 19505 16875 19545 16915
rect 19555 16875 19595 16915
rect 19605 16875 19645 16915
rect 19655 16875 19695 16915
rect 19705 16875 19745 16915
rect 19755 16875 19795 16915
rect 19805 16875 19845 16915
rect 19855 16875 19895 16915
rect 19905 16875 19945 16915
rect 19955 16875 19995 16915
rect 20005 16875 20045 16915
rect 20055 16875 20095 16915
rect 20105 16875 20145 16915
rect 20155 16875 20195 16915
rect 20205 16875 20245 16915
rect 20255 16875 20295 16915
rect 20305 16875 20345 16915
rect 20355 16875 20395 16915
rect 20405 16875 20445 16915
rect 20455 16875 20495 16915
rect 20505 16875 20545 16915
rect 20555 16875 20595 16915
rect 20605 16875 20645 16915
rect 20655 16875 20695 16915
rect 20705 16875 20745 16915
rect 20755 16875 20795 16915
rect 20805 16875 20845 16915
rect 20855 16875 20895 16915
rect 20905 16875 20945 16915
rect 20955 16875 20995 16915
rect 21005 16875 21045 16915
rect 21055 16875 21095 16915
rect 21105 16875 21145 16915
rect 21155 16875 21195 16915
rect 21205 16875 21245 16915
rect 21255 16875 21295 16915
rect 21305 16875 21345 16915
rect 21355 16875 21395 16915
rect 21405 16875 21445 16915
rect 21455 16875 21495 16915
rect 21505 16875 21545 16915
rect 21555 16875 21595 16915
rect 21605 16875 21645 16915
rect 21655 16875 21695 16915
rect 21705 16875 21745 16915
rect 21755 16875 21795 16915
rect 21805 16875 21845 16915
rect 21855 16875 21895 16915
rect 21905 16875 21945 16915
rect 21955 16875 21995 16915
rect 22005 16875 22045 16915
rect 22055 16875 22095 16915
rect 22105 16875 22145 16915
rect 22155 16875 22195 16915
rect 22205 16875 22245 16915
rect 22255 16875 22295 16915
rect 22305 16875 22345 16915
rect 22355 16875 22395 16915
rect 22405 16875 22445 16915
rect 22455 16875 22495 16915
rect 22505 16875 22545 16915
rect 22555 16875 22595 16915
rect 22605 16875 22645 16915
rect 22655 16875 22695 16915
rect 22705 16875 22745 16915
rect 22755 16875 22795 16915
rect 22805 16875 22845 16915
rect 22855 16875 22895 16915
rect 22905 16875 22945 16915
rect 22955 16875 22995 16915
rect 23005 16875 23045 16915
rect 23055 16875 23095 16915
rect 23105 16875 23145 16915
rect 23155 16875 23195 16915
rect 23205 16875 23245 16915
rect 23255 16875 23295 16915
rect 23305 16875 23345 16915
rect 23355 16875 23395 16915
rect 23405 16875 23445 16915
rect 23455 16875 23495 16915
rect 23505 16875 23545 16915
rect 23555 16875 23595 16915
rect 23605 16875 23645 16915
rect 23655 16875 23695 16915
rect 23705 16875 23745 16915
rect 23755 16875 23795 16915
rect 23805 16875 23845 16915
rect 23855 16875 23895 16915
rect 23905 16875 23945 16915
rect 23955 16875 23995 16915
rect 24005 16875 24045 16915
rect 24055 16875 24095 16915
rect 24105 16875 24145 16915
rect 24155 16875 24195 16915
rect 24205 16875 24245 16915
rect 24255 16875 24295 16915
rect 24305 16875 24345 16915
rect 24355 16875 24395 16915
rect 24405 16875 24445 16915
rect 24455 16875 24495 16915
rect 24505 16875 24545 16915
rect 24555 16875 24595 16915
rect 24605 16875 24645 16915
rect 24655 16875 24695 16915
rect 24705 16875 24745 16915
rect 24755 16875 24795 16915
rect 24805 16875 24845 16915
rect 24855 16875 24895 16915
rect 24905 16875 24945 16915
rect 24955 16875 24995 16915
rect 25005 16875 25045 16915
rect 25055 16875 25095 16915
rect 25105 16875 25145 16915
rect 25155 16875 25195 16915
rect 25205 16875 25245 16915
rect 25255 16875 25295 16915
rect 25305 16875 25345 16915
rect 25355 16875 25395 16915
rect 25405 16875 25445 16915
rect 25455 16875 25495 16915
rect 25505 16875 25545 16915
rect 25555 16875 25595 16915
rect 25605 16875 25645 16915
rect 25655 16875 25695 16915
rect 25705 16875 25745 16915
rect 25755 16875 25795 16915
rect 25805 16875 25845 16915
rect 25855 16875 25895 16915
rect 25905 16875 25945 16915
rect 25955 16875 25995 16915
rect 26005 16875 26045 16915
rect 26055 16875 26095 16915
rect 26105 16875 26145 16915
rect 26155 16875 26195 16915
rect 26205 16875 26245 16915
rect 26255 16875 26295 16915
rect 26305 16875 26345 16915
rect 26355 16875 26395 16915
rect 26405 16875 26445 16915
rect 26455 16875 26495 16915
rect 26505 16875 26545 16915
rect 26555 16875 26595 16915
rect 26605 16875 26645 16915
rect 26655 16875 26695 16915
rect 26705 16875 26745 16915
rect 26755 16875 26795 16915
rect 26805 16875 26845 16915
rect 26855 16875 26895 16915
rect 26905 16875 26945 16915
rect 26955 16875 26995 16915
rect 27005 16875 27045 16915
rect 27055 16875 27095 16915
rect 27105 16875 27145 16915
rect 27155 16875 27195 16915
rect 27205 16875 27245 16915
rect 27255 16875 27295 16915
rect 27305 16875 27345 16915
rect 27355 16875 27395 16915
rect 27405 16875 27445 16915
rect 27455 16875 27495 16915
rect 27505 16875 27545 16915
rect 27555 16875 27595 16915
rect 27605 16875 27645 16915
rect 27655 16875 27695 16915
rect 27705 16875 27745 16915
rect 27755 16875 27795 16915
rect 27805 16875 27845 16915
rect 27855 16875 27895 16915
rect 27905 16875 27945 16915
rect 27955 16875 27995 16915
rect 28005 16875 28045 16915
rect 28055 16875 28095 16915
rect 28105 16875 28145 16915
rect 28155 16875 28195 16915
rect 28205 16875 28245 16915
rect 28255 16875 28295 16915
rect 28305 16875 28345 16915
rect 28355 16875 28395 16915
rect 28405 16875 28445 16915
rect 28455 16875 28495 16915
rect 28505 16875 28545 16915
rect 28555 16875 28595 16915
rect 28605 16875 28645 16915
rect 28655 16875 28695 16915
rect 28705 16875 28745 16915
rect 28755 16875 28795 16915
rect 28805 16875 28845 16915
rect 28855 16875 28895 16915
rect 28905 16875 28945 16915
rect 28955 16875 28995 16915
rect 29005 16875 29045 16915
rect 29055 16875 29095 16915
rect 29105 16875 29145 16915
rect 29155 16875 29195 16915
rect 29205 16875 29245 16915
rect 29255 16875 29295 16915
rect 29305 16875 29345 16915
rect 29355 16875 29395 16915
rect 29405 16875 29445 16915
rect 29455 16875 29495 16915
rect 29505 16875 29545 16915
rect 29555 16875 29595 16915
rect 29605 16875 29645 16915
rect 29655 16875 29695 16915
rect 29705 16875 29745 16915
rect 29755 16875 29795 16915
rect 29805 16875 29845 16915
rect 29855 16875 29895 16915
rect 29905 16875 29945 16915
rect 29955 16875 29995 16915
rect 30005 16875 30045 16915
rect 30055 16875 30095 16915
rect 30105 16875 30145 16915
rect 30155 16875 30195 16915
rect 30205 16875 30245 16915
rect 30255 16875 30295 16915
rect 30305 16875 30345 16915
rect 30355 16875 30395 16915
rect 30405 16875 30445 16915
rect 30455 16875 30495 16915
rect 30505 16875 30545 16915
rect 30555 16875 30595 16915
rect 30605 16875 30645 16915
rect 30655 16875 30695 16915
rect 30705 16875 30745 16915
rect 30755 16875 30795 16915
rect 30805 16875 30845 16915
rect 30855 16875 30895 16915
rect 30905 16875 30945 16915
rect 30955 16875 30995 16915
rect 31005 16875 31045 16915
rect 31055 16875 31095 16915
rect 31105 16875 31145 16915
rect 31155 16875 31195 16915
rect 31205 16875 31245 16915
rect 31255 16875 31295 16915
rect 31305 16875 31345 16915
rect 31355 16875 31395 16915
rect 31405 16875 31445 16915
rect 31455 16875 31495 16915
rect 31505 16875 31545 16915
rect 31555 16875 31595 16915
rect 31605 16875 31645 16915
rect 31655 16875 31695 16915
rect 31705 16875 31745 16915
rect 31755 16875 31795 16915
rect 31805 16875 31845 16915
rect 31855 16875 31895 16915
rect 31905 16875 31945 16915
rect 31955 16875 31995 16915
rect 32005 16875 32045 16915
rect 32055 16875 32095 16915
rect 32105 16875 32145 16915
rect 32155 16875 32195 16915
rect 32205 16875 32245 16915
rect 32255 16875 32295 16915
rect 32305 16875 32345 16915
rect 32355 16875 32395 16915
rect 32405 16875 32445 16915
rect 32455 16875 32495 16915
rect 32505 16875 32545 16915
rect 32555 16875 32595 16915
rect 32605 16875 32645 16915
rect 32655 16875 32695 16915
rect 32705 16875 32745 16915
rect 32755 16875 32795 16915
rect 32805 16875 32845 16915
rect 32855 16875 32895 16915
rect 32905 16875 32945 16915
rect 32955 16875 32995 16915
rect 33005 16875 33045 16915
rect 33055 16875 33095 16915
rect 33105 16875 33145 16915
rect 33155 16875 33195 16915
rect 33205 16875 33245 16915
rect 33255 16875 33295 16915
rect 33305 16875 33345 16915
rect 33355 16875 33395 16915
rect 33405 16875 33445 16915
rect 33455 16875 33495 16915
rect 33505 16875 33545 16915
rect 33555 16875 33595 16915
rect 33605 16875 33645 16915
rect 33655 16875 33695 16915
rect 33705 16875 33745 16915
rect 33755 16875 33795 16915
rect 33805 16875 33845 16915
rect 33855 16875 33895 16915
rect 33905 16875 33945 16915
rect 33955 16875 33995 16915
rect 34005 16875 34045 16915
rect 34055 16875 34095 16915
rect 34105 16875 34145 16915
rect 34155 16875 34195 16915
rect 34205 16875 34245 16915
rect 34255 16875 34295 16915
rect 34305 16875 34345 16915
rect 34355 16875 34395 16915
rect 34405 16875 34445 16915
rect 34455 16875 34495 16915
rect 34505 16875 34545 16915
rect 34555 16875 34595 16915
rect 34605 16875 34645 16915
rect 34655 16875 34695 16915
rect 34705 16875 34745 16915
rect 34755 16875 34795 16915
rect 34805 16875 34845 16915
rect 34855 16875 34895 16915
rect 34905 16875 34945 16915
rect 34955 16875 34995 16915
rect 35005 16875 35045 16915
rect 35055 16875 35095 16915
rect 35105 16875 35145 16915
rect 35155 16875 35195 16915
rect 35205 16875 35245 16915
rect 35255 16875 35295 16915
rect 35305 16875 35345 16915
rect 35355 16875 35395 16915
rect 35405 16875 35445 16915
rect 35455 16875 35495 16915
rect 35505 16875 35545 16915
rect 35555 16875 35595 16915
rect 35605 16875 35645 16915
rect 35655 16875 35695 16915
rect 35705 16875 35745 16915
rect 35755 16875 35795 16915
rect 35805 16875 35845 16915
rect 35855 16875 35895 16915
rect 35905 16875 35945 16915
rect 35955 16875 35995 16915
rect 36005 16875 36045 16915
rect 36055 16875 36095 16915
rect 36105 16875 36145 16915
rect 36155 16875 36195 16915
rect 36205 16875 36245 16915
rect 36255 16875 36295 16915
rect 36305 16875 36345 16915
rect 36355 16875 36395 16915
rect 36405 16875 36445 16915
rect 36455 16875 36495 16915
rect 36505 16875 36545 16915
rect 36555 16875 36595 16915
rect 36605 16875 36645 16915
rect 36655 16875 36695 16915
rect 36705 16875 36745 16915
rect 36755 16875 36795 16915
rect 36805 16875 36845 16915
rect 36855 16875 36895 16915
rect 36905 16875 36945 16915
rect 36955 16875 36995 16915
rect 37005 16875 37045 16915
rect 37055 16875 37095 16915
rect 37105 16875 37145 16915
rect 37155 16875 37195 16915
rect 37205 16875 37245 16915
rect 37255 16875 37295 16915
rect 37305 16875 37345 16915
rect 37355 16875 37395 16915
rect 37405 16875 37445 16915
rect 37455 16875 37495 16915
rect 37505 16875 37545 16915
rect 37555 16875 37595 16915
rect 37605 16875 37645 16915
rect 37655 16875 37695 16915
rect 37705 16875 37745 16915
rect 37755 16875 37795 16915
rect 37805 16875 37845 16915
rect 37855 16875 37895 16915
rect 37905 16875 37945 16915
rect 37955 16875 37995 16915
rect 38005 16875 38045 16915
rect 38055 16875 38095 16915
rect 38105 16875 38145 16915
rect 38155 16875 38195 16915
rect 38205 16875 38245 16915
rect 38255 16875 38295 16915
rect 38305 16875 38345 16915
rect 38355 16875 38395 16915
rect 38405 16875 38445 16915
rect 38455 16875 38495 16915
rect 38505 16875 38545 16915
rect 38555 16875 38595 16915
rect 38605 16875 38645 16915
rect 38655 16875 38695 16915
rect 38705 16875 38745 16915
rect 38755 16875 38795 16915
rect 38805 16875 38845 16915
rect 38855 16875 38895 16915
rect 38905 16875 38945 16915
rect 38955 16875 38995 16915
rect 39005 16875 39045 16915
rect 39055 16875 39095 16915
rect 39105 16875 39145 16915
rect 39155 16875 39195 16915
rect 39205 16875 39245 16915
rect 39255 16875 39295 16915
rect 39305 16875 39345 16915
rect 39355 16875 39395 16915
rect 39405 16875 39445 16915
rect 39455 16875 39495 16915
rect 39505 16875 39545 16915
rect 39555 16875 39595 16915
rect 39605 16875 39645 16915
rect 39655 16875 39695 16915
rect 39705 16875 39745 16915
rect 5 15805 45 15845
rect 55 15805 95 15845
rect 105 15805 145 15845
rect 155 15805 195 15845
rect 205 15805 245 15845
rect 255 15805 295 15845
rect 305 15805 345 15845
rect 355 15805 395 15845
rect 405 15805 445 15845
rect 455 15805 495 15845
rect 505 15805 545 15845
rect 555 15805 595 15845
rect 605 15805 645 15845
rect 655 15805 695 15845
rect 705 15805 745 15845
rect 755 15805 795 15845
rect 805 15805 845 15845
rect 855 15805 895 15845
rect 905 15805 945 15845
rect 955 15805 995 15845
rect 1005 15805 1045 15845
rect 1055 15805 1095 15845
rect 1105 15805 1145 15845
rect 1155 15805 1195 15845
rect 1205 15805 1245 15845
rect 1255 15805 1295 15845
rect 1305 15805 1345 15845
rect 1355 15805 1395 15845
rect 1405 15805 1445 15845
rect 1455 15805 1495 15845
rect 1505 15805 1545 15845
rect 1555 15805 1595 15845
rect 1605 15805 1645 15845
rect 1655 15805 1695 15845
rect 1705 15805 1745 15845
rect 1755 15805 1795 15845
rect 1805 15805 1845 15845
rect 1855 15805 1895 15845
rect 1905 15805 1945 15845
rect 1955 15805 1995 15845
rect 2005 15805 2045 15845
rect 2055 15805 2095 15845
rect 2105 15805 2145 15845
rect 2155 15805 2195 15845
rect 2205 15805 2245 15845
rect 2255 15805 2295 15845
rect 2305 15805 2345 15845
rect 2355 15805 2395 15845
rect 2405 15805 2445 15845
rect 2455 15805 2495 15845
rect 2505 15805 2545 15845
rect 2555 15805 2595 15845
rect 2605 15805 2645 15845
rect 2655 15805 2695 15845
rect 2705 15805 2745 15845
rect 2755 15805 2795 15845
rect 2805 15805 2845 15845
rect 2855 15805 2895 15845
rect 2905 15805 2945 15845
rect 2955 15805 2995 15845
rect 3005 15805 3045 15845
rect 3055 15805 3095 15845
rect 3105 15805 3145 15845
rect 3155 15805 3195 15845
rect 3205 15805 3245 15845
rect 3255 15805 3295 15845
rect 3305 15805 3345 15845
rect 3355 15805 3395 15845
rect 3405 15805 3445 15845
rect 3455 15805 3495 15845
rect 3505 15805 3545 15845
rect 3555 15805 3595 15845
rect 3605 15805 3645 15845
rect 3655 15805 3695 15845
rect 3705 15805 3745 15845
rect 3755 15805 3795 15845
rect 3805 15805 3845 15845
rect 3855 15805 3895 15845
rect 3905 15805 3945 15845
rect 3955 15805 3995 15845
rect 4005 15805 4045 15845
rect 4055 15805 4095 15845
rect 4105 15805 4145 15845
rect 4155 15805 4195 15845
rect 4205 15805 4245 15845
rect 4255 15805 4295 15845
rect 4305 15805 4345 15845
rect 4355 15805 4395 15845
rect 4405 15805 4445 15845
rect 4455 15805 4495 15845
rect 4505 15805 4545 15845
rect 4555 15805 4595 15845
rect 4605 15805 4645 15845
rect 4655 15805 4695 15845
rect 4705 15805 4745 15845
rect 4755 15805 4795 15845
rect 4805 15805 4845 15845
rect 4855 15805 4895 15845
rect 4905 15805 4945 15845
rect 4955 15805 4995 15845
rect 5005 15805 5045 15845
rect 5055 15805 5095 15845
rect 5105 15805 5145 15845
rect 5155 15805 5195 15845
rect 5205 15805 5245 15845
rect 5255 15805 5295 15845
rect 5305 15805 5345 15845
rect 5355 15805 5395 15845
rect 5405 15805 5445 15845
rect 5455 15805 5495 15845
rect 5505 15805 5545 15845
rect 5555 15805 5595 15845
rect 5605 15805 5645 15845
rect 5655 15805 5695 15845
rect 5705 15805 5745 15845
rect 5755 15805 5795 15845
rect 5805 15805 5845 15845
rect 5855 15805 5895 15845
rect 5905 15805 5945 15845
rect 5955 15805 5995 15845
rect 6005 15805 6045 15845
rect 6055 15805 6095 15845
rect 6105 15805 6145 15845
rect 6155 15805 6195 15845
rect 6205 15805 6245 15845
rect 6255 15805 6295 15845
rect 6305 15805 6345 15845
rect 6355 15805 6395 15845
rect 6405 15805 6445 15845
rect 6455 15805 6495 15845
rect 6505 15805 6545 15845
rect 6555 15805 6595 15845
rect 6605 15805 6645 15845
rect 6655 15805 6695 15845
rect 6705 15805 6745 15845
rect 6755 15805 6795 15845
rect 6805 15805 6845 15845
rect 6855 15805 6895 15845
rect 6905 15805 6945 15845
rect 6955 15805 6995 15845
rect 7005 15805 7045 15845
rect 7055 15805 7095 15845
rect 7105 15805 7145 15845
rect 7155 15805 7195 15845
rect 7205 15805 7245 15845
rect 7255 15805 7295 15845
rect 7305 15805 7345 15845
rect 7355 15805 7395 15845
rect 7405 15805 7445 15845
rect 7455 15805 7495 15845
rect 7505 15805 7545 15845
rect 7555 15805 7595 15845
rect 7605 15805 7645 15845
rect 7655 15805 7695 15845
rect 7705 15805 7745 15845
rect 7755 15805 7795 15845
rect 7805 15805 7845 15845
rect 7855 15805 7895 15845
rect 7905 15805 7945 15845
rect 7955 15805 7995 15845
rect 8005 15805 8045 15845
rect 8055 15805 8095 15845
rect 8105 15805 8145 15845
rect 8155 15805 8195 15845
rect 8205 15805 8245 15845
rect 8255 15805 8295 15845
rect 8305 15805 8345 15845
rect 8355 15805 8395 15845
rect 8405 15805 8445 15845
rect 8455 15805 8495 15845
rect 8505 15805 8545 15845
rect 8555 15805 8595 15845
rect 8605 15805 8645 15845
rect 8655 15805 8695 15845
rect 8705 15805 8745 15845
rect 8755 15805 8795 15845
rect 8805 15805 8845 15845
rect 8855 15805 8895 15845
rect 8905 15805 8945 15845
rect 8955 15805 8995 15845
rect 9005 15805 9045 15845
rect 9055 15805 9095 15845
rect 9105 15805 9145 15845
rect 9155 15805 9195 15845
rect 9205 15805 9245 15845
rect 9255 15805 9295 15845
rect 9305 15805 9345 15845
rect 9355 15805 9395 15845
rect 9405 15805 9445 15845
rect 9455 15805 9495 15845
rect 9505 15805 9545 15845
rect 9555 15805 9595 15845
rect 9605 15805 9645 15845
rect 9655 15805 9695 15845
rect 9705 15805 9745 15845
rect 9755 15805 9795 15845
rect 9805 15805 9845 15845
rect 9855 15805 9895 15845
rect 9905 15805 9945 15845
rect 9955 15805 9995 15845
rect 10005 15805 10045 15845
rect 10055 15805 10095 15845
rect 10105 15805 10145 15845
rect 10155 15805 10195 15845
rect 10205 15805 10245 15845
rect 10255 15805 10295 15845
rect 10305 15805 10345 15845
rect 10355 15805 10395 15845
rect 10405 15805 10445 15845
rect 10455 15805 10495 15845
rect 10505 15805 10545 15845
rect 10555 15805 10595 15845
rect 10605 15805 10645 15845
rect 10655 15805 10695 15845
rect 10705 15805 10745 15845
rect 10755 15805 10795 15845
rect 10805 15805 10845 15845
rect 10855 15805 10895 15845
rect 10905 15805 10945 15845
rect 10955 15805 10995 15845
rect 11005 15805 11045 15845
rect 11055 15805 11095 15845
rect 11105 15805 11145 15845
rect 11155 15805 11195 15845
rect 11205 15805 11245 15845
rect 11255 15805 11295 15845
rect 11305 15805 11345 15845
rect 11355 15805 11395 15845
rect 11405 15805 11445 15845
rect 11455 15805 11495 15845
rect 11505 15805 11545 15845
rect 11555 15805 11595 15845
rect 11605 15805 11645 15845
rect 11655 15805 11695 15845
rect 11705 15805 11745 15845
rect 11755 15805 11795 15845
rect 11805 15805 11845 15845
rect 11855 15805 11895 15845
rect 11905 15805 11945 15845
rect 11955 15805 11995 15845
rect 12005 15805 12045 15845
rect 12055 15805 12095 15845
rect 12105 15805 12145 15845
rect 12155 15805 12195 15845
rect 12205 15805 12245 15845
rect 12255 15805 12295 15845
rect 12305 15805 12345 15845
rect 12355 15805 12395 15845
rect 12405 15805 12445 15845
rect 12455 15805 12495 15845
rect 12505 15805 12545 15845
rect 12555 15805 12595 15845
rect 12605 15805 12645 15845
rect 12655 15805 12695 15845
rect 12705 15805 12745 15845
rect 12755 15805 12795 15845
rect 12805 15805 12845 15845
rect 12855 15805 12895 15845
rect 12905 15805 12945 15845
rect 12955 15805 12995 15845
rect 13005 15805 13045 15845
rect 13055 15805 13095 15845
rect 13105 15805 13145 15845
rect 13155 15805 13195 15845
rect 13205 15805 13245 15845
rect 13255 15805 13295 15845
rect 13305 15805 13345 15845
rect 13355 15805 13395 15845
rect 13405 15805 13445 15845
rect 13455 15805 13495 15845
rect 13505 15805 13545 15845
rect 13555 15805 13595 15845
rect 13605 15805 13645 15845
rect 13655 15805 13695 15845
rect 13705 15805 13745 15845
rect 13755 15805 13795 15845
rect 13805 15805 13845 15845
rect 13855 15805 13895 15845
rect 13905 15805 13945 15845
rect 13955 15805 13995 15845
rect 14005 15805 14045 15845
rect 14055 15805 14095 15845
rect 14105 15805 14145 15845
rect 14155 15805 14195 15845
rect 14205 15805 14245 15845
rect 14255 15805 14295 15845
rect 14305 15805 14345 15845
rect 14355 15805 14395 15845
rect 14405 15805 14445 15845
rect 14455 15805 14495 15845
rect 14505 15805 14545 15845
rect 14555 15805 14595 15845
rect 14605 15805 14645 15845
rect 14655 15805 14695 15845
rect 14705 15805 14745 15845
rect 14755 15805 14795 15845
rect 14805 15805 14845 15845
rect 14855 15805 14895 15845
rect 14905 15805 14945 15845
rect 14955 15805 14995 15845
rect 15005 15805 15045 15845
rect 15055 15805 15095 15845
rect 15105 15805 15145 15845
rect 15155 15805 15195 15845
rect 15205 15805 15245 15845
rect 15255 15805 15295 15845
rect 15305 15805 15345 15845
rect 15355 15805 15395 15845
rect 15405 15805 15445 15845
rect 15455 15805 15495 15845
rect 15505 15805 15545 15845
rect 15555 15805 15595 15845
rect 15605 15805 15645 15845
rect 15655 15805 15695 15845
rect 15705 15805 15745 15845
rect 15755 15805 15795 15845
rect 15805 15805 15845 15845
rect 15855 15805 15895 15845
rect 15905 15805 15945 15845
rect 15955 15805 15995 15845
rect 16005 15805 16045 15845
rect 16055 15805 16095 15845
rect 16105 15805 16145 15845
rect 16155 15805 16195 15845
rect 16205 15805 16245 15845
rect 16255 15805 16295 15845
rect 16305 15805 16345 15845
rect 16355 15805 16395 15845
rect 16405 15805 16445 15845
rect 16455 15805 16495 15845
rect 16505 15805 16545 15845
rect 16555 15805 16595 15845
rect 16605 15805 16645 15845
rect 16655 15805 16695 15845
rect 16705 15805 16745 15845
rect 16755 15805 16795 15845
rect 16805 15805 16845 15845
rect 16855 15805 16895 15845
rect 16905 15805 16945 15845
rect 16955 15805 16995 15845
rect 17005 15805 17045 15845
rect 17055 15805 17095 15845
rect 17105 15805 17145 15845
rect 17155 15805 17195 15845
rect 17205 15805 17245 15845
rect 17255 15805 17295 15845
rect 17305 15805 17345 15845
rect 17355 15805 17395 15845
rect 17405 15805 17445 15845
rect 17455 15805 17495 15845
rect 17505 15805 17545 15845
rect 17555 15805 17595 15845
rect 17605 15805 17645 15845
rect 17655 15805 17695 15845
rect 17705 15805 17745 15845
rect 17755 15805 17795 15845
rect 17805 15805 17845 15845
rect 17855 15805 17895 15845
rect 17905 15805 17945 15845
rect 17955 15805 17995 15845
rect 18005 15805 18045 15845
rect 18055 15805 18095 15845
rect 18105 15805 18145 15845
rect 18155 15805 18195 15845
rect 18205 15805 18245 15845
rect 18255 15805 18295 15845
rect 18305 15805 18345 15845
rect 18355 15805 18395 15845
rect 18405 15805 18445 15845
rect 18455 15805 18495 15845
rect 18505 15805 18545 15845
rect 18555 15805 18595 15845
rect 18605 15805 18645 15845
rect 18655 15805 18695 15845
rect 18705 15805 18745 15845
rect 18755 15805 18795 15845
rect 18805 15805 18845 15845
rect 18855 15805 18895 15845
rect 18905 15805 18945 15845
rect 18955 15805 18995 15845
rect 19005 15805 19045 15845
rect 19055 15805 19095 15845
rect 19105 15805 19145 15845
rect 19155 15805 19195 15845
rect 19205 15805 19245 15845
rect 19255 15805 19295 15845
rect 19305 15805 19345 15845
rect 19355 15805 19395 15845
rect 19405 15805 19445 15845
rect 19455 15805 19495 15845
rect 19505 15805 19545 15845
rect 19555 15805 19595 15845
rect 19605 15805 19645 15845
rect 19655 15805 19695 15845
rect 19705 15805 19745 15845
rect 19755 15805 19795 15845
rect 19805 15805 19845 15845
rect 19855 15805 19895 15845
rect 19905 15805 19945 15845
rect 19955 15805 19995 15845
rect 20005 15805 20045 15845
rect 20055 15805 20095 15845
rect 20105 15805 20145 15845
rect 20155 15805 20195 15845
rect 20205 15805 20245 15845
rect 20255 15805 20295 15845
rect 20305 15805 20345 15845
rect 20355 15805 20395 15845
rect 20405 15805 20445 15845
rect 20455 15805 20495 15845
rect 20505 15805 20545 15845
rect 20555 15805 20595 15845
rect 20605 15805 20645 15845
rect 20655 15805 20695 15845
rect 20705 15805 20745 15845
rect 20755 15805 20795 15845
rect 20805 15805 20845 15845
rect 20855 15805 20895 15845
rect 20905 15805 20945 15845
rect 20955 15805 20995 15845
rect 21005 15805 21045 15845
rect 21055 15805 21095 15845
rect 21105 15805 21145 15845
rect 21155 15805 21195 15845
rect 21205 15805 21245 15845
rect 21255 15805 21295 15845
rect 21305 15805 21345 15845
rect 21355 15805 21395 15845
rect 21405 15805 21445 15845
rect 21455 15805 21495 15845
rect 21505 15805 21545 15845
rect 21555 15805 21595 15845
rect 21605 15805 21645 15845
rect 21655 15805 21695 15845
rect 21705 15805 21745 15845
rect 21755 15805 21795 15845
rect 21805 15805 21845 15845
rect 21855 15805 21895 15845
rect 21905 15805 21945 15845
rect 21955 15805 21995 15845
rect 22005 15805 22045 15845
rect 22055 15805 22095 15845
rect 22105 15805 22145 15845
rect 22155 15805 22195 15845
rect 22205 15805 22245 15845
rect 22255 15805 22295 15845
rect 22305 15805 22345 15845
rect 22355 15805 22395 15845
rect 22405 15805 22445 15845
rect 22455 15805 22495 15845
rect 22505 15805 22545 15845
rect 22555 15805 22595 15845
rect 22605 15805 22645 15845
rect 22655 15805 22695 15845
rect 22705 15805 22745 15845
rect 22755 15805 22795 15845
rect 22805 15805 22845 15845
rect 22855 15805 22895 15845
rect 22905 15805 22945 15845
rect 22955 15805 22995 15845
rect 23005 15805 23045 15845
rect 23055 15805 23095 15845
rect 23105 15805 23145 15845
rect 23155 15805 23195 15845
rect 23205 15805 23245 15845
rect 23255 15805 23295 15845
rect 23305 15805 23345 15845
rect 23355 15805 23395 15845
rect 23405 15805 23445 15845
rect 23455 15805 23495 15845
rect 23505 15805 23545 15845
rect 23555 15805 23595 15845
rect 23605 15805 23645 15845
rect 23655 15805 23695 15845
rect 23705 15805 23745 15845
rect 23755 15805 23795 15845
rect 23805 15805 23845 15845
rect 23855 15805 23895 15845
rect 23905 15805 23945 15845
rect 23955 15805 23995 15845
rect 24005 15805 24045 15845
rect 24055 15805 24095 15845
rect 24105 15805 24145 15845
rect 24155 15805 24195 15845
rect 24205 15805 24245 15845
rect 24255 15805 24295 15845
rect 24305 15805 24345 15845
rect 24355 15805 24395 15845
rect 24405 15805 24445 15845
rect 24455 15805 24495 15845
rect 24505 15805 24545 15845
rect 24555 15805 24595 15845
rect 24605 15805 24645 15845
rect 24655 15805 24695 15845
rect 24705 15805 24745 15845
rect 24755 15805 24795 15845
rect 24805 15805 24845 15845
rect 24855 15805 24895 15845
rect 24905 15805 24945 15845
rect 24955 15805 24995 15845
rect 25005 15805 25045 15845
rect 25055 15805 25095 15845
rect 25105 15805 25145 15845
rect 25155 15805 25195 15845
rect 25205 15805 25245 15845
rect 25255 15805 25295 15845
rect 25305 15805 25345 15845
rect 25355 15805 25395 15845
rect 25405 15805 25445 15845
rect 25455 15805 25495 15845
rect 25505 15805 25545 15845
rect 25555 15805 25595 15845
rect 25605 15805 25645 15845
rect 25655 15805 25695 15845
rect 25705 15805 25745 15845
rect 25755 15805 25795 15845
rect 25805 15805 25845 15845
rect 25855 15805 25895 15845
rect 25905 15805 25945 15845
rect 25955 15805 25995 15845
rect 26005 15805 26045 15845
rect 26055 15805 26095 15845
rect 26105 15805 26145 15845
rect 26155 15805 26195 15845
rect 26205 15805 26245 15845
rect 26255 15805 26295 15845
rect 26305 15805 26345 15845
rect 26355 15805 26395 15845
rect 26405 15805 26445 15845
rect 26455 15805 26495 15845
rect 26505 15805 26545 15845
rect 26555 15805 26595 15845
rect 26605 15805 26645 15845
rect 26655 15805 26695 15845
rect 26705 15805 26745 15845
rect 26755 15805 26795 15845
rect 26805 15805 26845 15845
rect 26855 15805 26895 15845
rect 26905 15805 26945 15845
rect 26955 15805 26995 15845
rect 27005 15805 27045 15845
rect 27055 15805 27095 15845
rect 27105 15805 27145 15845
rect 27155 15805 27195 15845
rect 27205 15805 27245 15845
rect 27255 15805 27295 15845
rect 27305 15805 27345 15845
rect 27355 15805 27395 15845
rect 27405 15805 27445 15845
rect 27455 15805 27495 15845
rect 27505 15805 27545 15845
rect 27555 15805 27595 15845
rect 27605 15805 27645 15845
rect 27655 15805 27695 15845
rect 27705 15805 27745 15845
rect 27755 15805 27795 15845
rect 27805 15805 27845 15845
rect 27855 15805 27895 15845
rect 27905 15805 27945 15845
rect 27955 15805 27995 15845
rect 28005 15805 28045 15845
rect 28055 15805 28095 15845
rect 28105 15805 28145 15845
rect 28155 15805 28195 15845
rect 28205 15805 28245 15845
rect 28255 15805 28295 15845
rect 28305 15805 28345 15845
rect 28355 15805 28395 15845
rect 28405 15805 28445 15845
rect 28455 15805 28495 15845
rect 28505 15805 28545 15845
rect 28555 15805 28595 15845
rect 28605 15805 28645 15845
rect 28655 15805 28695 15845
rect 28705 15805 28745 15845
rect 28755 15805 28795 15845
rect 28805 15805 28845 15845
rect 28855 15805 28895 15845
rect 28905 15805 28945 15845
rect 28955 15805 28995 15845
rect 29005 15805 29045 15845
rect 29055 15805 29095 15845
rect 29105 15805 29145 15845
rect 29155 15805 29195 15845
rect 29205 15805 29245 15845
rect 29255 15805 29295 15845
rect 29305 15805 29345 15845
rect 29355 15805 29395 15845
rect 29405 15805 29445 15845
rect 29455 15805 29495 15845
rect 29505 15805 29545 15845
rect 29555 15805 29595 15845
rect 29605 15805 29645 15845
rect 29655 15805 29695 15845
rect 29705 15805 29745 15845
rect 29755 15805 29795 15845
rect 29805 15805 29845 15845
rect 29855 15805 29895 15845
rect 29905 15805 29945 15845
rect 29955 15805 29995 15845
rect 30005 15805 30045 15845
rect 30055 15805 30095 15845
rect 30105 15805 30145 15845
rect 30155 15805 30195 15845
rect 30205 15805 30245 15845
rect 30255 15805 30295 15845
rect 30305 15805 30345 15845
rect 30355 15805 30395 15845
rect 30405 15805 30445 15845
rect 30455 15805 30495 15845
rect 30505 15805 30545 15845
rect 30555 15805 30595 15845
rect 30605 15805 30645 15845
rect 30655 15805 30695 15845
rect 30705 15805 30745 15845
rect 30755 15805 30795 15845
rect 30805 15805 30845 15845
rect 30855 15805 30895 15845
rect 30905 15805 30945 15845
rect 30955 15805 30995 15845
rect 31005 15805 31045 15845
rect 31055 15805 31095 15845
rect 31105 15805 31145 15845
rect 31155 15805 31195 15845
rect 31205 15805 31245 15845
rect 31255 15805 31295 15845
rect 31305 15805 31345 15845
rect 31355 15805 31395 15845
rect 31405 15805 31445 15845
rect 31455 15805 31495 15845
rect 31505 15805 31545 15845
rect 31555 15805 31595 15845
rect 31605 15805 31645 15845
rect 31655 15805 31695 15845
rect 31705 15805 31745 15845
rect 31755 15805 31795 15845
rect 31805 15805 31845 15845
rect 31855 15805 31895 15845
rect 31905 15805 31945 15845
rect 31955 15805 31995 15845
rect 32005 15805 32045 15845
rect 32055 15805 32095 15845
rect 32105 15805 32145 15845
rect 32155 15805 32195 15845
rect 32205 15805 32245 15845
rect 32255 15805 32295 15845
rect 32305 15805 32345 15845
rect 32355 15805 32395 15845
rect 32405 15805 32445 15845
rect 32455 15805 32495 15845
rect 32505 15805 32545 15845
rect 32555 15805 32595 15845
rect 32605 15805 32645 15845
rect 32655 15805 32695 15845
rect 32705 15805 32745 15845
rect 32755 15805 32795 15845
rect 32805 15805 32845 15845
rect 32855 15805 32895 15845
rect 32905 15805 32945 15845
rect 32955 15805 32995 15845
rect 33005 15805 33045 15845
rect 33055 15805 33095 15845
rect 33105 15805 33145 15845
rect 33155 15805 33195 15845
rect 33205 15805 33245 15845
rect 33255 15805 33295 15845
rect 33305 15805 33345 15845
rect 33355 15805 33395 15845
rect 33405 15805 33445 15845
rect 33455 15805 33495 15845
rect 33505 15805 33545 15845
rect 33555 15805 33595 15845
rect 33605 15805 33645 15845
rect 33655 15805 33695 15845
rect 33705 15805 33745 15845
rect 33755 15805 33795 15845
rect 33805 15805 33845 15845
rect 33855 15805 33895 15845
rect 33905 15805 33945 15845
rect 33955 15805 33995 15845
rect 34005 15805 34045 15845
rect 34055 15805 34095 15845
rect 34105 15805 34145 15845
rect 34155 15805 34195 15845
rect 34205 15805 34245 15845
rect 34255 15805 34295 15845
rect 34305 15805 34345 15845
rect 34355 15805 34395 15845
rect 34405 15805 34445 15845
rect 34455 15805 34495 15845
rect 34505 15805 34545 15845
rect 34555 15805 34595 15845
rect 34605 15805 34645 15845
rect 34655 15805 34695 15845
rect 34705 15805 34745 15845
rect 34755 15805 34795 15845
rect 34805 15805 34845 15845
rect 34855 15805 34895 15845
rect 34905 15805 34945 15845
rect 34955 15805 34995 15845
rect 35005 15805 35045 15845
rect 35055 15805 35095 15845
rect 35105 15805 35145 15845
rect 35155 15805 35195 15845
rect 35205 15805 35245 15845
rect 35255 15805 35295 15845
rect 35305 15805 35345 15845
rect 35355 15805 35395 15845
rect 35405 15805 35445 15845
rect 35455 15805 35495 15845
rect 35505 15805 35545 15845
rect 35555 15805 35595 15845
rect 35605 15805 35645 15845
rect 35655 15805 35695 15845
rect 35705 15805 35745 15845
rect 35755 15805 35795 15845
rect 35805 15805 35845 15845
rect 35855 15805 35895 15845
rect 35905 15805 35945 15845
rect 35955 15805 35995 15845
rect 36005 15805 36045 15845
rect 36055 15805 36095 15845
rect 36105 15805 36145 15845
rect 36155 15805 36195 15845
rect 36205 15805 36245 15845
rect 36255 15805 36295 15845
rect 36305 15805 36345 15845
rect 36355 15805 36395 15845
rect 36405 15805 36445 15845
rect 36455 15805 36495 15845
rect 36505 15805 36545 15845
rect 36555 15805 36595 15845
rect 36605 15805 36645 15845
rect 36655 15805 36695 15845
rect 36705 15805 36745 15845
rect 36755 15805 36795 15845
rect 36805 15805 36845 15845
rect 36855 15805 36895 15845
rect 36905 15805 36945 15845
rect 36955 15805 36995 15845
rect 37005 15805 37045 15845
rect 37055 15805 37095 15845
rect 37105 15805 37145 15845
rect 37155 15805 37195 15845
rect 37205 15805 37245 15845
rect 37255 15805 37295 15845
rect 37305 15805 37345 15845
rect 37355 15805 37395 15845
rect 37405 15805 37445 15845
rect 37455 15805 37495 15845
rect 37505 15805 37545 15845
rect 37555 15805 37595 15845
rect 37605 15805 37645 15845
rect 37655 15805 37695 15845
rect 37705 15805 37745 15845
rect 37755 15805 37795 15845
rect 37805 15805 37845 15845
rect 37855 15805 37895 15845
rect 37905 15805 37945 15845
rect 37955 15805 37995 15845
rect 38005 15805 38045 15845
rect 38055 15805 38095 15845
rect 38105 15805 38145 15845
rect 38155 15805 38195 15845
rect 38205 15805 38245 15845
rect 38255 15805 38295 15845
rect 38305 15805 38345 15845
rect 38355 15805 38395 15845
rect 38405 15805 38445 15845
rect 38455 15805 38495 15845
rect 38505 15805 38545 15845
rect 38555 15805 38595 15845
rect 38605 15805 38645 15845
rect 38655 15805 38695 15845
rect 38705 15805 38745 15845
rect 38755 15805 38795 15845
rect 38805 15805 38845 15845
rect 38855 15805 38895 15845
rect 38905 15805 38945 15845
rect 38955 15805 38995 15845
rect 39005 15805 39045 15845
rect 39055 15805 39095 15845
rect 39105 15805 39145 15845
rect 39155 15805 39195 15845
rect 39205 15805 39245 15845
rect 39255 15805 39295 15845
rect 39305 15805 39345 15845
rect 39355 15805 39395 15845
rect 39405 15805 39445 15845
rect 39455 15805 39495 15845
rect 39505 15805 39545 15845
rect 39555 15805 39595 15845
rect 39605 15805 39645 15845
rect 39655 15805 39695 15845
rect 39705 15805 39745 15845
rect -3495 15740 -3455 15745
rect -3495 15710 -3490 15740
rect -3490 15710 -3460 15740
rect -3460 15710 -3455 15740
rect -3495 15705 -3455 15710
rect -3295 15740 -3255 15745
rect -3295 15710 -3290 15740
rect -3290 15710 -3260 15740
rect -3260 15710 -3255 15740
rect -3295 15705 -3255 15710
rect -3095 15740 -3055 15745
rect -3095 15710 -3090 15740
rect -3090 15710 -3060 15740
rect -3060 15710 -3055 15740
rect -3095 15705 -3055 15710
rect -1595 15740 -1555 15745
rect -1595 15710 -1590 15740
rect -1590 15710 -1560 15740
rect -1560 15710 -1555 15740
rect -1595 15705 -1555 15710
rect -1195 15740 -1155 15745
rect -1195 15710 -1190 15740
rect -1190 15710 -1160 15740
rect -1160 15710 -1155 15740
rect -1195 15705 -1155 15710
rect -1095 15740 -1055 15745
rect -1095 15710 -1090 15740
rect -1090 15710 -1060 15740
rect -1060 15710 -1055 15740
rect -1095 15705 -1055 15710
rect -995 15740 -955 15745
rect -995 15710 -990 15740
rect -990 15710 -960 15740
rect -960 15710 -955 15740
rect -995 15705 -955 15710
rect -895 15740 -855 15745
rect -895 15710 -890 15740
rect -890 15710 -860 15740
rect -860 15710 -855 15740
rect -895 15705 -855 15710
rect -695 15740 -655 15745
rect -695 15710 -690 15740
rect -690 15710 -660 15740
rect -660 15710 -655 15740
rect -695 15705 -655 15710
rect -595 15740 -555 15745
rect -595 15710 -590 15740
rect -590 15710 -560 15740
rect -560 15710 -555 15740
rect -595 15705 -555 15710
rect -495 15740 -455 15745
rect -495 15710 -490 15740
rect -490 15710 -460 15740
rect -460 15710 -455 15740
rect -495 15705 -455 15710
rect -295 15740 -255 15745
rect -295 15710 -290 15740
rect -290 15710 -260 15740
rect -260 15710 -255 15740
rect -295 15705 -255 15710
rect -195 15740 -155 15745
rect -195 15710 -190 15740
rect -190 15710 -160 15740
rect -160 15710 -155 15740
rect -195 15705 -155 15710
rect -95 15740 -55 15745
rect -95 15710 -90 15740
rect -90 15710 -60 15740
rect -60 15710 -55 15740
rect -95 15705 -55 15710
rect 5 15705 45 15745
rect 55 15705 95 15745
rect 105 15705 145 15745
rect 155 15705 195 15745
rect 205 15705 245 15745
rect 255 15705 295 15745
rect 305 15705 345 15745
rect 355 15705 395 15745
rect 405 15705 445 15745
rect 455 15705 495 15745
rect 505 15705 545 15745
rect 555 15705 595 15745
rect 605 15705 645 15745
rect 655 15705 695 15745
rect 705 15705 745 15745
rect 755 15705 795 15745
rect 805 15705 845 15745
rect 855 15705 895 15745
rect 905 15705 945 15745
rect 955 15705 995 15745
rect 1005 15705 1045 15745
rect 1055 15705 1095 15745
rect 1105 15705 1145 15745
rect 1155 15705 1195 15745
rect 1205 15705 1245 15745
rect 1255 15705 1295 15745
rect 1305 15705 1345 15745
rect 1355 15705 1395 15745
rect 1405 15705 1445 15745
rect 1455 15705 1495 15745
rect 1505 15705 1545 15745
rect 1555 15705 1595 15745
rect 1605 15705 1645 15745
rect 1655 15705 1695 15745
rect 1705 15705 1745 15745
rect 1755 15705 1795 15745
rect 1805 15705 1845 15745
rect 1855 15705 1895 15745
rect 1905 15705 1945 15745
rect 1955 15705 1995 15745
rect 2005 15705 2045 15745
rect 2055 15705 2095 15745
rect 2105 15705 2145 15745
rect 2155 15705 2195 15745
rect 2205 15705 2245 15745
rect 2255 15705 2295 15745
rect 2305 15705 2345 15745
rect 2355 15705 2395 15745
rect 2405 15705 2445 15745
rect 2455 15705 2495 15745
rect 2505 15705 2545 15745
rect 2555 15705 2595 15745
rect 2605 15705 2645 15745
rect 2655 15705 2695 15745
rect 2705 15705 2745 15745
rect 2755 15705 2795 15745
rect 2805 15705 2845 15745
rect 2855 15705 2895 15745
rect 2905 15705 2945 15745
rect 2955 15705 2995 15745
rect 3005 15705 3045 15745
rect 3055 15705 3095 15745
rect 3105 15705 3145 15745
rect 3155 15705 3195 15745
rect 3205 15705 3245 15745
rect 3255 15705 3295 15745
rect 3305 15705 3345 15745
rect 3355 15705 3395 15745
rect 3405 15705 3445 15745
rect 3455 15705 3495 15745
rect 3505 15705 3545 15745
rect 3555 15705 3595 15745
rect 3605 15705 3645 15745
rect 3655 15705 3695 15745
rect 3705 15705 3745 15745
rect 3755 15705 3795 15745
rect 3805 15705 3845 15745
rect 3855 15705 3895 15745
rect 3905 15705 3945 15745
rect 3955 15705 3995 15745
rect 4005 15705 4045 15745
rect 4055 15705 4095 15745
rect 4105 15705 4145 15745
rect 4155 15705 4195 15745
rect 4205 15705 4245 15745
rect 4255 15705 4295 15745
rect 4305 15705 4345 15745
rect 4355 15705 4395 15745
rect 4405 15705 4445 15745
rect 4455 15705 4495 15745
rect 4505 15705 4545 15745
rect 4555 15705 4595 15745
rect 4605 15705 4645 15745
rect 4655 15705 4695 15745
rect 4705 15705 4745 15745
rect 4755 15705 4795 15745
rect 4805 15705 4845 15745
rect 4855 15705 4895 15745
rect 4905 15705 4945 15745
rect 4955 15705 4995 15745
rect 5005 15705 5045 15745
rect 5055 15705 5095 15745
rect 5105 15705 5145 15745
rect 5155 15705 5195 15745
rect 5205 15705 5245 15745
rect 5255 15705 5295 15745
rect 5305 15705 5345 15745
rect 5355 15705 5395 15745
rect 5405 15705 5445 15745
rect 5455 15705 5495 15745
rect 5505 15705 5545 15745
rect 5555 15705 5595 15745
rect 5605 15705 5645 15745
rect 5655 15705 5695 15745
rect 5705 15705 5745 15745
rect 5755 15705 5795 15745
rect 5805 15705 5845 15745
rect 5855 15705 5895 15745
rect 5905 15705 5945 15745
rect 5955 15705 5995 15745
rect 6005 15705 6045 15745
rect 6055 15705 6095 15745
rect 6105 15705 6145 15745
rect 6155 15705 6195 15745
rect 6205 15705 6245 15745
rect 6255 15705 6295 15745
rect 6305 15705 6345 15745
rect 6355 15705 6395 15745
rect 6405 15705 6445 15745
rect 6455 15705 6495 15745
rect 6505 15705 6545 15745
rect 6555 15705 6595 15745
rect 6605 15705 6645 15745
rect 6655 15705 6695 15745
rect 6705 15705 6745 15745
rect 6755 15705 6795 15745
rect 6805 15705 6845 15745
rect 6855 15705 6895 15745
rect 6905 15705 6945 15745
rect 6955 15705 6995 15745
rect 7005 15705 7045 15745
rect 7055 15705 7095 15745
rect 7105 15705 7145 15745
rect 7155 15705 7195 15745
rect 7205 15705 7245 15745
rect 7255 15705 7295 15745
rect 7305 15705 7345 15745
rect 7355 15705 7395 15745
rect 7405 15705 7445 15745
rect 7455 15705 7495 15745
rect 7505 15705 7545 15745
rect 7555 15705 7595 15745
rect 7605 15705 7645 15745
rect 7655 15705 7695 15745
rect 7705 15705 7745 15745
rect 7755 15705 7795 15745
rect 7805 15705 7845 15745
rect 7855 15705 7895 15745
rect 7905 15705 7945 15745
rect 7955 15705 7995 15745
rect 8005 15705 8045 15745
rect 8055 15705 8095 15745
rect 8105 15705 8145 15745
rect 8155 15705 8195 15745
rect 8205 15705 8245 15745
rect 8255 15705 8295 15745
rect 8305 15705 8345 15745
rect 8355 15705 8395 15745
rect 8405 15705 8445 15745
rect 8455 15705 8495 15745
rect 8505 15705 8545 15745
rect 8555 15705 8595 15745
rect 8605 15705 8645 15745
rect 8655 15705 8695 15745
rect 8705 15705 8745 15745
rect 8755 15705 8795 15745
rect 8805 15705 8845 15745
rect 8855 15705 8895 15745
rect 8905 15705 8945 15745
rect 8955 15705 8995 15745
rect 9005 15705 9045 15745
rect 9055 15705 9095 15745
rect 9105 15705 9145 15745
rect 9155 15705 9195 15745
rect 9205 15705 9245 15745
rect 9255 15705 9295 15745
rect 9305 15705 9345 15745
rect 9355 15705 9395 15745
rect 9405 15705 9445 15745
rect 9455 15705 9495 15745
rect 9505 15705 9545 15745
rect 9555 15705 9595 15745
rect 9605 15705 9645 15745
rect 9655 15705 9695 15745
rect 9705 15705 9745 15745
rect 9755 15705 9795 15745
rect 9805 15705 9845 15745
rect 9855 15705 9895 15745
rect 9905 15705 9945 15745
rect 9955 15705 9995 15745
rect 10005 15705 10045 15745
rect 10055 15705 10095 15745
rect 10105 15705 10145 15745
rect 10155 15705 10195 15745
rect 10205 15705 10245 15745
rect 10255 15705 10295 15745
rect 10305 15705 10345 15745
rect 10355 15705 10395 15745
rect 10405 15705 10445 15745
rect 10455 15705 10495 15745
rect 10505 15705 10545 15745
rect 10555 15705 10595 15745
rect 10605 15705 10645 15745
rect 10655 15705 10695 15745
rect 10705 15705 10745 15745
rect 10755 15705 10795 15745
rect 10805 15705 10845 15745
rect 10855 15705 10895 15745
rect 10905 15705 10945 15745
rect 10955 15705 10995 15745
rect 11005 15705 11045 15745
rect 11055 15705 11095 15745
rect 11105 15705 11145 15745
rect 11155 15705 11195 15745
rect 11205 15705 11245 15745
rect 11255 15705 11295 15745
rect 11305 15705 11345 15745
rect 11355 15705 11395 15745
rect 11405 15705 11445 15745
rect 11455 15705 11495 15745
rect 11505 15705 11545 15745
rect 11555 15705 11595 15745
rect 11605 15705 11645 15745
rect 11655 15705 11695 15745
rect 11705 15705 11745 15745
rect 11755 15705 11795 15745
rect 11805 15705 11845 15745
rect 11855 15705 11895 15745
rect 11905 15705 11945 15745
rect 11955 15705 11995 15745
rect 12005 15705 12045 15745
rect 12055 15705 12095 15745
rect 12105 15705 12145 15745
rect 12155 15705 12195 15745
rect 12205 15705 12245 15745
rect 12255 15705 12295 15745
rect 12305 15705 12345 15745
rect 12355 15705 12395 15745
rect 12405 15705 12445 15745
rect 12455 15705 12495 15745
rect 12505 15705 12545 15745
rect 12555 15705 12595 15745
rect 12605 15705 12645 15745
rect 12655 15705 12695 15745
rect 12705 15705 12745 15745
rect 12755 15705 12795 15745
rect 12805 15705 12845 15745
rect 12855 15705 12895 15745
rect 12905 15705 12945 15745
rect 12955 15705 12995 15745
rect 13005 15705 13045 15745
rect 13055 15705 13095 15745
rect 13105 15705 13145 15745
rect 13155 15705 13195 15745
rect 13205 15705 13245 15745
rect 13255 15705 13295 15745
rect 13305 15705 13345 15745
rect 13355 15705 13395 15745
rect 13405 15705 13445 15745
rect 13455 15705 13495 15745
rect 13505 15705 13545 15745
rect 13555 15705 13595 15745
rect 13605 15705 13645 15745
rect 13655 15705 13695 15745
rect 13705 15705 13745 15745
rect 13755 15705 13795 15745
rect 13805 15705 13845 15745
rect 13855 15705 13895 15745
rect 13905 15705 13945 15745
rect 13955 15705 13995 15745
rect 14005 15705 14045 15745
rect 14055 15705 14095 15745
rect 14105 15705 14145 15745
rect 14155 15705 14195 15745
rect 14205 15705 14245 15745
rect 14255 15705 14295 15745
rect 14305 15705 14345 15745
rect 14355 15705 14395 15745
rect 14405 15705 14445 15745
rect 14455 15705 14495 15745
rect 14505 15705 14545 15745
rect 14555 15705 14595 15745
rect 14605 15705 14645 15745
rect 14655 15705 14695 15745
rect 14705 15705 14745 15745
rect 14755 15705 14795 15745
rect 14805 15705 14845 15745
rect 14855 15705 14895 15745
rect 14905 15705 14945 15745
rect 14955 15705 14995 15745
rect 15005 15705 15045 15745
rect 15055 15705 15095 15745
rect 15105 15705 15145 15745
rect 15155 15705 15195 15745
rect 15205 15705 15245 15745
rect 15255 15705 15295 15745
rect 15305 15705 15345 15745
rect 15355 15705 15395 15745
rect 15405 15705 15445 15745
rect 15455 15705 15495 15745
rect 15505 15705 15545 15745
rect 15555 15705 15595 15745
rect 15605 15705 15645 15745
rect 15655 15705 15695 15745
rect 15705 15705 15745 15745
rect 15755 15705 15795 15745
rect 15805 15705 15845 15745
rect 15855 15705 15895 15745
rect 15905 15705 15945 15745
rect 15955 15705 15995 15745
rect 16005 15705 16045 15745
rect 16055 15705 16095 15745
rect 16105 15705 16145 15745
rect 16155 15705 16195 15745
rect 16205 15705 16245 15745
rect 16255 15705 16295 15745
rect 16305 15705 16345 15745
rect 16355 15705 16395 15745
rect 16405 15705 16445 15745
rect 16455 15705 16495 15745
rect 16505 15705 16545 15745
rect 16555 15705 16595 15745
rect 16605 15705 16645 15745
rect 16655 15705 16695 15745
rect 16705 15705 16745 15745
rect 16755 15705 16795 15745
rect 16805 15705 16845 15745
rect 16855 15705 16895 15745
rect 16905 15705 16945 15745
rect 16955 15705 16995 15745
rect 17005 15705 17045 15745
rect 17055 15705 17095 15745
rect 17105 15705 17145 15745
rect 17155 15705 17195 15745
rect 17205 15705 17245 15745
rect 17255 15705 17295 15745
rect 17305 15705 17345 15745
rect 17355 15705 17395 15745
rect 17405 15705 17445 15745
rect 17455 15705 17495 15745
rect 17505 15705 17545 15745
rect 17555 15705 17595 15745
rect 17605 15705 17645 15745
rect 17655 15705 17695 15745
rect 17705 15705 17745 15745
rect 17755 15705 17795 15745
rect 17805 15705 17845 15745
rect 17855 15705 17895 15745
rect 17905 15705 17945 15745
rect 17955 15705 17995 15745
rect 18005 15705 18045 15745
rect 18055 15705 18095 15745
rect 18105 15705 18145 15745
rect 18155 15705 18195 15745
rect 18205 15705 18245 15745
rect 18255 15705 18295 15745
rect 18305 15705 18345 15745
rect 18355 15705 18395 15745
rect 18405 15705 18445 15745
rect 18455 15705 18495 15745
rect 18505 15705 18545 15745
rect 18555 15705 18595 15745
rect 18605 15705 18645 15745
rect 18655 15705 18695 15745
rect 18705 15705 18745 15745
rect 18755 15705 18795 15745
rect 18805 15705 18845 15745
rect 18855 15705 18895 15745
rect 18905 15705 18945 15745
rect 18955 15705 18995 15745
rect 19005 15705 19045 15745
rect 19055 15705 19095 15745
rect 19105 15705 19145 15745
rect 19155 15705 19195 15745
rect 19205 15705 19245 15745
rect 19255 15705 19295 15745
rect 19305 15705 19345 15745
rect 19355 15705 19395 15745
rect 19405 15705 19445 15745
rect 19455 15705 19495 15745
rect 19505 15705 19545 15745
rect 19555 15705 19595 15745
rect 19605 15705 19645 15745
rect 19655 15705 19695 15745
rect 19705 15705 19745 15745
rect 19755 15705 19795 15745
rect 19805 15705 19845 15745
rect 19855 15705 19895 15745
rect 19905 15705 19945 15745
rect 19955 15705 19995 15745
rect 20005 15705 20045 15745
rect 20055 15705 20095 15745
rect 20105 15705 20145 15745
rect 20155 15705 20195 15745
rect 20205 15705 20245 15745
rect 20255 15705 20295 15745
rect 20305 15705 20345 15745
rect 20355 15705 20395 15745
rect 20405 15705 20445 15745
rect 20455 15705 20495 15745
rect 20505 15705 20545 15745
rect 20555 15705 20595 15745
rect 20605 15705 20645 15745
rect 20655 15705 20695 15745
rect 20705 15705 20745 15745
rect 20755 15705 20795 15745
rect 20805 15705 20845 15745
rect 20855 15705 20895 15745
rect 20905 15705 20945 15745
rect 20955 15705 20995 15745
rect 21005 15705 21045 15745
rect 21055 15705 21095 15745
rect 21105 15705 21145 15745
rect 21155 15705 21195 15745
rect 21205 15705 21245 15745
rect 21255 15705 21295 15745
rect 21305 15705 21345 15745
rect 21355 15705 21395 15745
rect 21405 15705 21445 15745
rect 21455 15705 21495 15745
rect 21505 15705 21545 15745
rect 21555 15705 21595 15745
rect 21605 15705 21645 15745
rect 21655 15705 21695 15745
rect 21705 15705 21745 15745
rect 21755 15705 21795 15745
rect 21805 15705 21845 15745
rect 21855 15705 21895 15745
rect 21905 15705 21945 15745
rect 21955 15705 21995 15745
rect 22005 15705 22045 15745
rect 22055 15705 22095 15745
rect 22105 15705 22145 15745
rect 22155 15705 22195 15745
rect 22205 15705 22245 15745
rect 22255 15705 22295 15745
rect 22305 15705 22345 15745
rect 22355 15705 22395 15745
rect 22405 15705 22445 15745
rect 22455 15705 22495 15745
rect 22505 15705 22545 15745
rect 22555 15705 22595 15745
rect 22605 15705 22645 15745
rect 22655 15705 22695 15745
rect 22705 15705 22745 15745
rect 22755 15705 22795 15745
rect 22805 15705 22845 15745
rect 22855 15705 22895 15745
rect 22905 15705 22945 15745
rect 22955 15705 22995 15745
rect 23005 15705 23045 15745
rect 23055 15705 23095 15745
rect 23105 15705 23145 15745
rect 23155 15705 23195 15745
rect 23205 15705 23245 15745
rect 23255 15705 23295 15745
rect 23305 15705 23345 15745
rect 23355 15705 23395 15745
rect 23405 15705 23445 15745
rect 23455 15705 23495 15745
rect 23505 15705 23545 15745
rect 23555 15705 23595 15745
rect 23605 15705 23645 15745
rect 23655 15705 23695 15745
rect 23705 15705 23745 15745
rect 23755 15705 23795 15745
rect 23805 15705 23845 15745
rect 23855 15705 23895 15745
rect 23905 15705 23945 15745
rect 23955 15705 23995 15745
rect 24005 15705 24045 15745
rect 24055 15705 24095 15745
rect 24105 15705 24145 15745
rect 24155 15705 24195 15745
rect 24205 15705 24245 15745
rect 24255 15705 24295 15745
rect 24305 15705 24345 15745
rect 24355 15705 24395 15745
rect 24405 15705 24445 15745
rect 24455 15705 24495 15745
rect 24505 15705 24545 15745
rect 24555 15705 24595 15745
rect 24605 15705 24645 15745
rect 24655 15705 24695 15745
rect 24705 15705 24745 15745
rect 24755 15705 24795 15745
rect 24805 15705 24845 15745
rect 24855 15705 24895 15745
rect 24905 15705 24945 15745
rect 24955 15705 24995 15745
rect 25005 15705 25045 15745
rect 25055 15705 25095 15745
rect 25105 15705 25145 15745
rect 25155 15705 25195 15745
rect 25205 15705 25245 15745
rect 25255 15705 25295 15745
rect 25305 15705 25345 15745
rect 25355 15705 25395 15745
rect 25405 15705 25445 15745
rect 25455 15705 25495 15745
rect 25505 15705 25545 15745
rect 25555 15705 25595 15745
rect 25605 15705 25645 15745
rect 25655 15705 25695 15745
rect 25705 15705 25745 15745
rect 25755 15705 25795 15745
rect 25805 15705 25845 15745
rect 25855 15705 25895 15745
rect 25905 15705 25945 15745
rect 25955 15705 25995 15745
rect 26005 15705 26045 15745
rect 26055 15705 26095 15745
rect 26105 15705 26145 15745
rect 26155 15705 26195 15745
rect 26205 15705 26245 15745
rect 26255 15705 26295 15745
rect 26305 15705 26345 15745
rect 26355 15705 26395 15745
rect 26405 15705 26445 15745
rect 26455 15705 26495 15745
rect 26505 15705 26545 15745
rect 26555 15705 26595 15745
rect 26605 15705 26645 15745
rect 26655 15705 26695 15745
rect 26705 15705 26745 15745
rect 26755 15705 26795 15745
rect 26805 15705 26845 15745
rect 26855 15705 26895 15745
rect 26905 15705 26945 15745
rect 26955 15705 26995 15745
rect 27005 15705 27045 15745
rect 27055 15705 27095 15745
rect 27105 15705 27145 15745
rect 27155 15705 27195 15745
rect 27205 15705 27245 15745
rect 27255 15705 27295 15745
rect 27305 15705 27345 15745
rect 27355 15705 27395 15745
rect 27405 15705 27445 15745
rect 27455 15705 27495 15745
rect 27505 15705 27545 15745
rect 27555 15705 27595 15745
rect 27605 15705 27645 15745
rect 27655 15705 27695 15745
rect 27705 15705 27745 15745
rect 27755 15705 27795 15745
rect 27805 15705 27845 15745
rect 27855 15705 27895 15745
rect 27905 15705 27945 15745
rect 27955 15705 27995 15745
rect 28005 15705 28045 15745
rect 28055 15705 28095 15745
rect 28105 15705 28145 15745
rect 28155 15705 28195 15745
rect 28205 15705 28245 15745
rect 28255 15705 28295 15745
rect 28305 15705 28345 15745
rect 28355 15705 28395 15745
rect 28405 15705 28445 15745
rect 28455 15705 28495 15745
rect 28505 15705 28545 15745
rect 28555 15705 28595 15745
rect 28605 15705 28645 15745
rect 28655 15705 28695 15745
rect 28705 15705 28745 15745
rect 28755 15705 28795 15745
rect 28805 15705 28845 15745
rect 28855 15705 28895 15745
rect 28905 15705 28945 15745
rect 28955 15705 28995 15745
rect 29005 15705 29045 15745
rect 29055 15705 29095 15745
rect 29105 15705 29145 15745
rect 29155 15705 29195 15745
rect 29205 15705 29245 15745
rect 29255 15705 29295 15745
rect 29305 15705 29345 15745
rect 29355 15705 29395 15745
rect 29405 15705 29445 15745
rect 29455 15705 29495 15745
rect 29505 15705 29545 15745
rect 29555 15705 29595 15745
rect 29605 15705 29645 15745
rect 29655 15705 29695 15745
rect 29705 15705 29745 15745
rect 29755 15705 29795 15745
rect 29805 15705 29845 15745
rect 29855 15705 29895 15745
rect 29905 15705 29945 15745
rect 29955 15705 29995 15745
rect 30005 15705 30045 15745
rect 30055 15705 30095 15745
rect 30105 15705 30145 15745
rect 30155 15705 30195 15745
rect 30205 15705 30245 15745
rect 30255 15705 30295 15745
rect 30305 15705 30345 15745
rect 30355 15705 30395 15745
rect 30405 15705 30445 15745
rect 30455 15705 30495 15745
rect 30505 15705 30545 15745
rect 30555 15705 30595 15745
rect 30605 15705 30645 15745
rect 30655 15705 30695 15745
rect 30705 15705 30745 15745
rect 30755 15705 30795 15745
rect 30805 15705 30845 15745
rect 30855 15705 30895 15745
rect 30905 15705 30945 15745
rect 30955 15705 30995 15745
rect 31005 15705 31045 15745
rect 31055 15705 31095 15745
rect 31105 15705 31145 15745
rect 31155 15705 31195 15745
rect 31205 15705 31245 15745
rect 31255 15705 31295 15745
rect 31305 15705 31345 15745
rect 31355 15705 31395 15745
rect 31405 15705 31445 15745
rect 31455 15705 31495 15745
rect 31505 15705 31545 15745
rect 31555 15705 31595 15745
rect 31605 15705 31645 15745
rect 31655 15705 31695 15745
rect 31705 15705 31745 15745
rect 31755 15705 31795 15745
rect 31805 15705 31845 15745
rect 31855 15705 31895 15745
rect 31905 15705 31945 15745
rect 31955 15705 31995 15745
rect 32005 15705 32045 15745
rect 32055 15705 32095 15745
rect 32105 15705 32145 15745
rect 32155 15705 32195 15745
rect 32205 15705 32245 15745
rect 32255 15705 32295 15745
rect 32305 15705 32345 15745
rect 32355 15705 32395 15745
rect 32405 15705 32445 15745
rect 32455 15705 32495 15745
rect 32505 15705 32545 15745
rect 32555 15705 32595 15745
rect 32605 15705 32645 15745
rect 32655 15705 32695 15745
rect 32705 15705 32745 15745
rect 32755 15705 32795 15745
rect 32805 15705 32845 15745
rect 32855 15705 32895 15745
rect 32905 15705 32945 15745
rect 32955 15705 32995 15745
rect 33005 15705 33045 15745
rect 33055 15705 33095 15745
rect 33105 15705 33145 15745
rect 33155 15705 33195 15745
rect 33205 15705 33245 15745
rect 33255 15705 33295 15745
rect 33305 15705 33345 15745
rect 33355 15705 33395 15745
rect 33405 15705 33445 15745
rect 33455 15705 33495 15745
rect 33505 15705 33545 15745
rect 33555 15705 33595 15745
rect 33605 15705 33645 15745
rect 33655 15705 33695 15745
rect 33705 15705 33745 15745
rect 33755 15705 33795 15745
rect 33805 15705 33845 15745
rect 33855 15705 33895 15745
rect 33905 15705 33945 15745
rect 33955 15705 33995 15745
rect 34005 15705 34045 15745
rect 34055 15705 34095 15745
rect 34105 15705 34145 15745
rect 34155 15705 34195 15745
rect 34205 15705 34245 15745
rect 34255 15705 34295 15745
rect 34305 15705 34345 15745
rect 34355 15705 34395 15745
rect 34405 15705 34445 15745
rect 34455 15705 34495 15745
rect 34505 15705 34545 15745
rect 34555 15705 34595 15745
rect 34605 15705 34645 15745
rect 34655 15705 34695 15745
rect 34705 15705 34745 15745
rect 34755 15705 34795 15745
rect 34805 15705 34845 15745
rect 34855 15705 34895 15745
rect 34905 15705 34945 15745
rect 34955 15705 34995 15745
rect 35005 15705 35045 15745
rect 35055 15705 35095 15745
rect 35105 15705 35145 15745
rect 35155 15705 35195 15745
rect 35205 15705 35245 15745
rect 35255 15705 35295 15745
rect 35305 15705 35345 15745
rect 35355 15705 35395 15745
rect 35405 15705 35445 15745
rect 35455 15705 35495 15745
rect 35505 15705 35545 15745
rect 35555 15705 35595 15745
rect 35605 15705 35645 15745
rect 35655 15705 35695 15745
rect 35705 15705 35745 15745
rect 35755 15705 35795 15745
rect 35805 15705 35845 15745
rect 35855 15705 35895 15745
rect 35905 15705 35945 15745
rect 35955 15705 35995 15745
rect 36005 15705 36045 15745
rect 36055 15705 36095 15745
rect 36105 15705 36145 15745
rect 36155 15705 36195 15745
rect 36205 15705 36245 15745
rect 36255 15705 36295 15745
rect 36305 15705 36345 15745
rect 36355 15705 36395 15745
rect 36405 15705 36445 15745
rect 36455 15705 36495 15745
rect 36505 15705 36545 15745
rect 36555 15705 36595 15745
rect 36605 15705 36645 15745
rect 36655 15705 36695 15745
rect 36705 15705 36745 15745
rect 36755 15705 36795 15745
rect 36805 15705 36845 15745
rect 36855 15705 36895 15745
rect 36905 15705 36945 15745
rect 36955 15705 36995 15745
rect 37005 15705 37045 15745
rect 37055 15705 37095 15745
rect 37105 15705 37145 15745
rect 37155 15705 37195 15745
rect 37205 15705 37245 15745
rect 37255 15705 37295 15745
rect 37305 15705 37345 15745
rect 37355 15705 37395 15745
rect 37405 15705 37445 15745
rect 37455 15705 37495 15745
rect 37505 15705 37545 15745
rect 37555 15705 37595 15745
rect 37605 15705 37645 15745
rect 37655 15705 37695 15745
rect 37705 15705 37745 15745
rect 37755 15705 37795 15745
rect 37805 15705 37845 15745
rect 37855 15705 37895 15745
rect 37905 15705 37945 15745
rect 37955 15705 37995 15745
rect 38005 15705 38045 15745
rect 38055 15705 38095 15745
rect 38105 15705 38145 15745
rect 38155 15705 38195 15745
rect 38205 15705 38245 15745
rect 38255 15705 38295 15745
rect 38305 15705 38345 15745
rect 38355 15705 38395 15745
rect 38405 15705 38445 15745
rect 38455 15705 38495 15745
rect 38505 15705 38545 15745
rect 38555 15705 38595 15745
rect 38605 15705 38645 15745
rect 38655 15705 38695 15745
rect 38705 15705 38745 15745
rect 38755 15705 38795 15745
rect 38805 15705 38845 15745
rect 38855 15705 38895 15745
rect 38905 15705 38945 15745
rect 38955 15705 38995 15745
rect 39005 15705 39045 15745
rect 39055 15705 39095 15745
rect 39105 15705 39145 15745
rect 39155 15705 39195 15745
rect 39205 15705 39245 15745
rect 39255 15705 39295 15745
rect 39305 15705 39345 15745
rect 39355 15705 39395 15745
rect 39405 15705 39445 15745
rect 39455 15705 39495 15745
rect 39505 15705 39545 15745
rect 39555 15705 39595 15745
rect 39605 15705 39645 15745
rect 39655 15705 39695 15745
rect 39705 15705 39745 15745
rect 39905 15705 39945 15745
rect 39955 15705 39995 15745
rect 40005 15705 40045 15745
rect 40055 15705 40095 15745
rect 40105 15705 40145 15745
rect 40155 15705 40195 15745
rect 40205 15705 40245 15745
rect 40255 15705 40295 15745
rect 40305 15705 40345 15745
rect 40355 15705 40395 15745
rect 40405 15705 40445 15745
rect 40455 15705 40495 15745
rect 40505 15705 40545 15745
rect 40555 15705 40595 15745
rect 40605 15705 40645 15745
rect 40655 15705 40695 15745
rect 40705 15705 40745 15745
rect 40755 15705 40795 15745
rect 40805 15705 40845 15745
rect 40855 15705 40895 15745
rect -3495 15340 -3455 15345
rect -3495 15310 -3490 15340
rect -3490 15310 -3460 15340
rect -3460 15310 -3455 15340
rect -3495 15305 -3455 15310
rect -3295 15340 -3255 15345
rect -3295 15310 -3290 15340
rect -3290 15310 -3260 15340
rect -3260 15310 -3255 15340
rect -3295 15305 -3255 15310
rect -3095 15340 -3055 15345
rect -3095 15310 -3090 15340
rect -3090 15310 -3060 15340
rect -3060 15310 -3055 15340
rect -3095 15305 -3055 15310
rect -1595 15340 -1555 15345
rect -1595 15310 -1590 15340
rect -1590 15310 -1560 15340
rect -1560 15310 -1555 15340
rect -1595 15305 -1555 15310
rect -1095 15340 -1055 15345
rect -1095 15310 -1090 15340
rect -1090 15310 -1060 15340
rect -1060 15310 -1055 15340
rect -1095 15305 -1055 15310
rect -895 15340 -855 15345
rect -895 15310 -890 15340
rect -890 15310 -860 15340
rect -860 15310 -855 15340
rect -895 15305 -855 15310
rect -695 15340 -655 15345
rect -695 15310 -690 15340
rect -690 15310 -660 15340
rect -660 15310 -655 15340
rect -695 15305 -655 15310
rect -495 15340 -455 15345
rect -495 15310 -490 15340
rect -490 15310 -460 15340
rect -460 15310 -455 15340
rect -495 15305 -455 15310
rect -295 15340 -255 15345
rect -295 15310 -290 15340
rect -290 15310 -260 15340
rect -260 15310 -255 15340
rect -295 15305 -255 15310
rect -95 15340 -55 15345
rect -95 15310 -90 15340
rect -90 15310 -60 15340
rect -60 15310 -55 15340
rect -95 15305 -55 15310
rect -3495 15290 -3455 15295
rect -3495 15260 -3490 15290
rect -3490 15260 -3460 15290
rect -3460 15260 -3455 15290
rect -3495 15255 -3455 15260
rect -3295 15290 -3255 15295
rect -3295 15260 -3290 15290
rect -3290 15260 -3260 15290
rect -3260 15260 -3255 15290
rect -3295 15255 -3255 15260
rect -3095 15290 -3055 15295
rect -3095 15260 -3090 15290
rect -3090 15260 -3060 15290
rect -3060 15260 -3055 15290
rect -3095 15255 -3055 15260
rect -1595 15290 -1555 15295
rect -1595 15260 -1590 15290
rect -1590 15260 -1560 15290
rect -1560 15260 -1555 15290
rect -1595 15255 -1555 15260
rect -1095 15290 -1055 15295
rect -1095 15260 -1090 15290
rect -1090 15260 -1060 15290
rect -1060 15260 -1055 15290
rect -1095 15255 -1055 15260
rect -895 15290 -855 15295
rect -895 15260 -890 15290
rect -890 15260 -860 15290
rect -860 15260 -855 15290
rect -895 15255 -855 15260
rect -695 15290 -655 15295
rect -695 15260 -690 15290
rect -690 15260 -660 15290
rect -660 15260 -655 15290
rect -695 15255 -655 15260
rect -495 15290 -455 15295
rect -495 15260 -490 15290
rect -490 15260 -460 15290
rect -460 15260 -455 15290
rect -495 15255 -455 15260
rect -295 15290 -255 15295
rect -295 15260 -290 15290
rect -290 15260 -260 15290
rect -260 15260 -255 15290
rect -295 15255 -255 15260
rect -95 15290 -55 15295
rect -95 15260 -90 15290
rect -90 15260 -60 15290
rect -60 15260 -55 15290
rect -95 15255 -55 15260
rect -3495 15240 -3455 15245
rect -3495 15210 -3490 15240
rect -3490 15210 -3460 15240
rect -3460 15210 -3455 15240
rect -3495 15205 -3455 15210
rect -3295 15240 -3255 15245
rect -3295 15210 -3290 15240
rect -3290 15210 -3260 15240
rect -3260 15210 -3255 15240
rect -3295 15205 -3255 15210
rect -3095 15240 -3055 15245
rect -3095 15210 -3090 15240
rect -3090 15210 -3060 15240
rect -3060 15210 -3055 15240
rect -3095 15205 -3055 15210
rect -1595 15240 -1555 15245
rect -1595 15210 -1590 15240
rect -1590 15210 -1560 15240
rect -1560 15210 -1555 15240
rect -1595 15205 -1555 15210
rect -1095 15240 -1055 15245
rect -1095 15210 -1090 15240
rect -1090 15210 -1060 15240
rect -1060 15210 -1055 15240
rect -1095 15205 -1055 15210
rect -895 15240 -855 15245
rect -895 15210 -890 15240
rect -890 15210 -860 15240
rect -860 15210 -855 15240
rect -895 15205 -855 15210
rect -695 15240 -655 15245
rect -695 15210 -690 15240
rect -690 15210 -660 15240
rect -660 15210 -655 15240
rect -695 15205 -655 15210
rect -495 15240 -455 15245
rect -495 15210 -490 15240
rect -490 15210 -460 15240
rect -460 15210 -455 15240
rect -495 15205 -455 15210
rect -295 15240 -255 15245
rect -295 15210 -290 15240
rect -290 15210 -260 15240
rect -260 15210 -255 15240
rect -295 15205 -255 15210
rect -95 15240 -55 15245
rect -95 15210 -90 15240
rect -90 15210 -60 15240
rect -60 15210 -55 15240
rect -95 15205 -55 15210
rect -195 14605 -155 14645
rect -395 14205 -355 14245
rect -595 14005 -555 14045
rect -3495 13640 -3455 13645
rect -3495 13610 -3490 13640
rect -3490 13610 -3460 13640
rect -3460 13610 -3455 13640
rect -3495 13605 -3455 13610
rect -3295 13640 -3255 13645
rect -3295 13610 -3290 13640
rect -3290 13610 -3260 13640
rect -3260 13610 -3255 13640
rect -3295 13605 -3255 13610
rect -3095 13640 -3055 13645
rect -3095 13610 -3090 13640
rect -3090 13610 -3060 13640
rect -3060 13610 -3055 13640
rect -3095 13605 -3055 13610
rect -1595 13640 -1555 13645
rect -1595 13610 -1590 13640
rect -1590 13610 -1560 13640
rect -1560 13610 -1555 13640
rect -1595 13605 -1555 13610
rect -1095 13640 -1055 13645
rect -1095 13610 -1090 13640
rect -1090 13610 -1060 13640
rect -1060 13610 -1055 13640
rect -1095 13605 -1055 13610
rect -895 13640 -855 13645
rect -895 13610 -890 13640
rect -890 13610 -860 13640
rect -860 13610 -855 13640
rect -895 13605 -855 13610
rect -695 13640 -655 13645
rect -695 13610 -690 13640
rect -690 13610 -660 13640
rect -660 13610 -655 13640
rect -695 13605 -655 13610
rect -495 13640 -455 13645
rect -495 13610 -490 13640
rect -490 13610 -460 13640
rect -460 13610 -455 13640
rect -495 13605 -455 13610
rect -295 13640 -255 13645
rect -295 13610 -290 13640
rect -290 13610 -260 13640
rect -260 13610 -255 13640
rect -295 13605 -255 13610
rect -95 13640 -55 13645
rect -95 13610 -90 13640
rect -90 13610 -60 13640
rect -60 13610 -55 13640
rect -95 13605 -55 13610
rect -3495 13590 -3455 13595
rect -3495 13560 -3490 13590
rect -3490 13560 -3460 13590
rect -3460 13560 -3455 13590
rect -3495 13555 -3455 13560
rect -3295 13590 -3255 13595
rect -3295 13560 -3290 13590
rect -3290 13560 -3260 13590
rect -3260 13560 -3255 13590
rect -3295 13555 -3255 13560
rect -3095 13590 -3055 13595
rect -3095 13560 -3090 13590
rect -3090 13560 -3060 13590
rect -3060 13560 -3055 13590
rect -3095 13555 -3055 13560
rect -1595 13590 -1555 13595
rect -1595 13560 -1590 13590
rect -1590 13560 -1560 13590
rect -1560 13560 -1555 13590
rect -1595 13555 -1555 13560
rect -1095 13590 -1055 13595
rect -1095 13560 -1090 13590
rect -1090 13560 -1060 13590
rect -1060 13560 -1055 13590
rect -1095 13555 -1055 13560
rect -895 13590 -855 13595
rect -895 13560 -890 13590
rect -890 13560 -860 13590
rect -860 13560 -855 13590
rect -895 13555 -855 13560
rect -695 13590 -655 13595
rect -695 13560 -690 13590
rect -690 13560 -660 13590
rect -660 13560 -655 13590
rect -695 13555 -655 13560
rect -495 13590 -455 13595
rect -495 13560 -490 13590
rect -490 13560 -460 13590
rect -460 13560 -455 13590
rect -495 13555 -455 13560
rect -295 13590 -255 13595
rect -295 13560 -290 13590
rect -290 13560 -260 13590
rect -260 13560 -255 13590
rect -295 13555 -255 13560
rect -95 13590 -55 13595
rect -95 13560 -90 13590
rect -90 13560 -60 13590
rect -60 13560 -55 13590
rect -95 13555 -55 13560
rect -3495 13540 -3455 13545
rect -3495 13510 -3490 13540
rect -3490 13510 -3460 13540
rect -3460 13510 -3455 13540
rect -3495 13505 -3455 13510
rect -3295 13540 -3255 13545
rect -3295 13510 -3290 13540
rect -3290 13510 -3260 13540
rect -3260 13510 -3255 13540
rect -3295 13505 -3255 13510
rect -3095 13540 -3055 13545
rect -3095 13510 -3090 13540
rect -3090 13510 -3060 13540
rect -3060 13510 -3055 13540
rect -3095 13505 -3055 13510
rect -1595 13540 -1555 13545
rect -1595 13510 -1590 13540
rect -1590 13510 -1560 13540
rect -1560 13510 -1555 13540
rect -1595 13505 -1555 13510
rect -1095 13540 -1055 13545
rect -1095 13510 -1090 13540
rect -1090 13510 -1060 13540
rect -1060 13510 -1055 13540
rect -1095 13505 -1055 13510
rect -895 13540 -855 13545
rect -895 13510 -890 13540
rect -890 13510 -860 13540
rect -860 13510 -855 13540
rect -895 13505 -855 13510
rect -695 13540 -655 13545
rect -695 13510 -690 13540
rect -690 13510 -660 13540
rect -660 13510 -655 13540
rect -695 13505 -655 13510
rect -495 13540 -455 13545
rect -495 13510 -490 13540
rect -490 13510 -460 13540
rect -460 13510 -455 13540
rect -495 13505 -455 13510
rect -295 13540 -255 13545
rect -295 13510 -290 13540
rect -290 13510 -260 13540
rect -260 13510 -255 13540
rect -295 13505 -255 13510
rect -95 13540 -55 13545
rect -95 13510 -90 13540
rect -90 13510 -60 13540
rect -60 13510 -55 13540
rect -95 13505 -55 13510
rect -795 13105 -755 13145
rect -995 12905 -955 12945
rect -1195 12505 -1155 12545
rect -1295 12405 -1255 12445
rect -1395 12305 -1355 12345
rect -1495 12205 -1455 12245
rect -3495 11940 -3455 11945
rect -3495 11910 -3490 11940
rect -3490 11910 -3460 11940
rect -3460 11910 -3455 11940
rect -3495 11905 -3455 11910
rect -3295 11940 -3255 11945
rect -3295 11910 -3290 11940
rect -3290 11910 -3260 11940
rect -3260 11910 -3255 11940
rect -3295 11905 -3255 11910
rect -3095 11940 -3055 11945
rect -3095 11910 -3090 11940
rect -3090 11910 -3060 11940
rect -3060 11910 -3055 11940
rect -3095 11905 -3055 11910
rect -1595 11940 -1555 11945
rect -1595 11910 -1590 11940
rect -1590 11910 -1560 11940
rect -1560 11910 -1555 11940
rect -1595 11905 -1555 11910
rect -1095 11940 -1055 11945
rect -1095 11910 -1090 11940
rect -1090 11910 -1060 11940
rect -1060 11910 -1055 11940
rect -1095 11905 -1055 11910
rect -895 11940 -855 11945
rect -895 11910 -890 11940
rect -890 11910 -860 11940
rect -860 11910 -855 11940
rect -895 11905 -855 11910
rect -695 11940 -655 11945
rect -695 11910 -690 11940
rect -690 11910 -660 11940
rect -660 11910 -655 11940
rect -695 11905 -655 11910
rect -495 11940 -455 11945
rect -495 11910 -490 11940
rect -490 11910 -460 11940
rect -460 11910 -455 11940
rect -495 11905 -455 11910
rect -295 11940 -255 11945
rect -295 11910 -290 11940
rect -290 11910 -260 11940
rect -260 11910 -255 11940
rect -295 11905 -255 11910
rect -95 11940 -55 11945
rect -95 11910 -90 11940
rect -90 11910 -60 11940
rect -60 11910 -55 11940
rect -95 11905 -55 11910
rect -3495 11890 -3455 11895
rect -3495 11860 -3490 11890
rect -3490 11860 -3460 11890
rect -3460 11860 -3455 11890
rect -3495 11855 -3455 11860
rect -3295 11890 -3255 11895
rect -3295 11860 -3290 11890
rect -3290 11860 -3260 11890
rect -3260 11860 -3255 11890
rect -3295 11855 -3255 11860
rect -3095 11890 -3055 11895
rect -3095 11860 -3090 11890
rect -3090 11860 -3060 11890
rect -3060 11860 -3055 11890
rect -3095 11855 -3055 11860
rect -1595 11890 -1555 11895
rect -1595 11860 -1590 11890
rect -1590 11860 -1560 11890
rect -1560 11860 -1555 11890
rect -1595 11855 -1555 11860
rect -1095 11890 -1055 11895
rect -1095 11860 -1090 11890
rect -1090 11860 -1060 11890
rect -1060 11860 -1055 11890
rect -1095 11855 -1055 11860
rect -895 11890 -855 11895
rect -895 11860 -890 11890
rect -890 11860 -860 11890
rect -860 11860 -855 11890
rect -895 11855 -855 11860
rect -695 11890 -655 11895
rect -695 11860 -690 11890
rect -690 11860 -660 11890
rect -660 11860 -655 11890
rect -695 11855 -655 11860
rect -495 11890 -455 11895
rect -495 11860 -490 11890
rect -490 11860 -460 11890
rect -460 11860 -455 11890
rect -495 11855 -455 11860
rect -295 11890 -255 11895
rect -295 11860 -290 11890
rect -290 11860 -260 11890
rect -260 11860 -255 11890
rect -295 11855 -255 11860
rect -95 11890 -55 11895
rect -95 11860 -90 11890
rect -90 11860 -60 11890
rect -60 11860 -55 11890
rect -95 11855 -55 11860
rect -3495 11840 -3455 11845
rect -3495 11810 -3490 11840
rect -3490 11810 -3460 11840
rect -3460 11810 -3455 11840
rect -3495 11805 -3455 11810
rect -3295 11840 -3255 11845
rect -3295 11810 -3290 11840
rect -3290 11810 -3260 11840
rect -3260 11810 -3255 11840
rect -3295 11805 -3255 11810
rect -3095 11840 -3055 11845
rect -3095 11810 -3090 11840
rect -3090 11810 -3060 11840
rect -3060 11810 -3055 11840
rect -3095 11805 -3055 11810
rect -1595 11840 -1555 11845
rect -1595 11810 -1590 11840
rect -1590 11810 -1560 11840
rect -1560 11810 -1555 11840
rect -1595 11805 -1555 11810
rect -1095 11840 -1055 11845
rect -1095 11810 -1090 11840
rect -1090 11810 -1060 11840
rect -1060 11810 -1055 11840
rect -1095 11805 -1055 11810
rect -895 11840 -855 11845
rect -895 11810 -890 11840
rect -890 11810 -860 11840
rect -860 11810 -855 11840
rect -895 11805 -855 11810
rect -695 11840 -655 11845
rect -695 11810 -690 11840
rect -690 11810 -660 11840
rect -660 11810 -655 11840
rect -695 11805 -655 11810
rect -495 11840 -455 11845
rect -495 11810 -490 11840
rect -490 11810 -460 11840
rect -460 11810 -455 11840
rect -495 11805 -455 11810
rect -295 11840 -255 11845
rect -295 11810 -290 11840
rect -290 11810 -260 11840
rect -260 11810 -255 11840
rect -295 11805 -255 11810
rect -95 11840 -55 11845
rect -95 11810 -90 11840
rect -90 11810 -60 11840
rect -60 11810 -55 11840
rect -95 11805 -55 11810
rect -3195 11405 -3155 11445
rect 39805 11340 39845 11345
rect 39805 11310 39810 11340
rect 39810 11310 39840 11340
rect 39840 11310 39845 11340
rect 39805 11305 39845 11310
rect 39905 11240 39945 11245
rect 39905 11210 39910 11240
rect 39910 11210 39940 11240
rect 39940 11210 39945 11240
rect 39905 11205 39945 11210
rect 39955 11240 39995 11245
rect 39955 11210 39960 11240
rect 39960 11210 39990 11240
rect 39990 11210 39995 11240
rect 39955 11205 39995 11210
rect 40005 11240 40045 11245
rect 40005 11210 40010 11240
rect 40010 11210 40040 11240
rect 40040 11210 40045 11240
rect 40005 11205 40045 11210
rect 40055 11240 40095 11245
rect 40055 11210 40060 11240
rect 40060 11210 40090 11240
rect 40090 11210 40095 11240
rect 40055 11205 40095 11210
rect 40105 11240 40145 11245
rect 40105 11210 40110 11240
rect 40110 11210 40140 11240
rect 40140 11210 40145 11240
rect 40105 11205 40145 11210
rect 40155 11240 40195 11245
rect 40155 11210 40160 11240
rect 40160 11210 40190 11240
rect 40190 11210 40195 11240
rect 40155 11205 40195 11210
rect 40205 11240 40245 11245
rect 40205 11210 40210 11240
rect 40210 11210 40240 11240
rect 40240 11210 40245 11240
rect 40205 11205 40245 11210
rect 40255 11240 40295 11245
rect 40255 11210 40260 11240
rect 40260 11210 40290 11240
rect 40290 11210 40295 11240
rect 40255 11205 40295 11210
rect 40305 11240 40345 11245
rect 40305 11210 40310 11240
rect 40310 11210 40340 11240
rect 40340 11210 40345 11240
rect 40305 11205 40345 11210
rect 40355 11240 40395 11245
rect 40355 11210 40360 11240
rect 40360 11210 40390 11240
rect 40390 11210 40395 11240
rect 40355 11205 40395 11210
rect 40405 11240 40445 11245
rect 40405 11210 40410 11240
rect 40410 11210 40440 11240
rect 40440 11210 40445 11240
rect 40405 11205 40445 11210
rect 40455 11240 40495 11245
rect 40455 11210 40460 11240
rect 40460 11210 40490 11240
rect 40490 11210 40495 11240
rect 40455 11205 40495 11210
rect 40505 11240 40545 11245
rect 40505 11210 40510 11240
rect 40510 11210 40540 11240
rect 40540 11210 40545 11240
rect 40505 11205 40545 11210
rect 40555 11240 40595 11245
rect 40555 11210 40560 11240
rect 40560 11210 40590 11240
rect 40590 11210 40595 11240
rect 40555 11205 40595 11210
rect 40605 11240 40645 11245
rect 40605 11210 40610 11240
rect 40610 11210 40640 11240
rect 40640 11210 40645 11240
rect 40605 11205 40645 11210
rect 40655 11240 40695 11245
rect 40655 11210 40660 11240
rect 40660 11210 40690 11240
rect 40690 11210 40695 11240
rect 40655 11205 40695 11210
rect 40705 11240 40745 11245
rect 40705 11210 40710 11240
rect 40710 11210 40740 11240
rect 40740 11210 40745 11240
rect 40705 11205 40745 11210
rect 40755 11240 40795 11245
rect 40755 11210 40760 11240
rect 40760 11210 40790 11240
rect 40790 11210 40795 11240
rect 40755 11205 40795 11210
rect 40805 11240 40845 11245
rect 40805 11210 40810 11240
rect 40810 11210 40840 11240
rect 40840 11210 40845 11240
rect 40805 11205 40845 11210
rect 40855 11240 40895 11245
rect 40855 11210 40860 11240
rect 40860 11210 40890 11240
rect 40890 11210 40895 11240
rect 40855 11205 40895 11210
rect 39905 11190 39945 11195
rect 39905 11160 39910 11190
rect 39910 11160 39940 11190
rect 39940 11160 39945 11190
rect 39905 11155 39945 11160
rect 39955 11190 39995 11195
rect 39955 11160 39960 11190
rect 39960 11160 39990 11190
rect 39990 11160 39995 11190
rect 39955 11155 39995 11160
rect 40005 11190 40045 11195
rect 40005 11160 40010 11190
rect 40010 11160 40040 11190
rect 40040 11160 40045 11190
rect 40005 11155 40045 11160
rect 40055 11190 40095 11195
rect 40055 11160 40060 11190
rect 40060 11160 40090 11190
rect 40090 11160 40095 11190
rect 40055 11155 40095 11160
rect 40105 11190 40145 11195
rect 40105 11160 40110 11190
rect 40110 11160 40140 11190
rect 40140 11160 40145 11190
rect 40105 11155 40145 11160
rect 40155 11190 40195 11195
rect 40155 11160 40160 11190
rect 40160 11160 40190 11190
rect 40190 11160 40195 11190
rect 40155 11155 40195 11160
rect 40205 11190 40245 11195
rect 40205 11160 40210 11190
rect 40210 11160 40240 11190
rect 40240 11160 40245 11190
rect 40205 11155 40245 11160
rect 40255 11190 40295 11195
rect 40255 11160 40260 11190
rect 40260 11160 40290 11190
rect 40290 11160 40295 11190
rect 40255 11155 40295 11160
rect 40305 11190 40345 11195
rect 40305 11160 40310 11190
rect 40310 11160 40340 11190
rect 40340 11160 40345 11190
rect 40305 11155 40345 11160
rect 40355 11190 40395 11195
rect 40355 11160 40360 11190
rect 40360 11160 40390 11190
rect 40390 11160 40395 11190
rect 40355 11155 40395 11160
rect 40405 11190 40445 11195
rect 40405 11160 40410 11190
rect 40410 11160 40440 11190
rect 40440 11160 40445 11190
rect 40405 11155 40445 11160
rect 40455 11190 40495 11195
rect 40455 11160 40460 11190
rect 40460 11160 40490 11190
rect 40490 11160 40495 11190
rect 40455 11155 40495 11160
rect 40505 11190 40545 11195
rect 40505 11160 40510 11190
rect 40510 11160 40540 11190
rect 40540 11160 40545 11190
rect 40505 11155 40545 11160
rect 40555 11190 40595 11195
rect 40555 11160 40560 11190
rect 40560 11160 40590 11190
rect 40590 11160 40595 11190
rect 40555 11155 40595 11160
rect 40605 11190 40645 11195
rect 40605 11160 40610 11190
rect 40610 11160 40640 11190
rect 40640 11160 40645 11190
rect 40605 11155 40645 11160
rect 40655 11190 40695 11195
rect 40655 11160 40660 11190
rect 40660 11160 40690 11190
rect 40690 11160 40695 11190
rect 40655 11155 40695 11160
rect 40705 11190 40745 11195
rect 40705 11160 40710 11190
rect 40710 11160 40740 11190
rect 40740 11160 40745 11190
rect 40705 11155 40745 11160
rect 40755 11190 40795 11195
rect 40755 11160 40760 11190
rect 40760 11160 40790 11190
rect 40790 11160 40795 11190
rect 40755 11155 40795 11160
rect 40805 11190 40845 11195
rect 40805 11160 40810 11190
rect 40810 11160 40840 11190
rect 40840 11160 40845 11190
rect 40805 11155 40845 11160
rect 40855 11190 40895 11195
rect 40855 11160 40860 11190
rect 40860 11160 40890 11190
rect 40890 11160 40895 11190
rect 40855 11155 40895 11160
rect 39905 11140 39945 11145
rect 39905 11110 39910 11140
rect 39910 11110 39940 11140
rect 39940 11110 39945 11140
rect 39905 11105 39945 11110
rect 39955 11140 39995 11145
rect 39955 11110 39960 11140
rect 39960 11110 39990 11140
rect 39990 11110 39995 11140
rect 39955 11105 39995 11110
rect 40005 11140 40045 11145
rect 40005 11110 40010 11140
rect 40010 11110 40040 11140
rect 40040 11110 40045 11140
rect 40005 11105 40045 11110
rect 40055 11140 40095 11145
rect 40055 11110 40060 11140
rect 40060 11110 40090 11140
rect 40090 11110 40095 11140
rect 40055 11105 40095 11110
rect 40105 11140 40145 11145
rect 40105 11110 40110 11140
rect 40110 11110 40140 11140
rect 40140 11110 40145 11140
rect 40105 11105 40145 11110
rect 40155 11140 40195 11145
rect 40155 11110 40160 11140
rect 40160 11110 40190 11140
rect 40190 11110 40195 11140
rect 40155 11105 40195 11110
rect 40205 11140 40245 11145
rect 40205 11110 40210 11140
rect 40210 11110 40240 11140
rect 40240 11110 40245 11140
rect 40205 11105 40245 11110
rect 40255 11140 40295 11145
rect 40255 11110 40260 11140
rect 40260 11110 40290 11140
rect 40290 11110 40295 11140
rect 40255 11105 40295 11110
rect 40305 11140 40345 11145
rect 40305 11110 40310 11140
rect 40310 11110 40340 11140
rect 40340 11110 40345 11140
rect 40305 11105 40345 11110
rect 40355 11140 40395 11145
rect 40355 11110 40360 11140
rect 40360 11110 40390 11140
rect 40390 11110 40395 11140
rect 40355 11105 40395 11110
rect 40405 11140 40445 11145
rect 40405 11110 40410 11140
rect 40410 11110 40440 11140
rect 40440 11110 40445 11140
rect 40405 11105 40445 11110
rect 40455 11140 40495 11145
rect 40455 11110 40460 11140
rect 40460 11110 40490 11140
rect 40490 11110 40495 11140
rect 40455 11105 40495 11110
rect 40505 11140 40545 11145
rect 40505 11110 40510 11140
rect 40510 11110 40540 11140
rect 40540 11110 40545 11140
rect 40505 11105 40545 11110
rect 40555 11140 40595 11145
rect 40555 11110 40560 11140
rect 40560 11110 40590 11140
rect 40590 11110 40595 11140
rect 40555 11105 40595 11110
rect 40605 11140 40645 11145
rect 40605 11110 40610 11140
rect 40610 11110 40640 11140
rect 40640 11110 40645 11140
rect 40605 11105 40645 11110
rect 40655 11140 40695 11145
rect 40655 11110 40660 11140
rect 40660 11110 40690 11140
rect 40690 11110 40695 11140
rect 40655 11105 40695 11110
rect 40705 11140 40745 11145
rect 40705 11110 40710 11140
rect 40710 11110 40740 11140
rect 40740 11110 40745 11140
rect 40705 11105 40745 11110
rect 40755 11140 40795 11145
rect 40755 11110 40760 11140
rect 40760 11110 40790 11140
rect 40790 11110 40795 11140
rect 40755 11105 40795 11110
rect 40805 11140 40845 11145
rect 40805 11110 40810 11140
rect 40810 11110 40840 11140
rect 40840 11110 40845 11140
rect 40805 11105 40845 11110
rect 40855 11140 40895 11145
rect 40855 11110 40860 11140
rect 40860 11110 40890 11140
rect 40890 11110 40895 11140
rect 40855 11105 40895 11110
rect 39905 11090 39945 11095
rect 39905 11060 39910 11090
rect 39910 11060 39940 11090
rect 39940 11060 39945 11090
rect 39905 11055 39945 11060
rect 39955 11090 39995 11095
rect 39955 11060 39960 11090
rect 39960 11060 39990 11090
rect 39990 11060 39995 11090
rect 39955 11055 39995 11060
rect 40005 11090 40045 11095
rect 40005 11060 40010 11090
rect 40010 11060 40040 11090
rect 40040 11060 40045 11090
rect 40005 11055 40045 11060
rect 40055 11090 40095 11095
rect 40055 11060 40060 11090
rect 40060 11060 40090 11090
rect 40090 11060 40095 11090
rect 40055 11055 40095 11060
rect 40105 11090 40145 11095
rect 40105 11060 40110 11090
rect 40110 11060 40140 11090
rect 40140 11060 40145 11090
rect 40105 11055 40145 11060
rect 40155 11090 40195 11095
rect 40155 11060 40160 11090
rect 40160 11060 40190 11090
rect 40190 11060 40195 11090
rect 40155 11055 40195 11060
rect 40205 11090 40245 11095
rect 40205 11060 40210 11090
rect 40210 11060 40240 11090
rect 40240 11060 40245 11090
rect 40205 11055 40245 11060
rect 40255 11090 40295 11095
rect 40255 11060 40260 11090
rect 40260 11060 40290 11090
rect 40290 11060 40295 11090
rect 40255 11055 40295 11060
rect 40305 11090 40345 11095
rect 40305 11060 40310 11090
rect 40310 11060 40340 11090
rect 40340 11060 40345 11090
rect 40305 11055 40345 11060
rect 40355 11090 40395 11095
rect 40355 11060 40360 11090
rect 40360 11060 40390 11090
rect 40390 11060 40395 11090
rect 40355 11055 40395 11060
rect 40405 11090 40445 11095
rect 40405 11060 40410 11090
rect 40410 11060 40440 11090
rect 40440 11060 40445 11090
rect 40405 11055 40445 11060
rect 40455 11090 40495 11095
rect 40455 11060 40460 11090
rect 40460 11060 40490 11090
rect 40490 11060 40495 11090
rect 40455 11055 40495 11060
rect 40505 11090 40545 11095
rect 40505 11060 40510 11090
rect 40510 11060 40540 11090
rect 40540 11060 40545 11090
rect 40505 11055 40545 11060
rect 40555 11090 40595 11095
rect 40555 11060 40560 11090
rect 40560 11060 40590 11090
rect 40590 11060 40595 11090
rect 40555 11055 40595 11060
rect 40605 11090 40645 11095
rect 40605 11060 40610 11090
rect 40610 11060 40640 11090
rect 40640 11060 40645 11090
rect 40605 11055 40645 11060
rect 40655 11090 40695 11095
rect 40655 11060 40660 11090
rect 40660 11060 40690 11090
rect 40690 11060 40695 11090
rect 40655 11055 40695 11060
rect 40705 11090 40745 11095
rect 40705 11060 40710 11090
rect 40710 11060 40740 11090
rect 40740 11060 40745 11090
rect 40705 11055 40745 11060
rect 40755 11090 40795 11095
rect 40755 11060 40760 11090
rect 40760 11060 40790 11090
rect 40790 11060 40795 11090
rect 40755 11055 40795 11060
rect 40805 11090 40845 11095
rect 40805 11060 40810 11090
rect 40810 11060 40840 11090
rect 40840 11060 40845 11090
rect 40805 11055 40845 11060
rect 40855 11090 40895 11095
rect 40855 11060 40860 11090
rect 40860 11060 40890 11090
rect 40890 11060 40895 11090
rect 40855 11055 40895 11060
rect 39905 11040 39945 11045
rect 39905 11010 39910 11040
rect 39910 11010 39940 11040
rect 39940 11010 39945 11040
rect 39905 11005 39945 11010
rect 39955 11040 39995 11045
rect 39955 11010 39960 11040
rect 39960 11010 39990 11040
rect 39990 11010 39995 11040
rect 39955 11005 39995 11010
rect 40005 11040 40045 11045
rect 40005 11010 40010 11040
rect 40010 11010 40040 11040
rect 40040 11010 40045 11040
rect 40005 11005 40045 11010
rect 40055 11040 40095 11045
rect 40055 11010 40060 11040
rect 40060 11010 40090 11040
rect 40090 11010 40095 11040
rect 40055 11005 40095 11010
rect 40105 11040 40145 11045
rect 40105 11010 40110 11040
rect 40110 11010 40140 11040
rect 40140 11010 40145 11040
rect 40105 11005 40145 11010
rect 40155 11040 40195 11045
rect 40155 11010 40160 11040
rect 40160 11010 40190 11040
rect 40190 11010 40195 11040
rect 40155 11005 40195 11010
rect 40205 11040 40245 11045
rect 40205 11010 40210 11040
rect 40210 11010 40240 11040
rect 40240 11010 40245 11040
rect 40205 11005 40245 11010
rect 40255 11040 40295 11045
rect 40255 11010 40260 11040
rect 40260 11010 40290 11040
rect 40290 11010 40295 11040
rect 40255 11005 40295 11010
rect 40305 11040 40345 11045
rect 40305 11010 40310 11040
rect 40310 11010 40340 11040
rect 40340 11010 40345 11040
rect 40305 11005 40345 11010
rect 40355 11040 40395 11045
rect 40355 11010 40360 11040
rect 40360 11010 40390 11040
rect 40390 11010 40395 11040
rect 40355 11005 40395 11010
rect 40405 11040 40445 11045
rect 40405 11010 40410 11040
rect 40410 11010 40440 11040
rect 40440 11010 40445 11040
rect 40405 11005 40445 11010
rect 40455 11040 40495 11045
rect 40455 11010 40460 11040
rect 40460 11010 40490 11040
rect 40490 11010 40495 11040
rect 40455 11005 40495 11010
rect 40505 11040 40545 11045
rect 40505 11010 40510 11040
rect 40510 11010 40540 11040
rect 40540 11010 40545 11040
rect 40505 11005 40545 11010
rect 40555 11040 40595 11045
rect 40555 11010 40560 11040
rect 40560 11010 40590 11040
rect 40590 11010 40595 11040
rect 40555 11005 40595 11010
rect 40605 11040 40645 11045
rect 40605 11010 40610 11040
rect 40610 11010 40640 11040
rect 40640 11010 40645 11040
rect 40605 11005 40645 11010
rect 40655 11040 40695 11045
rect 40655 11010 40660 11040
rect 40660 11010 40690 11040
rect 40690 11010 40695 11040
rect 40655 11005 40695 11010
rect 40705 11040 40745 11045
rect 40705 11010 40710 11040
rect 40710 11010 40740 11040
rect 40740 11010 40745 11040
rect 40705 11005 40745 11010
rect 40755 11040 40795 11045
rect 40755 11010 40760 11040
rect 40760 11010 40790 11040
rect 40790 11010 40795 11040
rect 40755 11005 40795 11010
rect 40805 11040 40845 11045
rect 40805 11010 40810 11040
rect 40810 11010 40840 11040
rect 40840 11010 40845 11040
rect 40805 11005 40845 11010
rect 40855 11040 40895 11045
rect 40855 11010 40860 11040
rect 40860 11010 40890 11040
rect 40890 11010 40895 11040
rect 40855 11005 40895 11010
rect 39805 10940 39845 10945
rect 39805 10910 39810 10940
rect 39810 10910 39840 10940
rect 39840 10910 39845 10940
rect 39805 10905 39845 10910
rect -3395 10805 -3355 10845
rect -2995 10640 -2955 10645
rect -2995 10610 -2990 10640
rect -2990 10610 -2960 10640
rect -2960 10610 -2955 10640
rect -2995 10605 -2955 10610
rect -2795 10640 -2755 10645
rect -2795 10610 -2790 10640
rect -2790 10610 -2760 10640
rect -2760 10610 -2755 10640
rect -2795 10605 -2755 10610
rect -2595 10640 -2555 10645
rect -2595 10610 -2590 10640
rect -2590 10610 -2560 10640
rect -2560 10610 -2555 10640
rect -2595 10605 -2555 10610
rect -2395 10640 -2355 10645
rect -2395 10610 -2390 10640
rect -2390 10610 -2360 10640
rect -2360 10610 -2355 10640
rect -2395 10605 -2355 10610
rect -2195 10640 -2155 10645
rect -2195 10610 -2190 10640
rect -2190 10610 -2160 10640
rect -2160 10610 -2155 10640
rect -2195 10605 -2155 10610
rect -1995 10640 -1955 10645
rect -1995 10610 -1990 10640
rect -1990 10610 -1960 10640
rect -1960 10610 -1955 10640
rect -1995 10605 -1955 10610
rect -1695 10640 -1655 10645
rect -1695 10610 -1690 10640
rect -1690 10610 -1660 10640
rect -1660 10610 -1655 10640
rect -1695 10605 -1655 10610
rect -2995 10590 -2955 10595
rect -2995 10560 -2990 10590
rect -2990 10560 -2960 10590
rect -2960 10560 -2955 10590
rect -2995 10555 -2955 10560
rect -2795 10590 -2755 10595
rect -2795 10560 -2790 10590
rect -2790 10560 -2760 10590
rect -2760 10560 -2755 10590
rect -2795 10555 -2755 10560
rect -2595 10590 -2555 10595
rect -2595 10560 -2590 10590
rect -2590 10560 -2560 10590
rect -2560 10560 -2555 10590
rect -2595 10555 -2555 10560
rect -2395 10590 -2355 10595
rect -2395 10560 -2390 10590
rect -2390 10560 -2360 10590
rect -2360 10560 -2355 10590
rect -2395 10555 -2355 10560
rect -2195 10590 -2155 10595
rect -2195 10560 -2190 10590
rect -2190 10560 -2160 10590
rect -2160 10560 -2155 10590
rect -2195 10555 -2155 10560
rect -1995 10590 -1955 10595
rect -1995 10560 -1990 10590
rect -1990 10560 -1960 10590
rect -1960 10560 -1955 10590
rect -1995 10555 -1955 10560
rect -1695 10590 -1655 10595
rect -1695 10560 -1690 10590
rect -1690 10560 -1660 10590
rect -1660 10560 -1655 10590
rect -1695 10555 -1655 10560
rect -2995 10540 -2955 10545
rect -2995 10510 -2990 10540
rect -2990 10510 -2960 10540
rect -2960 10510 -2955 10540
rect -2995 10505 -2955 10510
rect -2795 10540 -2755 10545
rect -2795 10510 -2790 10540
rect -2790 10510 -2760 10540
rect -2760 10510 -2755 10540
rect -2795 10505 -2755 10510
rect -2595 10540 -2555 10545
rect -2595 10510 -2590 10540
rect -2590 10510 -2560 10540
rect -2560 10510 -2555 10540
rect -2595 10505 -2555 10510
rect -2395 10540 -2355 10545
rect -2395 10510 -2390 10540
rect -2390 10510 -2360 10540
rect -2360 10510 -2355 10540
rect -2395 10505 -2355 10510
rect -2195 10540 -2155 10545
rect -2195 10510 -2190 10540
rect -2190 10510 -2160 10540
rect -2160 10510 -2155 10540
rect -2195 10505 -2155 10510
rect -1995 10540 -1955 10545
rect -1995 10510 -1990 10540
rect -1990 10510 -1960 10540
rect -1960 10510 -1955 10540
rect -1995 10505 -1955 10510
rect -1695 10540 -1655 10545
rect -1695 10510 -1690 10540
rect -1690 10510 -1660 10540
rect -1660 10510 -1655 10540
rect -1695 10505 -1655 10510
rect -1795 10205 -1755 10245
rect -1895 10105 -1855 10145
rect -2095 9705 -2055 9745
rect -2295 9505 -2255 9545
rect -2995 9340 -2955 9345
rect -2995 9310 -2990 9340
rect -2990 9310 -2960 9340
rect -2960 9310 -2955 9340
rect -2995 9305 -2955 9310
rect -2795 9340 -2755 9345
rect -2795 9310 -2790 9340
rect -2790 9310 -2760 9340
rect -2760 9310 -2755 9340
rect -2795 9305 -2755 9310
rect -2595 9340 -2555 9345
rect -2595 9310 -2590 9340
rect -2590 9310 -2560 9340
rect -2560 9310 -2555 9340
rect -2595 9305 -2555 9310
rect -2395 9340 -2355 9345
rect -2395 9310 -2390 9340
rect -2390 9310 -2360 9340
rect -2360 9310 -2355 9340
rect -2395 9305 -2355 9310
rect -2195 9340 -2155 9345
rect -2195 9310 -2190 9340
rect -2190 9310 -2160 9340
rect -2160 9310 -2155 9340
rect -2195 9305 -2155 9310
rect -1995 9340 -1955 9345
rect -1995 9310 -1990 9340
rect -1990 9310 -1960 9340
rect -1960 9310 -1955 9340
rect -1995 9305 -1955 9310
rect -1695 9340 -1655 9345
rect -1695 9310 -1690 9340
rect -1690 9310 -1660 9340
rect -1660 9310 -1655 9340
rect -1695 9305 -1655 9310
rect -2995 9290 -2955 9295
rect -2995 9260 -2990 9290
rect -2990 9260 -2960 9290
rect -2960 9260 -2955 9290
rect -2995 9255 -2955 9260
rect -2795 9290 -2755 9295
rect -2795 9260 -2790 9290
rect -2790 9260 -2760 9290
rect -2760 9260 -2755 9290
rect -2795 9255 -2755 9260
rect -2595 9290 -2555 9295
rect -2595 9260 -2590 9290
rect -2590 9260 -2560 9290
rect -2560 9260 -2555 9290
rect -2595 9255 -2555 9260
rect -2395 9290 -2355 9295
rect -2395 9260 -2390 9290
rect -2390 9260 -2360 9290
rect -2360 9260 -2355 9290
rect -2395 9255 -2355 9260
rect -2195 9290 -2155 9295
rect -2195 9260 -2190 9290
rect -2190 9260 -2160 9290
rect -2160 9260 -2155 9290
rect -2195 9255 -2155 9260
rect -1995 9290 -1955 9295
rect -1995 9260 -1990 9290
rect -1990 9260 -1960 9290
rect -1960 9260 -1955 9290
rect -1995 9255 -1955 9260
rect -1695 9290 -1655 9295
rect -1695 9260 -1690 9290
rect -1690 9260 -1660 9290
rect -1660 9260 -1655 9290
rect -1695 9255 -1655 9260
rect -2995 9240 -2955 9245
rect -2995 9210 -2990 9240
rect -2990 9210 -2960 9240
rect -2960 9210 -2955 9240
rect -2995 9205 -2955 9210
rect -2795 9240 -2755 9245
rect -2795 9210 -2790 9240
rect -2790 9210 -2760 9240
rect -2760 9210 -2755 9240
rect -2795 9205 -2755 9210
rect -2595 9240 -2555 9245
rect -2595 9210 -2590 9240
rect -2590 9210 -2560 9240
rect -2560 9210 -2555 9240
rect -2595 9205 -2555 9210
rect -2395 9240 -2355 9245
rect -2395 9210 -2390 9240
rect -2390 9210 -2360 9240
rect -2360 9210 -2355 9240
rect -2395 9205 -2355 9210
rect -2195 9240 -2155 9245
rect -2195 9210 -2190 9240
rect -2190 9210 -2160 9240
rect -2160 9210 -2155 9240
rect -2195 9205 -2155 9210
rect -1995 9240 -1955 9245
rect -1995 9210 -1990 9240
rect -1990 9210 -1960 9240
rect -1960 9210 -1955 9240
rect -1995 9205 -1955 9210
rect -1695 9240 -1655 9245
rect -1695 9210 -1690 9240
rect -1690 9210 -1660 9240
rect -1660 9210 -1655 9240
rect -1695 9205 -1655 9210
rect -2495 9005 -2455 9045
rect -2695 8805 -2655 8845
rect -2895 8405 -2855 8445
rect -2995 8040 -2955 8045
rect -2995 8010 -2990 8040
rect -2990 8010 -2960 8040
rect -2960 8010 -2955 8040
rect -2995 8005 -2955 8010
rect -2795 8040 -2755 8045
rect -2795 8010 -2790 8040
rect -2790 8010 -2760 8040
rect -2760 8010 -2755 8040
rect -2795 8005 -2755 8010
rect -2595 8040 -2555 8045
rect -2595 8010 -2590 8040
rect -2590 8010 -2560 8040
rect -2560 8010 -2555 8040
rect -2595 8005 -2555 8010
rect -2395 8040 -2355 8045
rect -2395 8010 -2390 8040
rect -2390 8010 -2360 8040
rect -2360 8010 -2355 8040
rect -2395 8005 -2355 8010
rect -2195 8040 -2155 8045
rect -2195 8010 -2190 8040
rect -2190 8010 -2160 8040
rect -2160 8010 -2155 8040
rect -2195 8005 -2155 8010
rect -1995 8040 -1955 8045
rect -1995 8010 -1990 8040
rect -1990 8010 -1960 8040
rect -1960 8010 -1955 8040
rect -1995 8005 -1955 8010
rect -1695 8040 -1655 8045
rect -1695 8010 -1690 8040
rect -1690 8010 -1660 8040
rect -1660 8010 -1655 8040
rect -1695 8005 -1655 8010
rect -2995 7990 -2955 7995
rect -2995 7960 -2990 7990
rect -2990 7960 -2960 7990
rect -2960 7960 -2955 7990
rect -2995 7955 -2955 7960
rect -2795 7990 -2755 7995
rect -2795 7960 -2790 7990
rect -2790 7960 -2760 7990
rect -2760 7960 -2755 7990
rect -2795 7955 -2755 7960
rect -2595 7990 -2555 7995
rect -2595 7960 -2590 7990
rect -2590 7960 -2560 7990
rect -2560 7960 -2555 7990
rect -2595 7955 -2555 7960
rect -2395 7990 -2355 7995
rect -2395 7960 -2390 7990
rect -2390 7960 -2360 7990
rect -2360 7960 -2355 7990
rect -2395 7955 -2355 7960
rect -2195 7990 -2155 7995
rect -2195 7960 -2190 7990
rect -2190 7960 -2160 7990
rect -2160 7960 -2155 7990
rect -2195 7955 -2155 7960
rect -1995 7990 -1955 7995
rect -1995 7960 -1990 7990
rect -1990 7960 -1960 7990
rect -1960 7960 -1955 7990
rect -1995 7955 -1955 7960
rect -1695 7990 -1655 7995
rect -1695 7960 -1690 7990
rect -1690 7960 -1660 7990
rect -1660 7960 -1655 7990
rect -1695 7955 -1655 7960
rect -2995 7940 -2955 7945
rect -2995 7910 -2990 7940
rect -2990 7910 -2960 7940
rect -2960 7910 -2955 7940
rect -2995 7905 -2955 7910
rect -2795 7940 -2755 7945
rect -2795 7910 -2790 7940
rect -2790 7910 -2760 7940
rect -2760 7910 -2755 7940
rect -2795 7905 -2755 7910
rect -2595 7940 -2555 7945
rect -2595 7910 -2590 7940
rect -2590 7910 -2560 7940
rect -2560 7910 -2555 7940
rect -2595 7905 -2555 7910
rect -2395 7940 -2355 7945
rect -2395 7910 -2390 7940
rect -2390 7910 -2360 7940
rect -2360 7910 -2355 7940
rect -2395 7905 -2355 7910
rect -2195 7940 -2155 7945
rect -2195 7910 -2190 7940
rect -2190 7910 -2160 7940
rect -2160 7910 -2155 7940
rect -2195 7905 -2155 7910
rect -1995 7940 -1955 7945
rect -1995 7910 -1990 7940
rect -1990 7910 -1960 7940
rect -1960 7910 -1955 7940
rect -1995 7905 -1955 7910
rect -1695 7940 -1655 7945
rect -1695 7910 -1690 7940
rect -1690 7910 -1660 7940
rect -1660 7910 -1655 7940
rect -1695 7905 -1655 7910
rect -2995 7740 -2955 7745
rect -2995 7710 -2990 7740
rect -2990 7710 -2960 7740
rect -2960 7710 -2955 7740
rect -2995 7705 -2955 7710
rect -2795 7740 -2755 7745
rect -2795 7710 -2790 7740
rect -2790 7710 -2760 7740
rect -2760 7710 -2755 7740
rect -2795 7705 -2755 7710
rect -2595 7740 -2555 7745
rect -2595 7710 -2590 7740
rect -2590 7710 -2560 7740
rect -2560 7710 -2555 7740
rect -2595 7705 -2555 7710
rect -2395 7740 -2355 7745
rect -2395 7710 -2390 7740
rect -2390 7710 -2360 7740
rect -2360 7710 -2355 7740
rect -2395 7705 -2355 7710
rect -2195 7740 -2155 7745
rect -2195 7710 -2190 7740
rect -2190 7710 -2160 7740
rect -2160 7710 -2155 7740
rect -2195 7705 -2155 7710
rect -1995 7740 -1955 7745
rect -1995 7710 -1990 7740
rect -1990 7710 -1960 7740
rect -1960 7710 -1955 7740
rect -1995 7705 -1955 7710
rect -1695 7740 -1655 7745
rect -1695 7710 -1690 7740
rect -1690 7710 -1660 7740
rect -1660 7710 -1655 7740
rect -1695 7705 -1655 7710
rect -2995 7690 -2955 7695
rect -2995 7660 -2990 7690
rect -2990 7660 -2960 7690
rect -2960 7660 -2955 7690
rect -2995 7655 -2955 7660
rect -2795 7690 -2755 7695
rect -2795 7660 -2790 7690
rect -2790 7660 -2760 7690
rect -2760 7660 -2755 7690
rect -2795 7655 -2755 7660
rect -2595 7690 -2555 7695
rect -2595 7660 -2590 7690
rect -2590 7660 -2560 7690
rect -2560 7660 -2555 7690
rect -2595 7655 -2555 7660
rect -2395 7690 -2355 7695
rect -2395 7660 -2390 7690
rect -2390 7660 -2360 7690
rect -2360 7660 -2355 7690
rect -2395 7655 -2355 7660
rect -2195 7690 -2155 7695
rect -2195 7660 -2190 7690
rect -2190 7660 -2160 7690
rect -2160 7660 -2155 7690
rect -2195 7655 -2155 7660
rect -1995 7690 -1955 7695
rect -1995 7660 -1990 7690
rect -1990 7660 -1960 7690
rect -1960 7660 -1955 7690
rect -1995 7655 -1955 7660
rect -1695 7690 -1655 7695
rect -1695 7660 -1690 7690
rect -1690 7660 -1660 7690
rect -1660 7660 -1655 7690
rect -1695 7655 -1655 7660
rect -2995 7640 -2955 7645
rect -2995 7610 -2990 7640
rect -2990 7610 -2960 7640
rect -2960 7610 -2955 7640
rect -2995 7605 -2955 7610
rect -2795 7640 -2755 7645
rect -2795 7610 -2790 7640
rect -2790 7610 -2760 7640
rect -2760 7610 -2755 7640
rect -2795 7605 -2755 7610
rect -2595 7640 -2555 7645
rect -2595 7610 -2590 7640
rect -2590 7610 -2560 7640
rect -2560 7610 -2555 7640
rect -2595 7605 -2555 7610
rect -2395 7640 -2355 7645
rect -2395 7610 -2390 7640
rect -2390 7610 -2360 7640
rect -2360 7610 -2355 7640
rect -2395 7605 -2355 7610
rect -2195 7640 -2155 7645
rect -2195 7610 -2190 7640
rect -2190 7610 -2160 7640
rect -2160 7610 -2155 7640
rect -2195 7605 -2155 7610
rect -1995 7640 -1955 7645
rect -1995 7610 -1990 7640
rect -1990 7610 -1960 7640
rect -1960 7610 -1955 7640
rect -1995 7605 -1955 7610
rect -1695 7640 -1655 7645
rect -1695 7610 -1690 7640
rect -1690 7610 -1660 7640
rect -1660 7610 -1655 7640
rect -1695 7605 -1655 7610
rect -2895 7205 -2855 7245
rect -2695 6805 -2655 6845
rect -2495 6605 -2455 6645
rect -2995 6440 -2955 6445
rect -2995 6410 -2990 6440
rect -2990 6410 -2960 6440
rect -2960 6410 -2955 6440
rect -2995 6405 -2955 6410
rect -2795 6440 -2755 6445
rect -2795 6410 -2790 6440
rect -2790 6410 -2760 6440
rect -2760 6410 -2755 6440
rect -2795 6405 -2755 6410
rect -2595 6440 -2555 6445
rect -2595 6410 -2590 6440
rect -2590 6410 -2560 6440
rect -2560 6410 -2555 6440
rect -2595 6405 -2555 6410
rect -2395 6440 -2355 6445
rect -2395 6410 -2390 6440
rect -2390 6410 -2360 6440
rect -2360 6410 -2355 6440
rect -2395 6405 -2355 6410
rect -2195 6440 -2155 6445
rect -2195 6410 -2190 6440
rect -2190 6410 -2160 6440
rect -2160 6410 -2155 6440
rect -2195 6405 -2155 6410
rect -1995 6440 -1955 6445
rect -1995 6410 -1990 6440
rect -1990 6410 -1960 6440
rect -1960 6410 -1955 6440
rect -1995 6405 -1955 6410
rect -1695 6440 -1655 6445
rect -1695 6410 -1690 6440
rect -1690 6410 -1660 6440
rect -1660 6410 -1655 6440
rect -1695 6405 -1655 6410
rect -2995 6390 -2955 6395
rect -2995 6360 -2990 6390
rect -2990 6360 -2960 6390
rect -2960 6360 -2955 6390
rect -2995 6355 -2955 6360
rect -2795 6390 -2755 6395
rect -2795 6360 -2790 6390
rect -2790 6360 -2760 6390
rect -2760 6360 -2755 6390
rect -2795 6355 -2755 6360
rect -2595 6390 -2555 6395
rect -2595 6360 -2590 6390
rect -2590 6360 -2560 6390
rect -2560 6360 -2555 6390
rect -2595 6355 -2555 6360
rect -2395 6390 -2355 6395
rect -2395 6360 -2390 6390
rect -2390 6360 -2360 6390
rect -2360 6360 -2355 6390
rect -2395 6355 -2355 6360
rect -2195 6390 -2155 6395
rect -2195 6360 -2190 6390
rect -2190 6360 -2160 6390
rect -2160 6360 -2155 6390
rect -2195 6355 -2155 6360
rect -1995 6390 -1955 6395
rect -1995 6360 -1990 6390
rect -1990 6360 -1960 6390
rect -1960 6360 -1955 6390
rect -1995 6355 -1955 6360
rect -1695 6390 -1655 6395
rect -1695 6360 -1690 6390
rect -1690 6360 -1660 6390
rect -1660 6360 -1655 6390
rect -1695 6355 -1655 6360
rect -2995 6340 -2955 6345
rect -2995 6310 -2990 6340
rect -2990 6310 -2960 6340
rect -2960 6310 -2955 6340
rect -2995 6305 -2955 6310
rect -2795 6340 -2755 6345
rect -2795 6310 -2790 6340
rect -2790 6310 -2760 6340
rect -2760 6310 -2755 6340
rect -2795 6305 -2755 6310
rect -2595 6340 -2555 6345
rect -2595 6310 -2590 6340
rect -2590 6310 -2560 6340
rect -2560 6310 -2555 6340
rect -2595 6305 -2555 6310
rect -2395 6340 -2355 6345
rect -2395 6310 -2390 6340
rect -2390 6310 -2360 6340
rect -2360 6310 -2355 6340
rect -2395 6305 -2355 6310
rect -2195 6340 -2155 6345
rect -2195 6310 -2190 6340
rect -2190 6310 -2160 6340
rect -2160 6310 -2155 6340
rect -2195 6305 -2155 6310
rect -1995 6340 -1955 6345
rect -1995 6310 -1990 6340
rect -1990 6310 -1960 6340
rect -1960 6310 -1955 6340
rect -1995 6305 -1955 6310
rect -1695 6340 -1655 6345
rect -1695 6310 -1690 6340
rect -1690 6310 -1660 6340
rect -1660 6310 -1655 6340
rect -1695 6305 -1655 6310
rect -2295 6105 -2255 6145
rect -2095 5905 -2055 5945
rect -1895 5505 -1855 5545
rect -1795 5405 -1755 5445
rect -2995 5140 -2955 5145
rect -2995 5110 -2990 5140
rect -2990 5110 -2960 5140
rect -2960 5110 -2955 5140
rect -2995 5105 -2955 5110
rect -2795 5140 -2755 5145
rect -2795 5110 -2790 5140
rect -2790 5110 -2760 5140
rect -2760 5110 -2755 5140
rect -2795 5105 -2755 5110
rect -2595 5140 -2555 5145
rect -2595 5110 -2590 5140
rect -2590 5110 -2560 5140
rect -2560 5110 -2555 5140
rect -2595 5105 -2555 5110
rect -2395 5140 -2355 5145
rect -2395 5110 -2390 5140
rect -2390 5110 -2360 5140
rect -2360 5110 -2355 5140
rect -2395 5105 -2355 5110
rect -2195 5140 -2155 5145
rect -2195 5110 -2190 5140
rect -2190 5110 -2160 5140
rect -2160 5110 -2155 5140
rect -2195 5105 -2155 5110
rect -1995 5140 -1955 5145
rect -1995 5110 -1990 5140
rect -1990 5110 -1960 5140
rect -1960 5110 -1955 5140
rect -1995 5105 -1955 5110
rect -1695 5140 -1655 5145
rect -1695 5110 -1690 5140
rect -1690 5110 -1660 5140
rect -1660 5110 -1655 5140
rect -1695 5105 -1655 5110
rect -2995 5090 -2955 5095
rect -2995 5060 -2990 5090
rect -2990 5060 -2960 5090
rect -2960 5060 -2955 5090
rect -2995 5055 -2955 5060
rect -2795 5090 -2755 5095
rect -2795 5060 -2790 5090
rect -2790 5060 -2760 5090
rect -2760 5060 -2755 5090
rect -2795 5055 -2755 5060
rect -2595 5090 -2555 5095
rect -2595 5060 -2590 5090
rect -2590 5060 -2560 5090
rect -2560 5060 -2555 5090
rect -2595 5055 -2555 5060
rect -2395 5090 -2355 5095
rect -2395 5060 -2390 5090
rect -2390 5060 -2360 5090
rect -2360 5060 -2355 5090
rect -2395 5055 -2355 5060
rect -2195 5090 -2155 5095
rect -2195 5060 -2190 5090
rect -2190 5060 -2160 5090
rect -2160 5060 -2155 5090
rect -2195 5055 -2155 5060
rect -1995 5090 -1955 5095
rect -1995 5060 -1990 5090
rect -1990 5060 -1960 5090
rect -1960 5060 -1955 5090
rect -1995 5055 -1955 5060
rect -1695 5090 -1655 5095
rect -1695 5060 -1690 5090
rect -1690 5060 -1660 5090
rect -1660 5060 -1655 5090
rect -1695 5055 -1655 5060
rect -2995 5040 -2955 5045
rect -2995 5010 -2990 5040
rect -2990 5010 -2960 5040
rect -2960 5010 -2955 5040
rect -2995 5005 -2955 5010
rect -2795 5040 -2755 5045
rect -2795 5010 -2790 5040
rect -2790 5010 -2760 5040
rect -2760 5010 -2755 5040
rect -2795 5005 -2755 5010
rect -2595 5040 -2555 5045
rect -2595 5010 -2590 5040
rect -2590 5010 -2560 5040
rect -2560 5010 -2555 5040
rect -2595 5005 -2555 5010
rect -2395 5040 -2355 5045
rect -2395 5010 -2390 5040
rect -2390 5010 -2360 5040
rect -2360 5010 -2355 5040
rect -2395 5005 -2355 5010
rect -2195 5040 -2155 5045
rect -2195 5010 -2190 5040
rect -2190 5010 -2160 5040
rect -2160 5010 -2155 5040
rect -2195 5005 -2155 5010
rect -1995 5040 -1955 5045
rect -1995 5010 -1990 5040
rect -1990 5010 -1960 5040
rect -1960 5010 -1955 5040
rect -1995 5005 -1955 5010
rect -1695 5040 -1655 5045
rect -1695 5010 -1690 5040
rect -1690 5010 -1660 5040
rect -1660 5010 -1655 5040
rect -1695 5005 -1655 5010
rect -3395 4805 -3355 4845
rect 39805 4740 39845 4745
rect 39805 4710 39810 4740
rect 39810 4710 39840 4740
rect 39840 4710 39845 4740
rect 39805 4705 39845 4710
rect 39905 4640 39945 4645
rect 39905 4610 39910 4640
rect 39910 4610 39940 4640
rect 39940 4610 39945 4640
rect 39905 4605 39945 4610
rect 39955 4640 39995 4645
rect 39955 4610 39960 4640
rect 39960 4610 39990 4640
rect 39990 4610 39995 4640
rect 39955 4605 39995 4610
rect 40005 4640 40045 4645
rect 40005 4610 40010 4640
rect 40010 4610 40040 4640
rect 40040 4610 40045 4640
rect 40005 4605 40045 4610
rect 40055 4640 40095 4645
rect 40055 4610 40060 4640
rect 40060 4610 40090 4640
rect 40090 4610 40095 4640
rect 40055 4605 40095 4610
rect 40105 4640 40145 4645
rect 40105 4610 40110 4640
rect 40110 4610 40140 4640
rect 40140 4610 40145 4640
rect 40105 4605 40145 4610
rect 40155 4640 40195 4645
rect 40155 4610 40160 4640
rect 40160 4610 40190 4640
rect 40190 4610 40195 4640
rect 40155 4605 40195 4610
rect 40205 4640 40245 4645
rect 40205 4610 40210 4640
rect 40210 4610 40240 4640
rect 40240 4610 40245 4640
rect 40205 4605 40245 4610
rect 40255 4640 40295 4645
rect 40255 4610 40260 4640
rect 40260 4610 40290 4640
rect 40290 4610 40295 4640
rect 40255 4605 40295 4610
rect 40305 4640 40345 4645
rect 40305 4610 40310 4640
rect 40310 4610 40340 4640
rect 40340 4610 40345 4640
rect 40305 4605 40345 4610
rect 40355 4640 40395 4645
rect 40355 4610 40360 4640
rect 40360 4610 40390 4640
rect 40390 4610 40395 4640
rect 40355 4605 40395 4610
rect 40405 4640 40445 4645
rect 40405 4610 40410 4640
rect 40410 4610 40440 4640
rect 40440 4610 40445 4640
rect 40405 4605 40445 4610
rect 40455 4640 40495 4645
rect 40455 4610 40460 4640
rect 40460 4610 40490 4640
rect 40490 4610 40495 4640
rect 40455 4605 40495 4610
rect 40505 4640 40545 4645
rect 40505 4610 40510 4640
rect 40510 4610 40540 4640
rect 40540 4610 40545 4640
rect 40505 4605 40545 4610
rect 40555 4640 40595 4645
rect 40555 4610 40560 4640
rect 40560 4610 40590 4640
rect 40590 4610 40595 4640
rect 40555 4605 40595 4610
rect 40605 4640 40645 4645
rect 40605 4610 40610 4640
rect 40610 4610 40640 4640
rect 40640 4610 40645 4640
rect 40605 4605 40645 4610
rect 40655 4640 40695 4645
rect 40655 4610 40660 4640
rect 40660 4610 40690 4640
rect 40690 4610 40695 4640
rect 40655 4605 40695 4610
rect 40705 4640 40745 4645
rect 40705 4610 40710 4640
rect 40710 4610 40740 4640
rect 40740 4610 40745 4640
rect 40705 4605 40745 4610
rect 40755 4640 40795 4645
rect 40755 4610 40760 4640
rect 40760 4610 40790 4640
rect 40790 4610 40795 4640
rect 40755 4605 40795 4610
rect 40805 4640 40845 4645
rect 40805 4610 40810 4640
rect 40810 4610 40840 4640
rect 40840 4610 40845 4640
rect 40805 4605 40845 4610
rect 40855 4640 40895 4645
rect 40855 4610 40860 4640
rect 40860 4610 40890 4640
rect 40890 4610 40895 4640
rect 40855 4605 40895 4610
rect 39905 4590 39945 4595
rect 39905 4560 39910 4590
rect 39910 4560 39940 4590
rect 39940 4560 39945 4590
rect 39905 4555 39945 4560
rect 39955 4590 39995 4595
rect 39955 4560 39960 4590
rect 39960 4560 39990 4590
rect 39990 4560 39995 4590
rect 39955 4555 39995 4560
rect 40005 4590 40045 4595
rect 40005 4560 40010 4590
rect 40010 4560 40040 4590
rect 40040 4560 40045 4590
rect 40005 4555 40045 4560
rect 40055 4590 40095 4595
rect 40055 4560 40060 4590
rect 40060 4560 40090 4590
rect 40090 4560 40095 4590
rect 40055 4555 40095 4560
rect 40105 4590 40145 4595
rect 40105 4560 40110 4590
rect 40110 4560 40140 4590
rect 40140 4560 40145 4590
rect 40105 4555 40145 4560
rect 40155 4590 40195 4595
rect 40155 4560 40160 4590
rect 40160 4560 40190 4590
rect 40190 4560 40195 4590
rect 40155 4555 40195 4560
rect 40205 4590 40245 4595
rect 40205 4560 40210 4590
rect 40210 4560 40240 4590
rect 40240 4560 40245 4590
rect 40205 4555 40245 4560
rect 40255 4590 40295 4595
rect 40255 4560 40260 4590
rect 40260 4560 40290 4590
rect 40290 4560 40295 4590
rect 40255 4555 40295 4560
rect 40305 4590 40345 4595
rect 40305 4560 40310 4590
rect 40310 4560 40340 4590
rect 40340 4560 40345 4590
rect 40305 4555 40345 4560
rect 40355 4590 40395 4595
rect 40355 4560 40360 4590
rect 40360 4560 40390 4590
rect 40390 4560 40395 4590
rect 40355 4555 40395 4560
rect 40405 4590 40445 4595
rect 40405 4560 40410 4590
rect 40410 4560 40440 4590
rect 40440 4560 40445 4590
rect 40405 4555 40445 4560
rect 40455 4590 40495 4595
rect 40455 4560 40460 4590
rect 40460 4560 40490 4590
rect 40490 4560 40495 4590
rect 40455 4555 40495 4560
rect 40505 4590 40545 4595
rect 40505 4560 40510 4590
rect 40510 4560 40540 4590
rect 40540 4560 40545 4590
rect 40505 4555 40545 4560
rect 40555 4590 40595 4595
rect 40555 4560 40560 4590
rect 40560 4560 40590 4590
rect 40590 4560 40595 4590
rect 40555 4555 40595 4560
rect 40605 4590 40645 4595
rect 40605 4560 40610 4590
rect 40610 4560 40640 4590
rect 40640 4560 40645 4590
rect 40605 4555 40645 4560
rect 40655 4590 40695 4595
rect 40655 4560 40660 4590
rect 40660 4560 40690 4590
rect 40690 4560 40695 4590
rect 40655 4555 40695 4560
rect 40705 4590 40745 4595
rect 40705 4560 40710 4590
rect 40710 4560 40740 4590
rect 40740 4560 40745 4590
rect 40705 4555 40745 4560
rect 40755 4590 40795 4595
rect 40755 4560 40760 4590
rect 40760 4560 40790 4590
rect 40790 4560 40795 4590
rect 40755 4555 40795 4560
rect 40805 4590 40845 4595
rect 40805 4560 40810 4590
rect 40810 4560 40840 4590
rect 40840 4560 40845 4590
rect 40805 4555 40845 4560
rect 40855 4590 40895 4595
rect 40855 4560 40860 4590
rect 40860 4560 40890 4590
rect 40890 4560 40895 4590
rect 40855 4555 40895 4560
rect 39905 4540 39945 4545
rect 39905 4510 39910 4540
rect 39910 4510 39940 4540
rect 39940 4510 39945 4540
rect 39905 4505 39945 4510
rect 39955 4540 39995 4545
rect 39955 4510 39960 4540
rect 39960 4510 39990 4540
rect 39990 4510 39995 4540
rect 39955 4505 39995 4510
rect 40005 4540 40045 4545
rect 40005 4510 40010 4540
rect 40010 4510 40040 4540
rect 40040 4510 40045 4540
rect 40005 4505 40045 4510
rect 40055 4540 40095 4545
rect 40055 4510 40060 4540
rect 40060 4510 40090 4540
rect 40090 4510 40095 4540
rect 40055 4505 40095 4510
rect 40105 4540 40145 4545
rect 40105 4510 40110 4540
rect 40110 4510 40140 4540
rect 40140 4510 40145 4540
rect 40105 4505 40145 4510
rect 40155 4540 40195 4545
rect 40155 4510 40160 4540
rect 40160 4510 40190 4540
rect 40190 4510 40195 4540
rect 40155 4505 40195 4510
rect 40205 4540 40245 4545
rect 40205 4510 40210 4540
rect 40210 4510 40240 4540
rect 40240 4510 40245 4540
rect 40205 4505 40245 4510
rect 40255 4540 40295 4545
rect 40255 4510 40260 4540
rect 40260 4510 40290 4540
rect 40290 4510 40295 4540
rect 40255 4505 40295 4510
rect 40305 4540 40345 4545
rect 40305 4510 40310 4540
rect 40310 4510 40340 4540
rect 40340 4510 40345 4540
rect 40305 4505 40345 4510
rect 40355 4540 40395 4545
rect 40355 4510 40360 4540
rect 40360 4510 40390 4540
rect 40390 4510 40395 4540
rect 40355 4505 40395 4510
rect 40405 4540 40445 4545
rect 40405 4510 40410 4540
rect 40410 4510 40440 4540
rect 40440 4510 40445 4540
rect 40405 4505 40445 4510
rect 40455 4540 40495 4545
rect 40455 4510 40460 4540
rect 40460 4510 40490 4540
rect 40490 4510 40495 4540
rect 40455 4505 40495 4510
rect 40505 4540 40545 4545
rect 40505 4510 40510 4540
rect 40510 4510 40540 4540
rect 40540 4510 40545 4540
rect 40505 4505 40545 4510
rect 40555 4540 40595 4545
rect 40555 4510 40560 4540
rect 40560 4510 40590 4540
rect 40590 4510 40595 4540
rect 40555 4505 40595 4510
rect 40605 4540 40645 4545
rect 40605 4510 40610 4540
rect 40610 4510 40640 4540
rect 40640 4510 40645 4540
rect 40605 4505 40645 4510
rect 40655 4540 40695 4545
rect 40655 4510 40660 4540
rect 40660 4510 40690 4540
rect 40690 4510 40695 4540
rect 40655 4505 40695 4510
rect 40705 4540 40745 4545
rect 40705 4510 40710 4540
rect 40710 4510 40740 4540
rect 40740 4510 40745 4540
rect 40705 4505 40745 4510
rect 40755 4540 40795 4545
rect 40755 4510 40760 4540
rect 40760 4510 40790 4540
rect 40790 4510 40795 4540
rect 40755 4505 40795 4510
rect 40805 4540 40845 4545
rect 40805 4510 40810 4540
rect 40810 4510 40840 4540
rect 40840 4510 40845 4540
rect 40805 4505 40845 4510
rect 40855 4540 40895 4545
rect 40855 4510 40860 4540
rect 40860 4510 40890 4540
rect 40890 4510 40895 4540
rect 40855 4505 40895 4510
rect 39905 4490 39945 4495
rect 39905 4460 39910 4490
rect 39910 4460 39940 4490
rect 39940 4460 39945 4490
rect 39905 4455 39945 4460
rect 39955 4490 39995 4495
rect 39955 4460 39960 4490
rect 39960 4460 39990 4490
rect 39990 4460 39995 4490
rect 39955 4455 39995 4460
rect 40005 4490 40045 4495
rect 40005 4460 40010 4490
rect 40010 4460 40040 4490
rect 40040 4460 40045 4490
rect 40005 4455 40045 4460
rect 40055 4490 40095 4495
rect 40055 4460 40060 4490
rect 40060 4460 40090 4490
rect 40090 4460 40095 4490
rect 40055 4455 40095 4460
rect 40105 4490 40145 4495
rect 40105 4460 40110 4490
rect 40110 4460 40140 4490
rect 40140 4460 40145 4490
rect 40105 4455 40145 4460
rect 40155 4490 40195 4495
rect 40155 4460 40160 4490
rect 40160 4460 40190 4490
rect 40190 4460 40195 4490
rect 40155 4455 40195 4460
rect 40205 4490 40245 4495
rect 40205 4460 40210 4490
rect 40210 4460 40240 4490
rect 40240 4460 40245 4490
rect 40205 4455 40245 4460
rect 40255 4490 40295 4495
rect 40255 4460 40260 4490
rect 40260 4460 40290 4490
rect 40290 4460 40295 4490
rect 40255 4455 40295 4460
rect 40305 4490 40345 4495
rect 40305 4460 40310 4490
rect 40310 4460 40340 4490
rect 40340 4460 40345 4490
rect 40305 4455 40345 4460
rect 40355 4490 40395 4495
rect 40355 4460 40360 4490
rect 40360 4460 40390 4490
rect 40390 4460 40395 4490
rect 40355 4455 40395 4460
rect 40405 4490 40445 4495
rect 40405 4460 40410 4490
rect 40410 4460 40440 4490
rect 40440 4460 40445 4490
rect 40405 4455 40445 4460
rect 40455 4490 40495 4495
rect 40455 4460 40460 4490
rect 40460 4460 40490 4490
rect 40490 4460 40495 4490
rect 40455 4455 40495 4460
rect 40505 4490 40545 4495
rect 40505 4460 40510 4490
rect 40510 4460 40540 4490
rect 40540 4460 40545 4490
rect 40505 4455 40545 4460
rect 40555 4490 40595 4495
rect 40555 4460 40560 4490
rect 40560 4460 40590 4490
rect 40590 4460 40595 4490
rect 40555 4455 40595 4460
rect 40605 4490 40645 4495
rect 40605 4460 40610 4490
rect 40610 4460 40640 4490
rect 40640 4460 40645 4490
rect 40605 4455 40645 4460
rect 40655 4490 40695 4495
rect 40655 4460 40660 4490
rect 40660 4460 40690 4490
rect 40690 4460 40695 4490
rect 40655 4455 40695 4460
rect 40705 4490 40745 4495
rect 40705 4460 40710 4490
rect 40710 4460 40740 4490
rect 40740 4460 40745 4490
rect 40705 4455 40745 4460
rect 40755 4490 40795 4495
rect 40755 4460 40760 4490
rect 40760 4460 40790 4490
rect 40790 4460 40795 4490
rect 40755 4455 40795 4460
rect 40805 4490 40845 4495
rect 40805 4460 40810 4490
rect 40810 4460 40840 4490
rect 40840 4460 40845 4490
rect 40805 4455 40845 4460
rect 40855 4490 40895 4495
rect 40855 4460 40860 4490
rect 40860 4460 40890 4490
rect 40890 4460 40895 4490
rect 40855 4455 40895 4460
rect 39905 4440 39945 4445
rect 39905 4410 39910 4440
rect 39910 4410 39940 4440
rect 39940 4410 39945 4440
rect 39905 4405 39945 4410
rect 39955 4440 39995 4445
rect 39955 4410 39960 4440
rect 39960 4410 39990 4440
rect 39990 4410 39995 4440
rect 39955 4405 39995 4410
rect 40005 4440 40045 4445
rect 40005 4410 40010 4440
rect 40010 4410 40040 4440
rect 40040 4410 40045 4440
rect 40005 4405 40045 4410
rect 40055 4440 40095 4445
rect 40055 4410 40060 4440
rect 40060 4410 40090 4440
rect 40090 4410 40095 4440
rect 40055 4405 40095 4410
rect 40105 4440 40145 4445
rect 40105 4410 40110 4440
rect 40110 4410 40140 4440
rect 40140 4410 40145 4440
rect 40105 4405 40145 4410
rect 40155 4440 40195 4445
rect 40155 4410 40160 4440
rect 40160 4410 40190 4440
rect 40190 4410 40195 4440
rect 40155 4405 40195 4410
rect 40205 4440 40245 4445
rect 40205 4410 40210 4440
rect 40210 4410 40240 4440
rect 40240 4410 40245 4440
rect 40205 4405 40245 4410
rect 40255 4440 40295 4445
rect 40255 4410 40260 4440
rect 40260 4410 40290 4440
rect 40290 4410 40295 4440
rect 40255 4405 40295 4410
rect 40305 4440 40345 4445
rect 40305 4410 40310 4440
rect 40310 4410 40340 4440
rect 40340 4410 40345 4440
rect 40305 4405 40345 4410
rect 40355 4440 40395 4445
rect 40355 4410 40360 4440
rect 40360 4410 40390 4440
rect 40390 4410 40395 4440
rect 40355 4405 40395 4410
rect 40405 4440 40445 4445
rect 40405 4410 40410 4440
rect 40410 4410 40440 4440
rect 40440 4410 40445 4440
rect 40405 4405 40445 4410
rect 40455 4440 40495 4445
rect 40455 4410 40460 4440
rect 40460 4410 40490 4440
rect 40490 4410 40495 4440
rect 40455 4405 40495 4410
rect 40505 4440 40545 4445
rect 40505 4410 40510 4440
rect 40510 4410 40540 4440
rect 40540 4410 40545 4440
rect 40505 4405 40545 4410
rect 40555 4440 40595 4445
rect 40555 4410 40560 4440
rect 40560 4410 40590 4440
rect 40590 4410 40595 4440
rect 40555 4405 40595 4410
rect 40605 4440 40645 4445
rect 40605 4410 40610 4440
rect 40610 4410 40640 4440
rect 40640 4410 40645 4440
rect 40605 4405 40645 4410
rect 40655 4440 40695 4445
rect 40655 4410 40660 4440
rect 40660 4410 40690 4440
rect 40690 4410 40695 4440
rect 40655 4405 40695 4410
rect 40705 4440 40745 4445
rect 40705 4410 40710 4440
rect 40710 4410 40740 4440
rect 40740 4410 40745 4440
rect 40705 4405 40745 4410
rect 40755 4440 40795 4445
rect 40755 4410 40760 4440
rect 40760 4410 40790 4440
rect 40790 4410 40795 4440
rect 40755 4405 40795 4410
rect 40805 4440 40845 4445
rect 40805 4410 40810 4440
rect 40810 4410 40840 4440
rect 40840 4410 40845 4440
rect 40805 4405 40845 4410
rect 40855 4440 40895 4445
rect 40855 4410 40860 4440
rect 40860 4410 40890 4440
rect 40890 4410 40895 4440
rect 40855 4405 40895 4410
rect 39805 4340 39845 4345
rect 39805 4310 39810 4340
rect 39810 4310 39840 4340
rect 39840 4310 39845 4340
rect 39805 4305 39845 4310
rect -3195 4205 -3155 4245
rect -3495 3840 -3455 3845
rect -3495 3810 -3490 3840
rect -3490 3810 -3460 3840
rect -3460 3810 -3455 3840
rect -3495 3805 -3455 3810
rect -3295 3840 -3255 3845
rect -3295 3810 -3290 3840
rect -3290 3810 -3260 3840
rect -3260 3810 -3255 3840
rect -3295 3805 -3255 3810
rect -3095 3840 -3055 3845
rect -3095 3810 -3090 3840
rect -3090 3810 -3060 3840
rect -3060 3810 -3055 3840
rect -3095 3805 -3055 3810
rect -1595 3840 -1555 3845
rect -1595 3810 -1590 3840
rect -1590 3810 -1560 3840
rect -1560 3810 -1555 3840
rect -1595 3805 -1555 3810
rect -1095 3840 -1055 3845
rect -1095 3810 -1090 3840
rect -1090 3810 -1060 3840
rect -1060 3810 -1055 3840
rect -1095 3805 -1055 3810
rect -895 3840 -855 3845
rect -895 3810 -890 3840
rect -890 3810 -860 3840
rect -860 3810 -855 3840
rect -895 3805 -855 3810
rect -695 3840 -655 3845
rect -695 3810 -690 3840
rect -690 3810 -660 3840
rect -660 3810 -655 3840
rect -695 3805 -655 3810
rect -495 3840 -455 3845
rect -495 3810 -490 3840
rect -490 3810 -460 3840
rect -460 3810 -455 3840
rect -495 3805 -455 3810
rect -295 3840 -255 3845
rect -295 3810 -290 3840
rect -290 3810 -260 3840
rect -260 3810 -255 3840
rect -295 3805 -255 3810
rect -95 3840 -55 3845
rect -95 3810 -90 3840
rect -90 3810 -60 3840
rect -60 3810 -55 3840
rect -95 3805 -55 3810
rect -3495 3790 -3455 3795
rect -3495 3760 -3490 3790
rect -3490 3760 -3460 3790
rect -3460 3760 -3455 3790
rect -3495 3755 -3455 3760
rect -3295 3790 -3255 3795
rect -3295 3760 -3290 3790
rect -3290 3760 -3260 3790
rect -3260 3760 -3255 3790
rect -3295 3755 -3255 3760
rect -3095 3790 -3055 3795
rect -3095 3760 -3090 3790
rect -3090 3760 -3060 3790
rect -3060 3760 -3055 3790
rect -3095 3755 -3055 3760
rect -1595 3790 -1555 3795
rect -1595 3760 -1590 3790
rect -1590 3760 -1560 3790
rect -1560 3760 -1555 3790
rect -1595 3755 -1555 3760
rect -1095 3790 -1055 3795
rect -1095 3760 -1090 3790
rect -1090 3760 -1060 3790
rect -1060 3760 -1055 3790
rect -1095 3755 -1055 3760
rect -895 3790 -855 3795
rect -895 3760 -890 3790
rect -890 3760 -860 3790
rect -860 3760 -855 3790
rect -895 3755 -855 3760
rect -695 3790 -655 3795
rect -695 3760 -690 3790
rect -690 3760 -660 3790
rect -660 3760 -655 3790
rect -695 3755 -655 3760
rect -495 3790 -455 3795
rect -495 3760 -490 3790
rect -490 3760 -460 3790
rect -460 3760 -455 3790
rect -495 3755 -455 3760
rect -295 3790 -255 3795
rect -295 3760 -290 3790
rect -290 3760 -260 3790
rect -260 3760 -255 3790
rect -295 3755 -255 3760
rect -95 3790 -55 3795
rect -95 3760 -90 3790
rect -90 3760 -60 3790
rect -60 3760 -55 3790
rect -95 3755 -55 3760
rect -3495 3740 -3455 3745
rect -3495 3710 -3490 3740
rect -3490 3710 -3460 3740
rect -3460 3710 -3455 3740
rect -3495 3705 -3455 3710
rect -3295 3740 -3255 3745
rect -3295 3710 -3290 3740
rect -3290 3710 -3260 3740
rect -3260 3710 -3255 3740
rect -3295 3705 -3255 3710
rect -3095 3740 -3055 3745
rect -3095 3710 -3090 3740
rect -3090 3710 -3060 3740
rect -3060 3710 -3055 3740
rect -3095 3705 -3055 3710
rect -1595 3740 -1555 3745
rect -1595 3710 -1590 3740
rect -1590 3710 -1560 3740
rect -1560 3710 -1555 3740
rect -1595 3705 -1555 3710
rect -1095 3740 -1055 3745
rect -1095 3710 -1090 3740
rect -1090 3710 -1060 3740
rect -1060 3710 -1055 3740
rect -1095 3705 -1055 3710
rect -895 3740 -855 3745
rect -895 3710 -890 3740
rect -890 3710 -860 3740
rect -860 3710 -855 3740
rect -895 3705 -855 3710
rect -695 3740 -655 3745
rect -695 3710 -690 3740
rect -690 3710 -660 3740
rect -660 3710 -655 3740
rect -695 3705 -655 3710
rect -495 3740 -455 3745
rect -495 3710 -490 3740
rect -490 3710 -460 3740
rect -460 3710 -455 3740
rect -495 3705 -455 3710
rect -295 3740 -255 3745
rect -295 3710 -290 3740
rect -290 3710 -260 3740
rect -260 3710 -255 3740
rect -295 3705 -255 3710
rect -95 3740 -55 3745
rect -95 3710 -90 3740
rect -90 3710 -60 3740
rect -60 3710 -55 3740
rect -95 3705 -55 3710
rect -1495 3405 -1455 3445
rect -1395 3305 -1355 3345
rect -1295 3205 -1255 3245
rect -1195 3105 -1155 3145
rect -995 2705 -955 2745
rect -795 2505 -755 2545
rect -3495 2140 -3455 2145
rect -3495 2110 -3490 2140
rect -3490 2110 -3460 2140
rect -3460 2110 -3455 2140
rect -3495 2105 -3455 2110
rect -3295 2140 -3255 2145
rect -3295 2110 -3290 2140
rect -3290 2110 -3260 2140
rect -3260 2110 -3255 2140
rect -3295 2105 -3255 2110
rect -3095 2140 -3055 2145
rect -3095 2110 -3090 2140
rect -3090 2110 -3060 2140
rect -3060 2110 -3055 2140
rect -3095 2105 -3055 2110
rect -1595 2140 -1555 2145
rect -1595 2110 -1590 2140
rect -1590 2110 -1560 2140
rect -1560 2110 -1555 2140
rect -1595 2105 -1555 2110
rect -1095 2140 -1055 2145
rect -1095 2110 -1090 2140
rect -1090 2110 -1060 2140
rect -1060 2110 -1055 2140
rect -1095 2105 -1055 2110
rect -895 2140 -855 2145
rect -895 2110 -890 2140
rect -890 2110 -860 2140
rect -860 2110 -855 2140
rect -895 2105 -855 2110
rect -695 2140 -655 2145
rect -695 2110 -690 2140
rect -690 2110 -660 2140
rect -660 2110 -655 2140
rect -695 2105 -655 2110
rect -495 2140 -455 2145
rect -495 2110 -490 2140
rect -490 2110 -460 2140
rect -460 2110 -455 2140
rect -495 2105 -455 2110
rect -295 2140 -255 2145
rect -295 2110 -290 2140
rect -290 2110 -260 2140
rect -260 2110 -255 2140
rect -295 2105 -255 2110
rect -95 2140 -55 2145
rect -95 2110 -90 2140
rect -90 2110 -60 2140
rect -60 2110 -55 2140
rect -95 2105 -55 2110
rect -3495 2090 -3455 2095
rect -3495 2060 -3490 2090
rect -3490 2060 -3460 2090
rect -3460 2060 -3455 2090
rect -3495 2055 -3455 2060
rect -3295 2090 -3255 2095
rect -3295 2060 -3290 2090
rect -3290 2060 -3260 2090
rect -3260 2060 -3255 2090
rect -3295 2055 -3255 2060
rect -3095 2090 -3055 2095
rect -3095 2060 -3090 2090
rect -3090 2060 -3060 2090
rect -3060 2060 -3055 2090
rect -3095 2055 -3055 2060
rect -1595 2090 -1555 2095
rect -1595 2060 -1590 2090
rect -1590 2060 -1560 2090
rect -1560 2060 -1555 2090
rect -1595 2055 -1555 2060
rect -1095 2090 -1055 2095
rect -1095 2060 -1090 2090
rect -1090 2060 -1060 2090
rect -1060 2060 -1055 2090
rect -1095 2055 -1055 2060
rect -895 2090 -855 2095
rect -895 2060 -890 2090
rect -890 2060 -860 2090
rect -860 2060 -855 2090
rect -895 2055 -855 2060
rect -695 2090 -655 2095
rect -695 2060 -690 2090
rect -690 2060 -660 2090
rect -660 2060 -655 2090
rect -695 2055 -655 2060
rect -495 2090 -455 2095
rect -495 2060 -490 2090
rect -490 2060 -460 2090
rect -460 2060 -455 2090
rect -495 2055 -455 2060
rect -295 2090 -255 2095
rect -295 2060 -290 2090
rect -290 2060 -260 2090
rect -260 2060 -255 2090
rect -295 2055 -255 2060
rect -95 2090 -55 2095
rect -95 2060 -90 2090
rect -90 2060 -60 2090
rect -60 2060 -55 2090
rect -95 2055 -55 2060
rect -3495 2040 -3455 2045
rect -3495 2010 -3490 2040
rect -3490 2010 -3460 2040
rect -3460 2010 -3455 2040
rect -3495 2005 -3455 2010
rect -3295 2040 -3255 2045
rect -3295 2010 -3290 2040
rect -3290 2010 -3260 2040
rect -3260 2010 -3255 2040
rect -3295 2005 -3255 2010
rect -3095 2040 -3055 2045
rect -3095 2010 -3090 2040
rect -3090 2010 -3060 2040
rect -3060 2010 -3055 2040
rect -3095 2005 -3055 2010
rect -1595 2040 -1555 2045
rect -1595 2010 -1590 2040
rect -1590 2010 -1560 2040
rect -1560 2010 -1555 2040
rect -1595 2005 -1555 2010
rect -1095 2040 -1055 2045
rect -1095 2010 -1090 2040
rect -1090 2010 -1060 2040
rect -1060 2010 -1055 2040
rect -1095 2005 -1055 2010
rect -895 2040 -855 2045
rect -895 2010 -890 2040
rect -890 2010 -860 2040
rect -860 2010 -855 2040
rect -895 2005 -855 2010
rect -695 2040 -655 2045
rect -695 2010 -690 2040
rect -690 2010 -660 2040
rect -660 2010 -655 2040
rect -695 2005 -655 2010
rect -495 2040 -455 2045
rect -495 2010 -490 2040
rect -490 2010 -460 2040
rect -460 2010 -455 2040
rect -495 2005 -455 2010
rect -295 2040 -255 2045
rect -295 2010 -290 2040
rect -290 2010 -260 2040
rect -260 2010 -255 2040
rect -295 2005 -255 2010
rect -95 2040 -55 2045
rect -95 2010 -90 2040
rect -90 2010 -60 2040
rect -60 2010 -55 2040
rect -95 2005 -55 2010
rect -595 1605 -555 1645
rect -395 1405 -355 1445
rect -195 1005 -155 1045
rect -3495 440 -3455 445
rect -3495 410 -3490 440
rect -3490 410 -3460 440
rect -3460 410 -3455 440
rect -3495 405 -3455 410
rect -3295 440 -3255 445
rect -3295 410 -3290 440
rect -3290 410 -3260 440
rect -3260 410 -3255 440
rect -3295 405 -3255 410
rect -3095 440 -3055 445
rect -3095 410 -3090 440
rect -3090 410 -3060 440
rect -3060 410 -3055 440
rect -3095 405 -3055 410
rect -1595 440 -1555 445
rect -1595 410 -1590 440
rect -1590 410 -1560 440
rect -1560 410 -1555 440
rect -1595 405 -1555 410
rect -1095 440 -1055 445
rect -1095 410 -1090 440
rect -1090 410 -1060 440
rect -1060 410 -1055 440
rect -1095 405 -1055 410
rect -895 440 -855 445
rect -895 410 -890 440
rect -890 410 -860 440
rect -860 410 -855 440
rect -895 405 -855 410
rect -695 440 -655 445
rect -695 410 -690 440
rect -690 410 -660 440
rect -660 410 -655 440
rect -695 405 -655 410
rect -495 440 -455 445
rect -495 410 -490 440
rect -490 410 -460 440
rect -460 410 -455 440
rect -495 405 -455 410
rect -295 440 -255 445
rect -295 410 -290 440
rect -290 410 -260 440
rect -260 410 -255 440
rect -295 405 -255 410
rect -95 440 -55 445
rect -95 410 -90 440
rect -90 410 -60 440
rect -60 410 -55 440
rect -95 405 -55 410
rect -3495 390 -3455 395
rect -3495 360 -3490 390
rect -3490 360 -3460 390
rect -3460 360 -3455 390
rect -3495 355 -3455 360
rect -3295 390 -3255 395
rect -3295 360 -3290 390
rect -3290 360 -3260 390
rect -3260 360 -3255 390
rect -3295 355 -3255 360
rect -3095 390 -3055 395
rect -3095 360 -3090 390
rect -3090 360 -3060 390
rect -3060 360 -3055 390
rect -3095 355 -3055 360
rect -1595 390 -1555 395
rect -1595 360 -1590 390
rect -1590 360 -1560 390
rect -1560 360 -1555 390
rect -1595 355 -1555 360
rect -1095 390 -1055 395
rect -1095 360 -1090 390
rect -1090 360 -1060 390
rect -1060 360 -1055 390
rect -1095 355 -1055 360
rect -895 390 -855 395
rect -895 360 -890 390
rect -890 360 -860 390
rect -860 360 -855 390
rect -895 355 -855 360
rect -695 390 -655 395
rect -695 360 -690 390
rect -690 360 -660 390
rect -660 360 -655 390
rect -695 355 -655 360
rect -495 390 -455 395
rect -495 360 -490 390
rect -490 360 -460 390
rect -460 360 -455 390
rect -495 355 -455 360
rect -295 390 -255 395
rect -295 360 -290 390
rect -290 360 -260 390
rect -260 360 -255 390
rect -295 355 -255 360
rect -95 390 -55 395
rect -95 360 -90 390
rect -90 360 -60 390
rect -60 360 -55 390
rect -95 355 -55 360
rect -3495 340 -3455 345
rect -3495 310 -3490 340
rect -3490 310 -3460 340
rect -3460 310 -3455 340
rect -3495 305 -3455 310
rect -3295 340 -3255 345
rect -3295 310 -3290 340
rect -3290 310 -3260 340
rect -3260 310 -3255 340
rect -3295 305 -3255 310
rect -3095 340 -3055 345
rect -3095 310 -3090 340
rect -3090 310 -3060 340
rect -3060 310 -3055 340
rect -3095 305 -3055 310
rect -1595 340 -1555 345
rect -1595 310 -1590 340
rect -1590 310 -1560 340
rect -1560 310 -1555 340
rect -1595 305 -1555 310
rect -1095 340 -1055 345
rect -1095 310 -1090 340
rect -1090 310 -1060 340
rect -1060 310 -1055 340
rect -1095 305 -1055 310
rect -895 340 -855 345
rect -895 310 -890 340
rect -890 310 -860 340
rect -860 310 -855 340
rect -895 305 -855 310
rect -695 340 -655 345
rect -695 310 -690 340
rect -690 310 -660 340
rect -660 310 -655 340
rect -695 305 -655 310
rect -495 340 -455 345
rect -495 310 -490 340
rect -490 310 -460 340
rect -460 310 -455 340
rect -495 305 -455 310
rect -295 340 -255 345
rect -295 310 -290 340
rect -290 310 -260 340
rect -260 310 -255 340
rect -295 305 -255 310
rect -95 340 -55 345
rect -95 310 -90 340
rect -90 310 -60 340
rect -60 310 -55 340
rect -95 305 -55 310
<< mimcap >>
rect 150 17990 3150 18040
rect 150 17340 200 17990
rect 3100 17340 3150 17990
rect 150 17290 3150 17340
rect 3400 17990 6400 18040
rect 3400 17340 3450 17990
rect 6350 17340 6400 17990
rect 3400 17290 6400 17340
rect 6650 17990 9650 18040
rect 6650 17340 6700 17990
rect 9600 17340 9650 17990
rect 6650 17290 9650 17340
rect 9900 17990 12900 18040
rect 9900 17340 9950 17990
rect 12850 17340 12900 17990
rect 9900 17290 12900 17340
rect 13150 17990 16150 18040
rect 13150 17340 13200 17990
rect 16100 17340 16150 17990
rect 13150 17290 16150 17340
rect 16400 17990 19400 18040
rect 16400 17340 16450 17990
rect 19350 17340 19400 17990
rect 16400 17290 19400 17340
rect 19650 17990 22650 18040
rect 19650 17340 19700 17990
rect 22600 17340 22650 17990
rect 19650 17290 22650 17340
rect 22900 17990 25900 18040
rect 22900 17340 22950 17990
rect 25850 17340 25900 17990
rect 22900 17290 25900 17340
rect 26150 17990 29150 18040
rect 26150 17340 26200 17990
rect 29100 17340 29150 17990
rect 26150 17290 29150 17340
rect 29400 17990 32400 18040
rect 29400 17340 29450 17990
rect 32350 17340 32400 17990
rect 29400 17290 32400 17340
rect 32650 17990 35650 18040
rect 32650 17340 32700 17990
rect 35600 17340 35650 17990
rect 32650 17290 35650 17340
rect 35900 17990 38900 18040
rect 35900 17340 35950 17990
rect 38850 17340 38900 17990
rect 35900 17290 38900 17340
rect 39150 17990 39700 18040
rect 39150 17340 39200 17990
rect 39650 17340 39700 17990
rect 39150 17290 39700 17340
rect 150 16650 3150 16700
rect 150 16000 200 16650
rect 3100 16000 3150 16650
rect 150 15950 3150 16000
rect 3400 16650 6400 16700
rect 3400 16000 3450 16650
rect 6350 16000 6400 16650
rect 3400 15950 6400 16000
rect 6650 16650 9650 16700
rect 6650 16000 6700 16650
rect 9600 16000 9650 16650
rect 6650 15950 9650 16000
rect 9900 16650 12900 16700
rect 9900 16000 9950 16650
rect 12850 16000 12900 16650
rect 9900 15950 12900 16000
rect 13150 16650 16150 16700
rect 13150 16000 13200 16650
rect 16100 16000 16150 16650
rect 13150 15950 16150 16000
rect 16400 16650 19400 16700
rect 16400 16000 16450 16650
rect 19350 16000 19400 16650
rect 16400 15950 19400 16000
rect 19650 16650 22650 16700
rect 19650 16000 19700 16650
rect 22600 16000 22650 16650
rect 19650 15950 22650 16000
rect 22900 16650 25900 16700
rect 22900 16000 22950 16650
rect 25850 16000 25900 16650
rect 22900 15950 25900 16000
rect 26150 16650 29150 16700
rect 26150 16000 26200 16650
rect 29100 16000 29150 16650
rect 26150 15950 29150 16000
rect 29400 16650 32400 16700
rect 29400 16000 29450 16650
rect 32350 16000 32400 16650
rect 29400 15950 32400 16000
rect 32650 16650 35650 16700
rect 32650 16000 32700 16650
rect 35600 16000 35650 16650
rect 32650 15950 35650 16000
rect 35900 16650 38900 16700
rect 35900 16000 35950 16650
rect 38850 16000 38900 16650
rect 35900 15950 38900 16000
rect 39150 16650 39700 16700
rect 39150 16000 39200 16650
rect 39650 16000 39700 16650
rect 39150 15950 39700 16000
<< mimcapcontact >>
rect 200 17340 3100 17990
rect 3450 17340 6350 17990
rect 6700 17340 9600 17990
rect 9950 17340 12850 17990
rect 13200 17340 16100 17990
rect 16450 17340 19350 17990
rect 19700 17340 22600 17990
rect 22950 17340 25850 17990
rect 26200 17340 29100 17990
rect 29450 17340 32350 17990
rect 32700 17340 35600 17990
rect 35950 17340 38850 17990
rect 39200 17340 39650 17990
rect 200 16000 3100 16650
rect 3450 16000 6350 16650
rect 6700 16000 9600 16650
rect 9950 16000 12850 16650
rect 13200 16000 16100 16650
rect 16450 16000 19350 16650
rect 19700 16000 22600 16650
rect 22950 16000 25850 16650
rect 26200 16000 29100 16650
rect 29450 16000 32350 16650
rect 32700 16000 35600 16650
rect 35950 16000 38850 16650
rect 39200 16000 39650 16650
<< metal4 >>
rect -3500 17015 -3450 18290
rect -3500 16975 -3495 17015
rect -3455 16975 -3450 17015
rect -3500 15745 -3450 16975
rect -3500 15705 -3495 15745
rect -3455 15705 -3450 15745
rect -3500 15345 -3450 15705
rect -3500 15305 -3495 15345
rect -3455 15305 -3450 15345
rect -3500 15295 -3450 15305
rect -3500 15255 -3495 15295
rect -3455 15255 -3450 15295
rect -3500 15245 -3450 15255
rect -3500 15205 -3495 15245
rect -3455 15205 -3450 15245
rect -3500 13645 -3450 15205
rect -3500 13605 -3495 13645
rect -3455 13605 -3450 13645
rect -3500 13595 -3450 13605
rect -3500 13555 -3495 13595
rect -3455 13555 -3450 13595
rect -3500 13545 -3450 13555
rect -3500 13505 -3495 13545
rect -3455 13505 -3450 13545
rect -3500 11945 -3450 13505
rect -3500 11905 -3495 11945
rect -3455 11905 -3450 11945
rect -3500 11895 -3450 11905
rect -3500 11855 -3495 11895
rect -3455 11855 -3450 11895
rect -3500 11845 -3450 11855
rect -3500 11805 -3495 11845
rect -3455 11805 -3450 11845
rect -3500 3845 -3450 11805
rect -3500 3805 -3495 3845
rect -3455 3805 -3450 3845
rect -3500 3795 -3450 3805
rect -3500 3755 -3495 3795
rect -3455 3755 -3450 3795
rect -3500 3745 -3450 3755
rect -3500 3705 -3495 3745
rect -3455 3705 -3450 3745
rect -3500 2145 -3450 3705
rect -3500 2105 -3495 2145
rect -3455 2105 -3450 2145
rect -3500 2095 -3450 2105
rect -3500 2055 -3495 2095
rect -3455 2055 -3450 2095
rect -3500 2045 -3450 2055
rect -3500 2005 -3495 2045
rect -3455 2005 -3450 2045
rect -3500 445 -3450 2005
rect -3500 405 -3495 445
rect -3455 405 -3450 445
rect -3500 395 -3450 405
rect -3500 355 -3495 395
rect -3455 355 -3450 395
rect -3500 345 -3450 355
rect -3500 305 -3495 345
rect -3455 305 -3450 345
rect -3500 0 -3450 305
rect -3400 10845 -3350 18290
rect -3400 10805 -3395 10845
rect -3355 10805 -3350 10845
rect -3400 4845 -3350 10805
rect -3400 4805 -3395 4845
rect -3355 4805 -3350 4845
rect -3400 0 -3350 4805
rect -3300 17015 -3250 18290
rect -3300 16975 -3295 17015
rect -3255 16975 -3250 17015
rect -3300 15745 -3250 16975
rect -3300 15705 -3295 15745
rect -3255 15705 -3250 15745
rect -3300 15345 -3250 15705
rect -3300 15305 -3295 15345
rect -3255 15305 -3250 15345
rect -3300 15295 -3250 15305
rect -3300 15255 -3295 15295
rect -3255 15255 -3250 15295
rect -3300 15245 -3250 15255
rect -3300 15205 -3295 15245
rect -3255 15205 -3250 15245
rect -3300 13645 -3250 15205
rect -3300 13605 -3295 13645
rect -3255 13605 -3250 13645
rect -3300 13595 -3250 13605
rect -3300 13555 -3295 13595
rect -3255 13555 -3250 13595
rect -3300 13545 -3250 13555
rect -3300 13505 -3295 13545
rect -3255 13505 -3250 13545
rect -3300 11945 -3250 13505
rect -3300 11905 -3295 11945
rect -3255 11905 -3250 11945
rect -3300 11895 -3250 11905
rect -3300 11855 -3295 11895
rect -3255 11855 -3250 11895
rect -3300 11845 -3250 11855
rect -3300 11805 -3295 11845
rect -3255 11805 -3250 11845
rect -3300 3845 -3250 11805
rect -3300 3805 -3295 3845
rect -3255 3805 -3250 3845
rect -3300 3795 -3250 3805
rect -3300 3755 -3295 3795
rect -3255 3755 -3250 3795
rect -3300 3745 -3250 3755
rect -3300 3705 -3295 3745
rect -3255 3705 -3250 3745
rect -3300 2145 -3250 3705
rect -3300 2105 -3295 2145
rect -3255 2105 -3250 2145
rect -3300 2095 -3250 2105
rect -3300 2055 -3295 2095
rect -3255 2055 -3250 2095
rect -3300 2045 -3250 2055
rect -3300 2005 -3295 2045
rect -3255 2005 -3250 2045
rect -3300 445 -3250 2005
rect -3300 405 -3295 445
rect -3255 405 -3250 445
rect -3300 395 -3250 405
rect -3300 355 -3295 395
rect -3255 355 -3250 395
rect -3300 345 -3250 355
rect -3300 305 -3295 345
rect -3255 305 -3250 345
rect -3300 0 -3250 305
rect -3200 11445 -3150 18290
rect -3200 11405 -3195 11445
rect -3155 11405 -3150 11445
rect -3200 4245 -3150 11405
rect -3200 4205 -3195 4245
rect -3155 4205 -3150 4245
rect -3200 0 -3150 4205
rect -3100 17015 -3050 18290
rect -3100 16975 -3095 17015
rect -3055 16975 -3050 17015
rect -3100 15745 -3050 16975
rect -3100 15705 -3095 15745
rect -3055 15705 -3050 15745
rect -3100 15345 -3050 15705
rect -3100 15305 -3095 15345
rect -3055 15305 -3050 15345
rect -3100 15295 -3050 15305
rect -3100 15255 -3095 15295
rect -3055 15255 -3050 15295
rect -3100 15245 -3050 15255
rect -3100 15205 -3095 15245
rect -3055 15205 -3050 15245
rect -3100 13645 -3050 15205
rect -3100 13605 -3095 13645
rect -3055 13605 -3050 13645
rect -3100 13595 -3050 13605
rect -3100 13555 -3095 13595
rect -3055 13555 -3050 13595
rect -3100 13545 -3050 13555
rect -3100 13505 -3095 13545
rect -3055 13505 -3050 13545
rect -3100 11945 -3050 13505
rect -3100 11905 -3095 11945
rect -3055 11905 -3050 11945
rect -3100 11895 -3050 11905
rect -3100 11855 -3095 11895
rect -3055 11855 -3050 11895
rect -3100 11845 -3050 11855
rect -3100 11805 -3095 11845
rect -3055 11805 -3050 11845
rect -3100 3845 -3050 11805
rect -3100 3805 -3095 3845
rect -3055 3805 -3050 3845
rect -3100 3795 -3050 3805
rect -3100 3755 -3095 3795
rect -3055 3755 -3050 3795
rect -3100 3745 -3050 3755
rect -3100 3705 -3095 3745
rect -3055 3705 -3050 3745
rect -3100 2145 -3050 3705
rect -3100 2105 -3095 2145
rect -3055 2105 -3050 2145
rect -3100 2095 -3050 2105
rect -3100 2055 -3095 2095
rect -3055 2055 -3050 2095
rect -3100 2045 -3050 2055
rect -3100 2005 -3095 2045
rect -3055 2005 -3050 2045
rect -3100 445 -3050 2005
rect -3100 405 -3095 445
rect -3055 405 -3050 445
rect -3100 395 -3050 405
rect -3100 355 -3095 395
rect -3055 355 -3050 395
rect -3100 345 -3050 355
rect -3100 305 -3095 345
rect -3055 305 -3050 345
rect -3100 0 -3050 305
rect -3000 18240 -1650 18290
rect -3000 17290 -2950 18240
rect -2900 17290 -2850 18240
rect -2800 17290 -2750 18240
rect -2700 17290 -2650 18240
rect -2600 17290 -2550 18240
rect -2500 17290 -2450 18240
rect -2400 17290 -2350 18240
rect -2300 17290 -2250 18240
rect -2200 17290 -2150 18240
rect -2100 17290 -2050 18240
rect -2000 17290 -1950 18240
rect -1900 17290 -1850 18240
rect -1800 17290 -1750 18240
rect -1700 17290 -1650 18240
rect -3000 17240 -1650 17290
rect -3000 15750 -2950 17240
rect -2900 15750 -2850 17240
rect -2800 15750 -2750 17240
rect -3000 15700 -2750 15750
rect -3000 10645 -2950 15700
rect -3000 10605 -2995 10645
rect -2955 10605 -2950 10645
rect -3000 10595 -2950 10605
rect -3000 10555 -2995 10595
rect -2955 10555 -2950 10595
rect -3000 10545 -2950 10555
rect -3000 10505 -2995 10545
rect -2955 10505 -2950 10545
rect -3000 9345 -2950 10505
rect -3000 9305 -2995 9345
rect -2955 9305 -2950 9345
rect -3000 9295 -2950 9305
rect -3000 9255 -2995 9295
rect -2955 9255 -2950 9295
rect -3000 9245 -2950 9255
rect -3000 9205 -2995 9245
rect -2955 9205 -2950 9245
rect -3000 8045 -2950 9205
rect -3000 8005 -2995 8045
rect -2955 8005 -2950 8045
rect -3000 7995 -2950 8005
rect -3000 7955 -2995 7995
rect -2955 7955 -2950 7995
rect -3000 7945 -2950 7955
rect -3000 7905 -2995 7945
rect -2955 7905 -2950 7945
rect -3000 7745 -2950 7905
rect -3000 7705 -2995 7745
rect -2955 7705 -2950 7745
rect -3000 7695 -2950 7705
rect -3000 7655 -2995 7695
rect -2955 7655 -2950 7695
rect -3000 7645 -2950 7655
rect -3000 7605 -2995 7645
rect -2955 7605 -2950 7645
rect -3000 6445 -2950 7605
rect -3000 6405 -2995 6445
rect -2955 6405 -2950 6445
rect -3000 6395 -2950 6405
rect -3000 6355 -2995 6395
rect -2955 6355 -2950 6395
rect -3000 6345 -2950 6355
rect -3000 6305 -2995 6345
rect -2955 6305 -2950 6345
rect -3000 5145 -2950 6305
rect -3000 5105 -2995 5145
rect -2955 5105 -2950 5145
rect -3000 5095 -2950 5105
rect -3000 5055 -2995 5095
rect -2955 5055 -2950 5095
rect -3000 5045 -2950 5055
rect -3000 5005 -2995 5045
rect -2955 5005 -2950 5045
rect -3000 0 -2950 5005
rect -2900 8445 -2850 15650
rect -2900 8405 -2895 8445
rect -2855 8405 -2850 8445
rect -2900 7245 -2850 8405
rect -2900 7205 -2895 7245
rect -2855 7205 -2850 7245
rect -2900 0 -2850 7205
rect -2800 10645 -2750 15700
rect -2800 10605 -2795 10645
rect -2755 10605 -2750 10645
rect -2800 10595 -2750 10605
rect -2800 10555 -2795 10595
rect -2755 10555 -2750 10595
rect -2800 10545 -2750 10555
rect -2800 10505 -2795 10545
rect -2755 10505 -2750 10545
rect -2800 9345 -2750 10505
rect -2800 9305 -2795 9345
rect -2755 9305 -2750 9345
rect -2800 9295 -2750 9305
rect -2800 9255 -2795 9295
rect -2755 9255 -2750 9295
rect -2800 9245 -2750 9255
rect -2800 9205 -2795 9245
rect -2755 9205 -2750 9245
rect -2800 8045 -2750 9205
rect -2800 8005 -2795 8045
rect -2755 8005 -2750 8045
rect -2800 7995 -2750 8005
rect -2800 7955 -2795 7995
rect -2755 7955 -2750 7995
rect -2800 7945 -2750 7955
rect -2800 7905 -2795 7945
rect -2755 7905 -2750 7945
rect -2800 7745 -2750 7905
rect -2800 7705 -2795 7745
rect -2755 7705 -2750 7745
rect -2800 7695 -2750 7705
rect -2800 7655 -2795 7695
rect -2755 7655 -2750 7695
rect -2800 7645 -2750 7655
rect -2800 7605 -2795 7645
rect -2755 7605 -2750 7645
rect -2800 6445 -2750 7605
rect -2800 6405 -2795 6445
rect -2755 6405 -2750 6445
rect -2800 6395 -2750 6405
rect -2800 6355 -2795 6395
rect -2755 6355 -2750 6395
rect -2800 6345 -2750 6355
rect -2800 6305 -2795 6345
rect -2755 6305 -2750 6345
rect -2800 5145 -2750 6305
rect -2800 5105 -2795 5145
rect -2755 5105 -2750 5145
rect -2800 5095 -2750 5105
rect -2800 5055 -2795 5095
rect -2755 5055 -2750 5095
rect -2800 5045 -2750 5055
rect -2800 5005 -2795 5045
rect -2755 5005 -2750 5045
rect -2800 0 -2750 5005
rect -2700 17115 -2650 17120
rect -2700 17075 -2695 17115
rect -2655 17075 -2650 17115
rect -2700 8845 -2650 17075
rect -2700 8805 -2695 8845
rect -2655 8805 -2650 8845
rect -2700 6845 -2650 8805
rect -2700 6805 -2695 6845
rect -2655 6805 -2650 6845
rect -2700 0 -2650 6805
rect -2600 15750 -2550 17240
rect -2500 15750 -2450 17240
rect -2400 15750 -2350 17240
rect -2300 15750 -2250 17240
rect -2200 15750 -2150 17240
rect -2100 15750 -2050 17240
rect -2000 15750 -1950 17240
rect -1900 15750 -1850 17240
rect -1800 15750 -1750 17240
rect -1700 15750 -1650 17240
rect -2600 15700 -1650 15750
rect -2600 10645 -2550 15700
rect -2600 10605 -2595 10645
rect -2555 10605 -2550 10645
rect -2600 10595 -2550 10605
rect -2600 10555 -2595 10595
rect -2555 10555 -2550 10595
rect -2600 10545 -2550 10555
rect -2600 10505 -2595 10545
rect -2555 10505 -2550 10545
rect -2600 9345 -2550 10505
rect -2600 9305 -2595 9345
rect -2555 9305 -2550 9345
rect -2600 9295 -2550 9305
rect -2600 9255 -2595 9295
rect -2555 9255 -2550 9295
rect -2600 9245 -2550 9255
rect -2600 9205 -2595 9245
rect -2555 9205 -2550 9245
rect -2600 8045 -2550 9205
rect -2600 8005 -2595 8045
rect -2555 8005 -2550 8045
rect -2600 7995 -2550 8005
rect -2600 7955 -2595 7995
rect -2555 7955 -2550 7995
rect -2600 7945 -2550 7955
rect -2600 7905 -2595 7945
rect -2555 7905 -2550 7945
rect -2600 7745 -2550 7905
rect -2600 7705 -2595 7745
rect -2555 7705 -2550 7745
rect -2600 7695 -2550 7705
rect -2600 7655 -2595 7695
rect -2555 7655 -2550 7695
rect -2600 7645 -2550 7655
rect -2600 7605 -2595 7645
rect -2555 7605 -2550 7645
rect -2600 6445 -2550 7605
rect -2600 6405 -2595 6445
rect -2555 6405 -2550 6445
rect -2600 6395 -2550 6405
rect -2600 6355 -2595 6395
rect -2555 6355 -2550 6395
rect -2600 6345 -2550 6355
rect -2600 6305 -2595 6345
rect -2555 6305 -2550 6345
rect -2600 5145 -2550 6305
rect -2600 5105 -2595 5145
rect -2555 5105 -2550 5145
rect -2600 5095 -2550 5105
rect -2600 5055 -2595 5095
rect -2555 5055 -2550 5095
rect -2600 5045 -2550 5055
rect -2600 5005 -2595 5045
rect -2555 5005 -2550 5045
rect -2600 0 -2550 5005
rect -2500 9045 -2450 15650
rect -2500 9005 -2495 9045
rect -2455 9005 -2450 9045
rect -2500 6645 -2450 9005
rect -2500 6605 -2495 6645
rect -2455 6605 -2450 6645
rect -2500 0 -2450 6605
rect -2400 10645 -2350 15700
rect -2400 10605 -2395 10645
rect -2355 10605 -2350 10645
rect -2400 10595 -2350 10605
rect -2400 10555 -2395 10595
rect -2355 10555 -2350 10595
rect -2400 10545 -2350 10555
rect -2400 10505 -2395 10545
rect -2355 10505 -2350 10545
rect -2400 9345 -2350 10505
rect -2400 9305 -2395 9345
rect -2355 9305 -2350 9345
rect -2400 9295 -2350 9305
rect -2400 9255 -2395 9295
rect -2355 9255 -2350 9295
rect -2400 9245 -2350 9255
rect -2400 9205 -2395 9245
rect -2355 9205 -2350 9245
rect -2400 8045 -2350 9205
rect -2400 8005 -2395 8045
rect -2355 8005 -2350 8045
rect -2400 7995 -2350 8005
rect -2400 7955 -2395 7995
rect -2355 7955 -2350 7995
rect -2400 7945 -2350 7955
rect -2400 7905 -2395 7945
rect -2355 7905 -2350 7945
rect -2400 7745 -2350 7905
rect -2400 7705 -2395 7745
rect -2355 7705 -2350 7745
rect -2400 7695 -2350 7705
rect -2400 7655 -2395 7695
rect -2355 7655 -2350 7695
rect -2400 7645 -2350 7655
rect -2400 7605 -2395 7645
rect -2355 7605 -2350 7645
rect -2400 6445 -2350 7605
rect -2400 6405 -2395 6445
rect -2355 6405 -2350 6445
rect -2400 6395 -2350 6405
rect -2400 6355 -2395 6395
rect -2355 6355 -2350 6395
rect -2400 6345 -2350 6355
rect -2400 6305 -2395 6345
rect -2355 6305 -2350 6345
rect -2400 5145 -2350 6305
rect -2400 5105 -2395 5145
rect -2355 5105 -2350 5145
rect -2400 5095 -2350 5105
rect -2400 5055 -2395 5095
rect -2355 5055 -2350 5095
rect -2400 5045 -2350 5055
rect -2400 5005 -2395 5045
rect -2355 5005 -2350 5045
rect -2400 0 -2350 5005
rect -2300 9545 -2250 15650
rect -2300 9505 -2295 9545
rect -2255 9505 -2250 9545
rect -2300 6145 -2250 9505
rect -2300 6105 -2295 6145
rect -2255 6105 -2250 6145
rect -2300 0 -2250 6105
rect -2200 10645 -2150 15700
rect -2200 10605 -2195 10645
rect -2155 10605 -2150 10645
rect -2200 10595 -2150 10605
rect -2200 10555 -2195 10595
rect -2155 10555 -2150 10595
rect -2200 10545 -2150 10555
rect -2200 10505 -2195 10545
rect -2155 10505 -2150 10545
rect -2200 9345 -2150 10505
rect -2200 9305 -2195 9345
rect -2155 9305 -2150 9345
rect -2200 9295 -2150 9305
rect -2200 9255 -2195 9295
rect -2155 9255 -2150 9295
rect -2200 9245 -2150 9255
rect -2200 9205 -2195 9245
rect -2155 9205 -2150 9245
rect -2200 8045 -2150 9205
rect -2200 8005 -2195 8045
rect -2155 8005 -2150 8045
rect -2200 7995 -2150 8005
rect -2200 7955 -2195 7995
rect -2155 7955 -2150 7995
rect -2200 7945 -2150 7955
rect -2200 7905 -2195 7945
rect -2155 7905 -2150 7945
rect -2200 7745 -2150 7905
rect -2200 7705 -2195 7745
rect -2155 7705 -2150 7745
rect -2200 7695 -2150 7705
rect -2200 7655 -2195 7695
rect -2155 7655 -2150 7695
rect -2200 7645 -2150 7655
rect -2200 7605 -2195 7645
rect -2155 7605 -2150 7645
rect -2200 6445 -2150 7605
rect -2200 6405 -2195 6445
rect -2155 6405 -2150 6445
rect -2200 6395 -2150 6405
rect -2200 6355 -2195 6395
rect -2155 6355 -2150 6395
rect -2200 6345 -2150 6355
rect -2200 6305 -2195 6345
rect -2155 6305 -2150 6345
rect -2200 5145 -2150 6305
rect -2200 5105 -2195 5145
rect -2155 5105 -2150 5145
rect -2200 5095 -2150 5105
rect -2200 5055 -2195 5095
rect -2155 5055 -2150 5095
rect -2200 5045 -2150 5055
rect -2200 5005 -2195 5045
rect -2155 5005 -2150 5045
rect -2200 0 -2150 5005
rect -2100 9745 -2050 15650
rect -2100 9705 -2095 9745
rect -2055 9705 -2050 9745
rect -2100 5945 -2050 9705
rect -2100 5905 -2095 5945
rect -2055 5905 -2050 5945
rect -2100 0 -2050 5905
rect -2000 10645 -1950 15700
rect -2000 10605 -1995 10645
rect -1955 10605 -1950 10645
rect -2000 10595 -1950 10605
rect -2000 10555 -1995 10595
rect -1955 10555 -1950 10595
rect -2000 10545 -1950 10555
rect -2000 10505 -1995 10545
rect -1955 10505 -1950 10545
rect -2000 9345 -1950 10505
rect -2000 9305 -1995 9345
rect -1955 9305 -1950 9345
rect -2000 9295 -1950 9305
rect -2000 9255 -1995 9295
rect -1955 9255 -1950 9295
rect -2000 9245 -1950 9255
rect -2000 9205 -1995 9245
rect -1955 9205 -1950 9245
rect -2000 8045 -1950 9205
rect -2000 8005 -1995 8045
rect -1955 8005 -1950 8045
rect -2000 7995 -1950 8005
rect -2000 7955 -1995 7995
rect -1955 7955 -1950 7995
rect -2000 7945 -1950 7955
rect -2000 7905 -1995 7945
rect -1955 7905 -1950 7945
rect -2000 7745 -1950 7905
rect -2000 7705 -1995 7745
rect -1955 7705 -1950 7745
rect -2000 7695 -1950 7705
rect -2000 7655 -1995 7695
rect -1955 7655 -1950 7695
rect -2000 7645 -1950 7655
rect -2000 7605 -1995 7645
rect -1955 7605 -1950 7645
rect -2000 6445 -1950 7605
rect -2000 6405 -1995 6445
rect -1955 6405 -1950 6445
rect -2000 6395 -1950 6405
rect -2000 6355 -1995 6395
rect -1955 6355 -1950 6395
rect -2000 6345 -1950 6355
rect -2000 6305 -1995 6345
rect -1955 6305 -1950 6345
rect -2000 5145 -1950 6305
rect -2000 5105 -1995 5145
rect -1955 5105 -1950 5145
rect -2000 5095 -1950 5105
rect -2000 5055 -1995 5095
rect -1955 5055 -1950 5095
rect -2000 5045 -1950 5055
rect -2000 5005 -1995 5045
rect -1955 5005 -1950 5045
rect -2000 0 -1950 5005
rect -1900 10145 -1850 15650
rect -1900 10105 -1895 10145
rect -1855 10105 -1850 10145
rect -1900 5545 -1850 10105
rect -1900 5505 -1895 5545
rect -1855 5505 -1850 5545
rect -1900 0 -1850 5505
rect -1800 10245 -1750 15650
rect -1800 10205 -1795 10245
rect -1755 10205 -1750 10245
rect -1800 5445 -1750 10205
rect -1800 5405 -1795 5445
rect -1755 5405 -1750 5445
rect -1800 0 -1750 5405
rect -1700 10645 -1650 15700
rect -1700 10605 -1695 10645
rect -1655 10605 -1650 10645
rect -1700 10595 -1650 10605
rect -1700 10555 -1695 10595
rect -1655 10555 -1650 10595
rect -1700 10545 -1650 10555
rect -1700 10505 -1695 10545
rect -1655 10505 -1650 10545
rect -1700 9345 -1650 10505
rect -1700 9305 -1695 9345
rect -1655 9305 -1650 9345
rect -1700 9295 -1650 9305
rect -1700 9255 -1695 9295
rect -1655 9255 -1650 9295
rect -1700 9245 -1650 9255
rect -1700 9205 -1695 9245
rect -1655 9205 -1650 9245
rect -1700 8045 -1650 9205
rect -1700 8005 -1695 8045
rect -1655 8005 -1650 8045
rect -1700 7995 -1650 8005
rect -1700 7955 -1695 7995
rect -1655 7955 -1650 7995
rect -1700 7945 -1650 7955
rect -1700 7905 -1695 7945
rect -1655 7905 -1650 7945
rect -1700 7745 -1650 7905
rect -1700 7705 -1695 7745
rect -1655 7705 -1650 7745
rect -1700 7695 -1650 7705
rect -1700 7655 -1695 7695
rect -1655 7655 -1650 7695
rect -1700 7645 -1650 7655
rect -1700 7605 -1695 7645
rect -1655 7605 -1650 7645
rect -1700 6445 -1650 7605
rect -1700 6405 -1695 6445
rect -1655 6405 -1650 6445
rect -1700 6395 -1650 6405
rect -1700 6355 -1695 6395
rect -1655 6355 -1650 6395
rect -1700 6345 -1650 6355
rect -1700 6305 -1695 6345
rect -1655 6305 -1650 6345
rect -1700 5145 -1650 6305
rect -1700 5105 -1695 5145
rect -1655 5105 -1650 5145
rect -1700 5095 -1650 5105
rect -1700 5055 -1695 5095
rect -1655 5055 -1650 5095
rect -1700 5045 -1650 5055
rect -1700 5005 -1695 5045
rect -1655 5005 -1650 5045
rect -1700 0 -1650 5005
rect -1600 17015 -1550 18290
rect -1600 16975 -1595 17015
rect -1555 16975 -1550 17015
rect -1600 15745 -1550 16975
rect -1600 15705 -1595 15745
rect -1555 15705 -1550 15745
rect -1600 15345 -1550 15705
rect -1600 15305 -1595 15345
rect -1555 15305 -1550 15345
rect -1600 15295 -1550 15305
rect -1600 15255 -1595 15295
rect -1555 15255 -1550 15295
rect -1600 15245 -1550 15255
rect -1600 15205 -1595 15245
rect -1555 15205 -1550 15245
rect -1600 13645 -1550 15205
rect -1600 13605 -1595 13645
rect -1555 13605 -1550 13645
rect -1600 13595 -1550 13605
rect -1600 13555 -1595 13595
rect -1555 13555 -1550 13595
rect -1600 13545 -1550 13555
rect -1600 13505 -1595 13545
rect -1555 13505 -1550 13545
rect -1600 11945 -1550 13505
rect -1600 11905 -1595 11945
rect -1555 11905 -1550 11945
rect -1600 11895 -1550 11905
rect -1600 11855 -1595 11895
rect -1555 11855 -1550 11895
rect -1600 11845 -1550 11855
rect -1600 11805 -1595 11845
rect -1555 11805 -1550 11845
rect -1600 3845 -1550 11805
rect -1600 3805 -1595 3845
rect -1555 3805 -1550 3845
rect -1600 3795 -1550 3805
rect -1600 3755 -1595 3795
rect -1555 3755 -1550 3795
rect -1600 3745 -1550 3755
rect -1600 3705 -1595 3745
rect -1555 3705 -1550 3745
rect -1600 2145 -1550 3705
rect -1600 2105 -1595 2145
rect -1555 2105 -1550 2145
rect -1600 2095 -1550 2105
rect -1600 2055 -1595 2095
rect -1555 2055 -1550 2095
rect -1600 2045 -1550 2055
rect -1600 2005 -1595 2045
rect -1555 2005 -1550 2045
rect -1600 445 -1550 2005
rect -1600 405 -1595 445
rect -1555 405 -1550 445
rect -1600 395 -1550 405
rect -1600 355 -1595 395
rect -1555 355 -1550 395
rect -1600 345 -1550 355
rect -1600 305 -1595 345
rect -1555 305 -1550 345
rect -1600 0 -1550 305
rect -1500 12245 -1450 18290
rect -1500 12205 -1495 12245
rect -1455 12205 -1450 12245
rect -1500 3445 -1450 12205
rect -1500 3405 -1495 3445
rect -1455 3405 -1450 3445
rect -1500 0 -1450 3405
rect -1400 12345 -1350 18290
rect -1400 12305 -1395 12345
rect -1355 12305 -1350 12345
rect -1400 3345 -1350 12305
rect -1400 3305 -1395 3345
rect -1355 3305 -1350 3345
rect -1400 0 -1350 3305
rect -1300 18240 -1250 18290
rect -1300 12445 -1250 18190
rect -1200 18240 -50 18290
rect -1200 17020 -1150 18240
rect -1100 17020 -1050 18240
rect -1000 17020 -950 18240
rect -900 17020 -850 18240
rect -800 17020 -750 18240
rect -700 17020 -650 18240
rect -600 17020 -550 18240
rect -500 17020 -450 18240
rect -400 17020 -350 18240
rect -300 17020 -250 18240
rect -200 17020 -150 18240
rect -100 17020 -50 18240
rect -1200 17015 -50 17020
rect -1200 16975 -1195 17015
rect -1155 16975 -1095 17015
rect -1055 16975 -995 17015
rect -955 16975 -895 17015
rect -855 16975 -795 17015
rect -755 16975 -695 17015
rect -655 16975 -595 17015
rect -555 16975 -495 17015
rect -455 16975 -395 17015
rect -355 16975 -295 17015
rect -255 16975 -195 17015
rect -155 16975 -95 17015
rect -55 16975 -50 17015
rect -1200 16970 -50 16975
rect -1200 15750 -1150 16970
rect -1100 15750 -1050 16970
rect -1000 15750 -950 16970
rect -900 15750 -850 16970
rect -800 15750 -750 16970
rect -700 15750 -650 16970
rect -600 15750 -550 16970
rect -500 15750 -450 16970
rect -1200 15745 -450 15750
rect -1200 15705 -1195 15745
rect -1155 15705 -1095 15745
rect -1055 15705 -995 15745
rect -955 15705 -895 15745
rect -855 15705 -695 15745
rect -655 15705 -595 15745
rect -555 15705 -495 15745
rect -455 15705 -450 15745
rect -1200 15700 -450 15705
rect -1300 12405 -1295 12445
rect -1255 12405 -1250 12445
rect -1300 3245 -1250 12405
rect -1300 3205 -1295 3245
rect -1255 3205 -1250 3245
rect -1300 0 -1250 3205
rect -1200 12545 -1150 15650
rect -1200 12505 -1195 12545
rect -1155 12505 -1150 12545
rect -1200 3145 -1150 12505
rect -1200 3105 -1195 3145
rect -1155 3105 -1150 3145
rect -1200 0 -1150 3105
rect -1100 15345 -1050 15700
rect -1100 15305 -1095 15345
rect -1055 15305 -1050 15345
rect -1100 15295 -1050 15305
rect -1100 15255 -1095 15295
rect -1055 15255 -1050 15295
rect -1100 15245 -1050 15255
rect -1100 15205 -1095 15245
rect -1055 15205 -1050 15245
rect -1100 13645 -1050 15205
rect -1100 13605 -1095 13645
rect -1055 13605 -1050 13645
rect -1100 13595 -1050 13605
rect -1100 13555 -1095 13595
rect -1055 13555 -1050 13595
rect -1100 13545 -1050 13555
rect -1100 13505 -1095 13545
rect -1055 13505 -1050 13545
rect -1100 11945 -1050 13505
rect -1100 11905 -1095 11945
rect -1055 11905 -1050 11945
rect -1100 11895 -1050 11905
rect -1100 11855 -1095 11895
rect -1055 11855 -1050 11895
rect -1100 11845 -1050 11855
rect -1100 11805 -1095 11845
rect -1055 11805 -1050 11845
rect -1100 3845 -1050 11805
rect -1100 3805 -1095 3845
rect -1055 3805 -1050 3845
rect -1100 3795 -1050 3805
rect -1100 3755 -1095 3795
rect -1055 3755 -1050 3795
rect -1100 3745 -1050 3755
rect -1100 3705 -1095 3745
rect -1055 3705 -1050 3745
rect -1100 2145 -1050 3705
rect -1100 2105 -1095 2145
rect -1055 2105 -1050 2145
rect -1100 2095 -1050 2105
rect -1100 2055 -1095 2095
rect -1055 2055 -1050 2095
rect -1100 2045 -1050 2055
rect -1100 2005 -1095 2045
rect -1055 2005 -1050 2045
rect -1100 445 -1050 2005
rect -1100 405 -1095 445
rect -1055 405 -1050 445
rect -1100 395 -1050 405
rect -1100 355 -1095 395
rect -1055 355 -1050 395
rect -1100 345 -1050 355
rect -1100 305 -1095 345
rect -1055 305 -1050 345
rect -1100 0 -1050 305
rect -1000 12945 -950 15650
rect -1000 12905 -995 12945
rect -955 12905 -950 12945
rect -1000 2745 -950 12905
rect -1000 2705 -995 2745
rect -955 2705 -950 2745
rect -1000 0 -950 2705
rect -900 15345 -850 15700
rect -900 15305 -895 15345
rect -855 15305 -850 15345
rect -900 15295 -850 15305
rect -900 15255 -895 15295
rect -855 15255 -850 15295
rect -900 15245 -850 15255
rect -900 15205 -895 15245
rect -855 15205 -850 15245
rect -900 13645 -850 15205
rect -900 13605 -895 13645
rect -855 13605 -850 13645
rect -900 13595 -850 13605
rect -900 13555 -895 13595
rect -855 13555 -850 13595
rect -900 13545 -850 13555
rect -900 13505 -895 13545
rect -855 13505 -850 13545
rect -900 11945 -850 13505
rect -900 11905 -895 11945
rect -855 11905 -850 11945
rect -900 11895 -850 11905
rect -900 11855 -895 11895
rect -855 11855 -850 11895
rect -900 11845 -850 11855
rect -900 11805 -895 11845
rect -855 11805 -850 11845
rect -900 3845 -850 11805
rect -900 3805 -895 3845
rect -855 3805 -850 3845
rect -900 3795 -850 3805
rect -900 3755 -895 3795
rect -855 3755 -850 3795
rect -900 3745 -850 3755
rect -900 3705 -895 3745
rect -855 3705 -850 3745
rect -900 2145 -850 3705
rect -900 2105 -895 2145
rect -855 2105 -850 2145
rect -900 2095 -850 2105
rect -900 2055 -895 2095
rect -855 2055 -850 2095
rect -900 2045 -850 2055
rect -900 2005 -895 2045
rect -855 2005 -850 2045
rect -900 445 -850 2005
rect -900 405 -895 445
rect -855 405 -850 445
rect -900 395 -850 405
rect -900 355 -895 395
rect -855 355 -850 395
rect -900 345 -850 355
rect -900 305 -895 345
rect -855 305 -850 345
rect -900 0 -850 305
rect -800 13145 -750 15650
rect -800 13105 -795 13145
rect -755 13105 -750 13145
rect -800 2545 -750 13105
rect -800 2505 -795 2545
rect -755 2505 -750 2545
rect -800 0 -750 2505
rect -700 15345 -650 15700
rect -700 15305 -695 15345
rect -655 15305 -650 15345
rect -700 15295 -650 15305
rect -700 15255 -695 15295
rect -655 15255 -650 15295
rect -700 15245 -650 15255
rect -700 15205 -695 15245
rect -655 15205 -650 15245
rect -700 13645 -650 15205
rect -700 13605 -695 13645
rect -655 13605 -650 13645
rect -700 13595 -650 13605
rect -700 13555 -695 13595
rect -655 13555 -650 13595
rect -700 13545 -650 13555
rect -700 13505 -695 13545
rect -655 13505 -650 13545
rect -700 11945 -650 13505
rect -700 11905 -695 11945
rect -655 11905 -650 11945
rect -700 11895 -650 11905
rect -700 11855 -695 11895
rect -655 11855 -650 11895
rect -700 11845 -650 11855
rect -700 11805 -695 11845
rect -655 11805 -650 11845
rect -700 3845 -650 11805
rect -700 3805 -695 3845
rect -655 3805 -650 3845
rect -700 3795 -650 3805
rect -700 3755 -695 3795
rect -655 3755 -650 3795
rect -700 3745 -650 3755
rect -700 3705 -695 3745
rect -655 3705 -650 3745
rect -700 2145 -650 3705
rect -700 2105 -695 2145
rect -655 2105 -650 2145
rect -700 2095 -650 2105
rect -700 2055 -695 2095
rect -655 2055 -650 2095
rect -700 2045 -650 2055
rect -700 2005 -695 2045
rect -655 2005 -650 2045
rect -700 445 -650 2005
rect -700 405 -695 445
rect -655 405 -650 445
rect -700 395 -650 405
rect -700 355 -695 395
rect -655 355 -650 395
rect -700 345 -650 355
rect -700 305 -695 345
rect -655 305 -650 345
rect -700 0 -650 305
rect -600 14045 -550 15650
rect -600 14005 -595 14045
rect -555 14005 -550 14045
rect -600 1645 -550 14005
rect -600 1605 -595 1645
rect -555 1605 -550 1645
rect -600 0 -550 1605
rect -500 15345 -450 15700
rect -500 15305 -495 15345
rect -455 15305 -450 15345
rect -500 15295 -450 15305
rect -500 15255 -495 15295
rect -455 15255 -450 15295
rect -500 15245 -450 15255
rect -500 15205 -495 15245
rect -455 15205 -450 15245
rect -500 13645 -450 15205
rect -500 13605 -495 13645
rect -455 13605 -450 13645
rect -500 13595 -450 13605
rect -500 13555 -495 13595
rect -455 13555 -450 13595
rect -500 13545 -450 13555
rect -500 13505 -495 13545
rect -455 13505 -450 13545
rect -500 11945 -450 13505
rect -500 11905 -495 11945
rect -455 11905 -450 11945
rect -500 11895 -450 11905
rect -500 11855 -495 11895
rect -455 11855 -450 11895
rect -500 11845 -450 11855
rect -500 11805 -495 11845
rect -455 11805 -450 11845
rect -500 3845 -450 11805
rect -500 3805 -495 3845
rect -455 3805 -450 3845
rect -500 3795 -450 3805
rect -500 3755 -495 3795
rect -455 3755 -450 3795
rect -500 3745 -450 3755
rect -500 3705 -495 3745
rect -455 3705 -450 3745
rect -500 2145 -450 3705
rect -500 2105 -495 2145
rect -455 2105 -450 2145
rect -500 2095 -450 2105
rect -500 2055 -495 2095
rect -455 2055 -450 2095
rect -500 2045 -450 2055
rect -500 2005 -495 2045
rect -455 2005 -450 2045
rect -500 445 -450 2005
rect -500 405 -495 445
rect -455 405 -450 445
rect -500 395 -450 405
rect -500 355 -495 395
rect -455 355 -450 395
rect -500 345 -450 355
rect -500 305 -495 345
rect -455 305 -450 345
rect -500 0 -450 305
rect -400 16915 -350 16920
rect -400 16875 -395 16915
rect -355 16875 -350 16915
rect -400 14245 -350 16875
rect -400 14205 -395 14245
rect -355 14205 -350 14245
rect -400 1445 -350 14205
rect -400 1405 -395 1445
rect -355 1405 -350 1445
rect -400 0 -350 1405
rect -300 15750 -250 16970
rect -200 15750 -150 16970
rect -100 15750 -50 16970
rect -300 15745 -50 15750
rect -300 15705 -295 15745
rect -255 15705 -195 15745
rect -155 15705 -95 15745
rect -55 15705 -50 15745
rect -300 15700 -50 15705
rect 0 18285 39750 18290
rect 0 18245 5 18285
rect 45 18245 55 18285
rect 95 18245 105 18285
rect 145 18245 155 18285
rect 195 18245 205 18285
rect 245 18245 255 18285
rect 295 18245 305 18285
rect 345 18245 355 18285
rect 395 18245 405 18285
rect 445 18245 455 18285
rect 495 18245 505 18285
rect 545 18245 555 18285
rect 595 18245 605 18285
rect 645 18245 655 18285
rect 695 18245 705 18285
rect 745 18245 755 18285
rect 795 18245 805 18285
rect 845 18245 855 18285
rect 895 18245 905 18285
rect 945 18245 955 18285
rect 995 18245 1005 18285
rect 1045 18245 1055 18285
rect 1095 18245 1105 18285
rect 1145 18245 1155 18285
rect 1195 18245 1205 18285
rect 1245 18245 1255 18285
rect 1295 18245 1305 18285
rect 1345 18245 1355 18285
rect 1395 18245 1405 18285
rect 1445 18245 1455 18285
rect 1495 18245 1505 18285
rect 1545 18245 1555 18285
rect 1595 18245 1605 18285
rect 1645 18245 1655 18285
rect 1695 18245 1705 18285
rect 1745 18245 1755 18285
rect 1795 18245 1805 18285
rect 1845 18245 1855 18285
rect 1895 18245 1905 18285
rect 1945 18245 1955 18285
rect 1995 18245 2005 18285
rect 2045 18245 2055 18285
rect 2095 18245 2105 18285
rect 2145 18245 2155 18285
rect 2195 18245 2205 18285
rect 2245 18245 2255 18285
rect 2295 18245 2305 18285
rect 2345 18245 2355 18285
rect 2395 18245 2405 18285
rect 2445 18245 2455 18285
rect 2495 18245 2505 18285
rect 2545 18245 2555 18285
rect 2595 18245 2605 18285
rect 2645 18245 2655 18285
rect 2695 18245 2705 18285
rect 2745 18245 2755 18285
rect 2795 18245 2805 18285
rect 2845 18245 2855 18285
rect 2895 18245 2905 18285
rect 2945 18245 2955 18285
rect 2995 18245 3005 18285
rect 3045 18245 3055 18285
rect 3095 18245 3105 18285
rect 3145 18245 3155 18285
rect 3195 18245 3205 18285
rect 3245 18245 3255 18285
rect 3295 18245 3305 18285
rect 3345 18245 3355 18285
rect 3395 18245 3405 18285
rect 3445 18245 3455 18285
rect 3495 18245 3505 18285
rect 3545 18245 3555 18285
rect 3595 18245 3605 18285
rect 3645 18245 3655 18285
rect 3695 18245 3705 18285
rect 3745 18245 3755 18285
rect 3795 18245 3805 18285
rect 3845 18245 3855 18285
rect 3895 18245 3905 18285
rect 3945 18245 3955 18285
rect 3995 18245 4005 18285
rect 4045 18245 4055 18285
rect 4095 18245 4105 18285
rect 4145 18245 4155 18285
rect 4195 18245 4205 18285
rect 4245 18245 4255 18285
rect 4295 18245 4305 18285
rect 4345 18245 4355 18285
rect 4395 18245 4405 18285
rect 4445 18245 4455 18285
rect 4495 18245 4505 18285
rect 4545 18245 4555 18285
rect 4595 18245 4605 18285
rect 4645 18245 4655 18285
rect 4695 18245 4705 18285
rect 4745 18245 4755 18285
rect 4795 18245 4805 18285
rect 4845 18245 4855 18285
rect 4895 18245 4905 18285
rect 4945 18245 4955 18285
rect 4995 18245 5005 18285
rect 5045 18245 5055 18285
rect 5095 18245 5105 18285
rect 5145 18245 5155 18285
rect 5195 18245 5205 18285
rect 5245 18245 5255 18285
rect 5295 18245 5305 18285
rect 5345 18245 5355 18285
rect 5395 18245 5405 18285
rect 5445 18245 5455 18285
rect 5495 18245 5505 18285
rect 5545 18245 5555 18285
rect 5595 18245 5605 18285
rect 5645 18245 5655 18285
rect 5695 18245 5705 18285
rect 5745 18245 5755 18285
rect 5795 18245 5805 18285
rect 5845 18245 5855 18285
rect 5895 18245 5905 18285
rect 5945 18245 5955 18285
rect 5995 18245 6005 18285
rect 6045 18245 6055 18285
rect 6095 18245 6105 18285
rect 6145 18245 6155 18285
rect 6195 18245 6205 18285
rect 6245 18245 6255 18285
rect 6295 18245 6305 18285
rect 6345 18245 6355 18285
rect 6395 18245 6405 18285
rect 6445 18245 6455 18285
rect 6495 18245 6505 18285
rect 6545 18245 6555 18285
rect 6595 18245 6605 18285
rect 6645 18245 6655 18285
rect 6695 18245 6705 18285
rect 6745 18245 6755 18285
rect 6795 18245 6805 18285
rect 6845 18245 6855 18285
rect 6895 18245 6905 18285
rect 6945 18245 6955 18285
rect 6995 18245 7005 18285
rect 7045 18245 7055 18285
rect 7095 18245 7105 18285
rect 7145 18245 7155 18285
rect 7195 18245 7205 18285
rect 7245 18245 7255 18285
rect 7295 18245 7305 18285
rect 7345 18245 7355 18285
rect 7395 18245 7405 18285
rect 7445 18245 7455 18285
rect 7495 18245 7505 18285
rect 7545 18245 7555 18285
rect 7595 18245 7605 18285
rect 7645 18245 7655 18285
rect 7695 18245 7705 18285
rect 7745 18245 7755 18285
rect 7795 18245 7805 18285
rect 7845 18245 7855 18285
rect 7895 18245 7905 18285
rect 7945 18245 7955 18285
rect 7995 18245 8005 18285
rect 8045 18245 8055 18285
rect 8095 18245 8105 18285
rect 8145 18245 8155 18285
rect 8195 18245 8205 18285
rect 8245 18245 8255 18285
rect 8295 18245 8305 18285
rect 8345 18245 8355 18285
rect 8395 18245 8405 18285
rect 8445 18245 8455 18285
rect 8495 18245 8505 18285
rect 8545 18245 8555 18285
rect 8595 18245 8605 18285
rect 8645 18245 8655 18285
rect 8695 18245 8705 18285
rect 8745 18245 8755 18285
rect 8795 18245 8805 18285
rect 8845 18245 8855 18285
rect 8895 18245 8905 18285
rect 8945 18245 8955 18285
rect 8995 18245 9005 18285
rect 9045 18245 9055 18285
rect 9095 18245 9105 18285
rect 9145 18245 9155 18285
rect 9195 18245 9205 18285
rect 9245 18245 9255 18285
rect 9295 18245 9305 18285
rect 9345 18245 9355 18285
rect 9395 18245 9405 18285
rect 9445 18245 9455 18285
rect 9495 18245 9505 18285
rect 9545 18245 9555 18285
rect 9595 18245 9605 18285
rect 9645 18245 9655 18285
rect 9695 18245 9705 18285
rect 9745 18245 9755 18285
rect 9795 18245 9805 18285
rect 9845 18245 9855 18285
rect 9895 18245 9905 18285
rect 9945 18245 9955 18285
rect 9995 18245 10005 18285
rect 10045 18245 10055 18285
rect 10095 18245 10105 18285
rect 10145 18245 10155 18285
rect 10195 18245 10205 18285
rect 10245 18245 10255 18285
rect 10295 18245 10305 18285
rect 10345 18245 10355 18285
rect 10395 18245 10405 18285
rect 10445 18245 10455 18285
rect 10495 18245 10505 18285
rect 10545 18245 10555 18285
rect 10595 18245 10605 18285
rect 10645 18245 10655 18285
rect 10695 18245 10705 18285
rect 10745 18245 10755 18285
rect 10795 18245 10805 18285
rect 10845 18245 10855 18285
rect 10895 18245 10905 18285
rect 10945 18245 10955 18285
rect 10995 18245 11005 18285
rect 11045 18245 11055 18285
rect 11095 18245 11105 18285
rect 11145 18245 11155 18285
rect 11195 18245 11205 18285
rect 11245 18245 11255 18285
rect 11295 18245 11305 18285
rect 11345 18245 11355 18285
rect 11395 18245 11405 18285
rect 11445 18245 11455 18285
rect 11495 18245 11505 18285
rect 11545 18245 11555 18285
rect 11595 18245 11605 18285
rect 11645 18245 11655 18285
rect 11695 18245 11705 18285
rect 11745 18245 11755 18285
rect 11795 18245 11805 18285
rect 11845 18245 11855 18285
rect 11895 18245 11905 18285
rect 11945 18245 11955 18285
rect 11995 18245 12005 18285
rect 12045 18245 12055 18285
rect 12095 18245 12105 18285
rect 12145 18245 12155 18285
rect 12195 18245 12205 18285
rect 12245 18245 12255 18285
rect 12295 18245 12305 18285
rect 12345 18245 12355 18285
rect 12395 18245 12405 18285
rect 12445 18245 12455 18285
rect 12495 18245 12505 18285
rect 12545 18245 12555 18285
rect 12595 18245 12605 18285
rect 12645 18245 12655 18285
rect 12695 18245 12705 18285
rect 12745 18245 12755 18285
rect 12795 18245 12805 18285
rect 12845 18245 12855 18285
rect 12895 18245 12905 18285
rect 12945 18245 12955 18285
rect 12995 18245 13005 18285
rect 13045 18245 13055 18285
rect 13095 18245 13105 18285
rect 13145 18245 13155 18285
rect 13195 18245 13205 18285
rect 13245 18245 13255 18285
rect 13295 18245 13305 18285
rect 13345 18245 13355 18285
rect 13395 18245 13405 18285
rect 13445 18245 13455 18285
rect 13495 18245 13505 18285
rect 13545 18245 13555 18285
rect 13595 18245 13605 18285
rect 13645 18245 13655 18285
rect 13695 18245 13705 18285
rect 13745 18245 13755 18285
rect 13795 18245 13805 18285
rect 13845 18245 13855 18285
rect 13895 18245 13905 18285
rect 13945 18245 13955 18285
rect 13995 18245 14005 18285
rect 14045 18245 14055 18285
rect 14095 18245 14105 18285
rect 14145 18245 14155 18285
rect 14195 18245 14205 18285
rect 14245 18245 14255 18285
rect 14295 18245 14305 18285
rect 14345 18245 14355 18285
rect 14395 18245 14405 18285
rect 14445 18245 14455 18285
rect 14495 18245 14505 18285
rect 14545 18245 14555 18285
rect 14595 18245 14605 18285
rect 14645 18245 14655 18285
rect 14695 18245 14705 18285
rect 14745 18245 14755 18285
rect 14795 18245 14805 18285
rect 14845 18245 14855 18285
rect 14895 18245 14905 18285
rect 14945 18245 14955 18285
rect 14995 18245 15005 18285
rect 15045 18245 15055 18285
rect 15095 18245 15105 18285
rect 15145 18245 15155 18285
rect 15195 18245 15205 18285
rect 15245 18245 15255 18285
rect 15295 18245 15305 18285
rect 15345 18245 15355 18285
rect 15395 18245 15405 18285
rect 15445 18245 15455 18285
rect 15495 18245 15505 18285
rect 15545 18245 15555 18285
rect 15595 18245 15605 18285
rect 15645 18245 15655 18285
rect 15695 18245 15705 18285
rect 15745 18245 15755 18285
rect 15795 18245 15805 18285
rect 15845 18245 15855 18285
rect 15895 18245 15905 18285
rect 15945 18245 15955 18285
rect 15995 18245 16005 18285
rect 16045 18245 16055 18285
rect 16095 18245 16105 18285
rect 16145 18245 16155 18285
rect 16195 18245 16205 18285
rect 16245 18245 16255 18285
rect 16295 18245 16305 18285
rect 16345 18245 16355 18285
rect 16395 18245 16405 18285
rect 16445 18245 16455 18285
rect 16495 18245 16505 18285
rect 16545 18245 16555 18285
rect 16595 18245 16605 18285
rect 16645 18245 16655 18285
rect 16695 18245 16705 18285
rect 16745 18245 16755 18285
rect 16795 18245 16805 18285
rect 16845 18245 16855 18285
rect 16895 18245 16905 18285
rect 16945 18245 16955 18285
rect 16995 18245 17005 18285
rect 17045 18245 17055 18285
rect 17095 18245 17105 18285
rect 17145 18245 17155 18285
rect 17195 18245 17205 18285
rect 17245 18245 17255 18285
rect 17295 18245 17305 18285
rect 17345 18245 17355 18285
rect 17395 18245 17405 18285
rect 17445 18245 17455 18285
rect 17495 18245 17505 18285
rect 17545 18245 17555 18285
rect 17595 18245 17605 18285
rect 17645 18245 17655 18285
rect 17695 18245 17705 18285
rect 17745 18245 17755 18285
rect 17795 18245 17805 18285
rect 17845 18245 17855 18285
rect 17895 18245 17905 18285
rect 17945 18245 17955 18285
rect 17995 18245 18005 18285
rect 18045 18245 18055 18285
rect 18095 18245 18105 18285
rect 18145 18245 18155 18285
rect 18195 18245 18205 18285
rect 18245 18245 18255 18285
rect 18295 18245 18305 18285
rect 18345 18245 18355 18285
rect 18395 18245 18405 18285
rect 18445 18245 18455 18285
rect 18495 18245 18505 18285
rect 18545 18245 18555 18285
rect 18595 18245 18605 18285
rect 18645 18245 18655 18285
rect 18695 18245 18705 18285
rect 18745 18245 18755 18285
rect 18795 18245 18805 18285
rect 18845 18245 18855 18285
rect 18895 18245 18905 18285
rect 18945 18245 18955 18285
rect 18995 18245 19005 18285
rect 19045 18245 19055 18285
rect 19095 18245 19105 18285
rect 19145 18245 19155 18285
rect 19195 18245 19205 18285
rect 19245 18245 19255 18285
rect 19295 18245 19305 18285
rect 19345 18245 19355 18285
rect 19395 18245 19405 18285
rect 19445 18245 19455 18285
rect 19495 18245 19505 18285
rect 19545 18245 19555 18285
rect 19595 18245 19605 18285
rect 19645 18245 19655 18285
rect 19695 18245 19705 18285
rect 19745 18245 19755 18285
rect 19795 18245 19805 18285
rect 19845 18245 19855 18285
rect 19895 18245 19905 18285
rect 19945 18245 19955 18285
rect 19995 18245 20005 18285
rect 20045 18245 20055 18285
rect 20095 18245 20105 18285
rect 20145 18245 20155 18285
rect 20195 18245 20205 18285
rect 20245 18245 20255 18285
rect 20295 18245 20305 18285
rect 20345 18245 20355 18285
rect 20395 18245 20405 18285
rect 20445 18245 20455 18285
rect 20495 18245 20505 18285
rect 20545 18245 20555 18285
rect 20595 18245 20605 18285
rect 20645 18245 20655 18285
rect 20695 18245 20705 18285
rect 20745 18245 20755 18285
rect 20795 18245 20805 18285
rect 20845 18245 20855 18285
rect 20895 18245 20905 18285
rect 20945 18245 20955 18285
rect 20995 18245 21005 18285
rect 21045 18245 21055 18285
rect 21095 18245 21105 18285
rect 21145 18245 21155 18285
rect 21195 18245 21205 18285
rect 21245 18245 21255 18285
rect 21295 18245 21305 18285
rect 21345 18245 21355 18285
rect 21395 18245 21405 18285
rect 21445 18245 21455 18285
rect 21495 18245 21505 18285
rect 21545 18245 21555 18285
rect 21595 18245 21605 18285
rect 21645 18245 21655 18285
rect 21695 18245 21705 18285
rect 21745 18245 21755 18285
rect 21795 18245 21805 18285
rect 21845 18245 21855 18285
rect 21895 18245 21905 18285
rect 21945 18245 21955 18285
rect 21995 18245 22005 18285
rect 22045 18245 22055 18285
rect 22095 18245 22105 18285
rect 22145 18245 22155 18285
rect 22195 18245 22205 18285
rect 22245 18245 22255 18285
rect 22295 18245 22305 18285
rect 22345 18245 22355 18285
rect 22395 18245 22405 18285
rect 22445 18245 22455 18285
rect 22495 18245 22505 18285
rect 22545 18245 22555 18285
rect 22595 18245 22605 18285
rect 22645 18245 22655 18285
rect 22695 18245 22705 18285
rect 22745 18245 22755 18285
rect 22795 18245 22805 18285
rect 22845 18245 22855 18285
rect 22895 18245 22905 18285
rect 22945 18245 22955 18285
rect 22995 18245 23005 18285
rect 23045 18245 23055 18285
rect 23095 18245 23105 18285
rect 23145 18245 23155 18285
rect 23195 18245 23205 18285
rect 23245 18245 23255 18285
rect 23295 18245 23305 18285
rect 23345 18245 23355 18285
rect 23395 18245 23405 18285
rect 23445 18245 23455 18285
rect 23495 18245 23505 18285
rect 23545 18245 23555 18285
rect 23595 18245 23605 18285
rect 23645 18245 23655 18285
rect 23695 18245 23705 18285
rect 23745 18245 23755 18285
rect 23795 18245 23805 18285
rect 23845 18245 23855 18285
rect 23895 18245 23905 18285
rect 23945 18245 23955 18285
rect 23995 18245 24005 18285
rect 24045 18245 24055 18285
rect 24095 18245 24105 18285
rect 24145 18245 24155 18285
rect 24195 18245 24205 18285
rect 24245 18245 24255 18285
rect 24295 18245 24305 18285
rect 24345 18245 24355 18285
rect 24395 18245 24405 18285
rect 24445 18245 24455 18285
rect 24495 18245 24505 18285
rect 24545 18245 24555 18285
rect 24595 18245 24605 18285
rect 24645 18245 24655 18285
rect 24695 18245 24705 18285
rect 24745 18245 24755 18285
rect 24795 18245 24805 18285
rect 24845 18245 24855 18285
rect 24895 18245 24905 18285
rect 24945 18245 24955 18285
rect 24995 18245 25005 18285
rect 25045 18245 25055 18285
rect 25095 18245 25105 18285
rect 25145 18245 25155 18285
rect 25195 18245 25205 18285
rect 25245 18245 25255 18285
rect 25295 18245 25305 18285
rect 25345 18245 25355 18285
rect 25395 18245 25405 18285
rect 25445 18245 25455 18285
rect 25495 18245 25505 18285
rect 25545 18245 25555 18285
rect 25595 18245 25605 18285
rect 25645 18245 25655 18285
rect 25695 18245 25705 18285
rect 25745 18245 25755 18285
rect 25795 18245 25805 18285
rect 25845 18245 25855 18285
rect 25895 18245 25905 18285
rect 25945 18245 25955 18285
rect 25995 18245 26005 18285
rect 26045 18245 26055 18285
rect 26095 18245 26105 18285
rect 26145 18245 26155 18285
rect 26195 18245 26205 18285
rect 26245 18245 26255 18285
rect 26295 18245 26305 18285
rect 26345 18245 26355 18285
rect 26395 18245 26405 18285
rect 26445 18245 26455 18285
rect 26495 18245 26505 18285
rect 26545 18245 26555 18285
rect 26595 18245 26605 18285
rect 26645 18245 26655 18285
rect 26695 18245 26705 18285
rect 26745 18245 26755 18285
rect 26795 18245 26805 18285
rect 26845 18245 26855 18285
rect 26895 18245 26905 18285
rect 26945 18245 26955 18285
rect 26995 18245 27005 18285
rect 27045 18245 27055 18285
rect 27095 18245 27105 18285
rect 27145 18245 27155 18285
rect 27195 18245 27205 18285
rect 27245 18245 27255 18285
rect 27295 18245 27305 18285
rect 27345 18245 27355 18285
rect 27395 18245 27405 18285
rect 27445 18245 27455 18285
rect 27495 18245 27505 18285
rect 27545 18245 27555 18285
rect 27595 18245 27605 18285
rect 27645 18245 27655 18285
rect 27695 18245 27705 18285
rect 27745 18245 27755 18285
rect 27795 18245 27805 18285
rect 27845 18245 27855 18285
rect 27895 18245 27905 18285
rect 27945 18245 27955 18285
rect 27995 18245 28005 18285
rect 28045 18245 28055 18285
rect 28095 18245 28105 18285
rect 28145 18245 28155 18285
rect 28195 18245 28205 18285
rect 28245 18245 28255 18285
rect 28295 18245 28305 18285
rect 28345 18245 28355 18285
rect 28395 18245 28405 18285
rect 28445 18245 28455 18285
rect 28495 18245 28505 18285
rect 28545 18245 28555 18285
rect 28595 18245 28605 18285
rect 28645 18245 28655 18285
rect 28695 18245 28705 18285
rect 28745 18245 28755 18285
rect 28795 18245 28805 18285
rect 28845 18245 28855 18285
rect 28895 18245 28905 18285
rect 28945 18245 28955 18285
rect 28995 18245 29005 18285
rect 29045 18245 29055 18285
rect 29095 18245 29105 18285
rect 29145 18245 29155 18285
rect 29195 18245 29205 18285
rect 29245 18245 29255 18285
rect 29295 18245 29305 18285
rect 29345 18245 29355 18285
rect 29395 18245 29405 18285
rect 29445 18245 29455 18285
rect 29495 18245 29505 18285
rect 29545 18245 29555 18285
rect 29595 18245 29605 18285
rect 29645 18245 29655 18285
rect 29695 18245 29705 18285
rect 29745 18245 29755 18285
rect 29795 18245 29805 18285
rect 29845 18245 29855 18285
rect 29895 18245 29905 18285
rect 29945 18245 29955 18285
rect 29995 18245 30005 18285
rect 30045 18245 30055 18285
rect 30095 18245 30105 18285
rect 30145 18245 30155 18285
rect 30195 18245 30205 18285
rect 30245 18245 30255 18285
rect 30295 18245 30305 18285
rect 30345 18245 30355 18285
rect 30395 18245 30405 18285
rect 30445 18245 30455 18285
rect 30495 18245 30505 18285
rect 30545 18245 30555 18285
rect 30595 18245 30605 18285
rect 30645 18245 30655 18285
rect 30695 18245 30705 18285
rect 30745 18245 30755 18285
rect 30795 18245 30805 18285
rect 30845 18245 30855 18285
rect 30895 18245 30905 18285
rect 30945 18245 30955 18285
rect 30995 18245 31005 18285
rect 31045 18245 31055 18285
rect 31095 18245 31105 18285
rect 31145 18245 31155 18285
rect 31195 18245 31205 18285
rect 31245 18245 31255 18285
rect 31295 18245 31305 18285
rect 31345 18245 31355 18285
rect 31395 18245 31405 18285
rect 31445 18245 31455 18285
rect 31495 18245 31505 18285
rect 31545 18245 31555 18285
rect 31595 18245 31605 18285
rect 31645 18245 31655 18285
rect 31695 18245 31705 18285
rect 31745 18245 31755 18285
rect 31795 18245 31805 18285
rect 31845 18245 31855 18285
rect 31895 18245 31905 18285
rect 31945 18245 31955 18285
rect 31995 18245 32005 18285
rect 32045 18245 32055 18285
rect 32095 18245 32105 18285
rect 32145 18245 32155 18285
rect 32195 18245 32205 18285
rect 32245 18245 32255 18285
rect 32295 18245 32305 18285
rect 32345 18245 32355 18285
rect 32395 18245 32405 18285
rect 32445 18245 32455 18285
rect 32495 18245 32505 18285
rect 32545 18245 32555 18285
rect 32595 18245 32605 18285
rect 32645 18245 32655 18285
rect 32695 18245 32705 18285
rect 32745 18245 32755 18285
rect 32795 18245 32805 18285
rect 32845 18245 32855 18285
rect 32895 18245 32905 18285
rect 32945 18245 32955 18285
rect 32995 18245 33005 18285
rect 33045 18245 33055 18285
rect 33095 18245 33105 18285
rect 33145 18245 33155 18285
rect 33195 18245 33205 18285
rect 33245 18245 33255 18285
rect 33295 18245 33305 18285
rect 33345 18245 33355 18285
rect 33395 18245 33405 18285
rect 33445 18245 33455 18285
rect 33495 18245 33505 18285
rect 33545 18245 33555 18285
rect 33595 18245 33605 18285
rect 33645 18245 33655 18285
rect 33695 18245 33705 18285
rect 33745 18245 33755 18285
rect 33795 18245 33805 18285
rect 33845 18245 33855 18285
rect 33895 18245 33905 18285
rect 33945 18245 33955 18285
rect 33995 18245 34005 18285
rect 34045 18245 34055 18285
rect 34095 18245 34105 18285
rect 34145 18245 34155 18285
rect 34195 18245 34205 18285
rect 34245 18245 34255 18285
rect 34295 18245 34305 18285
rect 34345 18245 34355 18285
rect 34395 18245 34405 18285
rect 34445 18245 34455 18285
rect 34495 18245 34505 18285
rect 34545 18245 34555 18285
rect 34595 18245 34605 18285
rect 34645 18245 34655 18285
rect 34695 18245 34705 18285
rect 34745 18245 34755 18285
rect 34795 18245 34805 18285
rect 34845 18245 34855 18285
rect 34895 18245 34905 18285
rect 34945 18245 34955 18285
rect 34995 18245 35005 18285
rect 35045 18245 35055 18285
rect 35095 18245 35105 18285
rect 35145 18245 35155 18285
rect 35195 18245 35205 18285
rect 35245 18245 35255 18285
rect 35295 18245 35305 18285
rect 35345 18245 35355 18285
rect 35395 18245 35405 18285
rect 35445 18245 35455 18285
rect 35495 18245 35505 18285
rect 35545 18245 35555 18285
rect 35595 18245 35605 18285
rect 35645 18245 35655 18285
rect 35695 18245 35705 18285
rect 35745 18245 35755 18285
rect 35795 18245 35805 18285
rect 35845 18245 35855 18285
rect 35895 18245 35905 18285
rect 35945 18245 35955 18285
rect 35995 18245 36005 18285
rect 36045 18245 36055 18285
rect 36095 18245 36105 18285
rect 36145 18245 36155 18285
rect 36195 18245 36205 18285
rect 36245 18245 36255 18285
rect 36295 18245 36305 18285
rect 36345 18245 36355 18285
rect 36395 18245 36405 18285
rect 36445 18245 36455 18285
rect 36495 18245 36505 18285
rect 36545 18245 36555 18285
rect 36595 18245 36605 18285
rect 36645 18245 36655 18285
rect 36695 18245 36705 18285
rect 36745 18245 36755 18285
rect 36795 18245 36805 18285
rect 36845 18245 36855 18285
rect 36895 18245 36905 18285
rect 36945 18245 36955 18285
rect 36995 18245 37005 18285
rect 37045 18245 37055 18285
rect 37095 18245 37105 18285
rect 37145 18245 37155 18285
rect 37195 18245 37205 18285
rect 37245 18245 37255 18285
rect 37295 18245 37305 18285
rect 37345 18245 37355 18285
rect 37395 18245 37405 18285
rect 37445 18245 37455 18285
rect 37495 18245 37505 18285
rect 37545 18245 37555 18285
rect 37595 18245 37605 18285
rect 37645 18245 37655 18285
rect 37695 18245 37705 18285
rect 37745 18245 37755 18285
rect 37795 18245 37805 18285
rect 37845 18245 37855 18285
rect 37895 18245 37905 18285
rect 37945 18245 37955 18285
rect 37995 18245 38005 18285
rect 38045 18245 38055 18285
rect 38095 18245 38105 18285
rect 38145 18245 38155 18285
rect 38195 18245 38205 18285
rect 38245 18245 38255 18285
rect 38295 18245 38305 18285
rect 38345 18245 38355 18285
rect 38395 18245 38405 18285
rect 38445 18245 38455 18285
rect 38495 18245 38505 18285
rect 38545 18245 38555 18285
rect 38595 18245 38605 18285
rect 38645 18245 38655 18285
rect 38695 18245 38705 18285
rect 38745 18245 38755 18285
rect 38795 18245 38805 18285
rect 38845 18245 38855 18285
rect 38895 18245 38905 18285
rect 38945 18245 38955 18285
rect 38995 18245 39005 18285
rect 39045 18245 39055 18285
rect 39095 18245 39105 18285
rect 39145 18245 39155 18285
rect 39195 18245 39205 18285
rect 39245 18245 39255 18285
rect 39295 18245 39305 18285
rect 39345 18245 39355 18285
rect 39395 18245 39405 18285
rect 39445 18245 39455 18285
rect 39495 18245 39505 18285
rect 39545 18245 39555 18285
rect 39595 18245 39605 18285
rect 39645 18245 39655 18285
rect 39695 18245 39705 18285
rect 39745 18245 39750 18285
rect 0 18185 39750 18245
rect 0 18145 5 18185
rect 45 18145 55 18185
rect 95 18145 105 18185
rect 145 18145 155 18185
rect 195 18145 205 18185
rect 245 18145 255 18185
rect 295 18145 305 18185
rect 345 18145 355 18185
rect 395 18145 405 18185
rect 445 18145 455 18185
rect 495 18145 505 18185
rect 545 18145 555 18185
rect 595 18145 605 18185
rect 645 18145 655 18185
rect 695 18145 705 18185
rect 745 18145 755 18185
rect 795 18145 805 18185
rect 845 18145 855 18185
rect 895 18145 905 18185
rect 945 18145 955 18185
rect 995 18145 1005 18185
rect 1045 18145 1055 18185
rect 1095 18145 1105 18185
rect 1145 18145 1155 18185
rect 1195 18145 1205 18185
rect 1245 18145 1255 18185
rect 1295 18145 1305 18185
rect 1345 18145 1355 18185
rect 1395 18145 1405 18185
rect 1445 18145 1455 18185
rect 1495 18145 1505 18185
rect 1545 18145 1555 18185
rect 1595 18145 1605 18185
rect 1645 18145 1655 18185
rect 1695 18145 1705 18185
rect 1745 18145 1755 18185
rect 1795 18145 1805 18185
rect 1845 18145 1855 18185
rect 1895 18145 1905 18185
rect 1945 18145 1955 18185
rect 1995 18145 2005 18185
rect 2045 18145 2055 18185
rect 2095 18145 2105 18185
rect 2145 18145 2155 18185
rect 2195 18145 2205 18185
rect 2245 18145 2255 18185
rect 2295 18145 2305 18185
rect 2345 18145 2355 18185
rect 2395 18145 2405 18185
rect 2445 18145 2455 18185
rect 2495 18145 2505 18185
rect 2545 18145 2555 18185
rect 2595 18145 2605 18185
rect 2645 18145 2655 18185
rect 2695 18145 2705 18185
rect 2745 18145 2755 18185
rect 2795 18145 2805 18185
rect 2845 18145 2855 18185
rect 2895 18145 2905 18185
rect 2945 18145 2955 18185
rect 2995 18145 3005 18185
rect 3045 18145 3055 18185
rect 3095 18145 3105 18185
rect 3145 18145 3155 18185
rect 3195 18145 3205 18185
rect 3245 18145 3255 18185
rect 3295 18145 3305 18185
rect 3345 18145 3355 18185
rect 3395 18145 3405 18185
rect 3445 18145 3455 18185
rect 3495 18145 3505 18185
rect 3545 18145 3555 18185
rect 3595 18145 3605 18185
rect 3645 18145 3655 18185
rect 3695 18145 3705 18185
rect 3745 18145 3755 18185
rect 3795 18145 3805 18185
rect 3845 18145 3855 18185
rect 3895 18145 3905 18185
rect 3945 18145 3955 18185
rect 3995 18145 4005 18185
rect 4045 18145 4055 18185
rect 4095 18145 4105 18185
rect 4145 18145 4155 18185
rect 4195 18145 4205 18185
rect 4245 18145 4255 18185
rect 4295 18145 4305 18185
rect 4345 18145 4355 18185
rect 4395 18145 4405 18185
rect 4445 18145 4455 18185
rect 4495 18145 4505 18185
rect 4545 18145 4555 18185
rect 4595 18145 4605 18185
rect 4645 18145 4655 18185
rect 4695 18145 4705 18185
rect 4745 18145 4755 18185
rect 4795 18145 4805 18185
rect 4845 18145 4855 18185
rect 4895 18145 4905 18185
rect 4945 18145 4955 18185
rect 4995 18145 5005 18185
rect 5045 18145 5055 18185
rect 5095 18145 5105 18185
rect 5145 18145 5155 18185
rect 5195 18145 5205 18185
rect 5245 18145 5255 18185
rect 5295 18145 5305 18185
rect 5345 18145 5355 18185
rect 5395 18145 5405 18185
rect 5445 18145 5455 18185
rect 5495 18145 5505 18185
rect 5545 18145 5555 18185
rect 5595 18145 5605 18185
rect 5645 18145 5655 18185
rect 5695 18145 5705 18185
rect 5745 18145 5755 18185
rect 5795 18145 5805 18185
rect 5845 18145 5855 18185
rect 5895 18145 5905 18185
rect 5945 18145 5955 18185
rect 5995 18145 6005 18185
rect 6045 18145 6055 18185
rect 6095 18145 6105 18185
rect 6145 18145 6155 18185
rect 6195 18145 6205 18185
rect 6245 18145 6255 18185
rect 6295 18145 6305 18185
rect 6345 18145 6355 18185
rect 6395 18145 6405 18185
rect 6445 18145 6455 18185
rect 6495 18145 6505 18185
rect 6545 18145 6555 18185
rect 6595 18145 6605 18185
rect 6645 18145 6655 18185
rect 6695 18145 6705 18185
rect 6745 18145 6755 18185
rect 6795 18145 6805 18185
rect 6845 18145 6855 18185
rect 6895 18145 6905 18185
rect 6945 18145 6955 18185
rect 6995 18145 7005 18185
rect 7045 18145 7055 18185
rect 7095 18145 7105 18185
rect 7145 18145 7155 18185
rect 7195 18145 7205 18185
rect 7245 18145 7255 18185
rect 7295 18145 7305 18185
rect 7345 18145 7355 18185
rect 7395 18145 7405 18185
rect 7445 18145 7455 18185
rect 7495 18145 7505 18185
rect 7545 18145 7555 18185
rect 7595 18145 7605 18185
rect 7645 18145 7655 18185
rect 7695 18145 7705 18185
rect 7745 18145 7755 18185
rect 7795 18145 7805 18185
rect 7845 18145 7855 18185
rect 7895 18145 7905 18185
rect 7945 18145 7955 18185
rect 7995 18145 8005 18185
rect 8045 18145 8055 18185
rect 8095 18145 8105 18185
rect 8145 18145 8155 18185
rect 8195 18145 8205 18185
rect 8245 18145 8255 18185
rect 8295 18145 8305 18185
rect 8345 18145 8355 18185
rect 8395 18145 8405 18185
rect 8445 18145 8455 18185
rect 8495 18145 8505 18185
rect 8545 18145 8555 18185
rect 8595 18145 8605 18185
rect 8645 18145 8655 18185
rect 8695 18145 8705 18185
rect 8745 18145 8755 18185
rect 8795 18145 8805 18185
rect 8845 18145 8855 18185
rect 8895 18145 8905 18185
rect 8945 18145 8955 18185
rect 8995 18145 9005 18185
rect 9045 18145 9055 18185
rect 9095 18145 9105 18185
rect 9145 18145 9155 18185
rect 9195 18145 9205 18185
rect 9245 18145 9255 18185
rect 9295 18145 9305 18185
rect 9345 18145 9355 18185
rect 9395 18145 9405 18185
rect 9445 18145 9455 18185
rect 9495 18145 9505 18185
rect 9545 18145 9555 18185
rect 9595 18145 9605 18185
rect 9645 18145 9655 18185
rect 9695 18145 9705 18185
rect 9745 18145 9755 18185
rect 9795 18145 9805 18185
rect 9845 18145 9855 18185
rect 9895 18145 9905 18185
rect 9945 18145 9955 18185
rect 9995 18145 10005 18185
rect 10045 18145 10055 18185
rect 10095 18145 10105 18185
rect 10145 18145 10155 18185
rect 10195 18145 10205 18185
rect 10245 18145 10255 18185
rect 10295 18145 10305 18185
rect 10345 18145 10355 18185
rect 10395 18145 10405 18185
rect 10445 18145 10455 18185
rect 10495 18145 10505 18185
rect 10545 18145 10555 18185
rect 10595 18145 10605 18185
rect 10645 18145 10655 18185
rect 10695 18145 10705 18185
rect 10745 18145 10755 18185
rect 10795 18145 10805 18185
rect 10845 18145 10855 18185
rect 10895 18145 10905 18185
rect 10945 18145 10955 18185
rect 10995 18145 11005 18185
rect 11045 18145 11055 18185
rect 11095 18145 11105 18185
rect 11145 18145 11155 18185
rect 11195 18145 11205 18185
rect 11245 18145 11255 18185
rect 11295 18145 11305 18185
rect 11345 18145 11355 18185
rect 11395 18145 11405 18185
rect 11445 18145 11455 18185
rect 11495 18145 11505 18185
rect 11545 18145 11555 18185
rect 11595 18145 11605 18185
rect 11645 18145 11655 18185
rect 11695 18145 11705 18185
rect 11745 18145 11755 18185
rect 11795 18145 11805 18185
rect 11845 18145 11855 18185
rect 11895 18145 11905 18185
rect 11945 18145 11955 18185
rect 11995 18145 12005 18185
rect 12045 18145 12055 18185
rect 12095 18145 12105 18185
rect 12145 18145 12155 18185
rect 12195 18145 12205 18185
rect 12245 18145 12255 18185
rect 12295 18145 12305 18185
rect 12345 18145 12355 18185
rect 12395 18145 12405 18185
rect 12445 18145 12455 18185
rect 12495 18145 12505 18185
rect 12545 18145 12555 18185
rect 12595 18145 12605 18185
rect 12645 18145 12655 18185
rect 12695 18145 12705 18185
rect 12745 18145 12755 18185
rect 12795 18145 12805 18185
rect 12845 18145 12855 18185
rect 12895 18145 12905 18185
rect 12945 18145 12955 18185
rect 12995 18145 13005 18185
rect 13045 18145 13055 18185
rect 13095 18145 13105 18185
rect 13145 18145 13155 18185
rect 13195 18145 13205 18185
rect 13245 18145 13255 18185
rect 13295 18145 13305 18185
rect 13345 18145 13355 18185
rect 13395 18145 13405 18185
rect 13445 18145 13455 18185
rect 13495 18145 13505 18185
rect 13545 18145 13555 18185
rect 13595 18145 13605 18185
rect 13645 18145 13655 18185
rect 13695 18145 13705 18185
rect 13745 18145 13755 18185
rect 13795 18145 13805 18185
rect 13845 18145 13855 18185
rect 13895 18145 13905 18185
rect 13945 18145 13955 18185
rect 13995 18145 14005 18185
rect 14045 18145 14055 18185
rect 14095 18145 14105 18185
rect 14145 18145 14155 18185
rect 14195 18145 14205 18185
rect 14245 18145 14255 18185
rect 14295 18145 14305 18185
rect 14345 18145 14355 18185
rect 14395 18145 14405 18185
rect 14445 18145 14455 18185
rect 14495 18145 14505 18185
rect 14545 18145 14555 18185
rect 14595 18145 14605 18185
rect 14645 18145 14655 18185
rect 14695 18145 14705 18185
rect 14745 18145 14755 18185
rect 14795 18145 14805 18185
rect 14845 18145 14855 18185
rect 14895 18145 14905 18185
rect 14945 18145 14955 18185
rect 14995 18145 15005 18185
rect 15045 18145 15055 18185
rect 15095 18145 15105 18185
rect 15145 18145 15155 18185
rect 15195 18145 15205 18185
rect 15245 18145 15255 18185
rect 15295 18145 15305 18185
rect 15345 18145 15355 18185
rect 15395 18145 15405 18185
rect 15445 18145 15455 18185
rect 15495 18145 15505 18185
rect 15545 18145 15555 18185
rect 15595 18145 15605 18185
rect 15645 18145 15655 18185
rect 15695 18145 15705 18185
rect 15745 18145 15755 18185
rect 15795 18145 15805 18185
rect 15845 18145 15855 18185
rect 15895 18145 15905 18185
rect 15945 18145 15955 18185
rect 15995 18145 16005 18185
rect 16045 18145 16055 18185
rect 16095 18145 16105 18185
rect 16145 18145 16155 18185
rect 16195 18145 16205 18185
rect 16245 18145 16255 18185
rect 16295 18145 16305 18185
rect 16345 18145 16355 18185
rect 16395 18145 16405 18185
rect 16445 18145 16455 18185
rect 16495 18145 16505 18185
rect 16545 18145 16555 18185
rect 16595 18145 16605 18185
rect 16645 18145 16655 18185
rect 16695 18145 16705 18185
rect 16745 18145 16755 18185
rect 16795 18145 16805 18185
rect 16845 18145 16855 18185
rect 16895 18145 16905 18185
rect 16945 18145 16955 18185
rect 16995 18145 17005 18185
rect 17045 18145 17055 18185
rect 17095 18145 17105 18185
rect 17145 18145 17155 18185
rect 17195 18145 17205 18185
rect 17245 18145 17255 18185
rect 17295 18145 17305 18185
rect 17345 18145 17355 18185
rect 17395 18145 17405 18185
rect 17445 18145 17455 18185
rect 17495 18145 17505 18185
rect 17545 18145 17555 18185
rect 17595 18145 17605 18185
rect 17645 18145 17655 18185
rect 17695 18145 17705 18185
rect 17745 18145 17755 18185
rect 17795 18145 17805 18185
rect 17845 18145 17855 18185
rect 17895 18145 17905 18185
rect 17945 18145 17955 18185
rect 17995 18145 18005 18185
rect 18045 18145 18055 18185
rect 18095 18145 18105 18185
rect 18145 18145 18155 18185
rect 18195 18145 18205 18185
rect 18245 18145 18255 18185
rect 18295 18145 18305 18185
rect 18345 18145 18355 18185
rect 18395 18145 18405 18185
rect 18445 18145 18455 18185
rect 18495 18145 18505 18185
rect 18545 18145 18555 18185
rect 18595 18145 18605 18185
rect 18645 18145 18655 18185
rect 18695 18145 18705 18185
rect 18745 18145 18755 18185
rect 18795 18145 18805 18185
rect 18845 18145 18855 18185
rect 18895 18145 18905 18185
rect 18945 18145 18955 18185
rect 18995 18145 19005 18185
rect 19045 18145 19055 18185
rect 19095 18145 19105 18185
rect 19145 18145 19155 18185
rect 19195 18145 19205 18185
rect 19245 18145 19255 18185
rect 19295 18145 19305 18185
rect 19345 18145 19355 18185
rect 19395 18145 19405 18185
rect 19445 18145 19455 18185
rect 19495 18145 19505 18185
rect 19545 18145 19555 18185
rect 19595 18145 19605 18185
rect 19645 18145 19655 18185
rect 19695 18145 19705 18185
rect 19745 18145 19755 18185
rect 19795 18145 19805 18185
rect 19845 18145 19855 18185
rect 19895 18145 19905 18185
rect 19945 18145 19955 18185
rect 19995 18145 20005 18185
rect 20045 18145 20055 18185
rect 20095 18145 20105 18185
rect 20145 18145 20155 18185
rect 20195 18145 20205 18185
rect 20245 18145 20255 18185
rect 20295 18145 20305 18185
rect 20345 18145 20355 18185
rect 20395 18145 20405 18185
rect 20445 18145 20455 18185
rect 20495 18145 20505 18185
rect 20545 18145 20555 18185
rect 20595 18145 20605 18185
rect 20645 18145 20655 18185
rect 20695 18145 20705 18185
rect 20745 18145 20755 18185
rect 20795 18145 20805 18185
rect 20845 18145 20855 18185
rect 20895 18145 20905 18185
rect 20945 18145 20955 18185
rect 20995 18145 21005 18185
rect 21045 18145 21055 18185
rect 21095 18145 21105 18185
rect 21145 18145 21155 18185
rect 21195 18145 21205 18185
rect 21245 18145 21255 18185
rect 21295 18145 21305 18185
rect 21345 18145 21355 18185
rect 21395 18145 21405 18185
rect 21445 18145 21455 18185
rect 21495 18145 21505 18185
rect 21545 18145 21555 18185
rect 21595 18145 21605 18185
rect 21645 18145 21655 18185
rect 21695 18145 21705 18185
rect 21745 18145 21755 18185
rect 21795 18145 21805 18185
rect 21845 18145 21855 18185
rect 21895 18145 21905 18185
rect 21945 18145 21955 18185
rect 21995 18145 22005 18185
rect 22045 18145 22055 18185
rect 22095 18145 22105 18185
rect 22145 18145 22155 18185
rect 22195 18145 22205 18185
rect 22245 18145 22255 18185
rect 22295 18145 22305 18185
rect 22345 18145 22355 18185
rect 22395 18145 22405 18185
rect 22445 18145 22455 18185
rect 22495 18145 22505 18185
rect 22545 18145 22555 18185
rect 22595 18145 22605 18185
rect 22645 18145 22655 18185
rect 22695 18145 22705 18185
rect 22745 18145 22755 18185
rect 22795 18145 22805 18185
rect 22845 18145 22855 18185
rect 22895 18145 22905 18185
rect 22945 18145 22955 18185
rect 22995 18145 23005 18185
rect 23045 18145 23055 18185
rect 23095 18145 23105 18185
rect 23145 18145 23155 18185
rect 23195 18145 23205 18185
rect 23245 18145 23255 18185
rect 23295 18145 23305 18185
rect 23345 18145 23355 18185
rect 23395 18145 23405 18185
rect 23445 18145 23455 18185
rect 23495 18145 23505 18185
rect 23545 18145 23555 18185
rect 23595 18145 23605 18185
rect 23645 18145 23655 18185
rect 23695 18145 23705 18185
rect 23745 18145 23755 18185
rect 23795 18145 23805 18185
rect 23845 18145 23855 18185
rect 23895 18145 23905 18185
rect 23945 18145 23955 18185
rect 23995 18145 24005 18185
rect 24045 18145 24055 18185
rect 24095 18145 24105 18185
rect 24145 18145 24155 18185
rect 24195 18145 24205 18185
rect 24245 18145 24255 18185
rect 24295 18145 24305 18185
rect 24345 18145 24355 18185
rect 24395 18145 24405 18185
rect 24445 18145 24455 18185
rect 24495 18145 24505 18185
rect 24545 18145 24555 18185
rect 24595 18145 24605 18185
rect 24645 18145 24655 18185
rect 24695 18145 24705 18185
rect 24745 18145 24755 18185
rect 24795 18145 24805 18185
rect 24845 18145 24855 18185
rect 24895 18145 24905 18185
rect 24945 18145 24955 18185
rect 24995 18145 25005 18185
rect 25045 18145 25055 18185
rect 25095 18145 25105 18185
rect 25145 18145 25155 18185
rect 25195 18145 25205 18185
rect 25245 18145 25255 18185
rect 25295 18145 25305 18185
rect 25345 18145 25355 18185
rect 25395 18145 25405 18185
rect 25445 18145 25455 18185
rect 25495 18145 25505 18185
rect 25545 18145 25555 18185
rect 25595 18145 25605 18185
rect 25645 18145 25655 18185
rect 25695 18145 25705 18185
rect 25745 18145 25755 18185
rect 25795 18145 25805 18185
rect 25845 18145 25855 18185
rect 25895 18145 25905 18185
rect 25945 18145 25955 18185
rect 25995 18145 26005 18185
rect 26045 18145 26055 18185
rect 26095 18145 26105 18185
rect 26145 18145 26155 18185
rect 26195 18145 26205 18185
rect 26245 18145 26255 18185
rect 26295 18145 26305 18185
rect 26345 18145 26355 18185
rect 26395 18145 26405 18185
rect 26445 18145 26455 18185
rect 26495 18145 26505 18185
rect 26545 18145 26555 18185
rect 26595 18145 26605 18185
rect 26645 18145 26655 18185
rect 26695 18145 26705 18185
rect 26745 18145 26755 18185
rect 26795 18145 26805 18185
rect 26845 18145 26855 18185
rect 26895 18145 26905 18185
rect 26945 18145 26955 18185
rect 26995 18145 27005 18185
rect 27045 18145 27055 18185
rect 27095 18145 27105 18185
rect 27145 18145 27155 18185
rect 27195 18145 27205 18185
rect 27245 18145 27255 18185
rect 27295 18145 27305 18185
rect 27345 18145 27355 18185
rect 27395 18145 27405 18185
rect 27445 18145 27455 18185
rect 27495 18145 27505 18185
rect 27545 18145 27555 18185
rect 27595 18145 27605 18185
rect 27645 18145 27655 18185
rect 27695 18145 27705 18185
rect 27745 18145 27755 18185
rect 27795 18145 27805 18185
rect 27845 18145 27855 18185
rect 27895 18145 27905 18185
rect 27945 18145 27955 18185
rect 27995 18145 28005 18185
rect 28045 18145 28055 18185
rect 28095 18145 28105 18185
rect 28145 18145 28155 18185
rect 28195 18145 28205 18185
rect 28245 18145 28255 18185
rect 28295 18145 28305 18185
rect 28345 18145 28355 18185
rect 28395 18145 28405 18185
rect 28445 18145 28455 18185
rect 28495 18145 28505 18185
rect 28545 18145 28555 18185
rect 28595 18145 28605 18185
rect 28645 18145 28655 18185
rect 28695 18145 28705 18185
rect 28745 18145 28755 18185
rect 28795 18145 28805 18185
rect 28845 18145 28855 18185
rect 28895 18145 28905 18185
rect 28945 18145 28955 18185
rect 28995 18145 29005 18185
rect 29045 18145 29055 18185
rect 29095 18145 29105 18185
rect 29145 18145 29155 18185
rect 29195 18145 29205 18185
rect 29245 18145 29255 18185
rect 29295 18145 29305 18185
rect 29345 18145 29355 18185
rect 29395 18145 29405 18185
rect 29445 18145 29455 18185
rect 29495 18145 29505 18185
rect 29545 18145 29555 18185
rect 29595 18145 29605 18185
rect 29645 18145 29655 18185
rect 29695 18145 29705 18185
rect 29745 18145 29755 18185
rect 29795 18145 29805 18185
rect 29845 18145 29855 18185
rect 29895 18145 29905 18185
rect 29945 18145 29955 18185
rect 29995 18145 30005 18185
rect 30045 18145 30055 18185
rect 30095 18145 30105 18185
rect 30145 18145 30155 18185
rect 30195 18145 30205 18185
rect 30245 18145 30255 18185
rect 30295 18145 30305 18185
rect 30345 18145 30355 18185
rect 30395 18145 30405 18185
rect 30445 18145 30455 18185
rect 30495 18145 30505 18185
rect 30545 18145 30555 18185
rect 30595 18145 30605 18185
rect 30645 18145 30655 18185
rect 30695 18145 30705 18185
rect 30745 18145 30755 18185
rect 30795 18145 30805 18185
rect 30845 18145 30855 18185
rect 30895 18145 30905 18185
rect 30945 18145 30955 18185
rect 30995 18145 31005 18185
rect 31045 18145 31055 18185
rect 31095 18145 31105 18185
rect 31145 18145 31155 18185
rect 31195 18145 31205 18185
rect 31245 18145 31255 18185
rect 31295 18145 31305 18185
rect 31345 18145 31355 18185
rect 31395 18145 31405 18185
rect 31445 18145 31455 18185
rect 31495 18145 31505 18185
rect 31545 18145 31555 18185
rect 31595 18145 31605 18185
rect 31645 18145 31655 18185
rect 31695 18145 31705 18185
rect 31745 18145 31755 18185
rect 31795 18145 31805 18185
rect 31845 18145 31855 18185
rect 31895 18145 31905 18185
rect 31945 18145 31955 18185
rect 31995 18145 32005 18185
rect 32045 18145 32055 18185
rect 32095 18145 32105 18185
rect 32145 18145 32155 18185
rect 32195 18145 32205 18185
rect 32245 18145 32255 18185
rect 32295 18145 32305 18185
rect 32345 18145 32355 18185
rect 32395 18145 32405 18185
rect 32445 18145 32455 18185
rect 32495 18145 32505 18185
rect 32545 18145 32555 18185
rect 32595 18145 32605 18185
rect 32645 18145 32655 18185
rect 32695 18145 32705 18185
rect 32745 18145 32755 18185
rect 32795 18145 32805 18185
rect 32845 18145 32855 18185
rect 32895 18145 32905 18185
rect 32945 18145 32955 18185
rect 32995 18145 33005 18185
rect 33045 18145 33055 18185
rect 33095 18145 33105 18185
rect 33145 18145 33155 18185
rect 33195 18145 33205 18185
rect 33245 18145 33255 18185
rect 33295 18145 33305 18185
rect 33345 18145 33355 18185
rect 33395 18145 33405 18185
rect 33445 18145 33455 18185
rect 33495 18145 33505 18185
rect 33545 18145 33555 18185
rect 33595 18145 33605 18185
rect 33645 18145 33655 18185
rect 33695 18145 33705 18185
rect 33745 18145 33755 18185
rect 33795 18145 33805 18185
rect 33845 18145 33855 18185
rect 33895 18145 33905 18185
rect 33945 18145 33955 18185
rect 33995 18145 34005 18185
rect 34045 18145 34055 18185
rect 34095 18145 34105 18185
rect 34145 18145 34155 18185
rect 34195 18145 34205 18185
rect 34245 18145 34255 18185
rect 34295 18145 34305 18185
rect 34345 18145 34355 18185
rect 34395 18145 34405 18185
rect 34445 18145 34455 18185
rect 34495 18145 34505 18185
rect 34545 18145 34555 18185
rect 34595 18145 34605 18185
rect 34645 18145 34655 18185
rect 34695 18145 34705 18185
rect 34745 18145 34755 18185
rect 34795 18145 34805 18185
rect 34845 18145 34855 18185
rect 34895 18145 34905 18185
rect 34945 18145 34955 18185
rect 34995 18145 35005 18185
rect 35045 18145 35055 18185
rect 35095 18145 35105 18185
rect 35145 18145 35155 18185
rect 35195 18145 35205 18185
rect 35245 18145 35255 18185
rect 35295 18145 35305 18185
rect 35345 18145 35355 18185
rect 35395 18145 35405 18185
rect 35445 18145 35455 18185
rect 35495 18145 35505 18185
rect 35545 18145 35555 18185
rect 35595 18145 35605 18185
rect 35645 18145 35655 18185
rect 35695 18145 35705 18185
rect 35745 18145 35755 18185
rect 35795 18145 35805 18185
rect 35845 18145 35855 18185
rect 35895 18145 35905 18185
rect 35945 18145 35955 18185
rect 35995 18145 36005 18185
rect 36045 18145 36055 18185
rect 36095 18145 36105 18185
rect 36145 18145 36155 18185
rect 36195 18145 36205 18185
rect 36245 18145 36255 18185
rect 36295 18145 36305 18185
rect 36345 18145 36355 18185
rect 36395 18145 36405 18185
rect 36445 18145 36455 18185
rect 36495 18145 36505 18185
rect 36545 18145 36555 18185
rect 36595 18145 36605 18185
rect 36645 18145 36655 18185
rect 36695 18145 36705 18185
rect 36745 18145 36755 18185
rect 36795 18145 36805 18185
rect 36845 18145 36855 18185
rect 36895 18145 36905 18185
rect 36945 18145 36955 18185
rect 36995 18145 37005 18185
rect 37045 18145 37055 18185
rect 37095 18145 37105 18185
rect 37145 18145 37155 18185
rect 37195 18145 37205 18185
rect 37245 18145 37255 18185
rect 37295 18145 37305 18185
rect 37345 18145 37355 18185
rect 37395 18145 37405 18185
rect 37445 18145 37455 18185
rect 37495 18145 37505 18185
rect 37545 18145 37555 18185
rect 37595 18145 37605 18185
rect 37645 18145 37655 18185
rect 37695 18145 37705 18185
rect 37745 18145 37755 18185
rect 37795 18145 37805 18185
rect 37845 18145 37855 18185
rect 37895 18145 37905 18185
rect 37945 18145 37955 18185
rect 37995 18145 38005 18185
rect 38045 18145 38055 18185
rect 38095 18145 38105 18185
rect 38145 18145 38155 18185
rect 38195 18145 38205 18185
rect 38245 18145 38255 18185
rect 38295 18145 38305 18185
rect 38345 18145 38355 18185
rect 38395 18145 38405 18185
rect 38445 18145 38455 18185
rect 38495 18145 38505 18185
rect 38545 18145 38555 18185
rect 38595 18145 38605 18185
rect 38645 18145 38655 18185
rect 38695 18145 38705 18185
rect 38745 18145 38755 18185
rect 38795 18145 38805 18185
rect 38845 18145 38855 18185
rect 38895 18145 38905 18185
rect 38945 18145 38955 18185
rect 38995 18145 39005 18185
rect 39045 18145 39055 18185
rect 39095 18145 39105 18185
rect 39145 18145 39155 18185
rect 39195 18145 39205 18185
rect 39245 18145 39255 18185
rect 39295 18145 39305 18185
rect 39345 18145 39355 18185
rect 39395 18145 39405 18185
rect 39445 18145 39455 18185
rect 39495 18145 39505 18185
rect 39545 18145 39555 18185
rect 39595 18145 39605 18185
rect 39645 18145 39655 18185
rect 39695 18145 39705 18185
rect 39745 18145 39750 18185
rect 0 18140 39750 18145
rect 0 17020 50 18140
rect 100 17990 3200 18090
rect 100 17340 200 17990
rect 3100 17340 3200 17990
rect 100 17120 3200 17340
rect 3350 17990 6450 18090
rect 3350 17340 3450 17990
rect 6350 17340 6450 17990
rect 3350 17120 6450 17340
rect 6600 17990 9700 18090
rect 6600 17340 6700 17990
rect 9600 17340 9700 17990
rect 6600 17120 9700 17340
rect 9850 17990 12950 18090
rect 9850 17340 9950 17990
rect 12850 17340 12950 17990
rect 9850 17120 12950 17340
rect 13100 17990 16200 18090
rect 13100 17340 13200 17990
rect 16100 17340 16200 17990
rect 13100 17120 16200 17340
rect 16350 17990 19450 18090
rect 16350 17340 16450 17990
rect 19350 17340 19450 17990
rect 16350 17120 19450 17340
rect 19600 17990 22700 18090
rect 19600 17340 19700 17990
rect 22600 17340 22700 17990
rect 19600 17120 22700 17340
rect 22850 17990 25950 18090
rect 22850 17340 22950 17990
rect 25850 17340 25950 17990
rect 22850 17120 25950 17340
rect 26100 17990 29200 18090
rect 26100 17340 26200 17990
rect 29100 17340 29200 17990
rect 26100 17120 29200 17340
rect 29350 17990 32450 18090
rect 29350 17340 29450 17990
rect 32350 17340 32450 17990
rect 29350 17120 32450 17340
rect 32600 17990 35700 18090
rect 32600 17340 32700 17990
rect 35600 17340 35700 17990
rect 32600 17120 35700 17340
rect 35850 17990 38950 18090
rect 35850 17340 35950 17990
rect 38850 17340 38950 17990
rect 35850 17120 38950 17340
rect 39100 17990 39750 18090
rect 39100 17340 39200 17990
rect 39650 17340 39750 17990
rect 39100 17120 39750 17340
rect 100 17115 39750 17120
rect 100 17075 105 17115
rect 145 17075 155 17115
rect 195 17075 205 17115
rect 245 17075 255 17115
rect 295 17075 305 17115
rect 345 17075 355 17115
rect 395 17075 405 17115
rect 445 17075 455 17115
rect 495 17075 505 17115
rect 545 17075 555 17115
rect 595 17075 605 17115
rect 645 17075 655 17115
rect 695 17075 705 17115
rect 745 17075 755 17115
rect 795 17075 805 17115
rect 845 17075 855 17115
rect 895 17075 905 17115
rect 945 17075 955 17115
rect 995 17075 1005 17115
rect 1045 17075 1055 17115
rect 1095 17075 1105 17115
rect 1145 17075 1155 17115
rect 1195 17075 1205 17115
rect 1245 17075 1255 17115
rect 1295 17075 1305 17115
rect 1345 17075 1355 17115
rect 1395 17075 1405 17115
rect 1445 17075 1455 17115
rect 1495 17075 1505 17115
rect 1545 17075 1555 17115
rect 1595 17075 1605 17115
rect 1645 17075 1655 17115
rect 1695 17075 1705 17115
rect 1745 17075 1755 17115
rect 1795 17075 1805 17115
rect 1845 17075 1855 17115
rect 1895 17075 1905 17115
rect 1945 17075 1955 17115
rect 1995 17075 2005 17115
rect 2045 17075 2055 17115
rect 2095 17075 2105 17115
rect 2145 17075 2155 17115
rect 2195 17075 2205 17115
rect 2245 17075 2255 17115
rect 2295 17075 2305 17115
rect 2345 17075 2355 17115
rect 2395 17075 2405 17115
rect 2445 17075 2455 17115
rect 2495 17075 2505 17115
rect 2545 17075 2555 17115
rect 2595 17075 2605 17115
rect 2645 17075 2655 17115
rect 2695 17075 2705 17115
rect 2745 17075 2755 17115
rect 2795 17075 2805 17115
rect 2845 17075 2855 17115
rect 2895 17075 2905 17115
rect 2945 17075 2955 17115
rect 2995 17075 3005 17115
rect 3045 17075 3055 17115
rect 3095 17075 3105 17115
rect 3145 17075 3155 17115
rect 3195 17075 3205 17115
rect 3245 17075 3255 17115
rect 3295 17075 3305 17115
rect 3345 17075 3355 17115
rect 3395 17075 3405 17115
rect 3445 17075 3455 17115
rect 3495 17075 3505 17115
rect 3545 17075 3555 17115
rect 3595 17075 3605 17115
rect 3645 17075 3655 17115
rect 3695 17075 3705 17115
rect 3745 17075 3755 17115
rect 3795 17075 3805 17115
rect 3845 17075 3855 17115
rect 3895 17075 3905 17115
rect 3945 17075 3955 17115
rect 3995 17075 4005 17115
rect 4045 17075 4055 17115
rect 4095 17075 4105 17115
rect 4145 17075 4155 17115
rect 4195 17075 4205 17115
rect 4245 17075 4255 17115
rect 4295 17075 4305 17115
rect 4345 17075 4355 17115
rect 4395 17075 4405 17115
rect 4445 17075 4455 17115
rect 4495 17075 4505 17115
rect 4545 17075 4555 17115
rect 4595 17075 4605 17115
rect 4645 17075 4655 17115
rect 4695 17075 4705 17115
rect 4745 17075 4755 17115
rect 4795 17075 4805 17115
rect 4845 17075 4855 17115
rect 4895 17075 4905 17115
rect 4945 17075 4955 17115
rect 4995 17075 5005 17115
rect 5045 17075 5055 17115
rect 5095 17075 5105 17115
rect 5145 17075 5155 17115
rect 5195 17075 5205 17115
rect 5245 17075 5255 17115
rect 5295 17075 5305 17115
rect 5345 17075 5355 17115
rect 5395 17075 5405 17115
rect 5445 17075 5455 17115
rect 5495 17075 5505 17115
rect 5545 17075 5555 17115
rect 5595 17075 5605 17115
rect 5645 17075 5655 17115
rect 5695 17075 5705 17115
rect 5745 17075 5755 17115
rect 5795 17075 5805 17115
rect 5845 17075 5855 17115
rect 5895 17075 5905 17115
rect 5945 17075 5955 17115
rect 5995 17075 6005 17115
rect 6045 17075 6055 17115
rect 6095 17075 6105 17115
rect 6145 17075 6155 17115
rect 6195 17075 6205 17115
rect 6245 17075 6255 17115
rect 6295 17075 6305 17115
rect 6345 17075 6355 17115
rect 6395 17075 6405 17115
rect 6445 17075 6455 17115
rect 6495 17075 6505 17115
rect 6545 17075 6555 17115
rect 6595 17075 6605 17115
rect 6645 17075 6655 17115
rect 6695 17075 6705 17115
rect 6745 17075 6755 17115
rect 6795 17075 6805 17115
rect 6845 17075 6855 17115
rect 6895 17075 6905 17115
rect 6945 17075 6955 17115
rect 6995 17075 7005 17115
rect 7045 17075 7055 17115
rect 7095 17075 7105 17115
rect 7145 17075 7155 17115
rect 7195 17075 7205 17115
rect 7245 17075 7255 17115
rect 7295 17075 7305 17115
rect 7345 17075 7355 17115
rect 7395 17075 7405 17115
rect 7445 17075 7455 17115
rect 7495 17075 7505 17115
rect 7545 17075 7555 17115
rect 7595 17075 7605 17115
rect 7645 17075 7655 17115
rect 7695 17075 7705 17115
rect 7745 17075 7755 17115
rect 7795 17075 7805 17115
rect 7845 17075 7855 17115
rect 7895 17075 7905 17115
rect 7945 17075 7955 17115
rect 7995 17075 8005 17115
rect 8045 17075 8055 17115
rect 8095 17075 8105 17115
rect 8145 17075 8155 17115
rect 8195 17075 8205 17115
rect 8245 17075 8255 17115
rect 8295 17075 8305 17115
rect 8345 17075 8355 17115
rect 8395 17075 8405 17115
rect 8445 17075 8455 17115
rect 8495 17075 8505 17115
rect 8545 17075 8555 17115
rect 8595 17075 8605 17115
rect 8645 17075 8655 17115
rect 8695 17075 8705 17115
rect 8745 17075 8755 17115
rect 8795 17075 8805 17115
rect 8845 17075 8855 17115
rect 8895 17075 8905 17115
rect 8945 17075 8955 17115
rect 8995 17075 9005 17115
rect 9045 17075 9055 17115
rect 9095 17075 9105 17115
rect 9145 17075 9155 17115
rect 9195 17075 9205 17115
rect 9245 17075 9255 17115
rect 9295 17075 9305 17115
rect 9345 17075 9355 17115
rect 9395 17075 9405 17115
rect 9445 17075 9455 17115
rect 9495 17075 9505 17115
rect 9545 17075 9555 17115
rect 9595 17075 9605 17115
rect 9645 17075 9655 17115
rect 9695 17075 9705 17115
rect 9745 17075 9755 17115
rect 9795 17075 9805 17115
rect 9845 17075 9855 17115
rect 9895 17075 9905 17115
rect 9945 17075 9955 17115
rect 9995 17075 10005 17115
rect 10045 17075 10055 17115
rect 10095 17075 10105 17115
rect 10145 17075 10155 17115
rect 10195 17075 10205 17115
rect 10245 17075 10255 17115
rect 10295 17075 10305 17115
rect 10345 17075 10355 17115
rect 10395 17075 10405 17115
rect 10445 17075 10455 17115
rect 10495 17075 10505 17115
rect 10545 17075 10555 17115
rect 10595 17075 10605 17115
rect 10645 17075 10655 17115
rect 10695 17075 10705 17115
rect 10745 17075 10755 17115
rect 10795 17075 10805 17115
rect 10845 17075 10855 17115
rect 10895 17075 10905 17115
rect 10945 17075 10955 17115
rect 10995 17075 11005 17115
rect 11045 17075 11055 17115
rect 11095 17075 11105 17115
rect 11145 17075 11155 17115
rect 11195 17075 11205 17115
rect 11245 17075 11255 17115
rect 11295 17075 11305 17115
rect 11345 17075 11355 17115
rect 11395 17075 11405 17115
rect 11445 17075 11455 17115
rect 11495 17075 11505 17115
rect 11545 17075 11555 17115
rect 11595 17075 11605 17115
rect 11645 17075 11655 17115
rect 11695 17075 11705 17115
rect 11745 17075 11755 17115
rect 11795 17075 11805 17115
rect 11845 17075 11855 17115
rect 11895 17075 11905 17115
rect 11945 17075 11955 17115
rect 11995 17075 12005 17115
rect 12045 17075 12055 17115
rect 12095 17075 12105 17115
rect 12145 17075 12155 17115
rect 12195 17075 12205 17115
rect 12245 17075 12255 17115
rect 12295 17075 12305 17115
rect 12345 17075 12355 17115
rect 12395 17075 12405 17115
rect 12445 17075 12455 17115
rect 12495 17075 12505 17115
rect 12545 17075 12555 17115
rect 12595 17075 12605 17115
rect 12645 17075 12655 17115
rect 12695 17075 12705 17115
rect 12745 17075 12755 17115
rect 12795 17075 12805 17115
rect 12845 17075 12855 17115
rect 12895 17075 12905 17115
rect 12945 17075 12955 17115
rect 12995 17075 13005 17115
rect 13045 17075 13055 17115
rect 13095 17075 13105 17115
rect 13145 17075 13155 17115
rect 13195 17075 13205 17115
rect 13245 17075 13255 17115
rect 13295 17075 13305 17115
rect 13345 17075 13355 17115
rect 13395 17075 13405 17115
rect 13445 17075 13455 17115
rect 13495 17075 13505 17115
rect 13545 17075 13555 17115
rect 13595 17075 13605 17115
rect 13645 17075 13655 17115
rect 13695 17075 13705 17115
rect 13745 17075 13755 17115
rect 13795 17075 13805 17115
rect 13845 17075 13855 17115
rect 13895 17075 13905 17115
rect 13945 17075 13955 17115
rect 13995 17075 14005 17115
rect 14045 17075 14055 17115
rect 14095 17075 14105 17115
rect 14145 17075 14155 17115
rect 14195 17075 14205 17115
rect 14245 17075 14255 17115
rect 14295 17075 14305 17115
rect 14345 17075 14355 17115
rect 14395 17075 14405 17115
rect 14445 17075 14455 17115
rect 14495 17075 14505 17115
rect 14545 17075 14555 17115
rect 14595 17075 14605 17115
rect 14645 17075 14655 17115
rect 14695 17075 14705 17115
rect 14745 17075 14755 17115
rect 14795 17075 14805 17115
rect 14845 17075 14855 17115
rect 14895 17075 14905 17115
rect 14945 17075 14955 17115
rect 14995 17075 15005 17115
rect 15045 17075 15055 17115
rect 15095 17075 15105 17115
rect 15145 17075 15155 17115
rect 15195 17075 15205 17115
rect 15245 17075 15255 17115
rect 15295 17075 15305 17115
rect 15345 17075 15355 17115
rect 15395 17075 15405 17115
rect 15445 17075 15455 17115
rect 15495 17075 15505 17115
rect 15545 17075 15555 17115
rect 15595 17075 15605 17115
rect 15645 17075 15655 17115
rect 15695 17075 15705 17115
rect 15745 17075 15755 17115
rect 15795 17075 15805 17115
rect 15845 17075 15855 17115
rect 15895 17075 15905 17115
rect 15945 17075 15955 17115
rect 15995 17075 16005 17115
rect 16045 17075 16055 17115
rect 16095 17075 16105 17115
rect 16145 17075 16155 17115
rect 16195 17075 16205 17115
rect 16245 17075 16255 17115
rect 16295 17075 16305 17115
rect 16345 17075 16355 17115
rect 16395 17075 16405 17115
rect 16445 17075 16455 17115
rect 16495 17075 16505 17115
rect 16545 17075 16555 17115
rect 16595 17075 16605 17115
rect 16645 17075 16655 17115
rect 16695 17075 16705 17115
rect 16745 17075 16755 17115
rect 16795 17075 16805 17115
rect 16845 17075 16855 17115
rect 16895 17075 16905 17115
rect 16945 17075 16955 17115
rect 16995 17075 17005 17115
rect 17045 17075 17055 17115
rect 17095 17075 17105 17115
rect 17145 17075 17155 17115
rect 17195 17075 17205 17115
rect 17245 17075 17255 17115
rect 17295 17075 17305 17115
rect 17345 17075 17355 17115
rect 17395 17075 17405 17115
rect 17445 17075 17455 17115
rect 17495 17075 17505 17115
rect 17545 17075 17555 17115
rect 17595 17075 17605 17115
rect 17645 17075 17655 17115
rect 17695 17075 17705 17115
rect 17745 17075 17755 17115
rect 17795 17075 17805 17115
rect 17845 17075 17855 17115
rect 17895 17075 17905 17115
rect 17945 17075 17955 17115
rect 17995 17075 18005 17115
rect 18045 17075 18055 17115
rect 18095 17075 18105 17115
rect 18145 17075 18155 17115
rect 18195 17075 18205 17115
rect 18245 17075 18255 17115
rect 18295 17075 18305 17115
rect 18345 17075 18355 17115
rect 18395 17075 18405 17115
rect 18445 17075 18455 17115
rect 18495 17075 18505 17115
rect 18545 17075 18555 17115
rect 18595 17075 18605 17115
rect 18645 17075 18655 17115
rect 18695 17075 18705 17115
rect 18745 17075 18755 17115
rect 18795 17075 18805 17115
rect 18845 17075 18855 17115
rect 18895 17075 18905 17115
rect 18945 17075 18955 17115
rect 18995 17075 19005 17115
rect 19045 17075 19055 17115
rect 19095 17075 19105 17115
rect 19145 17075 19155 17115
rect 19195 17075 19205 17115
rect 19245 17075 19255 17115
rect 19295 17075 19305 17115
rect 19345 17075 19355 17115
rect 19395 17075 19405 17115
rect 19445 17075 19455 17115
rect 19495 17075 19505 17115
rect 19545 17075 19555 17115
rect 19595 17075 19605 17115
rect 19645 17075 19655 17115
rect 19695 17075 19705 17115
rect 19745 17075 19755 17115
rect 19795 17075 19805 17115
rect 19845 17075 19855 17115
rect 19895 17075 19905 17115
rect 19945 17075 19955 17115
rect 19995 17075 20005 17115
rect 20045 17075 20055 17115
rect 20095 17075 20105 17115
rect 20145 17075 20155 17115
rect 20195 17075 20205 17115
rect 20245 17075 20255 17115
rect 20295 17075 20305 17115
rect 20345 17075 20355 17115
rect 20395 17075 20405 17115
rect 20445 17075 20455 17115
rect 20495 17075 20505 17115
rect 20545 17075 20555 17115
rect 20595 17075 20605 17115
rect 20645 17075 20655 17115
rect 20695 17075 20705 17115
rect 20745 17075 20755 17115
rect 20795 17075 20805 17115
rect 20845 17075 20855 17115
rect 20895 17075 20905 17115
rect 20945 17075 20955 17115
rect 20995 17075 21005 17115
rect 21045 17075 21055 17115
rect 21095 17075 21105 17115
rect 21145 17075 21155 17115
rect 21195 17075 21205 17115
rect 21245 17075 21255 17115
rect 21295 17075 21305 17115
rect 21345 17075 21355 17115
rect 21395 17075 21405 17115
rect 21445 17075 21455 17115
rect 21495 17075 21505 17115
rect 21545 17075 21555 17115
rect 21595 17075 21605 17115
rect 21645 17075 21655 17115
rect 21695 17075 21705 17115
rect 21745 17075 21755 17115
rect 21795 17075 21805 17115
rect 21845 17075 21855 17115
rect 21895 17075 21905 17115
rect 21945 17075 21955 17115
rect 21995 17075 22005 17115
rect 22045 17075 22055 17115
rect 22095 17075 22105 17115
rect 22145 17075 22155 17115
rect 22195 17075 22205 17115
rect 22245 17075 22255 17115
rect 22295 17075 22305 17115
rect 22345 17075 22355 17115
rect 22395 17075 22405 17115
rect 22445 17075 22455 17115
rect 22495 17075 22505 17115
rect 22545 17075 22555 17115
rect 22595 17075 22605 17115
rect 22645 17075 22655 17115
rect 22695 17075 22705 17115
rect 22745 17075 22755 17115
rect 22795 17075 22805 17115
rect 22845 17075 22855 17115
rect 22895 17075 22905 17115
rect 22945 17075 22955 17115
rect 22995 17075 23005 17115
rect 23045 17075 23055 17115
rect 23095 17075 23105 17115
rect 23145 17075 23155 17115
rect 23195 17075 23205 17115
rect 23245 17075 23255 17115
rect 23295 17075 23305 17115
rect 23345 17075 23355 17115
rect 23395 17075 23405 17115
rect 23445 17075 23455 17115
rect 23495 17075 23505 17115
rect 23545 17075 23555 17115
rect 23595 17075 23605 17115
rect 23645 17075 23655 17115
rect 23695 17075 23705 17115
rect 23745 17075 23755 17115
rect 23795 17075 23805 17115
rect 23845 17075 23855 17115
rect 23895 17075 23905 17115
rect 23945 17075 23955 17115
rect 23995 17075 24005 17115
rect 24045 17075 24055 17115
rect 24095 17075 24105 17115
rect 24145 17075 24155 17115
rect 24195 17075 24205 17115
rect 24245 17075 24255 17115
rect 24295 17075 24305 17115
rect 24345 17075 24355 17115
rect 24395 17075 24405 17115
rect 24445 17075 24455 17115
rect 24495 17075 24505 17115
rect 24545 17075 24555 17115
rect 24595 17075 24605 17115
rect 24645 17075 24655 17115
rect 24695 17075 24705 17115
rect 24745 17075 24755 17115
rect 24795 17075 24805 17115
rect 24845 17075 24855 17115
rect 24895 17075 24905 17115
rect 24945 17075 24955 17115
rect 24995 17075 25005 17115
rect 25045 17075 25055 17115
rect 25095 17075 25105 17115
rect 25145 17075 25155 17115
rect 25195 17075 25205 17115
rect 25245 17075 25255 17115
rect 25295 17075 25305 17115
rect 25345 17075 25355 17115
rect 25395 17075 25405 17115
rect 25445 17075 25455 17115
rect 25495 17075 25505 17115
rect 25545 17075 25555 17115
rect 25595 17075 25605 17115
rect 25645 17075 25655 17115
rect 25695 17075 25705 17115
rect 25745 17075 25755 17115
rect 25795 17075 25805 17115
rect 25845 17075 25855 17115
rect 25895 17075 25905 17115
rect 25945 17075 25955 17115
rect 25995 17075 26005 17115
rect 26045 17075 26055 17115
rect 26095 17075 26105 17115
rect 26145 17075 26155 17115
rect 26195 17075 26205 17115
rect 26245 17075 26255 17115
rect 26295 17075 26305 17115
rect 26345 17075 26355 17115
rect 26395 17075 26405 17115
rect 26445 17075 26455 17115
rect 26495 17075 26505 17115
rect 26545 17075 26555 17115
rect 26595 17075 26605 17115
rect 26645 17075 26655 17115
rect 26695 17075 26705 17115
rect 26745 17075 26755 17115
rect 26795 17075 26805 17115
rect 26845 17075 26855 17115
rect 26895 17075 26905 17115
rect 26945 17075 26955 17115
rect 26995 17075 27005 17115
rect 27045 17075 27055 17115
rect 27095 17075 27105 17115
rect 27145 17075 27155 17115
rect 27195 17075 27205 17115
rect 27245 17075 27255 17115
rect 27295 17075 27305 17115
rect 27345 17075 27355 17115
rect 27395 17075 27405 17115
rect 27445 17075 27455 17115
rect 27495 17075 27505 17115
rect 27545 17075 27555 17115
rect 27595 17075 27605 17115
rect 27645 17075 27655 17115
rect 27695 17075 27705 17115
rect 27745 17075 27755 17115
rect 27795 17075 27805 17115
rect 27845 17075 27855 17115
rect 27895 17075 27905 17115
rect 27945 17075 27955 17115
rect 27995 17075 28005 17115
rect 28045 17075 28055 17115
rect 28095 17075 28105 17115
rect 28145 17075 28155 17115
rect 28195 17075 28205 17115
rect 28245 17075 28255 17115
rect 28295 17075 28305 17115
rect 28345 17075 28355 17115
rect 28395 17075 28405 17115
rect 28445 17075 28455 17115
rect 28495 17075 28505 17115
rect 28545 17075 28555 17115
rect 28595 17075 28605 17115
rect 28645 17075 28655 17115
rect 28695 17075 28705 17115
rect 28745 17075 28755 17115
rect 28795 17075 28805 17115
rect 28845 17075 28855 17115
rect 28895 17075 28905 17115
rect 28945 17075 28955 17115
rect 28995 17075 29005 17115
rect 29045 17075 29055 17115
rect 29095 17075 29105 17115
rect 29145 17075 29155 17115
rect 29195 17075 29205 17115
rect 29245 17075 29255 17115
rect 29295 17075 29305 17115
rect 29345 17075 29355 17115
rect 29395 17075 29405 17115
rect 29445 17075 29455 17115
rect 29495 17075 29505 17115
rect 29545 17075 29555 17115
rect 29595 17075 29605 17115
rect 29645 17075 29655 17115
rect 29695 17075 29705 17115
rect 29745 17075 29755 17115
rect 29795 17075 29805 17115
rect 29845 17075 29855 17115
rect 29895 17075 29905 17115
rect 29945 17075 29955 17115
rect 29995 17075 30005 17115
rect 30045 17075 30055 17115
rect 30095 17075 30105 17115
rect 30145 17075 30155 17115
rect 30195 17075 30205 17115
rect 30245 17075 30255 17115
rect 30295 17075 30305 17115
rect 30345 17075 30355 17115
rect 30395 17075 30405 17115
rect 30445 17075 30455 17115
rect 30495 17075 30505 17115
rect 30545 17075 30555 17115
rect 30595 17075 30605 17115
rect 30645 17075 30655 17115
rect 30695 17075 30705 17115
rect 30745 17075 30755 17115
rect 30795 17075 30805 17115
rect 30845 17075 30855 17115
rect 30895 17075 30905 17115
rect 30945 17075 30955 17115
rect 30995 17075 31005 17115
rect 31045 17075 31055 17115
rect 31095 17075 31105 17115
rect 31145 17075 31155 17115
rect 31195 17075 31205 17115
rect 31245 17075 31255 17115
rect 31295 17075 31305 17115
rect 31345 17075 31355 17115
rect 31395 17075 31405 17115
rect 31445 17075 31455 17115
rect 31495 17075 31505 17115
rect 31545 17075 31555 17115
rect 31595 17075 31605 17115
rect 31645 17075 31655 17115
rect 31695 17075 31705 17115
rect 31745 17075 31755 17115
rect 31795 17075 31805 17115
rect 31845 17075 31855 17115
rect 31895 17075 31905 17115
rect 31945 17075 31955 17115
rect 31995 17075 32005 17115
rect 32045 17075 32055 17115
rect 32095 17075 32105 17115
rect 32145 17075 32155 17115
rect 32195 17075 32205 17115
rect 32245 17075 32255 17115
rect 32295 17075 32305 17115
rect 32345 17075 32355 17115
rect 32395 17075 32405 17115
rect 32445 17075 32455 17115
rect 32495 17075 32505 17115
rect 32545 17075 32555 17115
rect 32595 17075 32605 17115
rect 32645 17075 32655 17115
rect 32695 17075 32705 17115
rect 32745 17075 32755 17115
rect 32795 17075 32805 17115
rect 32845 17075 32855 17115
rect 32895 17075 32905 17115
rect 32945 17075 32955 17115
rect 32995 17075 33005 17115
rect 33045 17075 33055 17115
rect 33095 17075 33105 17115
rect 33145 17075 33155 17115
rect 33195 17075 33205 17115
rect 33245 17075 33255 17115
rect 33295 17075 33305 17115
rect 33345 17075 33355 17115
rect 33395 17075 33405 17115
rect 33445 17075 33455 17115
rect 33495 17075 33505 17115
rect 33545 17075 33555 17115
rect 33595 17075 33605 17115
rect 33645 17075 33655 17115
rect 33695 17075 33705 17115
rect 33745 17075 33755 17115
rect 33795 17075 33805 17115
rect 33845 17075 33855 17115
rect 33895 17075 33905 17115
rect 33945 17075 33955 17115
rect 33995 17075 34005 17115
rect 34045 17075 34055 17115
rect 34095 17075 34105 17115
rect 34145 17075 34155 17115
rect 34195 17075 34205 17115
rect 34245 17075 34255 17115
rect 34295 17075 34305 17115
rect 34345 17075 34355 17115
rect 34395 17075 34405 17115
rect 34445 17075 34455 17115
rect 34495 17075 34505 17115
rect 34545 17075 34555 17115
rect 34595 17075 34605 17115
rect 34645 17075 34655 17115
rect 34695 17075 34705 17115
rect 34745 17075 34755 17115
rect 34795 17075 34805 17115
rect 34845 17075 34855 17115
rect 34895 17075 34905 17115
rect 34945 17075 34955 17115
rect 34995 17075 35005 17115
rect 35045 17075 35055 17115
rect 35095 17075 35105 17115
rect 35145 17075 35155 17115
rect 35195 17075 35205 17115
rect 35245 17075 35255 17115
rect 35295 17075 35305 17115
rect 35345 17075 35355 17115
rect 35395 17075 35405 17115
rect 35445 17075 35455 17115
rect 35495 17075 35505 17115
rect 35545 17075 35555 17115
rect 35595 17075 35605 17115
rect 35645 17075 35655 17115
rect 35695 17075 35705 17115
rect 35745 17075 35755 17115
rect 35795 17075 35805 17115
rect 35845 17075 35855 17115
rect 35895 17075 35905 17115
rect 35945 17075 35955 17115
rect 35995 17075 36005 17115
rect 36045 17075 36055 17115
rect 36095 17075 36105 17115
rect 36145 17075 36155 17115
rect 36195 17075 36205 17115
rect 36245 17075 36255 17115
rect 36295 17075 36305 17115
rect 36345 17075 36355 17115
rect 36395 17075 36405 17115
rect 36445 17075 36455 17115
rect 36495 17075 36505 17115
rect 36545 17075 36555 17115
rect 36595 17075 36605 17115
rect 36645 17075 36655 17115
rect 36695 17075 36705 17115
rect 36745 17075 36755 17115
rect 36795 17075 36805 17115
rect 36845 17075 36855 17115
rect 36895 17075 36905 17115
rect 36945 17075 36955 17115
rect 36995 17075 37005 17115
rect 37045 17075 37055 17115
rect 37095 17075 37105 17115
rect 37145 17075 37155 17115
rect 37195 17075 37205 17115
rect 37245 17075 37255 17115
rect 37295 17075 37305 17115
rect 37345 17075 37355 17115
rect 37395 17075 37405 17115
rect 37445 17075 37455 17115
rect 37495 17075 37505 17115
rect 37545 17075 37555 17115
rect 37595 17075 37605 17115
rect 37645 17075 37655 17115
rect 37695 17075 37705 17115
rect 37745 17075 37755 17115
rect 37795 17075 37805 17115
rect 37845 17075 37855 17115
rect 37895 17075 37905 17115
rect 37945 17075 37955 17115
rect 37995 17075 38005 17115
rect 38045 17075 38055 17115
rect 38095 17075 38105 17115
rect 38145 17075 38155 17115
rect 38195 17075 38205 17115
rect 38245 17075 38255 17115
rect 38295 17075 38305 17115
rect 38345 17075 38355 17115
rect 38395 17075 38405 17115
rect 38445 17075 38455 17115
rect 38495 17075 38505 17115
rect 38545 17075 38555 17115
rect 38595 17075 38605 17115
rect 38645 17075 38655 17115
rect 38695 17075 38705 17115
rect 38745 17075 38755 17115
rect 38795 17075 38805 17115
rect 38845 17075 38855 17115
rect 38895 17075 38905 17115
rect 38945 17075 38955 17115
rect 38995 17075 39005 17115
rect 39045 17075 39055 17115
rect 39095 17075 39105 17115
rect 39145 17075 39155 17115
rect 39195 17075 39205 17115
rect 39245 17075 39255 17115
rect 39295 17075 39305 17115
rect 39345 17075 39355 17115
rect 39395 17075 39405 17115
rect 39445 17075 39455 17115
rect 39495 17075 39505 17115
rect 39545 17075 39555 17115
rect 39595 17075 39605 17115
rect 39645 17075 39655 17115
rect 39695 17075 39705 17115
rect 39745 17075 39750 17115
rect 100 17070 39750 17075
rect 0 17015 39750 17020
rect 0 16975 5 17015
rect 45 16975 55 17015
rect 95 16975 105 17015
rect 145 16975 155 17015
rect 195 16975 205 17015
rect 245 16975 255 17015
rect 295 16975 305 17015
rect 345 16975 355 17015
rect 395 16975 405 17015
rect 445 16975 455 17015
rect 495 16975 505 17015
rect 545 16975 555 17015
rect 595 16975 605 17015
rect 645 16975 655 17015
rect 695 16975 705 17015
rect 745 16975 755 17015
rect 795 16975 805 17015
rect 845 16975 855 17015
rect 895 16975 905 17015
rect 945 16975 955 17015
rect 995 16975 1005 17015
rect 1045 16975 1055 17015
rect 1095 16975 1105 17015
rect 1145 16975 1155 17015
rect 1195 16975 1205 17015
rect 1245 16975 1255 17015
rect 1295 16975 1305 17015
rect 1345 16975 1355 17015
rect 1395 16975 1405 17015
rect 1445 16975 1455 17015
rect 1495 16975 1505 17015
rect 1545 16975 1555 17015
rect 1595 16975 1605 17015
rect 1645 16975 1655 17015
rect 1695 16975 1705 17015
rect 1745 16975 1755 17015
rect 1795 16975 1805 17015
rect 1845 16975 1855 17015
rect 1895 16975 1905 17015
rect 1945 16975 1955 17015
rect 1995 16975 2005 17015
rect 2045 16975 2055 17015
rect 2095 16975 2105 17015
rect 2145 16975 2155 17015
rect 2195 16975 2205 17015
rect 2245 16975 2255 17015
rect 2295 16975 2305 17015
rect 2345 16975 2355 17015
rect 2395 16975 2405 17015
rect 2445 16975 2455 17015
rect 2495 16975 2505 17015
rect 2545 16975 2555 17015
rect 2595 16975 2605 17015
rect 2645 16975 2655 17015
rect 2695 16975 2705 17015
rect 2745 16975 2755 17015
rect 2795 16975 2805 17015
rect 2845 16975 2855 17015
rect 2895 16975 2905 17015
rect 2945 16975 2955 17015
rect 2995 16975 3005 17015
rect 3045 16975 3055 17015
rect 3095 16975 3105 17015
rect 3145 16975 3155 17015
rect 3195 16975 3205 17015
rect 3245 16975 3255 17015
rect 3295 16975 3305 17015
rect 3345 16975 3355 17015
rect 3395 16975 3405 17015
rect 3445 16975 3455 17015
rect 3495 16975 3505 17015
rect 3545 16975 3555 17015
rect 3595 16975 3605 17015
rect 3645 16975 3655 17015
rect 3695 16975 3705 17015
rect 3745 16975 3755 17015
rect 3795 16975 3805 17015
rect 3845 16975 3855 17015
rect 3895 16975 3905 17015
rect 3945 16975 3955 17015
rect 3995 16975 4005 17015
rect 4045 16975 4055 17015
rect 4095 16975 4105 17015
rect 4145 16975 4155 17015
rect 4195 16975 4205 17015
rect 4245 16975 4255 17015
rect 4295 16975 4305 17015
rect 4345 16975 4355 17015
rect 4395 16975 4405 17015
rect 4445 16975 4455 17015
rect 4495 16975 4505 17015
rect 4545 16975 4555 17015
rect 4595 16975 4605 17015
rect 4645 16975 4655 17015
rect 4695 16975 4705 17015
rect 4745 16975 4755 17015
rect 4795 16975 4805 17015
rect 4845 16975 4855 17015
rect 4895 16975 4905 17015
rect 4945 16975 4955 17015
rect 4995 16975 5005 17015
rect 5045 16975 5055 17015
rect 5095 16975 5105 17015
rect 5145 16975 5155 17015
rect 5195 16975 5205 17015
rect 5245 16975 5255 17015
rect 5295 16975 5305 17015
rect 5345 16975 5355 17015
rect 5395 16975 5405 17015
rect 5445 16975 5455 17015
rect 5495 16975 5505 17015
rect 5545 16975 5555 17015
rect 5595 16975 5605 17015
rect 5645 16975 5655 17015
rect 5695 16975 5705 17015
rect 5745 16975 5755 17015
rect 5795 16975 5805 17015
rect 5845 16975 5855 17015
rect 5895 16975 5905 17015
rect 5945 16975 5955 17015
rect 5995 16975 6005 17015
rect 6045 16975 6055 17015
rect 6095 16975 6105 17015
rect 6145 16975 6155 17015
rect 6195 16975 6205 17015
rect 6245 16975 6255 17015
rect 6295 16975 6305 17015
rect 6345 16975 6355 17015
rect 6395 16975 6405 17015
rect 6445 16975 6455 17015
rect 6495 16975 6505 17015
rect 6545 16975 6555 17015
rect 6595 16975 6605 17015
rect 6645 16975 6655 17015
rect 6695 16975 6705 17015
rect 6745 16975 6755 17015
rect 6795 16975 6805 17015
rect 6845 16975 6855 17015
rect 6895 16975 6905 17015
rect 6945 16975 6955 17015
rect 6995 16975 7005 17015
rect 7045 16975 7055 17015
rect 7095 16975 7105 17015
rect 7145 16975 7155 17015
rect 7195 16975 7205 17015
rect 7245 16975 7255 17015
rect 7295 16975 7305 17015
rect 7345 16975 7355 17015
rect 7395 16975 7405 17015
rect 7445 16975 7455 17015
rect 7495 16975 7505 17015
rect 7545 16975 7555 17015
rect 7595 16975 7605 17015
rect 7645 16975 7655 17015
rect 7695 16975 7705 17015
rect 7745 16975 7755 17015
rect 7795 16975 7805 17015
rect 7845 16975 7855 17015
rect 7895 16975 7905 17015
rect 7945 16975 7955 17015
rect 7995 16975 8005 17015
rect 8045 16975 8055 17015
rect 8095 16975 8105 17015
rect 8145 16975 8155 17015
rect 8195 16975 8205 17015
rect 8245 16975 8255 17015
rect 8295 16975 8305 17015
rect 8345 16975 8355 17015
rect 8395 16975 8405 17015
rect 8445 16975 8455 17015
rect 8495 16975 8505 17015
rect 8545 16975 8555 17015
rect 8595 16975 8605 17015
rect 8645 16975 8655 17015
rect 8695 16975 8705 17015
rect 8745 16975 8755 17015
rect 8795 16975 8805 17015
rect 8845 16975 8855 17015
rect 8895 16975 8905 17015
rect 8945 16975 8955 17015
rect 8995 16975 9005 17015
rect 9045 16975 9055 17015
rect 9095 16975 9105 17015
rect 9145 16975 9155 17015
rect 9195 16975 9205 17015
rect 9245 16975 9255 17015
rect 9295 16975 9305 17015
rect 9345 16975 9355 17015
rect 9395 16975 9405 17015
rect 9445 16975 9455 17015
rect 9495 16975 9505 17015
rect 9545 16975 9555 17015
rect 9595 16975 9605 17015
rect 9645 16975 9655 17015
rect 9695 16975 9705 17015
rect 9745 16975 9755 17015
rect 9795 16975 9805 17015
rect 9845 16975 9855 17015
rect 9895 16975 9905 17015
rect 9945 16975 9955 17015
rect 9995 16975 10005 17015
rect 10045 16975 10055 17015
rect 10095 16975 10105 17015
rect 10145 16975 10155 17015
rect 10195 16975 10205 17015
rect 10245 16975 10255 17015
rect 10295 16975 10305 17015
rect 10345 16975 10355 17015
rect 10395 16975 10405 17015
rect 10445 16975 10455 17015
rect 10495 16975 10505 17015
rect 10545 16975 10555 17015
rect 10595 16975 10605 17015
rect 10645 16975 10655 17015
rect 10695 16975 10705 17015
rect 10745 16975 10755 17015
rect 10795 16975 10805 17015
rect 10845 16975 10855 17015
rect 10895 16975 10905 17015
rect 10945 16975 10955 17015
rect 10995 16975 11005 17015
rect 11045 16975 11055 17015
rect 11095 16975 11105 17015
rect 11145 16975 11155 17015
rect 11195 16975 11205 17015
rect 11245 16975 11255 17015
rect 11295 16975 11305 17015
rect 11345 16975 11355 17015
rect 11395 16975 11405 17015
rect 11445 16975 11455 17015
rect 11495 16975 11505 17015
rect 11545 16975 11555 17015
rect 11595 16975 11605 17015
rect 11645 16975 11655 17015
rect 11695 16975 11705 17015
rect 11745 16975 11755 17015
rect 11795 16975 11805 17015
rect 11845 16975 11855 17015
rect 11895 16975 11905 17015
rect 11945 16975 11955 17015
rect 11995 16975 12005 17015
rect 12045 16975 12055 17015
rect 12095 16975 12105 17015
rect 12145 16975 12155 17015
rect 12195 16975 12205 17015
rect 12245 16975 12255 17015
rect 12295 16975 12305 17015
rect 12345 16975 12355 17015
rect 12395 16975 12405 17015
rect 12445 16975 12455 17015
rect 12495 16975 12505 17015
rect 12545 16975 12555 17015
rect 12595 16975 12605 17015
rect 12645 16975 12655 17015
rect 12695 16975 12705 17015
rect 12745 16975 12755 17015
rect 12795 16975 12805 17015
rect 12845 16975 12855 17015
rect 12895 16975 12905 17015
rect 12945 16975 12955 17015
rect 12995 16975 13005 17015
rect 13045 16975 13055 17015
rect 13095 16975 13105 17015
rect 13145 16975 13155 17015
rect 13195 16975 13205 17015
rect 13245 16975 13255 17015
rect 13295 16975 13305 17015
rect 13345 16975 13355 17015
rect 13395 16975 13405 17015
rect 13445 16975 13455 17015
rect 13495 16975 13505 17015
rect 13545 16975 13555 17015
rect 13595 16975 13605 17015
rect 13645 16975 13655 17015
rect 13695 16975 13705 17015
rect 13745 16975 13755 17015
rect 13795 16975 13805 17015
rect 13845 16975 13855 17015
rect 13895 16975 13905 17015
rect 13945 16975 13955 17015
rect 13995 16975 14005 17015
rect 14045 16975 14055 17015
rect 14095 16975 14105 17015
rect 14145 16975 14155 17015
rect 14195 16975 14205 17015
rect 14245 16975 14255 17015
rect 14295 16975 14305 17015
rect 14345 16975 14355 17015
rect 14395 16975 14405 17015
rect 14445 16975 14455 17015
rect 14495 16975 14505 17015
rect 14545 16975 14555 17015
rect 14595 16975 14605 17015
rect 14645 16975 14655 17015
rect 14695 16975 14705 17015
rect 14745 16975 14755 17015
rect 14795 16975 14805 17015
rect 14845 16975 14855 17015
rect 14895 16975 14905 17015
rect 14945 16975 14955 17015
rect 14995 16975 15005 17015
rect 15045 16975 15055 17015
rect 15095 16975 15105 17015
rect 15145 16975 15155 17015
rect 15195 16975 15205 17015
rect 15245 16975 15255 17015
rect 15295 16975 15305 17015
rect 15345 16975 15355 17015
rect 15395 16975 15405 17015
rect 15445 16975 15455 17015
rect 15495 16975 15505 17015
rect 15545 16975 15555 17015
rect 15595 16975 15605 17015
rect 15645 16975 15655 17015
rect 15695 16975 15705 17015
rect 15745 16975 15755 17015
rect 15795 16975 15805 17015
rect 15845 16975 15855 17015
rect 15895 16975 15905 17015
rect 15945 16975 15955 17015
rect 15995 16975 16005 17015
rect 16045 16975 16055 17015
rect 16095 16975 16105 17015
rect 16145 16975 16155 17015
rect 16195 16975 16205 17015
rect 16245 16975 16255 17015
rect 16295 16975 16305 17015
rect 16345 16975 16355 17015
rect 16395 16975 16405 17015
rect 16445 16975 16455 17015
rect 16495 16975 16505 17015
rect 16545 16975 16555 17015
rect 16595 16975 16605 17015
rect 16645 16975 16655 17015
rect 16695 16975 16705 17015
rect 16745 16975 16755 17015
rect 16795 16975 16805 17015
rect 16845 16975 16855 17015
rect 16895 16975 16905 17015
rect 16945 16975 16955 17015
rect 16995 16975 17005 17015
rect 17045 16975 17055 17015
rect 17095 16975 17105 17015
rect 17145 16975 17155 17015
rect 17195 16975 17205 17015
rect 17245 16975 17255 17015
rect 17295 16975 17305 17015
rect 17345 16975 17355 17015
rect 17395 16975 17405 17015
rect 17445 16975 17455 17015
rect 17495 16975 17505 17015
rect 17545 16975 17555 17015
rect 17595 16975 17605 17015
rect 17645 16975 17655 17015
rect 17695 16975 17705 17015
rect 17745 16975 17755 17015
rect 17795 16975 17805 17015
rect 17845 16975 17855 17015
rect 17895 16975 17905 17015
rect 17945 16975 17955 17015
rect 17995 16975 18005 17015
rect 18045 16975 18055 17015
rect 18095 16975 18105 17015
rect 18145 16975 18155 17015
rect 18195 16975 18205 17015
rect 18245 16975 18255 17015
rect 18295 16975 18305 17015
rect 18345 16975 18355 17015
rect 18395 16975 18405 17015
rect 18445 16975 18455 17015
rect 18495 16975 18505 17015
rect 18545 16975 18555 17015
rect 18595 16975 18605 17015
rect 18645 16975 18655 17015
rect 18695 16975 18705 17015
rect 18745 16975 18755 17015
rect 18795 16975 18805 17015
rect 18845 16975 18855 17015
rect 18895 16975 18905 17015
rect 18945 16975 18955 17015
rect 18995 16975 19005 17015
rect 19045 16975 19055 17015
rect 19095 16975 19105 17015
rect 19145 16975 19155 17015
rect 19195 16975 19205 17015
rect 19245 16975 19255 17015
rect 19295 16975 19305 17015
rect 19345 16975 19355 17015
rect 19395 16975 19405 17015
rect 19445 16975 19455 17015
rect 19495 16975 19505 17015
rect 19545 16975 19555 17015
rect 19595 16975 19605 17015
rect 19645 16975 19655 17015
rect 19695 16975 19705 17015
rect 19745 16975 19755 17015
rect 19795 16975 19805 17015
rect 19845 16975 19855 17015
rect 19895 16975 19905 17015
rect 19945 16975 19955 17015
rect 19995 16975 20005 17015
rect 20045 16975 20055 17015
rect 20095 16975 20105 17015
rect 20145 16975 20155 17015
rect 20195 16975 20205 17015
rect 20245 16975 20255 17015
rect 20295 16975 20305 17015
rect 20345 16975 20355 17015
rect 20395 16975 20405 17015
rect 20445 16975 20455 17015
rect 20495 16975 20505 17015
rect 20545 16975 20555 17015
rect 20595 16975 20605 17015
rect 20645 16975 20655 17015
rect 20695 16975 20705 17015
rect 20745 16975 20755 17015
rect 20795 16975 20805 17015
rect 20845 16975 20855 17015
rect 20895 16975 20905 17015
rect 20945 16975 20955 17015
rect 20995 16975 21005 17015
rect 21045 16975 21055 17015
rect 21095 16975 21105 17015
rect 21145 16975 21155 17015
rect 21195 16975 21205 17015
rect 21245 16975 21255 17015
rect 21295 16975 21305 17015
rect 21345 16975 21355 17015
rect 21395 16975 21405 17015
rect 21445 16975 21455 17015
rect 21495 16975 21505 17015
rect 21545 16975 21555 17015
rect 21595 16975 21605 17015
rect 21645 16975 21655 17015
rect 21695 16975 21705 17015
rect 21745 16975 21755 17015
rect 21795 16975 21805 17015
rect 21845 16975 21855 17015
rect 21895 16975 21905 17015
rect 21945 16975 21955 17015
rect 21995 16975 22005 17015
rect 22045 16975 22055 17015
rect 22095 16975 22105 17015
rect 22145 16975 22155 17015
rect 22195 16975 22205 17015
rect 22245 16975 22255 17015
rect 22295 16975 22305 17015
rect 22345 16975 22355 17015
rect 22395 16975 22405 17015
rect 22445 16975 22455 17015
rect 22495 16975 22505 17015
rect 22545 16975 22555 17015
rect 22595 16975 22605 17015
rect 22645 16975 22655 17015
rect 22695 16975 22705 17015
rect 22745 16975 22755 17015
rect 22795 16975 22805 17015
rect 22845 16975 22855 17015
rect 22895 16975 22905 17015
rect 22945 16975 22955 17015
rect 22995 16975 23005 17015
rect 23045 16975 23055 17015
rect 23095 16975 23105 17015
rect 23145 16975 23155 17015
rect 23195 16975 23205 17015
rect 23245 16975 23255 17015
rect 23295 16975 23305 17015
rect 23345 16975 23355 17015
rect 23395 16975 23405 17015
rect 23445 16975 23455 17015
rect 23495 16975 23505 17015
rect 23545 16975 23555 17015
rect 23595 16975 23605 17015
rect 23645 16975 23655 17015
rect 23695 16975 23705 17015
rect 23745 16975 23755 17015
rect 23795 16975 23805 17015
rect 23845 16975 23855 17015
rect 23895 16975 23905 17015
rect 23945 16975 23955 17015
rect 23995 16975 24005 17015
rect 24045 16975 24055 17015
rect 24095 16975 24105 17015
rect 24145 16975 24155 17015
rect 24195 16975 24205 17015
rect 24245 16975 24255 17015
rect 24295 16975 24305 17015
rect 24345 16975 24355 17015
rect 24395 16975 24405 17015
rect 24445 16975 24455 17015
rect 24495 16975 24505 17015
rect 24545 16975 24555 17015
rect 24595 16975 24605 17015
rect 24645 16975 24655 17015
rect 24695 16975 24705 17015
rect 24745 16975 24755 17015
rect 24795 16975 24805 17015
rect 24845 16975 24855 17015
rect 24895 16975 24905 17015
rect 24945 16975 24955 17015
rect 24995 16975 25005 17015
rect 25045 16975 25055 17015
rect 25095 16975 25105 17015
rect 25145 16975 25155 17015
rect 25195 16975 25205 17015
rect 25245 16975 25255 17015
rect 25295 16975 25305 17015
rect 25345 16975 25355 17015
rect 25395 16975 25405 17015
rect 25445 16975 25455 17015
rect 25495 16975 25505 17015
rect 25545 16975 25555 17015
rect 25595 16975 25605 17015
rect 25645 16975 25655 17015
rect 25695 16975 25705 17015
rect 25745 16975 25755 17015
rect 25795 16975 25805 17015
rect 25845 16975 25855 17015
rect 25895 16975 25905 17015
rect 25945 16975 25955 17015
rect 25995 16975 26005 17015
rect 26045 16975 26055 17015
rect 26095 16975 26105 17015
rect 26145 16975 26155 17015
rect 26195 16975 26205 17015
rect 26245 16975 26255 17015
rect 26295 16975 26305 17015
rect 26345 16975 26355 17015
rect 26395 16975 26405 17015
rect 26445 16975 26455 17015
rect 26495 16975 26505 17015
rect 26545 16975 26555 17015
rect 26595 16975 26605 17015
rect 26645 16975 26655 17015
rect 26695 16975 26705 17015
rect 26745 16975 26755 17015
rect 26795 16975 26805 17015
rect 26845 16975 26855 17015
rect 26895 16975 26905 17015
rect 26945 16975 26955 17015
rect 26995 16975 27005 17015
rect 27045 16975 27055 17015
rect 27095 16975 27105 17015
rect 27145 16975 27155 17015
rect 27195 16975 27205 17015
rect 27245 16975 27255 17015
rect 27295 16975 27305 17015
rect 27345 16975 27355 17015
rect 27395 16975 27405 17015
rect 27445 16975 27455 17015
rect 27495 16975 27505 17015
rect 27545 16975 27555 17015
rect 27595 16975 27605 17015
rect 27645 16975 27655 17015
rect 27695 16975 27705 17015
rect 27745 16975 27755 17015
rect 27795 16975 27805 17015
rect 27845 16975 27855 17015
rect 27895 16975 27905 17015
rect 27945 16975 27955 17015
rect 27995 16975 28005 17015
rect 28045 16975 28055 17015
rect 28095 16975 28105 17015
rect 28145 16975 28155 17015
rect 28195 16975 28205 17015
rect 28245 16975 28255 17015
rect 28295 16975 28305 17015
rect 28345 16975 28355 17015
rect 28395 16975 28405 17015
rect 28445 16975 28455 17015
rect 28495 16975 28505 17015
rect 28545 16975 28555 17015
rect 28595 16975 28605 17015
rect 28645 16975 28655 17015
rect 28695 16975 28705 17015
rect 28745 16975 28755 17015
rect 28795 16975 28805 17015
rect 28845 16975 28855 17015
rect 28895 16975 28905 17015
rect 28945 16975 28955 17015
rect 28995 16975 29005 17015
rect 29045 16975 29055 17015
rect 29095 16975 29105 17015
rect 29145 16975 29155 17015
rect 29195 16975 29205 17015
rect 29245 16975 29255 17015
rect 29295 16975 29305 17015
rect 29345 16975 29355 17015
rect 29395 16975 29405 17015
rect 29445 16975 29455 17015
rect 29495 16975 29505 17015
rect 29545 16975 29555 17015
rect 29595 16975 29605 17015
rect 29645 16975 29655 17015
rect 29695 16975 29705 17015
rect 29745 16975 29755 17015
rect 29795 16975 29805 17015
rect 29845 16975 29855 17015
rect 29895 16975 29905 17015
rect 29945 16975 29955 17015
rect 29995 16975 30005 17015
rect 30045 16975 30055 17015
rect 30095 16975 30105 17015
rect 30145 16975 30155 17015
rect 30195 16975 30205 17015
rect 30245 16975 30255 17015
rect 30295 16975 30305 17015
rect 30345 16975 30355 17015
rect 30395 16975 30405 17015
rect 30445 16975 30455 17015
rect 30495 16975 30505 17015
rect 30545 16975 30555 17015
rect 30595 16975 30605 17015
rect 30645 16975 30655 17015
rect 30695 16975 30705 17015
rect 30745 16975 30755 17015
rect 30795 16975 30805 17015
rect 30845 16975 30855 17015
rect 30895 16975 30905 17015
rect 30945 16975 30955 17015
rect 30995 16975 31005 17015
rect 31045 16975 31055 17015
rect 31095 16975 31105 17015
rect 31145 16975 31155 17015
rect 31195 16975 31205 17015
rect 31245 16975 31255 17015
rect 31295 16975 31305 17015
rect 31345 16975 31355 17015
rect 31395 16975 31405 17015
rect 31445 16975 31455 17015
rect 31495 16975 31505 17015
rect 31545 16975 31555 17015
rect 31595 16975 31605 17015
rect 31645 16975 31655 17015
rect 31695 16975 31705 17015
rect 31745 16975 31755 17015
rect 31795 16975 31805 17015
rect 31845 16975 31855 17015
rect 31895 16975 31905 17015
rect 31945 16975 31955 17015
rect 31995 16975 32005 17015
rect 32045 16975 32055 17015
rect 32095 16975 32105 17015
rect 32145 16975 32155 17015
rect 32195 16975 32205 17015
rect 32245 16975 32255 17015
rect 32295 16975 32305 17015
rect 32345 16975 32355 17015
rect 32395 16975 32405 17015
rect 32445 16975 32455 17015
rect 32495 16975 32505 17015
rect 32545 16975 32555 17015
rect 32595 16975 32605 17015
rect 32645 16975 32655 17015
rect 32695 16975 32705 17015
rect 32745 16975 32755 17015
rect 32795 16975 32805 17015
rect 32845 16975 32855 17015
rect 32895 16975 32905 17015
rect 32945 16975 32955 17015
rect 32995 16975 33005 17015
rect 33045 16975 33055 17015
rect 33095 16975 33105 17015
rect 33145 16975 33155 17015
rect 33195 16975 33205 17015
rect 33245 16975 33255 17015
rect 33295 16975 33305 17015
rect 33345 16975 33355 17015
rect 33395 16975 33405 17015
rect 33445 16975 33455 17015
rect 33495 16975 33505 17015
rect 33545 16975 33555 17015
rect 33595 16975 33605 17015
rect 33645 16975 33655 17015
rect 33695 16975 33705 17015
rect 33745 16975 33755 17015
rect 33795 16975 33805 17015
rect 33845 16975 33855 17015
rect 33895 16975 33905 17015
rect 33945 16975 33955 17015
rect 33995 16975 34005 17015
rect 34045 16975 34055 17015
rect 34095 16975 34105 17015
rect 34145 16975 34155 17015
rect 34195 16975 34205 17015
rect 34245 16975 34255 17015
rect 34295 16975 34305 17015
rect 34345 16975 34355 17015
rect 34395 16975 34405 17015
rect 34445 16975 34455 17015
rect 34495 16975 34505 17015
rect 34545 16975 34555 17015
rect 34595 16975 34605 17015
rect 34645 16975 34655 17015
rect 34695 16975 34705 17015
rect 34745 16975 34755 17015
rect 34795 16975 34805 17015
rect 34845 16975 34855 17015
rect 34895 16975 34905 17015
rect 34945 16975 34955 17015
rect 34995 16975 35005 17015
rect 35045 16975 35055 17015
rect 35095 16975 35105 17015
rect 35145 16975 35155 17015
rect 35195 16975 35205 17015
rect 35245 16975 35255 17015
rect 35295 16975 35305 17015
rect 35345 16975 35355 17015
rect 35395 16975 35405 17015
rect 35445 16975 35455 17015
rect 35495 16975 35505 17015
rect 35545 16975 35555 17015
rect 35595 16975 35605 17015
rect 35645 16975 35655 17015
rect 35695 16975 35705 17015
rect 35745 16975 35755 17015
rect 35795 16975 35805 17015
rect 35845 16975 35855 17015
rect 35895 16975 35905 17015
rect 35945 16975 35955 17015
rect 35995 16975 36005 17015
rect 36045 16975 36055 17015
rect 36095 16975 36105 17015
rect 36145 16975 36155 17015
rect 36195 16975 36205 17015
rect 36245 16975 36255 17015
rect 36295 16975 36305 17015
rect 36345 16975 36355 17015
rect 36395 16975 36405 17015
rect 36445 16975 36455 17015
rect 36495 16975 36505 17015
rect 36545 16975 36555 17015
rect 36595 16975 36605 17015
rect 36645 16975 36655 17015
rect 36695 16975 36705 17015
rect 36745 16975 36755 17015
rect 36795 16975 36805 17015
rect 36845 16975 36855 17015
rect 36895 16975 36905 17015
rect 36945 16975 36955 17015
rect 36995 16975 37005 17015
rect 37045 16975 37055 17015
rect 37095 16975 37105 17015
rect 37145 16975 37155 17015
rect 37195 16975 37205 17015
rect 37245 16975 37255 17015
rect 37295 16975 37305 17015
rect 37345 16975 37355 17015
rect 37395 16975 37405 17015
rect 37445 16975 37455 17015
rect 37495 16975 37505 17015
rect 37545 16975 37555 17015
rect 37595 16975 37605 17015
rect 37645 16975 37655 17015
rect 37695 16975 37705 17015
rect 37745 16975 37755 17015
rect 37795 16975 37805 17015
rect 37845 16975 37855 17015
rect 37895 16975 37905 17015
rect 37945 16975 37955 17015
rect 37995 16975 38005 17015
rect 38045 16975 38055 17015
rect 38095 16975 38105 17015
rect 38145 16975 38155 17015
rect 38195 16975 38205 17015
rect 38245 16975 38255 17015
rect 38295 16975 38305 17015
rect 38345 16975 38355 17015
rect 38395 16975 38405 17015
rect 38445 16975 38455 17015
rect 38495 16975 38505 17015
rect 38545 16975 38555 17015
rect 38595 16975 38605 17015
rect 38645 16975 38655 17015
rect 38695 16975 38705 17015
rect 38745 16975 38755 17015
rect 38795 16975 38805 17015
rect 38845 16975 38855 17015
rect 38895 16975 38905 17015
rect 38945 16975 38955 17015
rect 38995 16975 39005 17015
rect 39045 16975 39055 17015
rect 39095 16975 39105 17015
rect 39145 16975 39155 17015
rect 39195 16975 39205 17015
rect 39245 16975 39255 17015
rect 39295 16975 39305 17015
rect 39345 16975 39355 17015
rect 39395 16975 39405 17015
rect 39445 16975 39455 17015
rect 39495 16975 39505 17015
rect 39545 16975 39555 17015
rect 39595 16975 39605 17015
rect 39645 16975 39655 17015
rect 39695 16975 39705 17015
rect 39745 16975 39750 17015
rect 0 16970 39750 16975
rect 0 15850 50 16970
rect 100 16915 39750 16920
rect 100 16875 105 16915
rect 145 16875 155 16915
rect 195 16875 205 16915
rect 245 16875 255 16915
rect 295 16875 305 16915
rect 345 16875 355 16915
rect 395 16875 405 16915
rect 445 16875 455 16915
rect 495 16875 505 16915
rect 545 16875 555 16915
rect 595 16875 605 16915
rect 645 16875 655 16915
rect 695 16875 705 16915
rect 745 16875 755 16915
rect 795 16875 805 16915
rect 845 16875 855 16915
rect 895 16875 905 16915
rect 945 16875 955 16915
rect 995 16875 1005 16915
rect 1045 16875 1055 16915
rect 1095 16875 1105 16915
rect 1145 16875 1155 16915
rect 1195 16875 1205 16915
rect 1245 16875 1255 16915
rect 1295 16875 1305 16915
rect 1345 16875 1355 16915
rect 1395 16875 1405 16915
rect 1445 16875 1455 16915
rect 1495 16875 1505 16915
rect 1545 16875 1555 16915
rect 1595 16875 1605 16915
rect 1645 16875 1655 16915
rect 1695 16875 1705 16915
rect 1745 16875 1755 16915
rect 1795 16875 1805 16915
rect 1845 16875 1855 16915
rect 1895 16875 1905 16915
rect 1945 16875 1955 16915
rect 1995 16875 2005 16915
rect 2045 16875 2055 16915
rect 2095 16875 2105 16915
rect 2145 16875 2155 16915
rect 2195 16875 2205 16915
rect 2245 16875 2255 16915
rect 2295 16875 2305 16915
rect 2345 16875 2355 16915
rect 2395 16875 2405 16915
rect 2445 16875 2455 16915
rect 2495 16875 2505 16915
rect 2545 16875 2555 16915
rect 2595 16875 2605 16915
rect 2645 16875 2655 16915
rect 2695 16875 2705 16915
rect 2745 16875 2755 16915
rect 2795 16875 2805 16915
rect 2845 16875 2855 16915
rect 2895 16875 2905 16915
rect 2945 16875 2955 16915
rect 2995 16875 3005 16915
rect 3045 16875 3055 16915
rect 3095 16875 3105 16915
rect 3145 16875 3155 16915
rect 3195 16875 3205 16915
rect 3245 16875 3255 16915
rect 3295 16875 3305 16915
rect 3345 16875 3355 16915
rect 3395 16875 3405 16915
rect 3445 16875 3455 16915
rect 3495 16875 3505 16915
rect 3545 16875 3555 16915
rect 3595 16875 3605 16915
rect 3645 16875 3655 16915
rect 3695 16875 3705 16915
rect 3745 16875 3755 16915
rect 3795 16875 3805 16915
rect 3845 16875 3855 16915
rect 3895 16875 3905 16915
rect 3945 16875 3955 16915
rect 3995 16875 4005 16915
rect 4045 16875 4055 16915
rect 4095 16875 4105 16915
rect 4145 16875 4155 16915
rect 4195 16875 4205 16915
rect 4245 16875 4255 16915
rect 4295 16875 4305 16915
rect 4345 16875 4355 16915
rect 4395 16875 4405 16915
rect 4445 16875 4455 16915
rect 4495 16875 4505 16915
rect 4545 16875 4555 16915
rect 4595 16875 4605 16915
rect 4645 16875 4655 16915
rect 4695 16875 4705 16915
rect 4745 16875 4755 16915
rect 4795 16875 4805 16915
rect 4845 16875 4855 16915
rect 4895 16875 4905 16915
rect 4945 16875 4955 16915
rect 4995 16875 5005 16915
rect 5045 16875 5055 16915
rect 5095 16875 5105 16915
rect 5145 16875 5155 16915
rect 5195 16875 5205 16915
rect 5245 16875 5255 16915
rect 5295 16875 5305 16915
rect 5345 16875 5355 16915
rect 5395 16875 5405 16915
rect 5445 16875 5455 16915
rect 5495 16875 5505 16915
rect 5545 16875 5555 16915
rect 5595 16875 5605 16915
rect 5645 16875 5655 16915
rect 5695 16875 5705 16915
rect 5745 16875 5755 16915
rect 5795 16875 5805 16915
rect 5845 16875 5855 16915
rect 5895 16875 5905 16915
rect 5945 16875 5955 16915
rect 5995 16875 6005 16915
rect 6045 16875 6055 16915
rect 6095 16875 6105 16915
rect 6145 16875 6155 16915
rect 6195 16875 6205 16915
rect 6245 16875 6255 16915
rect 6295 16875 6305 16915
rect 6345 16875 6355 16915
rect 6395 16875 6405 16915
rect 6445 16875 6455 16915
rect 6495 16875 6505 16915
rect 6545 16875 6555 16915
rect 6595 16875 6605 16915
rect 6645 16875 6655 16915
rect 6695 16875 6705 16915
rect 6745 16875 6755 16915
rect 6795 16875 6805 16915
rect 6845 16875 6855 16915
rect 6895 16875 6905 16915
rect 6945 16875 6955 16915
rect 6995 16875 7005 16915
rect 7045 16875 7055 16915
rect 7095 16875 7105 16915
rect 7145 16875 7155 16915
rect 7195 16875 7205 16915
rect 7245 16875 7255 16915
rect 7295 16875 7305 16915
rect 7345 16875 7355 16915
rect 7395 16875 7405 16915
rect 7445 16875 7455 16915
rect 7495 16875 7505 16915
rect 7545 16875 7555 16915
rect 7595 16875 7605 16915
rect 7645 16875 7655 16915
rect 7695 16875 7705 16915
rect 7745 16875 7755 16915
rect 7795 16875 7805 16915
rect 7845 16875 7855 16915
rect 7895 16875 7905 16915
rect 7945 16875 7955 16915
rect 7995 16875 8005 16915
rect 8045 16875 8055 16915
rect 8095 16875 8105 16915
rect 8145 16875 8155 16915
rect 8195 16875 8205 16915
rect 8245 16875 8255 16915
rect 8295 16875 8305 16915
rect 8345 16875 8355 16915
rect 8395 16875 8405 16915
rect 8445 16875 8455 16915
rect 8495 16875 8505 16915
rect 8545 16875 8555 16915
rect 8595 16875 8605 16915
rect 8645 16875 8655 16915
rect 8695 16875 8705 16915
rect 8745 16875 8755 16915
rect 8795 16875 8805 16915
rect 8845 16875 8855 16915
rect 8895 16875 8905 16915
rect 8945 16875 8955 16915
rect 8995 16875 9005 16915
rect 9045 16875 9055 16915
rect 9095 16875 9105 16915
rect 9145 16875 9155 16915
rect 9195 16875 9205 16915
rect 9245 16875 9255 16915
rect 9295 16875 9305 16915
rect 9345 16875 9355 16915
rect 9395 16875 9405 16915
rect 9445 16875 9455 16915
rect 9495 16875 9505 16915
rect 9545 16875 9555 16915
rect 9595 16875 9605 16915
rect 9645 16875 9655 16915
rect 9695 16875 9705 16915
rect 9745 16875 9755 16915
rect 9795 16875 9805 16915
rect 9845 16875 9855 16915
rect 9895 16875 9905 16915
rect 9945 16875 9955 16915
rect 9995 16875 10005 16915
rect 10045 16875 10055 16915
rect 10095 16875 10105 16915
rect 10145 16875 10155 16915
rect 10195 16875 10205 16915
rect 10245 16875 10255 16915
rect 10295 16875 10305 16915
rect 10345 16875 10355 16915
rect 10395 16875 10405 16915
rect 10445 16875 10455 16915
rect 10495 16875 10505 16915
rect 10545 16875 10555 16915
rect 10595 16875 10605 16915
rect 10645 16875 10655 16915
rect 10695 16875 10705 16915
rect 10745 16875 10755 16915
rect 10795 16875 10805 16915
rect 10845 16875 10855 16915
rect 10895 16875 10905 16915
rect 10945 16875 10955 16915
rect 10995 16875 11005 16915
rect 11045 16875 11055 16915
rect 11095 16875 11105 16915
rect 11145 16875 11155 16915
rect 11195 16875 11205 16915
rect 11245 16875 11255 16915
rect 11295 16875 11305 16915
rect 11345 16875 11355 16915
rect 11395 16875 11405 16915
rect 11445 16875 11455 16915
rect 11495 16875 11505 16915
rect 11545 16875 11555 16915
rect 11595 16875 11605 16915
rect 11645 16875 11655 16915
rect 11695 16875 11705 16915
rect 11745 16875 11755 16915
rect 11795 16875 11805 16915
rect 11845 16875 11855 16915
rect 11895 16875 11905 16915
rect 11945 16875 11955 16915
rect 11995 16875 12005 16915
rect 12045 16875 12055 16915
rect 12095 16875 12105 16915
rect 12145 16875 12155 16915
rect 12195 16875 12205 16915
rect 12245 16875 12255 16915
rect 12295 16875 12305 16915
rect 12345 16875 12355 16915
rect 12395 16875 12405 16915
rect 12445 16875 12455 16915
rect 12495 16875 12505 16915
rect 12545 16875 12555 16915
rect 12595 16875 12605 16915
rect 12645 16875 12655 16915
rect 12695 16875 12705 16915
rect 12745 16875 12755 16915
rect 12795 16875 12805 16915
rect 12845 16875 12855 16915
rect 12895 16875 12905 16915
rect 12945 16875 12955 16915
rect 12995 16875 13005 16915
rect 13045 16875 13055 16915
rect 13095 16875 13105 16915
rect 13145 16875 13155 16915
rect 13195 16875 13205 16915
rect 13245 16875 13255 16915
rect 13295 16875 13305 16915
rect 13345 16875 13355 16915
rect 13395 16875 13405 16915
rect 13445 16875 13455 16915
rect 13495 16875 13505 16915
rect 13545 16875 13555 16915
rect 13595 16875 13605 16915
rect 13645 16875 13655 16915
rect 13695 16875 13705 16915
rect 13745 16875 13755 16915
rect 13795 16875 13805 16915
rect 13845 16875 13855 16915
rect 13895 16875 13905 16915
rect 13945 16875 13955 16915
rect 13995 16875 14005 16915
rect 14045 16875 14055 16915
rect 14095 16875 14105 16915
rect 14145 16875 14155 16915
rect 14195 16875 14205 16915
rect 14245 16875 14255 16915
rect 14295 16875 14305 16915
rect 14345 16875 14355 16915
rect 14395 16875 14405 16915
rect 14445 16875 14455 16915
rect 14495 16875 14505 16915
rect 14545 16875 14555 16915
rect 14595 16875 14605 16915
rect 14645 16875 14655 16915
rect 14695 16875 14705 16915
rect 14745 16875 14755 16915
rect 14795 16875 14805 16915
rect 14845 16875 14855 16915
rect 14895 16875 14905 16915
rect 14945 16875 14955 16915
rect 14995 16875 15005 16915
rect 15045 16875 15055 16915
rect 15095 16875 15105 16915
rect 15145 16875 15155 16915
rect 15195 16875 15205 16915
rect 15245 16875 15255 16915
rect 15295 16875 15305 16915
rect 15345 16875 15355 16915
rect 15395 16875 15405 16915
rect 15445 16875 15455 16915
rect 15495 16875 15505 16915
rect 15545 16875 15555 16915
rect 15595 16875 15605 16915
rect 15645 16875 15655 16915
rect 15695 16875 15705 16915
rect 15745 16875 15755 16915
rect 15795 16875 15805 16915
rect 15845 16875 15855 16915
rect 15895 16875 15905 16915
rect 15945 16875 15955 16915
rect 15995 16875 16005 16915
rect 16045 16875 16055 16915
rect 16095 16875 16105 16915
rect 16145 16875 16155 16915
rect 16195 16875 16205 16915
rect 16245 16875 16255 16915
rect 16295 16875 16305 16915
rect 16345 16875 16355 16915
rect 16395 16875 16405 16915
rect 16445 16875 16455 16915
rect 16495 16875 16505 16915
rect 16545 16875 16555 16915
rect 16595 16875 16605 16915
rect 16645 16875 16655 16915
rect 16695 16875 16705 16915
rect 16745 16875 16755 16915
rect 16795 16875 16805 16915
rect 16845 16875 16855 16915
rect 16895 16875 16905 16915
rect 16945 16875 16955 16915
rect 16995 16875 17005 16915
rect 17045 16875 17055 16915
rect 17095 16875 17105 16915
rect 17145 16875 17155 16915
rect 17195 16875 17205 16915
rect 17245 16875 17255 16915
rect 17295 16875 17305 16915
rect 17345 16875 17355 16915
rect 17395 16875 17405 16915
rect 17445 16875 17455 16915
rect 17495 16875 17505 16915
rect 17545 16875 17555 16915
rect 17595 16875 17605 16915
rect 17645 16875 17655 16915
rect 17695 16875 17705 16915
rect 17745 16875 17755 16915
rect 17795 16875 17805 16915
rect 17845 16875 17855 16915
rect 17895 16875 17905 16915
rect 17945 16875 17955 16915
rect 17995 16875 18005 16915
rect 18045 16875 18055 16915
rect 18095 16875 18105 16915
rect 18145 16875 18155 16915
rect 18195 16875 18205 16915
rect 18245 16875 18255 16915
rect 18295 16875 18305 16915
rect 18345 16875 18355 16915
rect 18395 16875 18405 16915
rect 18445 16875 18455 16915
rect 18495 16875 18505 16915
rect 18545 16875 18555 16915
rect 18595 16875 18605 16915
rect 18645 16875 18655 16915
rect 18695 16875 18705 16915
rect 18745 16875 18755 16915
rect 18795 16875 18805 16915
rect 18845 16875 18855 16915
rect 18895 16875 18905 16915
rect 18945 16875 18955 16915
rect 18995 16875 19005 16915
rect 19045 16875 19055 16915
rect 19095 16875 19105 16915
rect 19145 16875 19155 16915
rect 19195 16875 19205 16915
rect 19245 16875 19255 16915
rect 19295 16875 19305 16915
rect 19345 16875 19355 16915
rect 19395 16875 19405 16915
rect 19445 16875 19455 16915
rect 19495 16875 19505 16915
rect 19545 16875 19555 16915
rect 19595 16875 19605 16915
rect 19645 16875 19655 16915
rect 19695 16875 19705 16915
rect 19745 16875 19755 16915
rect 19795 16875 19805 16915
rect 19845 16875 19855 16915
rect 19895 16875 19905 16915
rect 19945 16875 19955 16915
rect 19995 16875 20005 16915
rect 20045 16875 20055 16915
rect 20095 16875 20105 16915
rect 20145 16875 20155 16915
rect 20195 16875 20205 16915
rect 20245 16875 20255 16915
rect 20295 16875 20305 16915
rect 20345 16875 20355 16915
rect 20395 16875 20405 16915
rect 20445 16875 20455 16915
rect 20495 16875 20505 16915
rect 20545 16875 20555 16915
rect 20595 16875 20605 16915
rect 20645 16875 20655 16915
rect 20695 16875 20705 16915
rect 20745 16875 20755 16915
rect 20795 16875 20805 16915
rect 20845 16875 20855 16915
rect 20895 16875 20905 16915
rect 20945 16875 20955 16915
rect 20995 16875 21005 16915
rect 21045 16875 21055 16915
rect 21095 16875 21105 16915
rect 21145 16875 21155 16915
rect 21195 16875 21205 16915
rect 21245 16875 21255 16915
rect 21295 16875 21305 16915
rect 21345 16875 21355 16915
rect 21395 16875 21405 16915
rect 21445 16875 21455 16915
rect 21495 16875 21505 16915
rect 21545 16875 21555 16915
rect 21595 16875 21605 16915
rect 21645 16875 21655 16915
rect 21695 16875 21705 16915
rect 21745 16875 21755 16915
rect 21795 16875 21805 16915
rect 21845 16875 21855 16915
rect 21895 16875 21905 16915
rect 21945 16875 21955 16915
rect 21995 16875 22005 16915
rect 22045 16875 22055 16915
rect 22095 16875 22105 16915
rect 22145 16875 22155 16915
rect 22195 16875 22205 16915
rect 22245 16875 22255 16915
rect 22295 16875 22305 16915
rect 22345 16875 22355 16915
rect 22395 16875 22405 16915
rect 22445 16875 22455 16915
rect 22495 16875 22505 16915
rect 22545 16875 22555 16915
rect 22595 16875 22605 16915
rect 22645 16875 22655 16915
rect 22695 16875 22705 16915
rect 22745 16875 22755 16915
rect 22795 16875 22805 16915
rect 22845 16875 22855 16915
rect 22895 16875 22905 16915
rect 22945 16875 22955 16915
rect 22995 16875 23005 16915
rect 23045 16875 23055 16915
rect 23095 16875 23105 16915
rect 23145 16875 23155 16915
rect 23195 16875 23205 16915
rect 23245 16875 23255 16915
rect 23295 16875 23305 16915
rect 23345 16875 23355 16915
rect 23395 16875 23405 16915
rect 23445 16875 23455 16915
rect 23495 16875 23505 16915
rect 23545 16875 23555 16915
rect 23595 16875 23605 16915
rect 23645 16875 23655 16915
rect 23695 16875 23705 16915
rect 23745 16875 23755 16915
rect 23795 16875 23805 16915
rect 23845 16875 23855 16915
rect 23895 16875 23905 16915
rect 23945 16875 23955 16915
rect 23995 16875 24005 16915
rect 24045 16875 24055 16915
rect 24095 16875 24105 16915
rect 24145 16875 24155 16915
rect 24195 16875 24205 16915
rect 24245 16875 24255 16915
rect 24295 16875 24305 16915
rect 24345 16875 24355 16915
rect 24395 16875 24405 16915
rect 24445 16875 24455 16915
rect 24495 16875 24505 16915
rect 24545 16875 24555 16915
rect 24595 16875 24605 16915
rect 24645 16875 24655 16915
rect 24695 16875 24705 16915
rect 24745 16875 24755 16915
rect 24795 16875 24805 16915
rect 24845 16875 24855 16915
rect 24895 16875 24905 16915
rect 24945 16875 24955 16915
rect 24995 16875 25005 16915
rect 25045 16875 25055 16915
rect 25095 16875 25105 16915
rect 25145 16875 25155 16915
rect 25195 16875 25205 16915
rect 25245 16875 25255 16915
rect 25295 16875 25305 16915
rect 25345 16875 25355 16915
rect 25395 16875 25405 16915
rect 25445 16875 25455 16915
rect 25495 16875 25505 16915
rect 25545 16875 25555 16915
rect 25595 16875 25605 16915
rect 25645 16875 25655 16915
rect 25695 16875 25705 16915
rect 25745 16875 25755 16915
rect 25795 16875 25805 16915
rect 25845 16875 25855 16915
rect 25895 16875 25905 16915
rect 25945 16875 25955 16915
rect 25995 16875 26005 16915
rect 26045 16875 26055 16915
rect 26095 16875 26105 16915
rect 26145 16875 26155 16915
rect 26195 16875 26205 16915
rect 26245 16875 26255 16915
rect 26295 16875 26305 16915
rect 26345 16875 26355 16915
rect 26395 16875 26405 16915
rect 26445 16875 26455 16915
rect 26495 16875 26505 16915
rect 26545 16875 26555 16915
rect 26595 16875 26605 16915
rect 26645 16875 26655 16915
rect 26695 16875 26705 16915
rect 26745 16875 26755 16915
rect 26795 16875 26805 16915
rect 26845 16875 26855 16915
rect 26895 16875 26905 16915
rect 26945 16875 26955 16915
rect 26995 16875 27005 16915
rect 27045 16875 27055 16915
rect 27095 16875 27105 16915
rect 27145 16875 27155 16915
rect 27195 16875 27205 16915
rect 27245 16875 27255 16915
rect 27295 16875 27305 16915
rect 27345 16875 27355 16915
rect 27395 16875 27405 16915
rect 27445 16875 27455 16915
rect 27495 16875 27505 16915
rect 27545 16875 27555 16915
rect 27595 16875 27605 16915
rect 27645 16875 27655 16915
rect 27695 16875 27705 16915
rect 27745 16875 27755 16915
rect 27795 16875 27805 16915
rect 27845 16875 27855 16915
rect 27895 16875 27905 16915
rect 27945 16875 27955 16915
rect 27995 16875 28005 16915
rect 28045 16875 28055 16915
rect 28095 16875 28105 16915
rect 28145 16875 28155 16915
rect 28195 16875 28205 16915
rect 28245 16875 28255 16915
rect 28295 16875 28305 16915
rect 28345 16875 28355 16915
rect 28395 16875 28405 16915
rect 28445 16875 28455 16915
rect 28495 16875 28505 16915
rect 28545 16875 28555 16915
rect 28595 16875 28605 16915
rect 28645 16875 28655 16915
rect 28695 16875 28705 16915
rect 28745 16875 28755 16915
rect 28795 16875 28805 16915
rect 28845 16875 28855 16915
rect 28895 16875 28905 16915
rect 28945 16875 28955 16915
rect 28995 16875 29005 16915
rect 29045 16875 29055 16915
rect 29095 16875 29105 16915
rect 29145 16875 29155 16915
rect 29195 16875 29205 16915
rect 29245 16875 29255 16915
rect 29295 16875 29305 16915
rect 29345 16875 29355 16915
rect 29395 16875 29405 16915
rect 29445 16875 29455 16915
rect 29495 16875 29505 16915
rect 29545 16875 29555 16915
rect 29595 16875 29605 16915
rect 29645 16875 29655 16915
rect 29695 16875 29705 16915
rect 29745 16875 29755 16915
rect 29795 16875 29805 16915
rect 29845 16875 29855 16915
rect 29895 16875 29905 16915
rect 29945 16875 29955 16915
rect 29995 16875 30005 16915
rect 30045 16875 30055 16915
rect 30095 16875 30105 16915
rect 30145 16875 30155 16915
rect 30195 16875 30205 16915
rect 30245 16875 30255 16915
rect 30295 16875 30305 16915
rect 30345 16875 30355 16915
rect 30395 16875 30405 16915
rect 30445 16875 30455 16915
rect 30495 16875 30505 16915
rect 30545 16875 30555 16915
rect 30595 16875 30605 16915
rect 30645 16875 30655 16915
rect 30695 16875 30705 16915
rect 30745 16875 30755 16915
rect 30795 16875 30805 16915
rect 30845 16875 30855 16915
rect 30895 16875 30905 16915
rect 30945 16875 30955 16915
rect 30995 16875 31005 16915
rect 31045 16875 31055 16915
rect 31095 16875 31105 16915
rect 31145 16875 31155 16915
rect 31195 16875 31205 16915
rect 31245 16875 31255 16915
rect 31295 16875 31305 16915
rect 31345 16875 31355 16915
rect 31395 16875 31405 16915
rect 31445 16875 31455 16915
rect 31495 16875 31505 16915
rect 31545 16875 31555 16915
rect 31595 16875 31605 16915
rect 31645 16875 31655 16915
rect 31695 16875 31705 16915
rect 31745 16875 31755 16915
rect 31795 16875 31805 16915
rect 31845 16875 31855 16915
rect 31895 16875 31905 16915
rect 31945 16875 31955 16915
rect 31995 16875 32005 16915
rect 32045 16875 32055 16915
rect 32095 16875 32105 16915
rect 32145 16875 32155 16915
rect 32195 16875 32205 16915
rect 32245 16875 32255 16915
rect 32295 16875 32305 16915
rect 32345 16875 32355 16915
rect 32395 16875 32405 16915
rect 32445 16875 32455 16915
rect 32495 16875 32505 16915
rect 32545 16875 32555 16915
rect 32595 16875 32605 16915
rect 32645 16875 32655 16915
rect 32695 16875 32705 16915
rect 32745 16875 32755 16915
rect 32795 16875 32805 16915
rect 32845 16875 32855 16915
rect 32895 16875 32905 16915
rect 32945 16875 32955 16915
rect 32995 16875 33005 16915
rect 33045 16875 33055 16915
rect 33095 16875 33105 16915
rect 33145 16875 33155 16915
rect 33195 16875 33205 16915
rect 33245 16875 33255 16915
rect 33295 16875 33305 16915
rect 33345 16875 33355 16915
rect 33395 16875 33405 16915
rect 33445 16875 33455 16915
rect 33495 16875 33505 16915
rect 33545 16875 33555 16915
rect 33595 16875 33605 16915
rect 33645 16875 33655 16915
rect 33695 16875 33705 16915
rect 33745 16875 33755 16915
rect 33795 16875 33805 16915
rect 33845 16875 33855 16915
rect 33895 16875 33905 16915
rect 33945 16875 33955 16915
rect 33995 16875 34005 16915
rect 34045 16875 34055 16915
rect 34095 16875 34105 16915
rect 34145 16875 34155 16915
rect 34195 16875 34205 16915
rect 34245 16875 34255 16915
rect 34295 16875 34305 16915
rect 34345 16875 34355 16915
rect 34395 16875 34405 16915
rect 34445 16875 34455 16915
rect 34495 16875 34505 16915
rect 34545 16875 34555 16915
rect 34595 16875 34605 16915
rect 34645 16875 34655 16915
rect 34695 16875 34705 16915
rect 34745 16875 34755 16915
rect 34795 16875 34805 16915
rect 34845 16875 34855 16915
rect 34895 16875 34905 16915
rect 34945 16875 34955 16915
rect 34995 16875 35005 16915
rect 35045 16875 35055 16915
rect 35095 16875 35105 16915
rect 35145 16875 35155 16915
rect 35195 16875 35205 16915
rect 35245 16875 35255 16915
rect 35295 16875 35305 16915
rect 35345 16875 35355 16915
rect 35395 16875 35405 16915
rect 35445 16875 35455 16915
rect 35495 16875 35505 16915
rect 35545 16875 35555 16915
rect 35595 16875 35605 16915
rect 35645 16875 35655 16915
rect 35695 16875 35705 16915
rect 35745 16875 35755 16915
rect 35795 16875 35805 16915
rect 35845 16875 35855 16915
rect 35895 16875 35905 16915
rect 35945 16875 35955 16915
rect 35995 16875 36005 16915
rect 36045 16875 36055 16915
rect 36095 16875 36105 16915
rect 36145 16875 36155 16915
rect 36195 16875 36205 16915
rect 36245 16875 36255 16915
rect 36295 16875 36305 16915
rect 36345 16875 36355 16915
rect 36395 16875 36405 16915
rect 36445 16875 36455 16915
rect 36495 16875 36505 16915
rect 36545 16875 36555 16915
rect 36595 16875 36605 16915
rect 36645 16875 36655 16915
rect 36695 16875 36705 16915
rect 36745 16875 36755 16915
rect 36795 16875 36805 16915
rect 36845 16875 36855 16915
rect 36895 16875 36905 16915
rect 36945 16875 36955 16915
rect 36995 16875 37005 16915
rect 37045 16875 37055 16915
rect 37095 16875 37105 16915
rect 37145 16875 37155 16915
rect 37195 16875 37205 16915
rect 37245 16875 37255 16915
rect 37295 16875 37305 16915
rect 37345 16875 37355 16915
rect 37395 16875 37405 16915
rect 37445 16875 37455 16915
rect 37495 16875 37505 16915
rect 37545 16875 37555 16915
rect 37595 16875 37605 16915
rect 37645 16875 37655 16915
rect 37695 16875 37705 16915
rect 37745 16875 37755 16915
rect 37795 16875 37805 16915
rect 37845 16875 37855 16915
rect 37895 16875 37905 16915
rect 37945 16875 37955 16915
rect 37995 16875 38005 16915
rect 38045 16875 38055 16915
rect 38095 16875 38105 16915
rect 38145 16875 38155 16915
rect 38195 16875 38205 16915
rect 38245 16875 38255 16915
rect 38295 16875 38305 16915
rect 38345 16875 38355 16915
rect 38395 16875 38405 16915
rect 38445 16875 38455 16915
rect 38495 16875 38505 16915
rect 38545 16875 38555 16915
rect 38595 16875 38605 16915
rect 38645 16875 38655 16915
rect 38695 16875 38705 16915
rect 38745 16875 38755 16915
rect 38795 16875 38805 16915
rect 38845 16875 38855 16915
rect 38895 16875 38905 16915
rect 38945 16875 38955 16915
rect 38995 16875 39005 16915
rect 39045 16875 39055 16915
rect 39095 16875 39105 16915
rect 39145 16875 39155 16915
rect 39195 16875 39205 16915
rect 39245 16875 39255 16915
rect 39295 16875 39305 16915
rect 39345 16875 39355 16915
rect 39395 16875 39405 16915
rect 39445 16875 39455 16915
rect 39495 16875 39505 16915
rect 39545 16875 39555 16915
rect 39595 16875 39605 16915
rect 39645 16875 39655 16915
rect 39695 16875 39705 16915
rect 39745 16875 39750 16915
rect 100 16870 39750 16875
rect 100 16650 3200 16870
rect 100 16000 200 16650
rect 3100 16000 3200 16650
rect 100 15900 3200 16000
rect 3350 16650 6450 16870
rect 3350 16000 3450 16650
rect 6350 16000 6450 16650
rect 3350 15900 6450 16000
rect 6600 16650 9700 16870
rect 6600 16000 6700 16650
rect 9600 16000 9700 16650
rect 6600 15900 9700 16000
rect 9850 16650 12950 16870
rect 9850 16000 9950 16650
rect 12850 16000 12950 16650
rect 9850 15900 12950 16000
rect 13100 16650 16200 16870
rect 13100 16000 13200 16650
rect 16100 16000 16200 16650
rect 13100 15900 16200 16000
rect 16350 16650 19450 16870
rect 16350 16000 16450 16650
rect 19350 16000 19450 16650
rect 16350 15900 19450 16000
rect 19600 16650 22700 16870
rect 19600 16000 19700 16650
rect 22600 16000 22700 16650
rect 19600 15900 22700 16000
rect 22850 16650 25950 16870
rect 22850 16000 22950 16650
rect 25850 16000 25950 16650
rect 22850 15900 25950 16000
rect 26100 16650 29200 16870
rect 26100 16000 26200 16650
rect 29100 16000 29200 16650
rect 26100 15900 29200 16000
rect 29350 16650 32450 16870
rect 29350 16000 29450 16650
rect 32350 16000 32450 16650
rect 29350 15900 32450 16000
rect 32600 16650 35700 16870
rect 32600 16000 32700 16650
rect 35600 16000 35700 16650
rect 32600 15900 35700 16000
rect 35850 16650 38950 16870
rect 35850 16000 35950 16650
rect 38850 16000 38950 16650
rect 35850 15900 38950 16000
rect 39100 16650 39750 16870
rect 39100 16000 39200 16650
rect 39650 16000 39750 16650
rect 39100 15900 39750 16000
rect 0 15845 39750 15850
rect 0 15805 5 15845
rect 45 15805 55 15845
rect 95 15805 105 15845
rect 145 15805 155 15845
rect 195 15805 205 15845
rect 245 15805 255 15845
rect 295 15805 305 15845
rect 345 15805 355 15845
rect 395 15805 405 15845
rect 445 15805 455 15845
rect 495 15805 505 15845
rect 545 15805 555 15845
rect 595 15805 605 15845
rect 645 15805 655 15845
rect 695 15805 705 15845
rect 745 15805 755 15845
rect 795 15805 805 15845
rect 845 15805 855 15845
rect 895 15805 905 15845
rect 945 15805 955 15845
rect 995 15805 1005 15845
rect 1045 15805 1055 15845
rect 1095 15805 1105 15845
rect 1145 15805 1155 15845
rect 1195 15805 1205 15845
rect 1245 15805 1255 15845
rect 1295 15805 1305 15845
rect 1345 15805 1355 15845
rect 1395 15805 1405 15845
rect 1445 15805 1455 15845
rect 1495 15805 1505 15845
rect 1545 15805 1555 15845
rect 1595 15805 1605 15845
rect 1645 15805 1655 15845
rect 1695 15805 1705 15845
rect 1745 15805 1755 15845
rect 1795 15805 1805 15845
rect 1845 15805 1855 15845
rect 1895 15805 1905 15845
rect 1945 15805 1955 15845
rect 1995 15805 2005 15845
rect 2045 15805 2055 15845
rect 2095 15805 2105 15845
rect 2145 15805 2155 15845
rect 2195 15805 2205 15845
rect 2245 15805 2255 15845
rect 2295 15805 2305 15845
rect 2345 15805 2355 15845
rect 2395 15805 2405 15845
rect 2445 15805 2455 15845
rect 2495 15805 2505 15845
rect 2545 15805 2555 15845
rect 2595 15805 2605 15845
rect 2645 15805 2655 15845
rect 2695 15805 2705 15845
rect 2745 15805 2755 15845
rect 2795 15805 2805 15845
rect 2845 15805 2855 15845
rect 2895 15805 2905 15845
rect 2945 15805 2955 15845
rect 2995 15805 3005 15845
rect 3045 15805 3055 15845
rect 3095 15805 3105 15845
rect 3145 15805 3155 15845
rect 3195 15805 3205 15845
rect 3245 15805 3255 15845
rect 3295 15805 3305 15845
rect 3345 15805 3355 15845
rect 3395 15805 3405 15845
rect 3445 15805 3455 15845
rect 3495 15805 3505 15845
rect 3545 15805 3555 15845
rect 3595 15805 3605 15845
rect 3645 15805 3655 15845
rect 3695 15805 3705 15845
rect 3745 15805 3755 15845
rect 3795 15805 3805 15845
rect 3845 15805 3855 15845
rect 3895 15805 3905 15845
rect 3945 15805 3955 15845
rect 3995 15805 4005 15845
rect 4045 15805 4055 15845
rect 4095 15805 4105 15845
rect 4145 15805 4155 15845
rect 4195 15805 4205 15845
rect 4245 15805 4255 15845
rect 4295 15805 4305 15845
rect 4345 15805 4355 15845
rect 4395 15805 4405 15845
rect 4445 15805 4455 15845
rect 4495 15805 4505 15845
rect 4545 15805 4555 15845
rect 4595 15805 4605 15845
rect 4645 15805 4655 15845
rect 4695 15805 4705 15845
rect 4745 15805 4755 15845
rect 4795 15805 4805 15845
rect 4845 15805 4855 15845
rect 4895 15805 4905 15845
rect 4945 15805 4955 15845
rect 4995 15805 5005 15845
rect 5045 15805 5055 15845
rect 5095 15805 5105 15845
rect 5145 15805 5155 15845
rect 5195 15805 5205 15845
rect 5245 15805 5255 15845
rect 5295 15805 5305 15845
rect 5345 15805 5355 15845
rect 5395 15805 5405 15845
rect 5445 15805 5455 15845
rect 5495 15805 5505 15845
rect 5545 15805 5555 15845
rect 5595 15805 5605 15845
rect 5645 15805 5655 15845
rect 5695 15805 5705 15845
rect 5745 15805 5755 15845
rect 5795 15805 5805 15845
rect 5845 15805 5855 15845
rect 5895 15805 5905 15845
rect 5945 15805 5955 15845
rect 5995 15805 6005 15845
rect 6045 15805 6055 15845
rect 6095 15805 6105 15845
rect 6145 15805 6155 15845
rect 6195 15805 6205 15845
rect 6245 15805 6255 15845
rect 6295 15805 6305 15845
rect 6345 15805 6355 15845
rect 6395 15805 6405 15845
rect 6445 15805 6455 15845
rect 6495 15805 6505 15845
rect 6545 15805 6555 15845
rect 6595 15805 6605 15845
rect 6645 15805 6655 15845
rect 6695 15805 6705 15845
rect 6745 15805 6755 15845
rect 6795 15805 6805 15845
rect 6845 15805 6855 15845
rect 6895 15805 6905 15845
rect 6945 15805 6955 15845
rect 6995 15805 7005 15845
rect 7045 15805 7055 15845
rect 7095 15805 7105 15845
rect 7145 15805 7155 15845
rect 7195 15805 7205 15845
rect 7245 15805 7255 15845
rect 7295 15805 7305 15845
rect 7345 15805 7355 15845
rect 7395 15805 7405 15845
rect 7445 15805 7455 15845
rect 7495 15805 7505 15845
rect 7545 15805 7555 15845
rect 7595 15805 7605 15845
rect 7645 15805 7655 15845
rect 7695 15805 7705 15845
rect 7745 15805 7755 15845
rect 7795 15805 7805 15845
rect 7845 15805 7855 15845
rect 7895 15805 7905 15845
rect 7945 15805 7955 15845
rect 7995 15805 8005 15845
rect 8045 15805 8055 15845
rect 8095 15805 8105 15845
rect 8145 15805 8155 15845
rect 8195 15805 8205 15845
rect 8245 15805 8255 15845
rect 8295 15805 8305 15845
rect 8345 15805 8355 15845
rect 8395 15805 8405 15845
rect 8445 15805 8455 15845
rect 8495 15805 8505 15845
rect 8545 15805 8555 15845
rect 8595 15805 8605 15845
rect 8645 15805 8655 15845
rect 8695 15805 8705 15845
rect 8745 15805 8755 15845
rect 8795 15805 8805 15845
rect 8845 15805 8855 15845
rect 8895 15805 8905 15845
rect 8945 15805 8955 15845
rect 8995 15805 9005 15845
rect 9045 15805 9055 15845
rect 9095 15805 9105 15845
rect 9145 15805 9155 15845
rect 9195 15805 9205 15845
rect 9245 15805 9255 15845
rect 9295 15805 9305 15845
rect 9345 15805 9355 15845
rect 9395 15805 9405 15845
rect 9445 15805 9455 15845
rect 9495 15805 9505 15845
rect 9545 15805 9555 15845
rect 9595 15805 9605 15845
rect 9645 15805 9655 15845
rect 9695 15805 9705 15845
rect 9745 15805 9755 15845
rect 9795 15805 9805 15845
rect 9845 15805 9855 15845
rect 9895 15805 9905 15845
rect 9945 15805 9955 15845
rect 9995 15805 10005 15845
rect 10045 15805 10055 15845
rect 10095 15805 10105 15845
rect 10145 15805 10155 15845
rect 10195 15805 10205 15845
rect 10245 15805 10255 15845
rect 10295 15805 10305 15845
rect 10345 15805 10355 15845
rect 10395 15805 10405 15845
rect 10445 15805 10455 15845
rect 10495 15805 10505 15845
rect 10545 15805 10555 15845
rect 10595 15805 10605 15845
rect 10645 15805 10655 15845
rect 10695 15805 10705 15845
rect 10745 15805 10755 15845
rect 10795 15805 10805 15845
rect 10845 15805 10855 15845
rect 10895 15805 10905 15845
rect 10945 15805 10955 15845
rect 10995 15805 11005 15845
rect 11045 15805 11055 15845
rect 11095 15805 11105 15845
rect 11145 15805 11155 15845
rect 11195 15805 11205 15845
rect 11245 15805 11255 15845
rect 11295 15805 11305 15845
rect 11345 15805 11355 15845
rect 11395 15805 11405 15845
rect 11445 15805 11455 15845
rect 11495 15805 11505 15845
rect 11545 15805 11555 15845
rect 11595 15805 11605 15845
rect 11645 15805 11655 15845
rect 11695 15805 11705 15845
rect 11745 15805 11755 15845
rect 11795 15805 11805 15845
rect 11845 15805 11855 15845
rect 11895 15805 11905 15845
rect 11945 15805 11955 15845
rect 11995 15805 12005 15845
rect 12045 15805 12055 15845
rect 12095 15805 12105 15845
rect 12145 15805 12155 15845
rect 12195 15805 12205 15845
rect 12245 15805 12255 15845
rect 12295 15805 12305 15845
rect 12345 15805 12355 15845
rect 12395 15805 12405 15845
rect 12445 15805 12455 15845
rect 12495 15805 12505 15845
rect 12545 15805 12555 15845
rect 12595 15805 12605 15845
rect 12645 15805 12655 15845
rect 12695 15805 12705 15845
rect 12745 15805 12755 15845
rect 12795 15805 12805 15845
rect 12845 15805 12855 15845
rect 12895 15805 12905 15845
rect 12945 15805 12955 15845
rect 12995 15805 13005 15845
rect 13045 15805 13055 15845
rect 13095 15805 13105 15845
rect 13145 15805 13155 15845
rect 13195 15805 13205 15845
rect 13245 15805 13255 15845
rect 13295 15805 13305 15845
rect 13345 15805 13355 15845
rect 13395 15805 13405 15845
rect 13445 15805 13455 15845
rect 13495 15805 13505 15845
rect 13545 15805 13555 15845
rect 13595 15805 13605 15845
rect 13645 15805 13655 15845
rect 13695 15805 13705 15845
rect 13745 15805 13755 15845
rect 13795 15805 13805 15845
rect 13845 15805 13855 15845
rect 13895 15805 13905 15845
rect 13945 15805 13955 15845
rect 13995 15805 14005 15845
rect 14045 15805 14055 15845
rect 14095 15805 14105 15845
rect 14145 15805 14155 15845
rect 14195 15805 14205 15845
rect 14245 15805 14255 15845
rect 14295 15805 14305 15845
rect 14345 15805 14355 15845
rect 14395 15805 14405 15845
rect 14445 15805 14455 15845
rect 14495 15805 14505 15845
rect 14545 15805 14555 15845
rect 14595 15805 14605 15845
rect 14645 15805 14655 15845
rect 14695 15805 14705 15845
rect 14745 15805 14755 15845
rect 14795 15805 14805 15845
rect 14845 15805 14855 15845
rect 14895 15805 14905 15845
rect 14945 15805 14955 15845
rect 14995 15805 15005 15845
rect 15045 15805 15055 15845
rect 15095 15805 15105 15845
rect 15145 15805 15155 15845
rect 15195 15805 15205 15845
rect 15245 15805 15255 15845
rect 15295 15805 15305 15845
rect 15345 15805 15355 15845
rect 15395 15805 15405 15845
rect 15445 15805 15455 15845
rect 15495 15805 15505 15845
rect 15545 15805 15555 15845
rect 15595 15805 15605 15845
rect 15645 15805 15655 15845
rect 15695 15805 15705 15845
rect 15745 15805 15755 15845
rect 15795 15805 15805 15845
rect 15845 15805 15855 15845
rect 15895 15805 15905 15845
rect 15945 15805 15955 15845
rect 15995 15805 16005 15845
rect 16045 15805 16055 15845
rect 16095 15805 16105 15845
rect 16145 15805 16155 15845
rect 16195 15805 16205 15845
rect 16245 15805 16255 15845
rect 16295 15805 16305 15845
rect 16345 15805 16355 15845
rect 16395 15805 16405 15845
rect 16445 15805 16455 15845
rect 16495 15805 16505 15845
rect 16545 15805 16555 15845
rect 16595 15805 16605 15845
rect 16645 15805 16655 15845
rect 16695 15805 16705 15845
rect 16745 15805 16755 15845
rect 16795 15805 16805 15845
rect 16845 15805 16855 15845
rect 16895 15805 16905 15845
rect 16945 15805 16955 15845
rect 16995 15805 17005 15845
rect 17045 15805 17055 15845
rect 17095 15805 17105 15845
rect 17145 15805 17155 15845
rect 17195 15805 17205 15845
rect 17245 15805 17255 15845
rect 17295 15805 17305 15845
rect 17345 15805 17355 15845
rect 17395 15805 17405 15845
rect 17445 15805 17455 15845
rect 17495 15805 17505 15845
rect 17545 15805 17555 15845
rect 17595 15805 17605 15845
rect 17645 15805 17655 15845
rect 17695 15805 17705 15845
rect 17745 15805 17755 15845
rect 17795 15805 17805 15845
rect 17845 15805 17855 15845
rect 17895 15805 17905 15845
rect 17945 15805 17955 15845
rect 17995 15805 18005 15845
rect 18045 15805 18055 15845
rect 18095 15805 18105 15845
rect 18145 15805 18155 15845
rect 18195 15805 18205 15845
rect 18245 15805 18255 15845
rect 18295 15805 18305 15845
rect 18345 15805 18355 15845
rect 18395 15805 18405 15845
rect 18445 15805 18455 15845
rect 18495 15805 18505 15845
rect 18545 15805 18555 15845
rect 18595 15805 18605 15845
rect 18645 15805 18655 15845
rect 18695 15805 18705 15845
rect 18745 15805 18755 15845
rect 18795 15805 18805 15845
rect 18845 15805 18855 15845
rect 18895 15805 18905 15845
rect 18945 15805 18955 15845
rect 18995 15805 19005 15845
rect 19045 15805 19055 15845
rect 19095 15805 19105 15845
rect 19145 15805 19155 15845
rect 19195 15805 19205 15845
rect 19245 15805 19255 15845
rect 19295 15805 19305 15845
rect 19345 15805 19355 15845
rect 19395 15805 19405 15845
rect 19445 15805 19455 15845
rect 19495 15805 19505 15845
rect 19545 15805 19555 15845
rect 19595 15805 19605 15845
rect 19645 15805 19655 15845
rect 19695 15805 19705 15845
rect 19745 15805 19755 15845
rect 19795 15805 19805 15845
rect 19845 15805 19855 15845
rect 19895 15805 19905 15845
rect 19945 15805 19955 15845
rect 19995 15805 20005 15845
rect 20045 15805 20055 15845
rect 20095 15805 20105 15845
rect 20145 15805 20155 15845
rect 20195 15805 20205 15845
rect 20245 15805 20255 15845
rect 20295 15805 20305 15845
rect 20345 15805 20355 15845
rect 20395 15805 20405 15845
rect 20445 15805 20455 15845
rect 20495 15805 20505 15845
rect 20545 15805 20555 15845
rect 20595 15805 20605 15845
rect 20645 15805 20655 15845
rect 20695 15805 20705 15845
rect 20745 15805 20755 15845
rect 20795 15805 20805 15845
rect 20845 15805 20855 15845
rect 20895 15805 20905 15845
rect 20945 15805 20955 15845
rect 20995 15805 21005 15845
rect 21045 15805 21055 15845
rect 21095 15805 21105 15845
rect 21145 15805 21155 15845
rect 21195 15805 21205 15845
rect 21245 15805 21255 15845
rect 21295 15805 21305 15845
rect 21345 15805 21355 15845
rect 21395 15805 21405 15845
rect 21445 15805 21455 15845
rect 21495 15805 21505 15845
rect 21545 15805 21555 15845
rect 21595 15805 21605 15845
rect 21645 15805 21655 15845
rect 21695 15805 21705 15845
rect 21745 15805 21755 15845
rect 21795 15805 21805 15845
rect 21845 15805 21855 15845
rect 21895 15805 21905 15845
rect 21945 15805 21955 15845
rect 21995 15805 22005 15845
rect 22045 15805 22055 15845
rect 22095 15805 22105 15845
rect 22145 15805 22155 15845
rect 22195 15805 22205 15845
rect 22245 15805 22255 15845
rect 22295 15805 22305 15845
rect 22345 15805 22355 15845
rect 22395 15805 22405 15845
rect 22445 15805 22455 15845
rect 22495 15805 22505 15845
rect 22545 15805 22555 15845
rect 22595 15805 22605 15845
rect 22645 15805 22655 15845
rect 22695 15805 22705 15845
rect 22745 15805 22755 15845
rect 22795 15805 22805 15845
rect 22845 15805 22855 15845
rect 22895 15805 22905 15845
rect 22945 15805 22955 15845
rect 22995 15805 23005 15845
rect 23045 15805 23055 15845
rect 23095 15805 23105 15845
rect 23145 15805 23155 15845
rect 23195 15805 23205 15845
rect 23245 15805 23255 15845
rect 23295 15805 23305 15845
rect 23345 15805 23355 15845
rect 23395 15805 23405 15845
rect 23445 15805 23455 15845
rect 23495 15805 23505 15845
rect 23545 15805 23555 15845
rect 23595 15805 23605 15845
rect 23645 15805 23655 15845
rect 23695 15805 23705 15845
rect 23745 15805 23755 15845
rect 23795 15805 23805 15845
rect 23845 15805 23855 15845
rect 23895 15805 23905 15845
rect 23945 15805 23955 15845
rect 23995 15805 24005 15845
rect 24045 15805 24055 15845
rect 24095 15805 24105 15845
rect 24145 15805 24155 15845
rect 24195 15805 24205 15845
rect 24245 15805 24255 15845
rect 24295 15805 24305 15845
rect 24345 15805 24355 15845
rect 24395 15805 24405 15845
rect 24445 15805 24455 15845
rect 24495 15805 24505 15845
rect 24545 15805 24555 15845
rect 24595 15805 24605 15845
rect 24645 15805 24655 15845
rect 24695 15805 24705 15845
rect 24745 15805 24755 15845
rect 24795 15805 24805 15845
rect 24845 15805 24855 15845
rect 24895 15805 24905 15845
rect 24945 15805 24955 15845
rect 24995 15805 25005 15845
rect 25045 15805 25055 15845
rect 25095 15805 25105 15845
rect 25145 15805 25155 15845
rect 25195 15805 25205 15845
rect 25245 15805 25255 15845
rect 25295 15805 25305 15845
rect 25345 15805 25355 15845
rect 25395 15805 25405 15845
rect 25445 15805 25455 15845
rect 25495 15805 25505 15845
rect 25545 15805 25555 15845
rect 25595 15805 25605 15845
rect 25645 15805 25655 15845
rect 25695 15805 25705 15845
rect 25745 15805 25755 15845
rect 25795 15805 25805 15845
rect 25845 15805 25855 15845
rect 25895 15805 25905 15845
rect 25945 15805 25955 15845
rect 25995 15805 26005 15845
rect 26045 15805 26055 15845
rect 26095 15805 26105 15845
rect 26145 15805 26155 15845
rect 26195 15805 26205 15845
rect 26245 15805 26255 15845
rect 26295 15805 26305 15845
rect 26345 15805 26355 15845
rect 26395 15805 26405 15845
rect 26445 15805 26455 15845
rect 26495 15805 26505 15845
rect 26545 15805 26555 15845
rect 26595 15805 26605 15845
rect 26645 15805 26655 15845
rect 26695 15805 26705 15845
rect 26745 15805 26755 15845
rect 26795 15805 26805 15845
rect 26845 15805 26855 15845
rect 26895 15805 26905 15845
rect 26945 15805 26955 15845
rect 26995 15805 27005 15845
rect 27045 15805 27055 15845
rect 27095 15805 27105 15845
rect 27145 15805 27155 15845
rect 27195 15805 27205 15845
rect 27245 15805 27255 15845
rect 27295 15805 27305 15845
rect 27345 15805 27355 15845
rect 27395 15805 27405 15845
rect 27445 15805 27455 15845
rect 27495 15805 27505 15845
rect 27545 15805 27555 15845
rect 27595 15805 27605 15845
rect 27645 15805 27655 15845
rect 27695 15805 27705 15845
rect 27745 15805 27755 15845
rect 27795 15805 27805 15845
rect 27845 15805 27855 15845
rect 27895 15805 27905 15845
rect 27945 15805 27955 15845
rect 27995 15805 28005 15845
rect 28045 15805 28055 15845
rect 28095 15805 28105 15845
rect 28145 15805 28155 15845
rect 28195 15805 28205 15845
rect 28245 15805 28255 15845
rect 28295 15805 28305 15845
rect 28345 15805 28355 15845
rect 28395 15805 28405 15845
rect 28445 15805 28455 15845
rect 28495 15805 28505 15845
rect 28545 15805 28555 15845
rect 28595 15805 28605 15845
rect 28645 15805 28655 15845
rect 28695 15805 28705 15845
rect 28745 15805 28755 15845
rect 28795 15805 28805 15845
rect 28845 15805 28855 15845
rect 28895 15805 28905 15845
rect 28945 15805 28955 15845
rect 28995 15805 29005 15845
rect 29045 15805 29055 15845
rect 29095 15805 29105 15845
rect 29145 15805 29155 15845
rect 29195 15805 29205 15845
rect 29245 15805 29255 15845
rect 29295 15805 29305 15845
rect 29345 15805 29355 15845
rect 29395 15805 29405 15845
rect 29445 15805 29455 15845
rect 29495 15805 29505 15845
rect 29545 15805 29555 15845
rect 29595 15805 29605 15845
rect 29645 15805 29655 15845
rect 29695 15805 29705 15845
rect 29745 15805 29755 15845
rect 29795 15805 29805 15845
rect 29845 15805 29855 15845
rect 29895 15805 29905 15845
rect 29945 15805 29955 15845
rect 29995 15805 30005 15845
rect 30045 15805 30055 15845
rect 30095 15805 30105 15845
rect 30145 15805 30155 15845
rect 30195 15805 30205 15845
rect 30245 15805 30255 15845
rect 30295 15805 30305 15845
rect 30345 15805 30355 15845
rect 30395 15805 30405 15845
rect 30445 15805 30455 15845
rect 30495 15805 30505 15845
rect 30545 15805 30555 15845
rect 30595 15805 30605 15845
rect 30645 15805 30655 15845
rect 30695 15805 30705 15845
rect 30745 15805 30755 15845
rect 30795 15805 30805 15845
rect 30845 15805 30855 15845
rect 30895 15805 30905 15845
rect 30945 15805 30955 15845
rect 30995 15805 31005 15845
rect 31045 15805 31055 15845
rect 31095 15805 31105 15845
rect 31145 15805 31155 15845
rect 31195 15805 31205 15845
rect 31245 15805 31255 15845
rect 31295 15805 31305 15845
rect 31345 15805 31355 15845
rect 31395 15805 31405 15845
rect 31445 15805 31455 15845
rect 31495 15805 31505 15845
rect 31545 15805 31555 15845
rect 31595 15805 31605 15845
rect 31645 15805 31655 15845
rect 31695 15805 31705 15845
rect 31745 15805 31755 15845
rect 31795 15805 31805 15845
rect 31845 15805 31855 15845
rect 31895 15805 31905 15845
rect 31945 15805 31955 15845
rect 31995 15805 32005 15845
rect 32045 15805 32055 15845
rect 32095 15805 32105 15845
rect 32145 15805 32155 15845
rect 32195 15805 32205 15845
rect 32245 15805 32255 15845
rect 32295 15805 32305 15845
rect 32345 15805 32355 15845
rect 32395 15805 32405 15845
rect 32445 15805 32455 15845
rect 32495 15805 32505 15845
rect 32545 15805 32555 15845
rect 32595 15805 32605 15845
rect 32645 15805 32655 15845
rect 32695 15805 32705 15845
rect 32745 15805 32755 15845
rect 32795 15805 32805 15845
rect 32845 15805 32855 15845
rect 32895 15805 32905 15845
rect 32945 15805 32955 15845
rect 32995 15805 33005 15845
rect 33045 15805 33055 15845
rect 33095 15805 33105 15845
rect 33145 15805 33155 15845
rect 33195 15805 33205 15845
rect 33245 15805 33255 15845
rect 33295 15805 33305 15845
rect 33345 15805 33355 15845
rect 33395 15805 33405 15845
rect 33445 15805 33455 15845
rect 33495 15805 33505 15845
rect 33545 15805 33555 15845
rect 33595 15805 33605 15845
rect 33645 15805 33655 15845
rect 33695 15805 33705 15845
rect 33745 15805 33755 15845
rect 33795 15805 33805 15845
rect 33845 15805 33855 15845
rect 33895 15805 33905 15845
rect 33945 15805 33955 15845
rect 33995 15805 34005 15845
rect 34045 15805 34055 15845
rect 34095 15805 34105 15845
rect 34145 15805 34155 15845
rect 34195 15805 34205 15845
rect 34245 15805 34255 15845
rect 34295 15805 34305 15845
rect 34345 15805 34355 15845
rect 34395 15805 34405 15845
rect 34445 15805 34455 15845
rect 34495 15805 34505 15845
rect 34545 15805 34555 15845
rect 34595 15805 34605 15845
rect 34645 15805 34655 15845
rect 34695 15805 34705 15845
rect 34745 15805 34755 15845
rect 34795 15805 34805 15845
rect 34845 15805 34855 15845
rect 34895 15805 34905 15845
rect 34945 15805 34955 15845
rect 34995 15805 35005 15845
rect 35045 15805 35055 15845
rect 35095 15805 35105 15845
rect 35145 15805 35155 15845
rect 35195 15805 35205 15845
rect 35245 15805 35255 15845
rect 35295 15805 35305 15845
rect 35345 15805 35355 15845
rect 35395 15805 35405 15845
rect 35445 15805 35455 15845
rect 35495 15805 35505 15845
rect 35545 15805 35555 15845
rect 35595 15805 35605 15845
rect 35645 15805 35655 15845
rect 35695 15805 35705 15845
rect 35745 15805 35755 15845
rect 35795 15805 35805 15845
rect 35845 15805 35855 15845
rect 35895 15805 35905 15845
rect 35945 15805 35955 15845
rect 35995 15805 36005 15845
rect 36045 15805 36055 15845
rect 36095 15805 36105 15845
rect 36145 15805 36155 15845
rect 36195 15805 36205 15845
rect 36245 15805 36255 15845
rect 36295 15805 36305 15845
rect 36345 15805 36355 15845
rect 36395 15805 36405 15845
rect 36445 15805 36455 15845
rect 36495 15805 36505 15845
rect 36545 15805 36555 15845
rect 36595 15805 36605 15845
rect 36645 15805 36655 15845
rect 36695 15805 36705 15845
rect 36745 15805 36755 15845
rect 36795 15805 36805 15845
rect 36845 15805 36855 15845
rect 36895 15805 36905 15845
rect 36945 15805 36955 15845
rect 36995 15805 37005 15845
rect 37045 15805 37055 15845
rect 37095 15805 37105 15845
rect 37145 15805 37155 15845
rect 37195 15805 37205 15845
rect 37245 15805 37255 15845
rect 37295 15805 37305 15845
rect 37345 15805 37355 15845
rect 37395 15805 37405 15845
rect 37445 15805 37455 15845
rect 37495 15805 37505 15845
rect 37545 15805 37555 15845
rect 37595 15805 37605 15845
rect 37645 15805 37655 15845
rect 37695 15805 37705 15845
rect 37745 15805 37755 15845
rect 37795 15805 37805 15845
rect 37845 15805 37855 15845
rect 37895 15805 37905 15845
rect 37945 15805 37955 15845
rect 37995 15805 38005 15845
rect 38045 15805 38055 15845
rect 38095 15805 38105 15845
rect 38145 15805 38155 15845
rect 38195 15805 38205 15845
rect 38245 15805 38255 15845
rect 38295 15805 38305 15845
rect 38345 15805 38355 15845
rect 38395 15805 38405 15845
rect 38445 15805 38455 15845
rect 38495 15805 38505 15845
rect 38545 15805 38555 15845
rect 38595 15805 38605 15845
rect 38645 15805 38655 15845
rect 38695 15805 38705 15845
rect 38745 15805 38755 15845
rect 38795 15805 38805 15845
rect 38845 15805 38855 15845
rect 38895 15805 38905 15845
rect 38945 15805 38955 15845
rect 38995 15805 39005 15845
rect 39045 15805 39055 15845
rect 39095 15805 39105 15845
rect 39145 15805 39155 15845
rect 39195 15805 39205 15845
rect 39245 15805 39255 15845
rect 39295 15805 39305 15845
rect 39345 15805 39355 15845
rect 39395 15805 39405 15845
rect 39445 15805 39455 15845
rect 39495 15805 39505 15845
rect 39545 15805 39555 15845
rect 39595 15805 39605 15845
rect 39645 15805 39655 15845
rect 39695 15805 39705 15845
rect 39745 15805 39750 15845
rect 0 15745 39750 15805
rect 0 15705 5 15745
rect 45 15705 55 15745
rect 95 15705 105 15745
rect 145 15705 155 15745
rect 195 15705 205 15745
rect 245 15705 255 15745
rect 295 15705 305 15745
rect 345 15705 355 15745
rect 395 15705 405 15745
rect 445 15705 455 15745
rect 495 15705 505 15745
rect 545 15705 555 15745
rect 595 15705 605 15745
rect 645 15705 655 15745
rect 695 15705 705 15745
rect 745 15705 755 15745
rect 795 15705 805 15745
rect 845 15705 855 15745
rect 895 15705 905 15745
rect 945 15705 955 15745
rect 995 15705 1005 15745
rect 1045 15705 1055 15745
rect 1095 15705 1105 15745
rect 1145 15705 1155 15745
rect 1195 15705 1205 15745
rect 1245 15705 1255 15745
rect 1295 15705 1305 15745
rect 1345 15705 1355 15745
rect 1395 15705 1405 15745
rect 1445 15705 1455 15745
rect 1495 15705 1505 15745
rect 1545 15705 1555 15745
rect 1595 15705 1605 15745
rect 1645 15705 1655 15745
rect 1695 15705 1705 15745
rect 1745 15705 1755 15745
rect 1795 15705 1805 15745
rect 1845 15705 1855 15745
rect 1895 15705 1905 15745
rect 1945 15705 1955 15745
rect 1995 15705 2005 15745
rect 2045 15705 2055 15745
rect 2095 15705 2105 15745
rect 2145 15705 2155 15745
rect 2195 15705 2205 15745
rect 2245 15705 2255 15745
rect 2295 15705 2305 15745
rect 2345 15705 2355 15745
rect 2395 15705 2405 15745
rect 2445 15705 2455 15745
rect 2495 15705 2505 15745
rect 2545 15705 2555 15745
rect 2595 15705 2605 15745
rect 2645 15705 2655 15745
rect 2695 15705 2705 15745
rect 2745 15705 2755 15745
rect 2795 15705 2805 15745
rect 2845 15705 2855 15745
rect 2895 15705 2905 15745
rect 2945 15705 2955 15745
rect 2995 15705 3005 15745
rect 3045 15705 3055 15745
rect 3095 15705 3105 15745
rect 3145 15705 3155 15745
rect 3195 15705 3205 15745
rect 3245 15705 3255 15745
rect 3295 15705 3305 15745
rect 3345 15705 3355 15745
rect 3395 15705 3405 15745
rect 3445 15705 3455 15745
rect 3495 15705 3505 15745
rect 3545 15705 3555 15745
rect 3595 15705 3605 15745
rect 3645 15705 3655 15745
rect 3695 15705 3705 15745
rect 3745 15705 3755 15745
rect 3795 15705 3805 15745
rect 3845 15705 3855 15745
rect 3895 15705 3905 15745
rect 3945 15705 3955 15745
rect 3995 15705 4005 15745
rect 4045 15705 4055 15745
rect 4095 15705 4105 15745
rect 4145 15705 4155 15745
rect 4195 15705 4205 15745
rect 4245 15705 4255 15745
rect 4295 15705 4305 15745
rect 4345 15705 4355 15745
rect 4395 15705 4405 15745
rect 4445 15705 4455 15745
rect 4495 15705 4505 15745
rect 4545 15705 4555 15745
rect 4595 15705 4605 15745
rect 4645 15705 4655 15745
rect 4695 15705 4705 15745
rect 4745 15705 4755 15745
rect 4795 15705 4805 15745
rect 4845 15705 4855 15745
rect 4895 15705 4905 15745
rect 4945 15705 4955 15745
rect 4995 15705 5005 15745
rect 5045 15705 5055 15745
rect 5095 15705 5105 15745
rect 5145 15705 5155 15745
rect 5195 15705 5205 15745
rect 5245 15705 5255 15745
rect 5295 15705 5305 15745
rect 5345 15705 5355 15745
rect 5395 15705 5405 15745
rect 5445 15705 5455 15745
rect 5495 15705 5505 15745
rect 5545 15705 5555 15745
rect 5595 15705 5605 15745
rect 5645 15705 5655 15745
rect 5695 15705 5705 15745
rect 5745 15705 5755 15745
rect 5795 15705 5805 15745
rect 5845 15705 5855 15745
rect 5895 15705 5905 15745
rect 5945 15705 5955 15745
rect 5995 15705 6005 15745
rect 6045 15705 6055 15745
rect 6095 15705 6105 15745
rect 6145 15705 6155 15745
rect 6195 15705 6205 15745
rect 6245 15705 6255 15745
rect 6295 15705 6305 15745
rect 6345 15705 6355 15745
rect 6395 15705 6405 15745
rect 6445 15705 6455 15745
rect 6495 15705 6505 15745
rect 6545 15705 6555 15745
rect 6595 15705 6605 15745
rect 6645 15705 6655 15745
rect 6695 15705 6705 15745
rect 6745 15705 6755 15745
rect 6795 15705 6805 15745
rect 6845 15705 6855 15745
rect 6895 15705 6905 15745
rect 6945 15705 6955 15745
rect 6995 15705 7005 15745
rect 7045 15705 7055 15745
rect 7095 15705 7105 15745
rect 7145 15705 7155 15745
rect 7195 15705 7205 15745
rect 7245 15705 7255 15745
rect 7295 15705 7305 15745
rect 7345 15705 7355 15745
rect 7395 15705 7405 15745
rect 7445 15705 7455 15745
rect 7495 15705 7505 15745
rect 7545 15705 7555 15745
rect 7595 15705 7605 15745
rect 7645 15705 7655 15745
rect 7695 15705 7705 15745
rect 7745 15705 7755 15745
rect 7795 15705 7805 15745
rect 7845 15705 7855 15745
rect 7895 15705 7905 15745
rect 7945 15705 7955 15745
rect 7995 15705 8005 15745
rect 8045 15705 8055 15745
rect 8095 15705 8105 15745
rect 8145 15705 8155 15745
rect 8195 15705 8205 15745
rect 8245 15705 8255 15745
rect 8295 15705 8305 15745
rect 8345 15705 8355 15745
rect 8395 15705 8405 15745
rect 8445 15705 8455 15745
rect 8495 15705 8505 15745
rect 8545 15705 8555 15745
rect 8595 15705 8605 15745
rect 8645 15705 8655 15745
rect 8695 15705 8705 15745
rect 8745 15705 8755 15745
rect 8795 15705 8805 15745
rect 8845 15705 8855 15745
rect 8895 15705 8905 15745
rect 8945 15705 8955 15745
rect 8995 15705 9005 15745
rect 9045 15705 9055 15745
rect 9095 15705 9105 15745
rect 9145 15705 9155 15745
rect 9195 15705 9205 15745
rect 9245 15705 9255 15745
rect 9295 15705 9305 15745
rect 9345 15705 9355 15745
rect 9395 15705 9405 15745
rect 9445 15705 9455 15745
rect 9495 15705 9505 15745
rect 9545 15705 9555 15745
rect 9595 15705 9605 15745
rect 9645 15705 9655 15745
rect 9695 15705 9705 15745
rect 9745 15705 9755 15745
rect 9795 15705 9805 15745
rect 9845 15705 9855 15745
rect 9895 15705 9905 15745
rect 9945 15705 9955 15745
rect 9995 15705 10005 15745
rect 10045 15705 10055 15745
rect 10095 15705 10105 15745
rect 10145 15705 10155 15745
rect 10195 15705 10205 15745
rect 10245 15705 10255 15745
rect 10295 15705 10305 15745
rect 10345 15705 10355 15745
rect 10395 15705 10405 15745
rect 10445 15705 10455 15745
rect 10495 15705 10505 15745
rect 10545 15705 10555 15745
rect 10595 15705 10605 15745
rect 10645 15705 10655 15745
rect 10695 15705 10705 15745
rect 10745 15705 10755 15745
rect 10795 15705 10805 15745
rect 10845 15705 10855 15745
rect 10895 15705 10905 15745
rect 10945 15705 10955 15745
rect 10995 15705 11005 15745
rect 11045 15705 11055 15745
rect 11095 15705 11105 15745
rect 11145 15705 11155 15745
rect 11195 15705 11205 15745
rect 11245 15705 11255 15745
rect 11295 15705 11305 15745
rect 11345 15705 11355 15745
rect 11395 15705 11405 15745
rect 11445 15705 11455 15745
rect 11495 15705 11505 15745
rect 11545 15705 11555 15745
rect 11595 15705 11605 15745
rect 11645 15705 11655 15745
rect 11695 15705 11705 15745
rect 11745 15705 11755 15745
rect 11795 15705 11805 15745
rect 11845 15705 11855 15745
rect 11895 15705 11905 15745
rect 11945 15705 11955 15745
rect 11995 15705 12005 15745
rect 12045 15705 12055 15745
rect 12095 15705 12105 15745
rect 12145 15705 12155 15745
rect 12195 15705 12205 15745
rect 12245 15705 12255 15745
rect 12295 15705 12305 15745
rect 12345 15705 12355 15745
rect 12395 15705 12405 15745
rect 12445 15705 12455 15745
rect 12495 15705 12505 15745
rect 12545 15705 12555 15745
rect 12595 15705 12605 15745
rect 12645 15705 12655 15745
rect 12695 15705 12705 15745
rect 12745 15705 12755 15745
rect 12795 15705 12805 15745
rect 12845 15705 12855 15745
rect 12895 15705 12905 15745
rect 12945 15705 12955 15745
rect 12995 15705 13005 15745
rect 13045 15705 13055 15745
rect 13095 15705 13105 15745
rect 13145 15705 13155 15745
rect 13195 15705 13205 15745
rect 13245 15705 13255 15745
rect 13295 15705 13305 15745
rect 13345 15705 13355 15745
rect 13395 15705 13405 15745
rect 13445 15705 13455 15745
rect 13495 15705 13505 15745
rect 13545 15705 13555 15745
rect 13595 15705 13605 15745
rect 13645 15705 13655 15745
rect 13695 15705 13705 15745
rect 13745 15705 13755 15745
rect 13795 15705 13805 15745
rect 13845 15705 13855 15745
rect 13895 15705 13905 15745
rect 13945 15705 13955 15745
rect 13995 15705 14005 15745
rect 14045 15705 14055 15745
rect 14095 15705 14105 15745
rect 14145 15705 14155 15745
rect 14195 15705 14205 15745
rect 14245 15705 14255 15745
rect 14295 15705 14305 15745
rect 14345 15705 14355 15745
rect 14395 15705 14405 15745
rect 14445 15705 14455 15745
rect 14495 15705 14505 15745
rect 14545 15705 14555 15745
rect 14595 15705 14605 15745
rect 14645 15705 14655 15745
rect 14695 15705 14705 15745
rect 14745 15705 14755 15745
rect 14795 15705 14805 15745
rect 14845 15705 14855 15745
rect 14895 15705 14905 15745
rect 14945 15705 14955 15745
rect 14995 15705 15005 15745
rect 15045 15705 15055 15745
rect 15095 15705 15105 15745
rect 15145 15705 15155 15745
rect 15195 15705 15205 15745
rect 15245 15705 15255 15745
rect 15295 15705 15305 15745
rect 15345 15705 15355 15745
rect 15395 15705 15405 15745
rect 15445 15705 15455 15745
rect 15495 15705 15505 15745
rect 15545 15705 15555 15745
rect 15595 15705 15605 15745
rect 15645 15705 15655 15745
rect 15695 15705 15705 15745
rect 15745 15705 15755 15745
rect 15795 15705 15805 15745
rect 15845 15705 15855 15745
rect 15895 15705 15905 15745
rect 15945 15705 15955 15745
rect 15995 15705 16005 15745
rect 16045 15705 16055 15745
rect 16095 15705 16105 15745
rect 16145 15705 16155 15745
rect 16195 15705 16205 15745
rect 16245 15705 16255 15745
rect 16295 15705 16305 15745
rect 16345 15705 16355 15745
rect 16395 15705 16405 15745
rect 16445 15705 16455 15745
rect 16495 15705 16505 15745
rect 16545 15705 16555 15745
rect 16595 15705 16605 15745
rect 16645 15705 16655 15745
rect 16695 15705 16705 15745
rect 16745 15705 16755 15745
rect 16795 15705 16805 15745
rect 16845 15705 16855 15745
rect 16895 15705 16905 15745
rect 16945 15705 16955 15745
rect 16995 15705 17005 15745
rect 17045 15705 17055 15745
rect 17095 15705 17105 15745
rect 17145 15705 17155 15745
rect 17195 15705 17205 15745
rect 17245 15705 17255 15745
rect 17295 15705 17305 15745
rect 17345 15705 17355 15745
rect 17395 15705 17405 15745
rect 17445 15705 17455 15745
rect 17495 15705 17505 15745
rect 17545 15705 17555 15745
rect 17595 15705 17605 15745
rect 17645 15705 17655 15745
rect 17695 15705 17705 15745
rect 17745 15705 17755 15745
rect 17795 15705 17805 15745
rect 17845 15705 17855 15745
rect 17895 15705 17905 15745
rect 17945 15705 17955 15745
rect 17995 15705 18005 15745
rect 18045 15705 18055 15745
rect 18095 15705 18105 15745
rect 18145 15705 18155 15745
rect 18195 15705 18205 15745
rect 18245 15705 18255 15745
rect 18295 15705 18305 15745
rect 18345 15705 18355 15745
rect 18395 15705 18405 15745
rect 18445 15705 18455 15745
rect 18495 15705 18505 15745
rect 18545 15705 18555 15745
rect 18595 15705 18605 15745
rect 18645 15705 18655 15745
rect 18695 15705 18705 15745
rect 18745 15705 18755 15745
rect 18795 15705 18805 15745
rect 18845 15705 18855 15745
rect 18895 15705 18905 15745
rect 18945 15705 18955 15745
rect 18995 15705 19005 15745
rect 19045 15705 19055 15745
rect 19095 15705 19105 15745
rect 19145 15705 19155 15745
rect 19195 15705 19205 15745
rect 19245 15705 19255 15745
rect 19295 15705 19305 15745
rect 19345 15705 19355 15745
rect 19395 15705 19405 15745
rect 19445 15705 19455 15745
rect 19495 15705 19505 15745
rect 19545 15705 19555 15745
rect 19595 15705 19605 15745
rect 19645 15705 19655 15745
rect 19695 15705 19705 15745
rect 19745 15705 19755 15745
rect 19795 15705 19805 15745
rect 19845 15705 19855 15745
rect 19895 15705 19905 15745
rect 19945 15705 19955 15745
rect 19995 15705 20005 15745
rect 20045 15705 20055 15745
rect 20095 15705 20105 15745
rect 20145 15705 20155 15745
rect 20195 15705 20205 15745
rect 20245 15705 20255 15745
rect 20295 15705 20305 15745
rect 20345 15705 20355 15745
rect 20395 15705 20405 15745
rect 20445 15705 20455 15745
rect 20495 15705 20505 15745
rect 20545 15705 20555 15745
rect 20595 15705 20605 15745
rect 20645 15705 20655 15745
rect 20695 15705 20705 15745
rect 20745 15705 20755 15745
rect 20795 15705 20805 15745
rect 20845 15705 20855 15745
rect 20895 15705 20905 15745
rect 20945 15705 20955 15745
rect 20995 15705 21005 15745
rect 21045 15705 21055 15745
rect 21095 15705 21105 15745
rect 21145 15705 21155 15745
rect 21195 15705 21205 15745
rect 21245 15705 21255 15745
rect 21295 15705 21305 15745
rect 21345 15705 21355 15745
rect 21395 15705 21405 15745
rect 21445 15705 21455 15745
rect 21495 15705 21505 15745
rect 21545 15705 21555 15745
rect 21595 15705 21605 15745
rect 21645 15705 21655 15745
rect 21695 15705 21705 15745
rect 21745 15705 21755 15745
rect 21795 15705 21805 15745
rect 21845 15705 21855 15745
rect 21895 15705 21905 15745
rect 21945 15705 21955 15745
rect 21995 15705 22005 15745
rect 22045 15705 22055 15745
rect 22095 15705 22105 15745
rect 22145 15705 22155 15745
rect 22195 15705 22205 15745
rect 22245 15705 22255 15745
rect 22295 15705 22305 15745
rect 22345 15705 22355 15745
rect 22395 15705 22405 15745
rect 22445 15705 22455 15745
rect 22495 15705 22505 15745
rect 22545 15705 22555 15745
rect 22595 15705 22605 15745
rect 22645 15705 22655 15745
rect 22695 15705 22705 15745
rect 22745 15705 22755 15745
rect 22795 15705 22805 15745
rect 22845 15705 22855 15745
rect 22895 15705 22905 15745
rect 22945 15705 22955 15745
rect 22995 15705 23005 15745
rect 23045 15705 23055 15745
rect 23095 15705 23105 15745
rect 23145 15705 23155 15745
rect 23195 15705 23205 15745
rect 23245 15705 23255 15745
rect 23295 15705 23305 15745
rect 23345 15705 23355 15745
rect 23395 15705 23405 15745
rect 23445 15705 23455 15745
rect 23495 15705 23505 15745
rect 23545 15705 23555 15745
rect 23595 15705 23605 15745
rect 23645 15705 23655 15745
rect 23695 15705 23705 15745
rect 23745 15705 23755 15745
rect 23795 15705 23805 15745
rect 23845 15705 23855 15745
rect 23895 15705 23905 15745
rect 23945 15705 23955 15745
rect 23995 15705 24005 15745
rect 24045 15705 24055 15745
rect 24095 15705 24105 15745
rect 24145 15705 24155 15745
rect 24195 15705 24205 15745
rect 24245 15705 24255 15745
rect 24295 15705 24305 15745
rect 24345 15705 24355 15745
rect 24395 15705 24405 15745
rect 24445 15705 24455 15745
rect 24495 15705 24505 15745
rect 24545 15705 24555 15745
rect 24595 15705 24605 15745
rect 24645 15705 24655 15745
rect 24695 15705 24705 15745
rect 24745 15705 24755 15745
rect 24795 15705 24805 15745
rect 24845 15705 24855 15745
rect 24895 15705 24905 15745
rect 24945 15705 24955 15745
rect 24995 15705 25005 15745
rect 25045 15705 25055 15745
rect 25095 15705 25105 15745
rect 25145 15705 25155 15745
rect 25195 15705 25205 15745
rect 25245 15705 25255 15745
rect 25295 15705 25305 15745
rect 25345 15705 25355 15745
rect 25395 15705 25405 15745
rect 25445 15705 25455 15745
rect 25495 15705 25505 15745
rect 25545 15705 25555 15745
rect 25595 15705 25605 15745
rect 25645 15705 25655 15745
rect 25695 15705 25705 15745
rect 25745 15705 25755 15745
rect 25795 15705 25805 15745
rect 25845 15705 25855 15745
rect 25895 15705 25905 15745
rect 25945 15705 25955 15745
rect 25995 15705 26005 15745
rect 26045 15705 26055 15745
rect 26095 15705 26105 15745
rect 26145 15705 26155 15745
rect 26195 15705 26205 15745
rect 26245 15705 26255 15745
rect 26295 15705 26305 15745
rect 26345 15705 26355 15745
rect 26395 15705 26405 15745
rect 26445 15705 26455 15745
rect 26495 15705 26505 15745
rect 26545 15705 26555 15745
rect 26595 15705 26605 15745
rect 26645 15705 26655 15745
rect 26695 15705 26705 15745
rect 26745 15705 26755 15745
rect 26795 15705 26805 15745
rect 26845 15705 26855 15745
rect 26895 15705 26905 15745
rect 26945 15705 26955 15745
rect 26995 15705 27005 15745
rect 27045 15705 27055 15745
rect 27095 15705 27105 15745
rect 27145 15705 27155 15745
rect 27195 15705 27205 15745
rect 27245 15705 27255 15745
rect 27295 15705 27305 15745
rect 27345 15705 27355 15745
rect 27395 15705 27405 15745
rect 27445 15705 27455 15745
rect 27495 15705 27505 15745
rect 27545 15705 27555 15745
rect 27595 15705 27605 15745
rect 27645 15705 27655 15745
rect 27695 15705 27705 15745
rect 27745 15705 27755 15745
rect 27795 15705 27805 15745
rect 27845 15705 27855 15745
rect 27895 15705 27905 15745
rect 27945 15705 27955 15745
rect 27995 15705 28005 15745
rect 28045 15705 28055 15745
rect 28095 15705 28105 15745
rect 28145 15705 28155 15745
rect 28195 15705 28205 15745
rect 28245 15705 28255 15745
rect 28295 15705 28305 15745
rect 28345 15705 28355 15745
rect 28395 15705 28405 15745
rect 28445 15705 28455 15745
rect 28495 15705 28505 15745
rect 28545 15705 28555 15745
rect 28595 15705 28605 15745
rect 28645 15705 28655 15745
rect 28695 15705 28705 15745
rect 28745 15705 28755 15745
rect 28795 15705 28805 15745
rect 28845 15705 28855 15745
rect 28895 15705 28905 15745
rect 28945 15705 28955 15745
rect 28995 15705 29005 15745
rect 29045 15705 29055 15745
rect 29095 15705 29105 15745
rect 29145 15705 29155 15745
rect 29195 15705 29205 15745
rect 29245 15705 29255 15745
rect 29295 15705 29305 15745
rect 29345 15705 29355 15745
rect 29395 15705 29405 15745
rect 29445 15705 29455 15745
rect 29495 15705 29505 15745
rect 29545 15705 29555 15745
rect 29595 15705 29605 15745
rect 29645 15705 29655 15745
rect 29695 15705 29705 15745
rect 29745 15705 29755 15745
rect 29795 15705 29805 15745
rect 29845 15705 29855 15745
rect 29895 15705 29905 15745
rect 29945 15705 29955 15745
rect 29995 15705 30005 15745
rect 30045 15705 30055 15745
rect 30095 15705 30105 15745
rect 30145 15705 30155 15745
rect 30195 15705 30205 15745
rect 30245 15705 30255 15745
rect 30295 15705 30305 15745
rect 30345 15705 30355 15745
rect 30395 15705 30405 15745
rect 30445 15705 30455 15745
rect 30495 15705 30505 15745
rect 30545 15705 30555 15745
rect 30595 15705 30605 15745
rect 30645 15705 30655 15745
rect 30695 15705 30705 15745
rect 30745 15705 30755 15745
rect 30795 15705 30805 15745
rect 30845 15705 30855 15745
rect 30895 15705 30905 15745
rect 30945 15705 30955 15745
rect 30995 15705 31005 15745
rect 31045 15705 31055 15745
rect 31095 15705 31105 15745
rect 31145 15705 31155 15745
rect 31195 15705 31205 15745
rect 31245 15705 31255 15745
rect 31295 15705 31305 15745
rect 31345 15705 31355 15745
rect 31395 15705 31405 15745
rect 31445 15705 31455 15745
rect 31495 15705 31505 15745
rect 31545 15705 31555 15745
rect 31595 15705 31605 15745
rect 31645 15705 31655 15745
rect 31695 15705 31705 15745
rect 31745 15705 31755 15745
rect 31795 15705 31805 15745
rect 31845 15705 31855 15745
rect 31895 15705 31905 15745
rect 31945 15705 31955 15745
rect 31995 15705 32005 15745
rect 32045 15705 32055 15745
rect 32095 15705 32105 15745
rect 32145 15705 32155 15745
rect 32195 15705 32205 15745
rect 32245 15705 32255 15745
rect 32295 15705 32305 15745
rect 32345 15705 32355 15745
rect 32395 15705 32405 15745
rect 32445 15705 32455 15745
rect 32495 15705 32505 15745
rect 32545 15705 32555 15745
rect 32595 15705 32605 15745
rect 32645 15705 32655 15745
rect 32695 15705 32705 15745
rect 32745 15705 32755 15745
rect 32795 15705 32805 15745
rect 32845 15705 32855 15745
rect 32895 15705 32905 15745
rect 32945 15705 32955 15745
rect 32995 15705 33005 15745
rect 33045 15705 33055 15745
rect 33095 15705 33105 15745
rect 33145 15705 33155 15745
rect 33195 15705 33205 15745
rect 33245 15705 33255 15745
rect 33295 15705 33305 15745
rect 33345 15705 33355 15745
rect 33395 15705 33405 15745
rect 33445 15705 33455 15745
rect 33495 15705 33505 15745
rect 33545 15705 33555 15745
rect 33595 15705 33605 15745
rect 33645 15705 33655 15745
rect 33695 15705 33705 15745
rect 33745 15705 33755 15745
rect 33795 15705 33805 15745
rect 33845 15705 33855 15745
rect 33895 15705 33905 15745
rect 33945 15705 33955 15745
rect 33995 15705 34005 15745
rect 34045 15705 34055 15745
rect 34095 15705 34105 15745
rect 34145 15705 34155 15745
rect 34195 15705 34205 15745
rect 34245 15705 34255 15745
rect 34295 15705 34305 15745
rect 34345 15705 34355 15745
rect 34395 15705 34405 15745
rect 34445 15705 34455 15745
rect 34495 15705 34505 15745
rect 34545 15705 34555 15745
rect 34595 15705 34605 15745
rect 34645 15705 34655 15745
rect 34695 15705 34705 15745
rect 34745 15705 34755 15745
rect 34795 15705 34805 15745
rect 34845 15705 34855 15745
rect 34895 15705 34905 15745
rect 34945 15705 34955 15745
rect 34995 15705 35005 15745
rect 35045 15705 35055 15745
rect 35095 15705 35105 15745
rect 35145 15705 35155 15745
rect 35195 15705 35205 15745
rect 35245 15705 35255 15745
rect 35295 15705 35305 15745
rect 35345 15705 35355 15745
rect 35395 15705 35405 15745
rect 35445 15705 35455 15745
rect 35495 15705 35505 15745
rect 35545 15705 35555 15745
rect 35595 15705 35605 15745
rect 35645 15705 35655 15745
rect 35695 15705 35705 15745
rect 35745 15705 35755 15745
rect 35795 15705 35805 15745
rect 35845 15705 35855 15745
rect 35895 15705 35905 15745
rect 35945 15705 35955 15745
rect 35995 15705 36005 15745
rect 36045 15705 36055 15745
rect 36095 15705 36105 15745
rect 36145 15705 36155 15745
rect 36195 15705 36205 15745
rect 36245 15705 36255 15745
rect 36295 15705 36305 15745
rect 36345 15705 36355 15745
rect 36395 15705 36405 15745
rect 36445 15705 36455 15745
rect 36495 15705 36505 15745
rect 36545 15705 36555 15745
rect 36595 15705 36605 15745
rect 36645 15705 36655 15745
rect 36695 15705 36705 15745
rect 36745 15705 36755 15745
rect 36795 15705 36805 15745
rect 36845 15705 36855 15745
rect 36895 15705 36905 15745
rect 36945 15705 36955 15745
rect 36995 15705 37005 15745
rect 37045 15705 37055 15745
rect 37095 15705 37105 15745
rect 37145 15705 37155 15745
rect 37195 15705 37205 15745
rect 37245 15705 37255 15745
rect 37295 15705 37305 15745
rect 37345 15705 37355 15745
rect 37395 15705 37405 15745
rect 37445 15705 37455 15745
rect 37495 15705 37505 15745
rect 37545 15705 37555 15745
rect 37595 15705 37605 15745
rect 37645 15705 37655 15745
rect 37695 15705 37705 15745
rect 37745 15705 37755 15745
rect 37795 15705 37805 15745
rect 37845 15705 37855 15745
rect 37895 15705 37905 15745
rect 37945 15705 37955 15745
rect 37995 15705 38005 15745
rect 38045 15705 38055 15745
rect 38095 15705 38105 15745
rect 38145 15705 38155 15745
rect 38195 15705 38205 15745
rect 38245 15705 38255 15745
rect 38295 15705 38305 15745
rect 38345 15705 38355 15745
rect 38395 15705 38405 15745
rect 38445 15705 38455 15745
rect 38495 15705 38505 15745
rect 38545 15705 38555 15745
rect 38595 15705 38605 15745
rect 38645 15705 38655 15745
rect 38695 15705 38705 15745
rect 38745 15705 38755 15745
rect 38795 15705 38805 15745
rect 38845 15705 38855 15745
rect 38895 15705 38905 15745
rect 38945 15705 38955 15745
rect 38995 15705 39005 15745
rect 39045 15705 39055 15745
rect 39095 15705 39105 15745
rect 39145 15705 39155 15745
rect 39195 15705 39205 15745
rect 39245 15705 39255 15745
rect 39295 15705 39305 15745
rect 39345 15705 39355 15745
rect 39395 15705 39405 15745
rect 39445 15705 39455 15745
rect 39495 15705 39505 15745
rect 39545 15705 39555 15745
rect 39595 15705 39605 15745
rect 39645 15705 39655 15745
rect 39695 15705 39705 15745
rect 39745 15705 39750 15745
rect 0 15700 39750 15705
rect -300 15345 -250 15700
rect -300 15305 -295 15345
rect -255 15305 -250 15345
rect -300 15295 -250 15305
rect -300 15255 -295 15295
rect -255 15255 -250 15295
rect -300 15245 -250 15255
rect -300 15205 -295 15245
rect -255 15205 -250 15245
rect -300 13645 -250 15205
rect -300 13605 -295 13645
rect -255 13605 -250 13645
rect -300 13595 -250 13605
rect -300 13555 -295 13595
rect -255 13555 -250 13595
rect -300 13545 -250 13555
rect -300 13505 -295 13545
rect -255 13505 -250 13545
rect -300 11945 -250 13505
rect -300 11905 -295 11945
rect -255 11905 -250 11945
rect -300 11895 -250 11905
rect -300 11855 -295 11895
rect -255 11855 -250 11895
rect -300 11845 -250 11855
rect -300 11805 -295 11845
rect -255 11805 -250 11845
rect -300 3845 -250 11805
rect -300 3805 -295 3845
rect -255 3805 -250 3845
rect -300 3795 -250 3805
rect -300 3755 -295 3795
rect -255 3755 -250 3795
rect -300 3745 -250 3755
rect -300 3705 -295 3745
rect -255 3705 -250 3745
rect -300 2145 -250 3705
rect -300 2105 -295 2145
rect -255 2105 -250 2145
rect -300 2095 -250 2105
rect -300 2055 -295 2095
rect -255 2055 -250 2095
rect -300 2045 -250 2055
rect -300 2005 -295 2045
rect -255 2005 -250 2045
rect -300 445 -250 2005
rect -300 405 -295 445
rect -255 405 -250 445
rect -300 395 -250 405
rect -300 355 -295 395
rect -255 355 -250 395
rect -300 345 -250 355
rect -300 305 -295 345
rect -255 305 -250 345
rect -300 0 -250 305
rect -200 14645 -150 15650
rect -200 14605 -195 14645
rect -155 14605 -150 14645
rect -200 1045 -150 14605
rect -200 1005 -195 1045
rect -155 1005 -150 1045
rect -200 0 -150 1005
rect -100 15345 -50 15700
rect -100 15305 -95 15345
rect -55 15305 -50 15345
rect -100 15295 -50 15305
rect -100 15255 -95 15295
rect -55 15255 -50 15295
rect -100 15245 -50 15255
rect -100 15205 -95 15245
rect -55 15205 -50 15245
rect -100 13645 -50 15205
rect -100 13605 -95 13645
rect -55 13605 -50 13645
rect -100 13595 -50 13605
rect -100 13555 -95 13595
rect -55 13555 -50 13595
rect -100 13545 -50 13555
rect -100 13505 -95 13545
rect -55 13505 -50 13545
rect -100 11945 -50 13505
rect -100 11905 -95 11945
rect -55 11905 -50 11945
rect -100 11895 -50 11905
rect -100 11855 -95 11895
rect -55 11855 -50 11895
rect -100 11845 -50 11855
rect -100 11805 -95 11845
rect -55 11805 -50 11845
rect -100 3845 -50 11805
rect -100 3805 -95 3845
rect -55 3805 -50 3845
rect -100 3795 -50 3805
rect -100 3755 -95 3795
rect -55 3755 -50 3795
rect -100 3745 -50 3755
rect -100 3705 -95 3745
rect -55 3705 -50 3745
rect -100 2145 -50 3705
rect -100 2105 -95 2145
rect -55 2105 -50 2145
rect -100 2095 -50 2105
rect -100 2055 -95 2095
rect -55 2055 -50 2095
rect -100 2045 -50 2055
rect -100 2005 -95 2045
rect -55 2005 -50 2045
rect -100 445 -50 2005
rect -100 405 -95 445
rect -55 405 -50 445
rect -100 395 -50 405
rect -100 355 -95 395
rect -55 355 -50 395
rect -100 345 -50 355
rect -100 305 -95 345
rect -55 305 -50 345
rect -100 0 -50 305
rect 39800 11345 39850 18290
rect 39800 11305 39805 11345
rect 39845 11305 39850 11345
rect 39800 10945 39850 11305
rect 39800 10905 39805 10945
rect 39845 10905 39850 10945
rect 39800 4745 39850 10905
rect 39800 4705 39805 4745
rect 39845 4705 39850 4745
rect 39800 4345 39850 4705
rect 39800 4305 39805 4345
rect 39845 4305 39850 4345
rect 39800 0 39850 4305
rect 39900 18285 40900 18290
rect 39900 18245 39905 18285
rect 39945 18245 39955 18285
rect 39995 18245 40005 18285
rect 40045 18245 40055 18285
rect 40095 18245 40105 18285
rect 40145 18245 40155 18285
rect 40195 18245 40205 18285
rect 40245 18245 40255 18285
rect 40295 18245 40305 18285
rect 40345 18245 40355 18285
rect 40395 18245 40405 18285
rect 40445 18245 40455 18285
rect 40495 18245 40505 18285
rect 40545 18245 40555 18285
rect 40595 18245 40605 18285
rect 40645 18245 40655 18285
rect 40695 18245 40705 18285
rect 40745 18245 40755 18285
rect 40795 18245 40805 18285
rect 40845 18245 40855 18285
rect 40895 18245 40900 18285
rect 39900 17015 40900 18245
rect 39900 16975 39905 17015
rect 39945 16975 39955 17015
rect 39995 16975 40005 17015
rect 40045 16975 40055 17015
rect 40095 16975 40105 17015
rect 40145 16975 40155 17015
rect 40195 16975 40205 17015
rect 40245 16975 40255 17015
rect 40295 16975 40305 17015
rect 40345 16975 40355 17015
rect 40395 16975 40405 17015
rect 40445 16975 40455 17015
rect 40495 16975 40505 17015
rect 40545 16975 40555 17015
rect 40595 16975 40605 17015
rect 40645 16975 40655 17015
rect 40695 16975 40705 17015
rect 40745 16975 40755 17015
rect 40795 16975 40805 17015
rect 40845 16975 40855 17015
rect 40895 16975 40900 17015
rect 39900 15745 40900 16975
rect 39900 15705 39905 15745
rect 39945 15705 39955 15745
rect 39995 15705 40005 15745
rect 40045 15705 40055 15745
rect 40095 15705 40105 15745
rect 40145 15705 40155 15745
rect 40195 15705 40205 15745
rect 40245 15705 40255 15745
rect 40295 15705 40305 15745
rect 40345 15705 40355 15745
rect 40395 15705 40405 15745
rect 40445 15705 40455 15745
rect 40495 15705 40505 15745
rect 40545 15705 40555 15745
rect 40595 15705 40605 15745
rect 40645 15705 40655 15745
rect 40695 15705 40705 15745
rect 40745 15705 40755 15745
rect 40795 15705 40805 15745
rect 40845 15705 40855 15745
rect 40895 15705 40900 15745
rect 39900 11245 40900 15705
rect 39900 11205 39905 11245
rect 39945 11205 39955 11245
rect 39995 11205 40005 11245
rect 40045 11205 40055 11245
rect 40095 11205 40105 11245
rect 40145 11205 40155 11245
rect 40195 11205 40205 11245
rect 40245 11205 40255 11245
rect 40295 11205 40305 11245
rect 40345 11205 40355 11245
rect 40395 11205 40405 11245
rect 40445 11205 40455 11245
rect 40495 11205 40505 11245
rect 40545 11205 40555 11245
rect 40595 11205 40605 11245
rect 40645 11205 40655 11245
rect 40695 11205 40705 11245
rect 40745 11205 40755 11245
rect 40795 11205 40805 11245
rect 40845 11205 40855 11245
rect 40895 11205 40900 11245
rect 39900 11195 40900 11205
rect 39900 11155 39905 11195
rect 39945 11155 39955 11195
rect 39995 11155 40005 11195
rect 40045 11155 40055 11195
rect 40095 11155 40105 11195
rect 40145 11155 40155 11195
rect 40195 11155 40205 11195
rect 40245 11155 40255 11195
rect 40295 11155 40305 11195
rect 40345 11155 40355 11195
rect 40395 11155 40405 11195
rect 40445 11155 40455 11195
rect 40495 11155 40505 11195
rect 40545 11155 40555 11195
rect 40595 11155 40605 11195
rect 40645 11155 40655 11195
rect 40695 11155 40705 11195
rect 40745 11155 40755 11195
rect 40795 11155 40805 11195
rect 40845 11155 40855 11195
rect 40895 11155 40900 11195
rect 39900 11145 40900 11155
rect 39900 11105 39905 11145
rect 39945 11105 39955 11145
rect 39995 11105 40005 11145
rect 40045 11105 40055 11145
rect 40095 11105 40105 11145
rect 40145 11105 40155 11145
rect 40195 11105 40205 11145
rect 40245 11105 40255 11145
rect 40295 11105 40305 11145
rect 40345 11105 40355 11145
rect 40395 11105 40405 11145
rect 40445 11105 40455 11145
rect 40495 11105 40505 11145
rect 40545 11105 40555 11145
rect 40595 11105 40605 11145
rect 40645 11105 40655 11145
rect 40695 11105 40705 11145
rect 40745 11105 40755 11145
rect 40795 11105 40805 11145
rect 40845 11105 40855 11145
rect 40895 11105 40900 11145
rect 39900 11095 40900 11105
rect 39900 11055 39905 11095
rect 39945 11055 39955 11095
rect 39995 11055 40005 11095
rect 40045 11055 40055 11095
rect 40095 11055 40105 11095
rect 40145 11055 40155 11095
rect 40195 11055 40205 11095
rect 40245 11055 40255 11095
rect 40295 11055 40305 11095
rect 40345 11055 40355 11095
rect 40395 11055 40405 11095
rect 40445 11055 40455 11095
rect 40495 11055 40505 11095
rect 40545 11055 40555 11095
rect 40595 11055 40605 11095
rect 40645 11055 40655 11095
rect 40695 11055 40705 11095
rect 40745 11055 40755 11095
rect 40795 11055 40805 11095
rect 40845 11055 40855 11095
rect 40895 11055 40900 11095
rect 39900 11045 40900 11055
rect 39900 11005 39905 11045
rect 39945 11005 39955 11045
rect 39995 11005 40005 11045
rect 40045 11005 40055 11045
rect 40095 11005 40105 11045
rect 40145 11005 40155 11045
rect 40195 11005 40205 11045
rect 40245 11005 40255 11045
rect 40295 11005 40305 11045
rect 40345 11005 40355 11045
rect 40395 11005 40405 11045
rect 40445 11005 40455 11045
rect 40495 11005 40505 11045
rect 40545 11005 40555 11045
rect 40595 11005 40605 11045
rect 40645 11005 40655 11045
rect 40695 11005 40705 11045
rect 40745 11005 40755 11045
rect 40795 11005 40805 11045
rect 40845 11005 40855 11045
rect 40895 11005 40900 11045
rect 39900 4645 40900 11005
rect 39900 4605 39905 4645
rect 39945 4605 39955 4645
rect 39995 4605 40005 4645
rect 40045 4605 40055 4645
rect 40095 4605 40105 4645
rect 40145 4605 40155 4645
rect 40195 4605 40205 4645
rect 40245 4605 40255 4645
rect 40295 4605 40305 4645
rect 40345 4605 40355 4645
rect 40395 4605 40405 4645
rect 40445 4605 40455 4645
rect 40495 4605 40505 4645
rect 40545 4605 40555 4645
rect 40595 4605 40605 4645
rect 40645 4605 40655 4645
rect 40695 4605 40705 4645
rect 40745 4605 40755 4645
rect 40795 4605 40805 4645
rect 40845 4605 40855 4645
rect 40895 4605 40900 4645
rect 39900 4595 40900 4605
rect 39900 4555 39905 4595
rect 39945 4555 39955 4595
rect 39995 4555 40005 4595
rect 40045 4555 40055 4595
rect 40095 4555 40105 4595
rect 40145 4555 40155 4595
rect 40195 4555 40205 4595
rect 40245 4555 40255 4595
rect 40295 4555 40305 4595
rect 40345 4555 40355 4595
rect 40395 4555 40405 4595
rect 40445 4555 40455 4595
rect 40495 4555 40505 4595
rect 40545 4555 40555 4595
rect 40595 4555 40605 4595
rect 40645 4555 40655 4595
rect 40695 4555 40705 4595
rect 40745 4555 40755 4595
rect 40795 4555 40805 4595
rect 40845 4555 40855 4595
rect 40895 4555 40900 4595
rect 39900 4545 40900 4555
rect 39900 4505 39905 4545
rect 39945 4505 39955 4545
rect 39995 4505 40005 4545
rect 40045 4505 40055 4545
rect 40095 4505 40105 4545
rect 40145 4505 40155 4545
rect 40195 4505 40205 4545
rect 40245 4505 40255 4545
rect 40295 4505 40305 4545
rect 40345 4505 40355 4545
rect 40395 4505 40405 4545
rect 40445 4505 40455 4545
rect 40495 4505 40505 4545
rect 40545 4505 40555 4545
rect 40595 4505 40605 4545
rect 40645 4505 40655 4545
rect 40695 4505 40705 4545
rect 40745 4505 40755 4545
rect 40795 4505 40805 4545
rect 40845 4505 40855 4545
rect 40895 4505 40900 4545
rect 39900 4495 40900 4505
rect 39900 4455 39905 4495
rect 39945 4455 39955 4495
rect 39995 4455 40005 4495
rect 40045 4455 40055 4495
rect 40095 4455 40105 4495
rect 40145 4455 40155 4495
rect 40195 4455 40205 4495
rect 40245 4455 40255 4495
rect 40295 4455 40305 4495
rect 40345 4455 40355 4495
rect 40395 4455 40405 4495
rect 40445 4455 40455 4495
rect 40495 4455 40505 4495
rect 40545 4455 40555 4495
rect 40595 4455 40605 4495
rect 40645 4455 40655 4495
rect 40695 4455 40705 4495
rect 40745 4455 40755 4495
rect 40795 4455 40805 4495
rect 40845 4455 40855 4495
rect 40895 4455 40900 4495
rect 39900 4445 40900 4455
rect 39900 4405 39905 4445
rect 39945 4405 39955 4445
rect 39995 4405 40005 4445
rect 40045 4405 40055 4445
rect 40095 4405 40105 4445
rect 40145 4405 40155 4445
rect 40195 4405 40205 4445
rect 40245 4405 40255 4445
rect 40295 4405 40305 4445
rect 40345 4405 40355 4445
rect 40395 4405 40405 4445
rect 40445 4405 40455 4445
rect 40495 4405 40505 4445
rect 40545 4405 40555 4445
rect 40595 4405 40605 4445
rect 40645 4405 40655 4445
rect 40695 4405 40705 4445
rect 40745 4405 40755 4445
rect 40795 4405 40805 4445
rect 40845 4405 40855 4445
rect 40895 4405 40900 4445
rect 39900 0 40900 4405
<< rmetal4 >>
rect -1300 18190 -1250 18240
use lpopamp_slice  slice0
timestamp 1713022628
transform -1 0 38750 0 -1 13550
box -1000 -2100 38750 5750
use lpopamp_slice  slice1
timestamp 1713022628
transform 1 0 1000 0 1 2100
box -1000 -2100 38750 5750
<< labels >>
rlabel metal3 -50 1000 0 1050 0 xn
rlabel metal3 -50 1400 0 1450 0 ynm
rlabel metal3 -50 1600 0 1650 0 ynp
rlabel metal3 -50 2500 0 2550 0 znm
rlabel metal3 -50 2700 0 2750 0 znp
rlabel metal3 -50 3100 0 3150 0 bna
rlabel metal3 -50 3200 0 3250 0 bnb
rlabel metal3 -50 5400 0 5450 0 bpb
rlabel metal3 -50 5500 0 5550 0 bpa
rlabel metal3 -50 5900 0 5950 0 zpp
rlabel metal3 -50 6100 0 6150 0 zpm
rlabel metal3 -50 6800 0 6850 0 ypm
rlabel metal3 -50 7200 0 7250 0 xp
rlabel metal3 -50 6600 0 6650 0 ypp
rlabel locali 0 0 50 50 0 vsub
port 9 nsew
rlabel metal4 -3400 18240 -3350 18290 0 im
port 1 nsew
rlabel metal4 -3200 18240 -3150 18290 0 ip
port 2 nsew
rlabel metal4 39900 18240 40900 18290 0 o
port 3 nsew
rlabel metal4 -1300 18240 -1250 18290 0 ib
port 4 nsew
rlabel metal4 -1400 18240 -1350 18290 0 en
port 5 nsew
rlabel metal4 -1500 18240 -1450 18290 0 enb
port 6 nsew
rlabel metal4 -3000 18240 -1650 18290 0 avdd
port 7 nsew
rlabel metal4 -1200 18240 -50 18290 0 avss
port 8 nsew
<< end >>
