magic
tech sky130A
timestamp 1711450593
<< error_p >>
rect 20400 1750 20450 1950
rect 20400 -1850 20433 -1817
rect 20367 -1900 20433 -1850
rect 20400 -1933 20433 -1900
rect 19950 -2000 20400 -1950
<< dnwell >>
rect -850 -1950 20400 1900
<< nwell >>
rect -700 2500 20450 5250
rect -900 1750 20450 1950
rect -900 -1800 -700 1750
rect -900 -2000 20400 -1800
<< mvnmos >>
rect -600 900 -500 1600
rect -450 900 -350 1600
rect -300 900 -200 1600
rect -150 900 -50 1600
rect 0 900 100 1600
rect 150 900 250 1600
rect 300 900 400 1600
rect 450 900 550 1600
rect 600 900 700 1600
rect 750 900 850 1600
rect 900 900 1000 1600
rect 1050 900 1150 1600
rect 1200 900 1300 1600
rect 1350 900 1450 1600
rect 1500 900 1600 1600
rect 1650 900 1750 1600
rect 1800 900 1900 1600
rect 1950 900 2050 1600
rect 2100 900 2200 1600
rect 2250 900 2350 1600
rect 2400 900 2500 1600
rect 2550 900 2650 1600
rect 2700 900 2800 1600
rect 2850 900 2950 1600
rect 3000 900 3100 1600
rect 3150 900 3250 1600
rect 3300 900 3400 1600
rect 3450 900 3550 1600
rect 3600 900 3700 1600
rect 3750 900 3850 1600
rect 3900 900 4000 1600
rect 4050 900 4150 1600
rect 4200 900 4300 1600
rect 4350 900 4450 1600
rect 4500 900 4600 1600
rect 4650 900 4750 1600
rect 4800 900 4900 1600
rect 4950 900 5050 1600
rect 5100 900 5200 1600
rect 5250 900 5350 1600
rect 5400 900 5500 1600
rect 5550 900 5650 1600
rect 5700 900 5800 1600
rect 5850 900 5950 1600
rect 6000 900 6100 1600
rect 6150 900 6250 1600
rect 6300 900 6400 1600
rect 6450 900 6550 1600
rect 6600 900 6700 1600
rect 6750 900 6850 1600
rect 6900 900 7000 1600
rect 7050 900 7150 1600
rect 7200 900 7300 1600
rect 7350 900 7450 1600
rect 7500 900 7600 1600
rect 7650 900 7750 1600
rect 7800 900 7900 1600
rect 7950 900 8050 1600
rect 8100 900 8200 1600
rect 8250 900 8350 1600
rect 8400 900 8500 1600
rect 8550 900 8650 1600
rect 8700 900 8800 1600
rect 8850 900 8950 1600
rect 9000 900 9100 1600
rect 9150 900 9250 1600
rect 9300 900 9400 1600
rect 9450 900 9550 1600
rect 9600 900 9700 1600
rect 9750 900 9850 1600
rect 9900 900 10000 1600
rect 10050 900 10150 1600
rect 10200 900 10300 1600
rect 10350 900 10450 1600
rect 10500 900 10600 1600
rect 10650 900 10750 1600
rect 10800 900 10900 1600
rect 10950 900 11050 1600
rect 11100 900 11200 1600
rect 11250 900 11350 1600
rect 11400 900 11500 1600
rect 11550 900 11650 1600
rect 11700 900 11800 1600
rect 11850 900 11950 1600
rect 12000 900 12100 1600
rect 12150 900 12250 1600
rect 12300 900 12400 1600
rect 12450 900 12550 1600
rect 12600 900 12700 1600
rect 12750 900 12850 1600
rect 12900 900 13000 1600
rect 13050 900 13150 1600
rect 13200 900 13300 1600
rect 13350 900 13450 1600
rect 13500 900 13600 1600
rect 13650 900 13750 1600
rect 13800 900 13900 1600
rect 13950 900 14050 1600
rect 14100 900 14200 1600
rect 14250 900 14350 1600
rect 14400 900 14500 1600
rect 14550 900 14650 1600
rect 14700 900 14800 1600
rect 14850 900 14950 1600
rect 15000 900 15100 1600
rect 15150 900 15250 1600
rect 15300 900 15400 1600
rect 15450 900 15550 1600
rect 15600 900 15700 1600
rect 15750 900 15850 1600
rect 15900 900 16000 1600
rect 16050 900 16150 1600
rect 16200 900 16300 1600
rect 16350 900 16450 1600
rect 16500 900 16600 1600
rect 16650 900 16750 1600
rect 16800 900 16900 1600
rect 16950 900 17050 1600
rect 17100 900 17200 1600
rect 17250 900 17350 1600
rect 17400 900 17500 1600
rect 17550 900 17650 1600
rect 17700 900 17800 1600
rect 17850 900 17950 1600
rect 18000 900 18100 1600
rect 18150 900 18250 1600
rect 18300 900 18400 1600
rect 18450 900 18550 1600
rect 18600 900 18700 1600
rect 18750 900 18850 1600
rect 18900 900 19000 1600
rect 19050 900 19150 1600
rect 19200 900 19300 1600
rect 19350 900 19450 1600
rect 19500 900 19600 1600
rect 19650 900 19750 1600
rect 19800 900 19900 1600
rect 19950 900 20050 1600
rect 20100 900 20200 1600
rect 20250 900 20350 1600
rect -600 50 -500 750
rect -450 50 -350 750
rect -300 50 -200 750
rect -150 50 -50 750
rect 0 50 100 750
rect 150 50 250 750
rect 300 50 400 750
rect 450 50 550 750
rect 600 50 700 750
rect 750 50 850 750
rect 900 50 1000 750
rect 1050 50 1150 750
rect 1200 50 1300 750
rect 1350 50 1450 750
rect 1500 50 1600 750
rect 1650 50 1750 750
rect 1800 50 1900 750
rect 1950 50 2050 750
rect 2100 50 2200 750
rect 2250 50 2350 750
rect 2400 50 2500 750
rect 2550 50 2650 750
rect 2700 50 2800 750
rect 2850 50 2950 750
rect 3000 50 3100 750
rect 3150 50 3250 750
rect 3300 50 3400 750
rect 3450 50 3550 750
rect 3600 50 3700 750
rect 3750 50 3850 750
rect 3900 50 4000 750
rect 4050 50 4150 750
rect 4200 50 4300 750
rect 4350 50 4450 750
rect 4500 50 4600 750
rect 4650 50 4750 750
rect 4800 50 4900 750
rect 4950 50 5050 750
rect 5100 50 5200 750
rect 5250 50 5350 750
rect 5400 50 5500 750
rect 5550 50 5650 750
rect 5700 50 5800 750
rect 5850 50 5950 750
rect 6000 50 6100 750
rect 6150 50 6250 750
rect 6300 50 6400 750
rect 6450 50 6550 750
rect 6600 50 6700 750
rect 6750 50 6850 750
rect 6900 50 7000 750
rect 7050 50 7150 750
rect 7200 50 7300 750
rect 7350 50 7450 750
rect 7500 50 7600 750
rect 7650 50 7750 750
rect 7800 50 7900 750
rect 7950 50 8050 750
rect 8100 50 8200 750
rect 8250 50 8350 750
rect 8400 50 8500 750
rect 8550 50 8650 750
rect 8700 50 8800 750
rect 8850 50 8950 750
rect 9000 50 9100 750
rect 9150 50 9250 750
rect 9300 50 9400 750
rect 9450 50 9550 750
rect 9600 50 9700 750
rect 9750 50 9850 750
rect 9900 50 10000 750
rect 10050 50 10150 750
rect 10200 50 10300 750
rect 10350 50 10450 750
rect 10500 50 10600 750
rect 10650 50 10750 750
rect 10800 50 10900 750
rect 10950 50 11050 750
rect 11100 50 11200 750
rect 11250 50 11350 750
rect 11400 50 11500 750
rect 11550 50 11650 750
rect 11700 50 11800 750
rect 11850 50 11950 750
rect 12000 50 12100 750
rect 12150 50 12250 750
rect 12300 50 12400 750
rect 12450 50 12550 750
rect 12600 50 12700 750
rect 12750 50 12850 750
rect 12900 50 13000 750
rect 13050 50 13150 750
rect 13200 50 13300 750
rect 13350 50 13450 750
rect 13500 50 13600 750
rect 13650 50 13750 750
rect 13800 50 13900 750
rect 13950 50 14050 750
rect 14100 50 14200 750
rect 14250 50 14350 750
rect 14400 50 14500 750
rect 14550 50 14650 750
rect 14700 50 14800 750
rect 14850 50 14950 750
rect 15000 50 15100 750
rect 15150 50 15250 750
rect 15300 50 15400 750
rect 15450 50 15550 750
rect 15600 50 15700 750
rect 15750 50 15850 750
rect 15900 50 16000 750
rect 16050 50 16150 750
rect 16200 50 16300 750
rect 16350 50 16450 750
rect 16500 50 16600 750
rect 16650 50 16750 750
rect 16800 50 16900 750
rect 16950 50 17050 750
rect 17100 50 17200 750
rect 17250 50 17350 750
rect 17400 50 17500 750
rect 17550 50 17650 750
rect 17700 50 17800 750
rect 17850 50 17950 750
rect 18000 50 18100 750
rect 18150 50 18250 750
rect 18300 50 18400 750
rect 18450 50 18550 750
rect 18600 50 18700 750
rect 18750 50 18850 750
rect 18900 50 19000 750
rect 19050 50 19150 750
rect 19200 50 19300 750
rect 19350 50 19450 750
rect 19500 50 19600 750
rect 19650 50 19750 750
rect 19800 50 19900 750
rect 19950 50 20050 750
rect 20100 50 20200 750
rect 20250 50 20350 750
rect -600 -800 -500 -100
rect -450 -800 -350 -100
rect -300 -800 -200 -100
rect -150 -800 -50 -100
rect 0 -800 100 -100
rect 150 -800 250 -100
rect 300 -800 400 -100
rect 450 -800 550 -100
rect 600 -800 700 -100
rect 750 -800 850 -100
rect 900 -800 1000 -100
rect 1050 -800 1150 -100
rect 1200 -800 1300 -100
rect 1350 -800 1450 -100
rect 1500 -800 1600 -100
rect 1650 -800 1750 -100
rect 1800 -800 1900 -100
rect 1950 -800 2050 -100
rect 2100 -800 2200 -100
rect 2250 -800 2350 -100
rect 2400 -800 2500 -100
rect 2550 -800 2650 -100
rect 2700 -800 2800 -100
rect 2850 -800 2950 -100
rect 3000 -800 3100 -100
rect 3150 -800 3250 -100
rect 3300 -800 3400 -100
rect 3450 -800 3550 -100
rect 3600 -800 3700 -100
rect 3750 -800 3850 -100
rect 3900 -800 4000 -100
rect 4050 -800 4150 -100
rect 4200 -800 4300 -100
rect 4350 -800 4450 -100
rect 4500 -800 4600 -100
rect 4650 -800 4750 -100
rect 4800 -800 4900 -100
rect 4950 -800 5050 -100
rect 5100 -800 5200 -100
rect 5250 -800 5350 -100
rect 5400 -800 5500 -100
rect 5550 -800 5650 -100
rect 5700 -800 5800 -100
rect 5850 -800 5950 -100
rect 6000 -800 6100 -100
rect 6150 -800 6250 -100
rect 6300 -800 6400 -100
rect 6450 -800 6550 -100
rect 6600 -800 6700 -100
rect 6750 -800 6850 -100
rect 6900 -800 7000 -100
rect 7050 -800 7150 -100
rect 7200 -800 7300 -100
rect 7350 -800 7450 -100
rect 7500 -800 7600 -100
rect 7650 -800 7750 -100
rect 7800 -800 7900 -100
rect 7950 -800 8050 -100
rect 8100 -800 8200 -100
rect 8250 -800 8350 -100
rect 8400 -800 8500 -100
rect 8550 -800 8650 -100
rect 8700 -800 8800 -100
rect 8850 -800 8950 -100
rect 9000 -800 9100 -100
rect 9150 -800 9250 -100
rect 9300 -800 9400 -100
rect 9450 -800 9550 -100
rect 9600 -800 9700 -100
rect 9750 -800 9850 -100
rect 9900 -800 10000 -100
rect 10050 -800 10150 -100
rect 10200 -800 10300 -100
rect 10350 -800 10450 -100
rect 10500 -800 10600 -100
rect 10650 -800 10750 -100
rect 10800 -800 10900 -100
rect 10950 -800 11050 -100
rect 11100 -800 11200 -100
rect 11250 -800 11350 -100
rect 11400 -800 11500 -100
rect 11550 -800 11650 -100
rect 11700 -800 11800 -100
rect 11850 -800 11950 -100
rect 12000 -800 12100 -100
rect 12150 -800 12250 -100
rect 12300 -800 12400 -100
rect 12450 -800 12550 -100
rect 12600 -800 12700 -100
rect 12750 -800 12850 -100
rect 12900 -800 13000 -100
rect 13050 -800 13150 -100
rect 13200 -800 13300 -100
rect 13350 -800 13450 -100
rect 13500 -800 13600 -100
rect 13650 -800 13750 -100
rect 13800 -800 13900 -100
rect 13950 -800 14050 -100
rect 14100 -800 14200 -100
rect 14250 -800 14350 -100
rect 14400 -800 14500 -100
rect 14550 -800 14650 -100
rect 14700 -800 14800 -100
rect 14850 -800 14950 -100
rect 15000 -800 15100 -100
rect 15150 -800 15250 -100
rect 15300 -800 15400 -100
rect 15450 -800 15550 -100
rect 15600 -800 15700 -100
rect 15750 -800 15850 -100
rect 15900 -800 16000 -100
rect 16050 -800 16150 -100
rect 16200 -800 16300 -100
rect 16350 -800 16450 -100
rect 16500 -800 16600 -100
rect 16650 -800 16750 -100
rect 16800 -800 16900 -100
rect 16950 -800 17050 -100
rect 17100 -800 17200 -100
rect 17250 -800 17350 -100
rect 17400 -800 17500 -100
rect 17550 -800 17650 -100
rect 17700 -800 17800 -100
rect 17850 -800 17950 -100
rect 18000 -800 18100 -100
rect 18150 -800 18250 -100
rect 18300 -800 18400 -100
rect 18450 -800 18550 -100
rect 18600 -800 18700 -100
rect 18750 -800 18850 -100
rect 18900 -800 19000 -100
rect 19050 -800 19150 -100
rect 19200 -800 19300 -100
rect 19350 -800 19450 -100
rect 19500 -800 19600 -100
rect 19650 -800 19750 -100
rect 19800 -800 19900 -100
rect 19950 -800 20050 -100
rect 20100 -800 20200 -100
rect 20250 -800 20350 -100
rect -600 -1650 -500 -950
rect -450 -1650 -350 -950
rect -300 -1650 -200 -950
rect -150 -1650 -50 -950
rect 0 -1650 100 -950
rect 150 -1650 250 -950
rect 300 -1650 400 -950
rect 450 -1650 550 -950
rect 600 -1650 700 -950
rect 750 -1650 850 -950
rect 900 -1650 1000 -950
rect 1050 -1650 1150 -950
rect 1200 -1650 1300 -950
rect 1350 -1650 1450 -950
rect 1500 -1650 1600 -950
rect 1650 -1650 1750 -950
rect 1800 -1650 1900 -950
rect 1950 -1650 2050 -950
rect 2100 -1650 2200 -950
rect 2250 -1650 2350 -950
rect 2400 -1650 2500 -950
rect 2550 -1650 2650 -950
rect 2700 -1650 2800 -950
rect 2850 -1650 2950 -950
rect 3000 -1650 3100 -950
rect 3150 -1650 3250 -950
rect 3300 -1650 3400 -950
rect 3450 -1650 3550 -950
rect 3600 -1650 3700 -950
rect 3750 -1650 3850 -950
rect 3900 -1650 4000 -950
rect 4050 -1650 4150 -950
rect 4200 -1650 4300 -950
rect 4350 -1650 4450 -950
rect 4500 -1650 4600 -950
rect 4650 -1650 4750 -950
rect 4800 -1650 4900 -950
rect 4950 -1650 5050 -950
rect 5100 -1650 5200 -950
rect 5250 -1650 5350 -950
rect 5400 -1650 5500 -950
rect 5550 -1650 5650 -950
rect 5700 -1650 5800 -950
rect 5850 -1650 5950 -950
rect 6000 -1650 6100 -950
rect 6150 -1650 6250 -950
rect 6300 -1650 6400 -950
rect 6450 -1650 6550 -950
rect 6600 -1650 6700 -950
rect 6750 -1650 6850 -950
rect 6900 -1650 7000 -950
rect 7050 -1650 7150 -950
rect 7200 -1650 7300 -950
rect 7350 -1650 7450 -950
rect 7500 -1650 7600 -950
rect 7650 -1650 7750 -950
rect 7800 -1650 7900 -950
rect 7950 -1650 8050 -950
rect 8100 -1650 8200 -950
rect 8250 -1650 8350 -950
rect 8400 -1650 8500 -950
rect 8550 -1650 8650 -950
rect 8700 -1650 8800 -950
rect 8850 -1650 8950 -950
rect 9000 -1650 9100 -950
rect 9150 -1650 9250 -950
rect 9300 -1650 9400 -950
rect 9450 -1650 9550 -950
rect 9600 -1650 9700 -950
rect 9750 -1650 9850 -950
rect 9900 -1650 10000 -950
rect 10050 -1650 10150 -950
rect 10200 -1650 10300 -950
rect 10350 -1650 10450 -950
rect 10500 -1650 10600 -950
rect 10650 -1650 10750 -950
rect 10800 -1650 10900 -950
rect 10950 -1650 11050 -950
rect 11100 -1650 11200 -950
rect 11250 -1650 11350 -950
rect 11400 -1650 11500 -950
rect 11550 -1650 11650 -950
rect 11700 -1650 11800 -950
rect 11850 -1650 11950 -950
rect 12000 -1650 12100 -950
rect 12150 -1650 12250 -950
rect 12300 -1650 12400 -950
rect 12450 -1650 12550 -950
rect 12600 -1650 12700 -950
rect 12750 -1650 12850 -950
rect 12900 -1650 13000 -950
rect 13050 -1650 13150 -950
rect 13200 -1650 13300 -950
rect 13350 -1650 13450 -950
rect 13500 -1650 13600 -950
rect 13650 -1650 13750 -950
rect 13800 -1650 13900 -950
rect 13950 -1650 14050 -950
rect 14100 -1650 14200 -950
rect 14250 -1650 14350 -950
rect 14400 -1650 14500 -950
rect 14550 -1650 14650 -950
rect 14700 -1650 14800 -950
rect 14850 -1650 14950 -950
rect 15000 -1650 15100 -950
rect 15150 -1650 15250 -950
rect 15300 -1650 15400 -950
rect 15450 -1650 15550 -950
rect 15600 -1650 15700 -950
rect 15750 -1650 15850 -950
rect 15900 -1650 16000 -950
rect 16050 -1650 16150 -950
rect 16200 -1650 16300 -950
rect 16350 -1650 16450 -950
rect 16500 -1650 16600 -950
rect 16650 -1650 16750 -950
rect 16800 -1650 16900 -950
rect 16950 -1650 17050 -950
rect 17100 -1650 17200 -950
rect 17250 -1650 17350 -950
rect 17400 -1650 17500 -950
rect 17550 -1650 17650 -950
rect 17700 -1650 17800 -950
rect 17850 -1650 17950 -950
rect 18000 -1650 18100 -950
rect 18150 -1650 18250 -950
rect 18300 -1650 18400 -950
rect 18450 -1650 18550 -950
rect 18600 -1650 18700 -950
rect 18750 -1650 18850 -950
rect 18900 -1650 19000 -950
rect 19050 -1650 19150 -950
rect 19200 -1650 19300 -950
rect 19350 -1650 19450 -950
rect 19500 -1650 19600 -950
rect 19650 -1650 19750 -950
rect 19800 -1650 19900 -950
rect 19950 -1650 20050 -950
rect 20100 -1650 20200 -950
rect 20250 -1650 20350 -950
<< mvpmos >>
rect -600 4600 -500 5100
rect -450 4600 -350 5100
rect -300 4600 -200 5100
rect -150 4600 -50 5100
rect 0 4600 100 5100
rect 150 4600 250 5100
rect 300 4600 400 5100
rect 450 4600 550 5100
rect 600 4600 700 5100
rect 750 4600 850 5100
rect 900 4600 1000 5100
rect 1050 4600 1150 5100
rect 1200 4600 1300 5100
rect 1350 4600 1450 5100
rect 1500 4600 1600 5100
rect 1650 4600 1750 5100
rect 1800 4600 1900 5100
rect 1950 4600 2050 5100
rect 2100 4600 2200 5100
rect 2250 4600 2350 5100
rect 2400 4600 2500 5100
rect 2550 4600 2650 5100
rect 2700 4600 2800 5100
rect 2850 4600 2950 5100
rect 3000 4600 3100 5100
rect 3150 4600 3250 5100
rect 3300 4600 3400 5100
rect 3450 4600 3550 5100
rect 3600 4600 3700 5100
rect 3750 4600 3850 5100
rect 3900 4600 4000 5100
rect 4050 4600 4150 5100
rect 4200 4600 4300 5100
rect 4350 4600 4450 5100
rect 4500 4600 4600 5100
rect 4650 4600 4750 5100
rect 4800 4600 4900 5100
rect 4950 4600 5050 5100
rect 5100 4600 5200 5100
rect 5250 4600 5350 5100
rect 5400 4600 5500 5100
rect 5550 4600 5650 5100
rect 5700 4600 5800 5100
rect 5850 4600 5950 5100
rect 6000 4600 6100 5100
rect 6150 4600 6250 5100
rect 6300 4600 6400 5100
rect 6450 4600 6550 5100
rect 6600 4600 6700 5100
rect 6750 4600 6850 5100
rect 6900 4600 7000 5100
rect 7050 4600 7150 5100
rect 7200 4600 7300 5100
rect 7350 4600 7450 5100
rect 7500 4600 7600 5100
rect 7650 4600 7750 5100
rect 7800 4600 7900 5100
rect 7950 4600 8050 5100
rect 8100 4600 8200 5100
rect 8250 4600 8350 5100
rect 8400 4600 8500 5100
rect 8550 4600 8650 5100
rect 8700 4600 8800 5100
rect 8850 4600 8950 5100
rect 9000 4600 9100 5100
rect 9150 4600 9250 5100
rect 9300 4600 9400 5100
rect 9450 4600 9550 5100
rect 9600 4600 9700 5100
rect 9750 4600 9850 5100
rect 9900 4600 10000 5100
rect 10050 4600 10150 5100
rect 10200 4600 10300 5100
rect 10350 4600 10450 5100
rect 10500 4600 10600 5100
rect 10650 4600 10750 5100
rect 10800 4600 10900 5100
rect 10950 4600 11050 5100
rect 11100 4600 11200 5100
rect 11250 4600 11350 5100
rect 11400 4600 11500 5100
rect 11550 4600 11650 5100
rect 11700 4600 11800 5100
rect 11850 4600 11950 5100
rect 12000 4600 12100 5100
rect 12150 4600 12250 5100
rect 12300 4600 12400 5100
rect 12450 4600 12550 5100
rect 12600 4600 12700 5100
rect 12750 4600 12850 5100
rect 12900 4600 13000 5100
rect 13050 4600 13150 5100
rect 13200 4600 13300 5100
rect 13350 4600 13450 5100
rect 13500 4600 13600 5100
rect 13650 4600 13750 5100
rect 13800 4600 13900 5100
rect 13950 4600 14050 5100
rect 14100 4600 14200 5100
rect 14250 4600 14350 5100
rect 14400 4600 14500 5100
rect 14550 4600 14650 5100
rect 14700 4600 14800 5100
rect 14850 4600 14950 5100
rect 15000 4600 15100 5100
rect 15150 4600 15250 5100
rect 15300 4600 15400 5100
rect 15450 4600 15550 5100
rect 15600 4600 15700 5100
rect 15750 4600 15850 5100
rect 15900 4600 16000 5100
rect 16050 4600 16150 5100
rect 16200 4600 16300 5100
rect 16350 4600 16450 5100
rect 16500 4600 16600 5100
rect 16650 4600 16750 5100
rect 16800 4600 16900 5100
rect 16950 4600 17050 5100
rect 17100 4600 17200 5100
rect 17250 4600 17350 5100
rect 17400 4600 17500 5100
rect 17550 4600 17650 5100
rect 17700 4600 17800 5100
rect 17850 4600 17950 5100
rect 18000 4600 18100 5100
rect 18150 4600 18250 5100
rect 18300 4600 18400 5100
rect 18450 4600 18550 5100
rect 18600 4600 18700 5100
rect 18750 4600 18850 5100
rect 18900 4600 19000 5100
rect 19050 4600 19150 5100
rect 19200 4600 19300 5100
rect 19350 4600 19450 5100
rect 19500 4600 19600 5100
rect 19650 4600 19750 5100
rect 19800 4600 19900 5100
rect 19950 4600 20050 5100
rect 20100 4600 20200 5100
rect 20250 4600 20350 5100
rect -600 3950 -500 4450
rect -450 3950 -350 4450
rect -300 3950 -200 4450
rect -150 3950 -50 4450
rect 0 3950 100 4450
rect 150 3950 250 4450
rect 300 3950 400 4450
rect 450 3950 550 4450
rect 600 3950 700 4450
rect 750 3950 850 4450
rect 900 3950 1000 4450
rect 1050 3950 1150 4450
rect 1200 3950 1300 4450
rect 1350 3950 1450 4450
rect 1500 3950 1600 4450
rect 1650 3950 1750 4450
rect 1800 3950 1900 4450
rect 1950 3950 2050 4450
rect 2100 3950 2200 4450
rect 2250 3950 2350 4450
rect 2400 3950 2500 4450
rect 2550 3950 2650 4450
rect 2700 3950 2800 4450
rect 2850 3950 2950 4450
rect 3000 3950 3100 4450
rect 3150 3950 3250 4450
rect 3300 3950 3400 4450
rect 3450 3950 3550 4450
rect 3600 3950 3700 4450
rect 3750 3950 3850 4450
rect 3900 3950 4000 4450
rect 4050 3950 4150 4450
rect 4200 3950 4300 4450
rect 4350 3950 4450 4450
rect 4500 3950 4600 4450
rect 4650 3950 4750 4450
rect 4800 3950 4900 4450
rect 4950 3950 5050 4450
rect 5100 3950 5200 4450
rect 5250 3950 5350 4450
rect 5400 3950 5500 4450
rect 5550 3950 5650 4450
rect 5700 3950 5800 4450
rect 5850 3950 5950 4450
rect 6000 3950 6100 4450
rect 6150 3950 6250 4450
rect 6300 3950 6400 4450
rect 6450 3950 6550 4450
rect 6600 3950 6700 4450
rect 6750 3950 6850 4450
rect 6900 3950 7000 4450
rect 7050 3950 7150 4450
rect 7200 3950 7300 4450
rect 7350 3950 7450 4450
rect 7500 3950 7600 4450
rect 7650 3950 7750 4450
rect 7800 3950 7900 4450
rect 7950 3950 8050 4450
rect 8100 3950 8200 4450
rect 8250 3950 8350 4450
rect 8400 3950 8500 4450
rect 8550 3950 8650 4450
rect 8700 3950 8800 4450
rect 8850 3950 8950 4450
rect 9000 3950 9100 4450
rect 9150 3950 9250 4450
rect 9300 3950 9400 4450
rect 9450 3950 9550 4450
rect 9600 3950 9700 4450
rect 9750 3950 9850 4450
rect 9900 3950 10000 4450
rect 10050 3950 10150 4450
rect 10200 3950 10300 4450
rect 10350 3950 10450 4450
rect 10500 3950 10600 4450
rect 10650 3950 10750 4450
rect 10800 3950 10900 4450
rect 10950 3950 11050 4450
rect 11100 3950 11200 4450
rect 11250 3950 11350 4450
rect 11400 3950 11500 4450
rect 11550 3950 11650 4450
rect 11700 3950 11800 4450
rect 11850 3950 11950 4450
rect 12000 3950 12100 4450
rect 12150 3950 12250 4450
rect 12300 3950 12400 4450
rect 12450 3950 12550 4450
rect 12600 3950 12700 4450
rect 12750 3950 12850 4450
rect 12900 3950 13000 4450
rect 13050 3950 13150 4450
rect 13200 3950 13300 4450
rect 13350 3950 13450 4450
rect 13500 3950 13600 4450
rect 13650 3950 13750 4450
rect 13800 3950 13900 4450
rect 13950 3950 14050 4450
rect 14100 3950 14200 4450
rect 14250 3950 14350 4450
rect 14400 3950 14500 4450
rect 14550 3950 14650 4450
rect 14700 3950 14800 4450
rect 14850 3950 14950 4450
rect 15000 3950 15100 4450
rect 15150 3950 15250 4450
rect 15300 3950 15400 4450
rect 15450 3950 15550 4450
rect 15600 3950 15700 4450
rect 15750 3950 15850 4450
rect 15900 3950 16000 4450
rect 16050 3950 16150 4450
rect 16200 3950 16300 4450
rect 16350 3950 16450 4450
rect 16500 3950 16600 4450
rect 16650 3950 16750 4450
rect 16800 3950 16900 4450
rect 16950 3950 17050 4450
rect 17100 3950 17200 4450
rect 17250 3950 17350 4450
rect 17400 3950 17500 4450
rect 17550 3950 17650 4450
rect 17700 3950 17800 4450
rect 17850 3950 17950 4450
rect 18000 3950 18100 4450
rect 18150 3950 18250 4450
rect 18300 3950 18400 4450
rect 18450 3950 18550 4450
rect 18600 3950 18700 4450
rect 18750 3950 18850 4450
rect 18900 3950 19000 4450
rect 19050 3950 19150 4450
rect 19200 3950 19300 4450
rect 19350 3950 19450 4450
rect 19500 3950 19600 4450
rect 19650 3950 19750 4450
rect 19800 3950 19900 4450
rect 19950 3950 20050 4450
rect 20100 3950 20200 4450
rect 20250 3950 20350 4450
rect -600 3300 -500 3800
rect -450 3300 -350 3800
rect -300 3300 -200 3800
rect -150 3300 -50 3800
rect 0 3300 100 3800
rect 150 3300 250 3800
rect 300 3300 400 3800
rect 450 3300 550 3800
rect 600 3300 700 3800
rect 750 3300 850 3800
rect 900 3300 1000 3800
rect 1050 3300 1150 3800
rect 1200 3300 1300 3800
rect 1350 3300 1450 3800
rect 1500 3300 1600 3800
rect 1650 3300 1750 3800
rect 1800 3300 1900 3800
rect 1950 3300 2050 3800
rect 2100 3300 2200 3800
rect 2250 3300 2350 3800
rect 2400 3300 2500 3800
rect 2550 3300 2650 3800
rect 2700 3300 2800 3800
rect 2850 3300 2950 3800
rect 3000 3300 3100 3800
rect 3150 3300 3250 3800
rect 3300 3300 3400 3800
rect 3450 3300 3550 3800
rect 3600 3300 3700 3800
rect 3750 3300 3850 3800
rect 3900 3300 4000 3800
rect 4050 3300 4150 3800
rect 4200 3300 4300 3800
rect 4350 3300 4450 3800
rect 4500 3300 4600 3800
rect 4650 3300 4750 3800
rect 4800 3300 4900 3800
rect 4950 3300 5050 3800
rect 5100 3300 5200 3800
rect 5250 3300 5350 3800
rect 5400 3300 5500 3800
rect 5550 3300 5650 3800
rect 5700 3300 5800 3800
rect 5850 3300 5950 3800
rect 6000 3300 6100 3800
rect 6150 3300 6250 3800
rect 6300 3300 6400 3800
rect 6450 3300 6550 3800
rect 6600 3300 6700 3800
rect 6750 3300 6850 3800
rect 6900 3300 7000 3800
rect 7050 3300 7150 3800
rect 7200 3300 7300 3800
rect 7350 3300 7450 3800
rect 7500 3300 7600 3800
rect 7650 3300 7750 3800
rect 7800 3300 7900 3800
rect 7950 3300 8050 3800
rect 8100 3300 8200 3800
rect 8250 3300 8350 3800
rect 8400 3300 8500 3800
rect 8550 3300 8650 3800
rect 8700 3300 8800 3800
rect 8850 3300 8950 3800
rect 9000 3300 9100 3800
rect 9150 3300 9250 3800
rect 9300 3300 9400 3800
rect 9450 3300 9550 3800
rect 9600 3300 9700 3800
rect 9750 3300 9850 3800
rect 9900 3300 10000 3800
rect 10050 3300 10150 3800
rect 10200 3300 10300 3800
rect 10350 3300 10450 3800
rect 10500 3300 10600 3800
rect 10650 3300 10750 3800
rect 10800 3300 10900 3800
rect 10950 3300 11050 3800
rect 11100 3300 11200 3800
rect 11250 3300 11350 3800
rect 11400 3300 11500 3800
rect 11550 3300 11650 3800
rect 11700 3300 11800 3800
rect 11850 3300 11950 3800
rect 12000 3300 12100 3800
rect 12150 3300 12250 3800
rect 12300 3300 12400 3800
rect 12450 3300 12550 3800
rect 12600 3300 12700 3800
rect 12750 3300 12850 3800
rect 12900 3300 13000 3800
rect 13050 3300 13150 3800
rect 13200 3300 13300 3800
rect 13350 3300 13450 3800
rect 13500 3300 13600 3800
rect 13650 3300 13750 3800
rect 13800 3300 13900 3800
rect 13950 3300 14050 3800
rect 14100 3300 14200 3800
rect 14250 3300 14350 3800
rect 14400 3300 14500 3800
rect 14550 3300 14650 3800
rect 14700 3300 14800 3800
rect 14850 3300 14950 3800
rect 15000 3300 15100 3800
rect 15150 3300 15250 3800
rect 15300 3300 15400 3800
rect 15450 3300 15550 3800
rect 15600 3300 15700 3800
rect 15750 3300 15850 3800
rect 15900 3300 16000 3800
rect 16050 3300 16150 3800
rect 16200 3300 16300 3800
rect 16350 3300 16450 3800
rect 16500 3300 16600 3800
rect 16650 3300 16750 3800
rect 16800 3300 16900 3800
rect 16950 3300 17050 3800
rect 17100 3300 17200 3800
rect 17250 3300 17350 3800
rect 17400 3300 17500 3800
rect 17550 3300 17650 3800
rect 17700 3300 17800 3800
rect 17850 3300 17950 3800
rect 18000 3300 18100 3800
rect 18150 3300 18250 3800
rect 18300 3300 18400 3800
rect 18450 3300 18550 3800
rect 18600 3300 18700 3800
rect 18750 3300 18850 3800
rect 18900 3300 19000 3800
rect 19050 3300 19150 3800
rect 19200 3300 19300 3800
rect 19350 3300 19450 3800
rect 19500 3300 19600 3800
rect 19650 3300 19750 3800
rect 19800 3300 19900 3800
rect 19950 3300 20050 3800
rect 20100 3300 20200 3800
rect 20250 3300 20350 3800
rect -600 2650 -500 3150
rect -450 2650 -350 3150
rect -300 2650 -200 3150
rect -150 2650 -50 3150
rect 0 2650 100 3150
rect 150 2650 250 3150
rect 300 2650 400 3150
rect 450 2650 550 3150
rect 600 2650 700 3150
rect 750 2650 850 3150
rect 900 2650 1000 3150
rect 1050 2650 1150 3150
rect 1200 2650 1300 3150
rect 1350 2650 1450 3150
rect 1500 2650 1600 3150
rect 1650 2650 1750 3150
rect 1800 2650 1900 3150
rect 1950 2650 2050 3150
rect 2100 2650 2200 3150
rect 2250 2650 2350 3150
rect 2400 2650 2500 3150
rect 2550 2650 2650 3150
rect 2700 2650 2800 3150
rect 2850 2650 2950 3150
rect 3000 2650 3100 3150
rect 3150 2650 3250 3150
rect 3300 2650 3400 3150
rect 3450 2650 3550 3150
rect 3600 2650 3700 3150
rect 3750 2650 3850 3150
rect 3900 2650 4000 3150
rect 4050 2650 4150 3150
rect 4200 2650 4300 3150
rect 4350 2650 4450 3150
rect 4500 2650 4600 3150
rect 4650 2650 4750 3150
rect 4800 2650 4900 3150
rect 4950 2650 5050 3150
rect 5100 2650 5200 3150
rect 5250 2650 5350 3150
rect 5400 2650 5500 3150
rect 5550 2650 5650 3150
rect 5700 2650 5800 3150
rect 5850 2650 5950 3150
rect 6000 2650 6100 3150
rect 6150 2650 6250 3150
rect 6300 2650 6400 3150
rect 6450 2650 6550 3150
rect 6600 2650 6700 3150
rect 6750 2650 6850 3150
rect 6900 2650 7000 3150
rect 7050 2650 7150 3150
rect 7200 2650 7300 3150
rect 7350 2650 7450 3150
rect 7500 2650 7600 3150
rect 7650 2650 7750 3150
rect 7800 2650 7900 3150
rect 7950 2650 8050 3150
rect 8100 2650 8200 3150
rect 8250 2650 8350 3150
rect 8400 2650 8500 3150
rect 8550 2650 8650 3150
rect 8700 2650 8800 3150
rect 8850 2650 8950 3150
rect 9000 2650 9100 3150
rect 9150 2650 9250 3150
rect 9300 2650 9400 3150
rect 9450 2650 9550 3150
rect 9600 2650 9700 3150
rect 9750 2650 9850 3150
rect 9900 2650 10000 3150
rect 10050 2650 10150 3150
rect 10200 2650 10300 3150
rect 10350 2650 10450 3150
rect 10500 2650 10600 3150
rect 10650 2650 10750 3150
rect 10800 2650 10900 3150
rect 10950 2650 11050 3150
rect 11100 2650 11200 3150
rect 11250 2650 11350 3150
rect 11400 2650 11500 3150
rect 11550 2650 11650 3150
rect 11700 2650 11800 3150
rect 11850 2650 11950 3150
rect 12000 2650 12100 3150
rect 12150 2650 12250 3150
rect 12300 2650 12400 3150
rect 12450 2650 12550 3150
rect 12600 2650 12700 3150
rect 12750 2650 12850 3150
rect 12900 2650 13000 3150
rect 13050 2650 13150 3150
rect 13200 2650 13300 3150
rect 13350 2650 13450 3150
rect 13500 2650 13600 3150
rect 13650 2650 13750 3150
rect 13800 2650 13900 3150
rect 13950 2650 14050 3150
rect 14100 2650 14200 3150
rect 14250 2650 14350 3150
rect 14400 2650 14500 3150
rect 14550 2650 14650 3150
rect 14700 2650 14800 3150
rect 14850 2650 14950 3150
rect 15000 2650 15100 3150
rect 15150 2650 15250 3150
rect 15300 2650 15400 3150
rect 15450 2650 15550 3150
rect 15600 2650 15700 3150
rect 15750 2650 15850 3150
rect 15900 2650 16000 3150
rect 16050 2650 16150 3150
rect 16200 2650 16300 3150
rect 16350 2650 16450 3150
rect 16500 2650 16600 3150
rect 16650 2650 16750 3150
rect 16800 2650 16900 3150
rect 16950 2650 17050 3150
rect 17100 2650 17200 3150
rect 17250 2650 17350 3150
rect 17400 2650 17500 3150
rect 17550 2650 17650 3150
rect 17700 2650 17800 3150
rect 17850 2650 17950 3150
rect 18000 2650 18100 3150
rect 18150 2650 18250 3150
rect 18300 2650 18400 3150
rect 18450 2650 18550 3150
rect 18600 2650 18700 3150
rect 18750 2650 18850 3150
rect 18900 2650 19000 3150
rect 19050 2650 19150 3150
rect 19200 2650 19300 3150
rect 19350 2650 19450 3150
rect 19500 2650 19600 3150
rect 19650 2650 19750 3150
rect 19800 2650 19900 3150
rect 19950 2650 20050 3150
rect 20100 2650 20200 3150
rect 20250 2650 20350 3150
<< mvndiff >>
rect -650 1585 -600 1600
rect -650 1565 -635 1585
rect -615 1565 -600 1585
rect -650 1535 -600 1565
rect -650 1515 -635 1535
rect -615 1515 -600 1535
rect -650 1485 -600 1515
rect -650 1465 -635 1485
rect -615 1465 -600 1485
rect -650 1435 -600 1465
rect -650 1415 -635 1435
rect -615 1415 -600 1435
rect -650 1385 -600 1415
rect -650 1365 -635 1385
rect -615 1365 -600 1385
rect -650 1335 -600 1365
rect -650 1315 -635 1335
rect -615 1315 -600 1335
rect -650 1285 -600 1315
rect -650 1265 -635 1285
rect -615 1265 -600 1285
rect -650 1235 -600 1265
rect -650 1215 -635 1235
rect -615 1215 -600 1235
rect -650 1185 -600 1215
rect -650 1165 -635 1185
rect -615 1165 -600 1185
rect -650 1135 -600 1165
rect -650 1115 -635 1135
rect -615 1115 -600 1135
rect -650 1085 -600 1115
rect -650 1065 -635 1085
rect -615 1065 -600 1085
rect -650 1035 -600 1065
rect -650 1015 -635 1035
rect -615 1015 -600 1035
rect -650 985 -600 1015
rect -650 965 -635 985
rect -615 965 -600 985
rect -650 935 -600 965
rect -650 915 -635 935
rect -615 915 -600 935
rect -650 900 -600 915
rect -500 1585 -450 1600
rect -500 1565 -485 1585
rect -465 1565 -450 1585
rect -500 1535 -450 1565
rect -500 1515 -485 1535
rect -465 1515 -450 1535
rect -500 1485 -450 1515
rect -500 1465 -485 1485
rect -465 1465 -450 1485
rect -500 1435 -450 1465
rect -500 1415 -485 1435
rect -465 1415 -450 1435
rect -500 1385 -450 1415
rect -500 1365 -485 1385
rect -465 1365 -450 1385
rect -500 1335 -450 1365
rect -500 1315 -485 1335
rect -465 1315 -450 1335
rect -500 1285 -450 1315
rect -500 1265 -485 1285
rect -465 1265 -450 1285
rect -500 1235 -450 1265
rect -500 1215 -485 1235
rect -465 1215 -450 1235
rect -500 1185 -450 1215
rect -500 1165 -485 1185
rect -465 1165 -450 1185
rect -500 1135 -450 1165
rect -500 1115 -485 1135
rect -465 1115 -450 1135
rect -500 1085 -450 1115
rect -500 1065 -485 1085
rect -465 1065 -450 1085
rect -500 1035 -450 1065
rect -500 1015 -485 1035
rect -465 1015 -450 1035
rect -500 985 -450 1015
rect -500 965 -485 985
rect -465 965 -450 985
rect -500 935 -450 965
rect -500 915 -485 935
rect -465 915 -450 935
rect -500 900 -450 915
rect -350 1585 -300 1600
rect -350 1565 -335 1585
rect -315 1565 -300 1585
rect -350 1535 -300 1565
rect -350 1515 -335 1535
rect -315 1515 -300 1535
rect -350 1485 -300 1515
rect -350 1465 -335 1485
rect -315 1465 -300 1485
rect -350 1435 -300 1465
rect -350 1415 -335 1435
rect -315 1415 -300 1435
rect -350 1385 -300 1415
rect -350 1365 -335 1385
rect -315 1365 -300 1385
rect -350 1335 -300 1365
rect -350 1315 -335 1335
rect -315 1315 -300 1335
rect -350 1285 -300 1315
rect -350 1265 -335 1285
rect -315 1265 -300 1285
rect -350 1235 -300 1265
rect -350 1215 -335 1235
rect -315 1215 -300 1235
rect -350 1185 -300 1215
rect -350 1165 -335 1185
rect -315 1165 -300 1185
rect -350 1135 -300 1165
rect -350 1115 -335 1135
rect -315 1115 -300 1135
rect -350 1085 -300 1115
rect -350 1065 -335 1085
rect -315 1065 -300 1085
rect -350 1035 -300 1065
rect -350 1015 -335 1035
rect -315 1015 -300 1035
rect -350 985 -300 1015
rect -350 965 -335 985
rect -315 965 -300 985
rect -350 935 -300 965
rect -350 915 -335 935
rect -315 915 -300 935
rect -350 900 -300 915
rect -200 1585 -150 1600
rect -200 1565 -185 1585
rect -165 1565 -150 1585
rect -200 1535 -150 1565
rect -200 1515 -185 1535
rect -165 1515 -150 1535
rect -200 1485 -150 1515
rect -200 1465 -185 1485
rect -165 1465 -150 1485
rect -200 1435 -150 1465
rect -200 1415 -185 1435
rect -165 1415 -150 1435
rect -200 1385 -150 1415
rect -200 1365 -185 1385
rect -165 1365 -150 1385
rect -200 1335 -150 1365
rect -200 1315 -185 1335
rect -165 1315 -150 1335
rect -200 1285 -150 1315
rect -200 1265 -185 1285
rect -165 1265 -150 1285
rect -200 1235 -150 1265
rect -200 1215 -185 1235
rect -165 1215 -150 1235
rect -200 1185 -150 1215
rect -200 1165 -185 1185
rect -165 1165 -150 1185
rect -200 1135 -150 1165
rect -200 1115 -185 1135
rect -165 1115 -150 1135
rect -200 1085 -150 1115
rect -200 1065 -185 1085
rect -165 1065 -150 1085
rect -200 1035 -150 1065
rect -200 1015 -185 1035
rect -165 1015 -150 1035
rect -200 985 -150 1015
rect -200 965 -185 985
rect -165 965 -150 985
rect -200 935 -150 965
rect -200 915 -185 935
rect -165 915 -150 935
rect -200 900 -150 915
rect -50 1585 0 1600
rect -50 1565 -35 1585
rect -15 1565 0 1585
rect -50 1535 0 1565
rect -50 1515 -35 1535
rect -15 1515 0 1535
rect -50 1485 0 1515
rect -50 1465 -35 1485
rect -15 1465 0 1485
rect -50 1435 0 1465
rect -50 1415 -35 1435
rect -15 1415 0 1435
rect -50 1385 0 1415
rect -50 1365 -35 1385
rect -15 1365 0 1385
rect -50 1335 0 1365
rect -50 1315 -35 1335
rect -15 1315 0 1335
rect -50 1285 0 1315
rect -50 1265 -35 1285
rect -15 1265 0 1285
rect -50 1235 0 1265
rect -50 1215 -35 1235
rect -15 1215 0 1235
rect -50 1185 0 1215
rect -50 1165 -35 1185
rect -15 1165 0 1185
rect -50 1135 0 1165
rect -50 1115 -35 1135
rect -15 1115 0 1135
rect -50 1085 0 1115
rect -50 1065 -35 1085
rect -15 1065 0 1085
rect -50 1035 0 1065
rect -50 1015 -35 1035
rect -15 1015 0 1035
rect -50 985 0 1015
rect -50 965 -35 985
rect -15 965 0 985
rect -50 935 0 965
rect -50 915 -35 935
rect -15 915 0 935
rect -50 900 0 915
rect 100 900 150 1600
rect 250 900 300 1600
rect 400 900 450 1600
rect 550 900 600 1600
rect 700 900 750 1600
rect 850 900 900 1600
rect 1000 900 1050 1600
rect 1150 1585 1200 1600
rect 1150 1565 1165 1585
rect 1185 1565 1200 1585
rect 1150 1535 1200 1565
rect 1150 1515 1165 1535
rect 1185 1515 1200 1535
rect 1150 1485 1200 1515
rect 1150 1465 1165 1485
rect 1185 1465 1200 1485
rect 1150 1435 1200 1465
rect 1150 1415 1165 1435
rect 1185 1415 1200 1435
rect 1150 1385 1200 1415
rect 1150 1365 1165 1385
rect 1185 1365 1200 1385
rect 1150 1335 1200 1365
rect 1150 1315 1165 1335
rect 1185 1315 1200 1335
rect 1150 1285 1200 1315
rect 1150 1265 1165 1285
rect 1185 1265 1200 1285
rect 1150 1235 1200 1265
rect 1150 1215 1165 1235
rect 1185 1215 1200 1235
rect 1150 1185 1200 1215
rect 1150 1165 1165 1185
rect 1185 1165 1200 1185
rect 1150 1135 1200 1165
rect 1150 1115 1165 1135
rect 1185 1115 1200 1135
rect 1150 1085 1200 1115
rect 1150 1065 1165 1085
rect 1185 1065 1200 1085
rect 1150 1035 1200 1065
rect 1150 1015 1165 1035
rect 1185 1015 1200 1035
rect 1150 985 1200 1015
rect 1150 965 1165 985
rect 1185 965 1200 985
rect 1150 935 1200 965
rect 1150 915 1165 935
rect 1185 915 1200 935
rect 1150 900 1200 915
rect 1300 900 1350 1600
rect 1450 1585 1500 1600
rect 1450 1565 1465 1585
rect 1485 1565 1500 1585
rect 1450 1535 1500 1565
rect 1450 1515 1465 1535
rect 1485 1515 1500 1535
rect 1450 1485 1500 1515
rect 1450 1465 1465 1485
rect 1485 1465 1500 1485
rect 1450 1435 1500 1465
rect 1450 1415 1465 1435
rect 1485 1415 1500 1435
rect 1450 1385 1500 1415
rect 1450 1365 1465 1385
rect 1485 1365 1500 1385
rect 1450 1335 1500 1365
rect 1450 1315 1465 1335
rect 1485 1315 1500 1335
rect 1450 1285 1500 1315
rect 1450 1265 1465 1285
rect 1485 1265 1500 1285
rect 1450 1235 1500 1265
rect 1450 1215 1465 1235
rect 1485 1215 1500 1235
rect 1450 1185 1500 1215
rect 1450 1165 1465 1185
rect 1485 1165 1500 1185
rect 1450 1135 1500 1165
rect 1450 1115 1465 1135
rect 1485 1115 1500 1135
rect 1450 1085 1500 1115
rect 1450 1065 1465 1085
rect 1485 1065 1500 1085
rect 1450 1035 1500 1065
rect 1450 1015 1465 1035
rect 1485 1015 1500 1035
rect 1450 985 1500 1015
rect 1450 965 1465 985
rect 1485 965 1500 985
rect 1450 935 1500 965
rect 1450 915 1465 935
rect 1485 915 1500 935
rect 1450 900 1500 915
rect 1600 900 1650 1600
rect 1750 1585 1800 1600
rect 1750 1565 1765 1585
rect 1785 1565 1800 1585
rect 1750 1535 1800 1565
rect 1750 1515 1765 1535
rect 1785 1515 1800 1535
rect 1750 1485 1800 1515
rect 1750 1465 1765 1485
rect 1785 1465 1800 1485
rect 1750 1435 1800 1465
rect 1750 1415 1765 1435
rect 1785 1415 1800 1435
rect 1750 1385 1800 1415
rect 1750 1365 1765 1385
rect 1785 1365 1800 1385
rect 1750 1335 1800 1365
rect 1750 1315 1765 1335
rect 1785 1315 1800 1335
rect 1750 1285 1800 1315
rect 1750 1265 1765 1285
rect 1785 1265 1800 1285
rect 1750 1235 1800 1265
rect 1750 1215 1765 1235
rect 1785 1215 1800 1235
rect 1750 1185 1800 1215
rect 1750 1165 1765 1185
rect 1785 1165 1800 1185
rect 1750 1135 1800 1165
rect 1750 1115 1765 1135
rect 1785 1115 1800 1135
rect 1750 1085 1800 1115
rect 1750 1065 1765 1085
rect 1785 1065 1800 1085
rect 1750 1035 1800 1065
rect 1750 1015 1765 1035
rect 1785 1015 1800 1035
rect 1750 985 1800 1015
rect 1750 965 1765 985
rect 1785 965 1800 985
rect 1750 935 1800 965
rect 1750 915 1765 935
rect 1785 915 1800 935
rect 1750 900 1800 915
rect 1900 900 1950 1600
rect 2050 1585 2100 1600
rect 2050 1565 2065 1585
rect 2085 1565 2100 1585
rect 2050 1535 2100 1565
rect 2050 1515 2065 1535
rect 2085 1515 2100 1535
rect 2050 1485 2100 1515
rect 2050 1465 2065 1485
rect 2085 1465 2100 1485
rect 2050 1435 2100 1465
rect 2050 1415 2065 1435
rect 2085 1415 2100 1435
rect 2050 1385 2100 1415
rect 2050 1365 2065 1385
rect 2085 1365 2100 1385
rect 2050 1335 2100 1365
rect 2050 1315 2065 1335
rect 2085 1315 2100 1335
rect 2050 1285 2100 1315
rect 2050 1265 2065 1285
rect 2085 1265 2100 1285
rect 2050 1235 2100 1265
rect 2050 1215 2065 1235
rect 2085 1215 2100 1235
rect 2050 1185 2100 1215
rect 2050 1165 2065 1185
rect 2085 1165 2100 1185
rect 2050 1135 2100 1165
rect 2050 1115 2065 1135
rect 2085 1115 2100 1135
rect 2050 1085 2100 1115
rect 2050 1065 2065 1085
rect 2085 1065 2100 1085
rect 2050 1035 2100 1065
rect 2050 1015 2065 1035
rect 2085 1015 2100 1035
rect 2050 985 2100 1015
rect 2050 965 2065 985
rect 2085 965 2100 985
rect 2050 935 2100 965
rect 2050 915 2065 935
rect 2085 915 2100 935
rect 2050 900 2100 915
rect 2200 900 2250 1600
rect 2350 1585 2400 1600
rect 2350 1565 2365 1585
rect 2385 1565 2400 1585
rect 2350 1535 2400 1565
rect 2350 1515 2365 1535
rect 2385 1515 2400 1535
rect 2350 1485 2400 1515
rect 2350 1465 2365 1485
rect 2385 1465 2400 1485
rect 2350 1435 2400 1465
rect 2350 1415 2365 1435
rect 2385 1415 2400 1435
rect 2350 1385 2400 1415
rect 2350 1365 2365 1385
rect 2385 1365 2400 1385
rect 2350 1335 2400 1365
rect 2350 1315 2365 1335
rect 2385 1315 2400 1335
rect 2350 1285 2400 1315
rect 2350 1265 2365 1285
rect 2385 1265 2400 1285
rect 2350 1235 2400 1265
rect 2350 1215 2365 1235
rect 2385 1215 2400 1235
rect 2350 1185 2400 1215
rect 2350 1165 2365 1185
rect 2385 1165 2400 1185
rect 2350 1135 2400 1165
rect 2350 1115 2365 1135
rect 2385 1115 2400 1135
rect 2350 1085 2400 1115
rect 2350 1065 2365 1085
rect 2385 1065 2400 1085
rect 2350 1035 2400 1065
rect 2350 1015 2365 1035
rect 2385 1015 2400 1035
rect 2350 985 2400 1015
rect 2350 965 2365 985
rect 2385 965 2400 985
rect 2350 935 2400 965
rect 2350 915 2365 935
rect 2385 915 2400 935
rect 2350 900 2400 915
rect 2500 900 2550 1600
rect 2650 1585 2700 1600
rect 2650 1565 2665 1585
rect 2685 1565 2700 1585
rect 2650 1535 2700 1565
rect 2650 1515 2665 1535
rect 2685 1515 2700 1535
rect 2650 1485 2700 1515
rect 2650 1465 2665 1485
rect 2685 1465 2700 1485
rect 2650 1435 2700 1465
rect 2650 1415 2665 1435
rect 2685 1415 2700 1435
rect 2650 1385 2700 1415
rect 2650 1365 2665 1385
rect 2685 1365 2700 1385
rect 2650 1335 2700 1365
rect 2650 1315 2665 1335
rect 2685 1315 2700 1335
rect 2650 1285 2700 1315
rect 2650 1265 2665 1285
rect 2685 1265 2700 1285
rect 2650 1235 2700 1265
rect 2650 1215 2665 1235
rect 2685 1215 2700 1235
rect 2650 1185 2700 1215
rect 2650 1165 2665 1185
rect 2685 1165 2700 1185
rect 2650 1135 2700 1165
rect 2650 1115 2665 1135
rect 2685 1115 2700 1135
rect 2650 1085 2700 1115
rect 2650 1065 2665 1085
rect 2685 1065 2700 1085
rect 2650 1035 2700 1065
rect 2650 1015 2665 1035
rect 2685 1015 2700 1035
rect 2650 985 2700 1015
rect 2650 965 2665 985
rect 2685 965 2700 985
rect 2650 935 2700 965
rect 2650 915 2665 935
rect 2685 915 2700 935
rect 2650 900 2700 915
rect 2800 900 2850 1600
rect 2950 1585 3000 1600
rect 2950 1565 2965 1585
rect 2985 1565 3000 1585
rect 2950 1535 3000 1565
rect 2950 1515 2965 1535
rect 2985 1515 3000 1535
rect 2950 1485 3000 1515
rect 2950 1465 2965 1485
rect 2985 1465 3000 1485
rect 2950 1435 3000 1465
rect 2950 1415 2965 1435
rect 2985 1415 3000 1435
rect 2950 1385 3000 1415
rect 2950 1365 2965 1385
rect 2985 1365 3000 1385
rect 2950 1335 3000 1365
rect 2950 1315 2965 1335
rect 2985 1315 3000 1335
rect 2950 1285 3000 1315
rect 2950 1265 2965 1285
rect 2985 1265 3000 1285
rect 2950 1235 3000 1265
rect 2950 1215 2965 1235
rect 2985 1215 3000 1235
rect 2950 1185 3000 1215
rect 2950 1165 2965 1185
rect 2985 1165 3000 1185
rect 2950 1135 3000 1165
rect 2950 1115 2965 1135
rect 2985 1115 3000 1135
rect 2950 1085 3000 1115
rect 2950 1065 2965 1085
rect 2985 1065 3000 1085
rect 2950 1035 3000 1065
rect 2950 1015 2965 1035
rect 2985 1015 3000 1035
rect 2950 985 3000 1015
rect 2950 965 2965 985
rect 2985 965 3000 985
rect 2950 935 3000 965
rect 2950 915 2965 935
rect 2985 915 3000 935
rect 2950 900 3000 915
rect 3100 900 3150 1600
rect 3250 1585 3300 1600
rect 3250 1565 3265 1585
rect 3285 1565 3300 1585
rect 3250 1535 3300 1565
rect 3250 1515 3265 1535
rect 3285 1515 3300 1535
rect 3250 1485 3300 1515
rect 3250 1465 3265 1485
rect 3285 1465 3300 1485
rect 3250 1435 3300 1465
rect 3250 1415 3265 1435
rect 3285 1415 3300 1435
rect 3250 1385 3300 1415
rect 3250 1365 3265 1385
rect 3285 1365 3300 1385
rect 3250 1335 3300 1365
rect 3250 1315 3265 1335
rect 3285 1315 3300 1335
rect 3250 1285 3300 1315
rect 3250 1265 3265 1285
rect 3285 1265 3300 1285
rect 3250 1235 3300 1265
rect 3250 1215 3265 1235
rect 3285 1215 3300 1235
rect 3250 1185 3300 1215
rect 3250 1165 3265 1185
rect 3285 1165 3300 1185
rect 3250 1135 3300 1165
rect 3250 1115 3265 1135
rect 3285 1115 3300 1135
rect 3250 1085 3300 1115
rect 3250 1065 3265 1085
rect 3285 1065 3300 1085
rect 3250 1035 3300 1065
rect 3250 1015 3265 1035
rect 3285 1015 3300 1035
rect 3250 985 3300 1015
rect 3250 965 3265 985
rect 3285 965 3300 985
rect 3250 935 3300 965
rect 3250 915 3265 935
rect 3285 915 3300 935
rect 3250 900 3300 915
rect 3400 900 3450 1600
rect 3550 1585 3600 1600
rect 3550 1565 3565 1585
rect 3585 1565 3600 1585
rect 3550 1535 3600 1565
rect 3550 1515 3565 1535
rect 3585 1515 3600 1535
rect 3550 1485 3600 1515
rect 3550 1465 3565 1485
rect 3585 1465 3600 1485
rect 3550 1435 3600 1465
rect 3550 1415 3565 1435
rect 3585 1415 3600 1435
rect 3550 1385 3600 1415
rect 3550 1365 3565 1385
rect 3585 1365 3600 1385
rect 3550 1335 3600 1365
rect 3550 1315 3565 1335
rect 3585 1315 3600 1335
rect 3550 1285 3600 1315
rect 3550 1265 3565 1285
rect 3585 1265 3600 1285
rect 3550 1235 3600 1265
rect 3550 1215 3565 1235
rect 3585 1215 3600 1235
rect 3550 1185 3600 1215
rect 3550 1165 3565 1185
rect 3585 1165 3600 1185
rect 3550 1135 3600 1165
rect 3550 1115 3565 1135
rect 3585 1115 3600 1135
rect 3550 1085 3600 1115
rect 3550 1065 3565 1085
rect 3585 1065 3600 1085
rect 3550 1035 3600 1065
rect 3550 1015 3565 1035
rect 3585 1015 3600 1035
rect 3550 985 3600 1015
rect 3550 965 3565 985
rect 3585 965 3600 985
rect 3550 935 3600 965
rect 3550 915 3565 935
rect 3585 915 3600 935
rect 3550 900 3600 915
rect 3700 1585 3750 1600
rect 3700 1565 3715 1585
rect 3735 1565 3750 1585
rect 3700 1535 3750 1565
rect 3700 1515 3715 1535
rect 3735 1515 3750 1535
rect 3700 1485 3750 1515
rect 3700 1465 3715 1485
rect 3735 1465 3750 1485
rect 3700 1435 3750 1465
rect 3700 1415 3715 1435
rect 3735 1415 3750 1435
rect 3700 1385 3750 1415
rect 3700 1365 3715 1385
rect 3735 1365 3750 1385
rect 3700 1335 3750 1365
rect 3700 1315 3715 1335
rect 3735 1315 3750 1335
rect 3700 1285 3750 1315
rect 3700 1265 3715 1285
rect 3735 1265 3750 1285
rect 3700 1235 3750 1265
rect 3700 1215 3715 1235
rect 3735 1215 3750 1235
rect 3700 1185 3750 1215
rect 3700 1165 3715 1185
rect 3735 1165 3750 1185
rect 3700 1135 3750 1165
rect 3700 1115 3715 1135
rect 3735 1115 3750 1135
rect 3700 1085 3750 1115
rect 3700 1065 3715 1085
rect 3735 1065 3750 1085
rect 3700 1035 3750 1065
rect 3700 1015 3715 1035
rect 3735 1015 3750 1035
rect 3700 985 3750 1015
rect 3700 965 3715 985
rect 3735 965 3750 985
rect 3700 935 3750 965
rect 3700 915 3715 935
rect 3735 915 3750 935
rect 3700 900 3750 915
rect 3850 1585 3900 1600
rect 3850 1565 3865 1585
rect 3885 1565 3900 1585
rect 3850 1535 3900 1565
rect 3850 1515 3865 1535
rect 3885 1515 3900 1535
rect 3850 1485 3900 1515
rect 3850 1465 3865 1485
rect 3885 1465 3900 1485
rect 3850 1435 3900 1465
rect 3850 1415 3865 1435
rect 3885 1415 3900 1435
rect 3850 1385 3900 1415
rect 3850 1365 3865 1385
rect 3885 1365 3900 1385
rect 3850 1335 3900 1365
rect 3850 1315 3865 1335
rect 3885 1315 3900 1335
rect 3850 1285 3900 1315
rect 3850 1265 3865 1285
rect 3885 1265 3900 1285
rect 3850 1235 3900 1265
rect 3850 1215 3865 1235
rect 3885 1215 3900 1235
rect 3850 1185 3900 1215
rect 3850 1165 3865 1185
rect 3885 1165 3900 1185
rect 3850 1135 3900 1165
rect 3850 1115 3865 1135
rect 3885 1115 3900 1135
rect 3850 1085 3900 1115
rect 3850 1065 3865 1085
rect 3885 1065 3900 1085
rect 3850 1035 3900 1065
rect 3850 1015 3865 1035
rect 3885 1015 3900 1035
rect 3850 985 3900 1015
rect 3850 965 3865 985
rect 3885 965 3900 985
rect 3850 935 3900 965
rect 3850 915 3865 935
rect 3885 915 3900 935
rect 3850 900 3900 915
rect 4000 1585 4050 1600
rect 4000 1565 4015 1585
rect 4035 1565 4050 1585
rect 4000 1535 4050 1565
rect 4000 1515 4015 1535
rect 4035 1515 4050 1535
rect 4000 1485 4050 1515
rect 4000 1465 4015 1485
rect 4035 1465 4050 1485
rect 4000 1435 4050 1465
rect 4000 1415 4015 1435
rect 4035 1415 4050 1435
rect 4000 1385 4050 1415
rect 4000 1365 4015 1385
rect 4035 1365 4050 1385
rect 4000 1335 4050 1365
rect 4000 1315 4015 1335
rect 4035 1315 4050 1335
rect 4000 1285 4050 1315
rect 4000 1265 4015 1285
rect 4035 1265 4050 1285
rect 4000 1235 4050 1265
rect 4000 1215 4015 1235
rect 4035 1215 4050 1235
rect 4000 1185 4050 1215
rect 4000 1165 4015 1185
rect 4035 1165 4050 1185
rect 4000 1135 4050 1165
rect 4000 1115 4015 1135
rect 4035 1115 4050 1135
rect 4000 1085 4050 1115
rect 4000 1065 4015 1085
rect 4035 1065 4050 1085
rect 4000 1035 4050 1065
rect 4000 1015 4015 1035
rect 4035 1015 4050 1035
rect 4000 985 4050 1015
rect 4000 965 4015 985
rect 4035 965 4050 985
rect 4000 935 4050 965
rect 4000 915 4015 935
rect 4035 915 4050 935
rect 4000 900 4050 915
rect 4150 1585 4200 1600
rect 4150 1565 4165 1585
rect 4185 1565 4200 1585
rect 4150 1535 4200 1565
rect 4150 1515 4165 1535
rect 4185 1515 4200 1535
rect 4150 1485 4200 1515
rect 4150 1465 4165 1485
rect 4185 1465 4200 1485
rect 4150 1435 4200 1465
rect 4150 1415 4165 1435
rect 4185 1415 4200 1435
rect 4150 1385 4200 1415
rect 4150 1365 4165 1385
rect 4185 1365 4200 1385
rect 4150 1335 4200 1365
rect 4150 1315 4165 1335
rect 4185 1315 4200 1335
rect 4150 1285 4200 1315
rect 4150 1265 4165 1285
rect 4185 1265 4200 1285
rect 4150 1235 4200 1265
rect 4150 1215 4165 1235
rect 4185 1215 4200 1235
rect 4150 1185 4200 1215
rect 4150 1165 4165 1185
rect 4185 1165 4200 1185
rect 4150 1135 4200 1165
rect 4150 1115 4165 1135
rect 4185 1115 4200 1135
rect 4150 1085 4200 1115
rect 4150 1065 4165 1085
rect 4185 1065 4200 1085
rect 4150 1035 4200 1065
rect 4150 1015 4165 1035
rect 4185 1015 4200 1035
rect 4150 985 4200 1015
rect 4150 965 4165 985
rect 4185 965 4200 985
rect 4150 935 4200 965
rect 4150 915 4165 935
rect 4185 915 4200 935
rect 4150 900 4200 915
rect 4300 1585 4350 1600
rect 4300 1565 4315 1585
rect 4335 1565 4350 1585
rect 4300 1535 4350 1565
rect 4300 1515 4315 1535
rect 4335 1515 4350 1535
rect 4300 1485 4350 1515
rect 4300 1465 4315 1485
rect 4335 1465 4350 1485
rect 4300 1435 4350 1465
rect 4300 1415 4315 1435
rect 4335 1415 4350 1435
rect 4300 1385 4350 1415
rect 4300 1365 4315 1385
rect 4335 1365 4350 1385
rect 4300 1335 4350 1365
rect 4300 1315 4315 1335
rect 4335 1315 4350 1335
rect 4300 1285 4350 1315
rect 4300 1265 4315 1285
rect 4335 1265 4350 1285
rect 4300 1235 4350 1265
rect 4300 1215 4315 1235
rect 4335 1215 4350 1235
rect 4300 1185 4350 1215
rect 4300 1165 4315 1185
rect 4335 1165 4350 1185
rect 4300 1135 4350 1165
rect 4300 1115 4315 1135
rect 4335 1115 4350 1135
rect 4300 1085 4350 1115
rect 4300 1065 4315 1085
rect 4335 1065 4350 1085
rect 4300 1035 4350 1065
rect 4300 1015 4315 1035
rect 4335 1015 4350 1035
rect 4300 985 4350 1015
rect 4300 965 4315 985
rect 4335 965 4350 985
rect 4300 935 4350 965
rect 4300 915 4315 935
rect 4335 915 4350 935
rect 4300 900 4350 915
rect 4450 1585 4500 1600
rect 4450 1565 4465 1585
rect 4485 1565 4500 1585
rect 4450 1535 4500 1565
rect 4450 1515 4465 1535
rect 4485 1515 4500 1535
rect 4450 1485 4500 1515
rect 4450 1465 4465 1485
rect 4485 1465 4500 1485
rect 4450 1435 4500 1465
rect 4450 1415 4465 1435
rect 4485 1415 4500 1435
rect 4450 1385 4500 1415
rect 4450 1365 4465 1385
rect 4485 1365 4500 1385
rect 4450 1335 4500 1365
rect 4450 1315 4465 1335
rect 4485 1315 4500 1335
rect 4450 1285 4500 1315
rect 4450 1265 4465 1285
rect 4485 1265 4500 1285
rect 4450 1235 4500 1265
rect 4450 1215 4465 1235
rect 4485 1215 4500 1235
rect 4450 1185 4500 1215
rect 4450 1165 4465 1185
rect 4485 1165 4500 1185
rect 4450 1135 4500 1165
rect 4450 1115 4465 1135
rect 4485 1115 4500 1135
rect 4450 1085 4500 1115
rect 4450 1065 4465 1085
rect 4485 1065 4500 1085
rect 4450 1035 4500 1065
rect 4450 1015 4465 1035
rect 4485 1015 4500 1035
rect 4450 985 4500 1015
rect 4450 965 4465 985
rect 4485 965 4500 985
rect 4450 935 4500 965
rect 4450 915 4465 935
rect 4485 915 4500 935
rect 4450 900 4500 915
rect 4600 1585 4650 1600
rect 4600 1565 4615 1585
rect 4635 1565 4650 1585
rect 4600 1535 4650 1565
rect 4600 1515 4615 1535
rect 4635 1515 4650 1535
rect 4600 1485 4650 1515
rect 4600 1465 4615 1485
rect 4635 1465 4650 1485
rect 4600 1435 4650 1465
rect 4600 1415 4615 1435
rect 4635 1415 4650 1435
rect 4600 1385 4650 1415
rect 4600 1365 4615 1385
rect 4635 1365 4650 1385
rect 4600 1335 4650 1365
rect 4600 1315 4615 1335
rect 4635 1315 4650 1335
rect 4600 1285 4650 1315
rect 4600 1265 4615 1285
rect 4635 1265 4650 1285
rect 4600 1235 4650 1265
rect 4600 1215 4615 1235
rect 4635 1215 4650 1235
rect 4600 1185 4650 1215
rect 4600 1165 4615 1185
rect 4635 1165 4650 1185
rect 4600 1135 4650 1165
rect 4600 1115 4615 1135
rect 4635 1115 4650 1135
rect 4600 1085 4650 1115
rect 4600 1065 4615 1085
rect 4635 1065 4650 1085
rect 4600 1035 4650 1065
rect 4600 1015 4615 1035
rect 4635 1015 4650 1035
rect 4600 985 4650 1015
rect 4600 965 4615 985
rect 4635 965 4650 985
rect 4600 935 4650 965
rect 4600 915 4615 935
rect 4635 915 4650 935
rect 4600 900 4650 915
rect 4750 1585 4800 1600
rect 4750 1565 4765 1585
rect 4785 1565 4800 1585
rect 4750 1535 4800 1565
rect 4750 1515 4765 1535
rect 4785 1515 4800 1535
rect 4750 1485 4800 1515
rect 4750 1465 4765 1485
rect 4785 1465 4800 1485
rect 4750 1435 4800 1465
rect 4750 1415 4765 1435
rect 4785 1415 4800 1435
rect 4750 1385 4800 1415
rect 4750 1365 4765 1385
rect 4785 1365 4800 1385
rect 4750 1335 4800 1365
rect 4750 1315 4765 1335
rect 4785 1315 4800 1335
rect 4750 1285 4800 1315
rect 4750 1265 4765 1285
rect 4785 1265 4800 1285
rect 4750 1235 4800 1265
rect 4750 1215 4765 1235
rect 4785 1215 4800 1235
rect 4750 1185 4800 1215
rect 4750 1165 4765 1185
rect 4785 1165 4800 1185
rect 4750 1135 4800 1165
rect 4750 1115 4765 1135
rect 4785 1115 4800 1135
rect 4750 1085 4800 1115
rect 4750 1065 4765 1085
rect 4785 1065 4800 1085
rect 4750 1035 4800 1065
rect 4750 1015 4765 1035
rect 4785 1015 4800 1035
rect 4750 985 4800 1015
rect 4750 965 4765 985
rect 4785 965 4800 985
rect 4750 935 4800 965
rect 4750 915 4765 935
rect 4785 915 4800 935
rect 4750 900 4800 915
rect 4900 900 4950 1600
rect 5050 1585 5100 1600
rect 5050 1565 5065 1585
rect 5085 1565 5100 1585
rect 5050 1535 5100 1565
rect 5050 1515 5065 1535
rect 5085 1515 5100 1535
rect 5050 1485 5100 1515
rect 5050 1465 5065 1485
rect 5085 1465 5100 1485
rect 5050 1435 5100 1465
rect 5050 1415 5065 1435
rect 5085 1415 5100 1435
rect 5050 1385 5100 1415
rect 5050 1365 5065 1385
rect 5085 1365 5100 1385
rect 5050 1335 5100 1365
rect 5050 1315 5065 1335
rect 5085 1315 5100 1335
rect 5050 1285 5100 1315
rect 5050 1265 5065 1285
rect 5085 1265 5100 1285
rect 5050 1235 5100 1265
rect 5050 1215 5065 1235
rect 5085 1215 5100 1235
rect 5050 1185 5100 1215
rect 5050 1165 5065 1185
rect 5085 1165 5100 1185
rect 5050 1135 5100 1165
rect 5050 1115 5065 1135
rect 5085 1115 5100 1135
rect 5050 1085 5100 1115
rect 5050 1065 5065 1085
rect 5085 1065 5100 1085
rect 5050 1035 5100 1065
rect 5050 1015 5065 1035
rect 5085 1015 5100 1035
rect 5050 985 5100 1015
rect 5050 965 5065 985
rect 5085 965 5100 985
rect 5050 935 5100 965
rect 5050 915 5065 935
rect 5085 915 5100 935
rect 5050 900 5100 915
rect 5200 900 5250 1600
rect 5350 1585 5400 1600
rect 5350 1565 5365 1585
rect 5385 1565 5400 1585
rect 5350 1535 5400 1565
rect 5350 1515 5365 1535
rect 5385 1515 5400 1535
rect 5350 1485 5400 1515
rect 5350 1465 5365 1485
rect 5385 1465 5400 1485
rect 5350 1435 5400 1465
rect 5350 1415 5365 1435
rect 5385 1415 5400 1435
rect 5350 1385 5400 1415
rect 5350 1365 5365 1385
rect 5385 1365 5400 1385
rect 5350 1335 5400 1365
rect 5350 1315 5365 1335
rect 5385 1315 5400 1335
rect 5350 1285 5400 1315
rect 5350 1265 5365 1285
rect 5385 1265 5400 1285
rect 5350 1235 5400 1265
rect 5350 1215 5365 1235
rect 5385 1215 5400 1235
rect 5350 1185 5400 1215
rect 5350 1165 5365 1185
rect 5385 1165 5400 1185
rect 5350 1135 5400 1165
rect 5350 1115 5365 1135
rect 5385 1115 5400 1135
rect 5350 1085 5400 1115
rect 5350 1065 5365 1085
rect 5385 1065 5400 1085
rect 5350 1035 5400 1065
rect 5350 1015 5365 1035
rect 5385 1015 5400 1035
rect 5350 985 5400 1015
rect 5350 965 5365 985
rect 5385 965 5400 985
rect 5350 935 5400 965
rect 5350 915 5365 935
rect 5385 915 5400 935
rect 5350 900 5400 915
rect 5500 900 5550 1600
rect 5650 1585 5700 1600
rect 5650 1565 5665 1585
rect 5685 1565 5700 1585
rect 5650 1535 5700 1565
rect 5650 1515 5665 1535
rect 5685 1515 5700 1535
rect 5650 1485 5700 1515
rect 5650 1465 5665 1485
rect 5685 1465 5700 1485
rect 5650 1435 5700 1465
rect 5650 1415 5665 1435
rect 5685 1415 5700 1435
rect 5650 1385 5700 1415
rect 5650 1365 5665 1385
rect 5685 1365 5700 1385
rect 5650 1335 5700 1365
rect 5650 1315 5665 1335
rect 5685 1315 5700 1335
rect 5650 1285 5700 1315
rect 5650 1265 5665 1285
rect 5685 1265 5700 1285
rect 5650 1235 5700 1265
rect 5650 1215 5665 1235
rect 5685 1215 5700 1235
rect 5650 1185 5700 1215
rect 5650 1165 5665 1185
rect 5685 1165 5700 1185
rect 5650 1135 5700 1165
rect 5650 1115 5665 1135
rect 5685 1115 5700 1135
rect 5650 1085 5700 1115
rect 5650 1065 5665 1085
rect 5685 1065 5700 1085
rect 5650 1035 5700 1065
rect 5650 1015 5665 1035
rect 5685 1015 5700 1035
rect 5650 985 5700 1015
rect 5650 965 5665 985
rect 5685 965 5700 985
rect 5650 935 5700 965
rect 5650 915 5665 935
rect 5685 915 5700 935
rect 5650 900 5700 915
rect 5800 900 5850 1600
rect 5950 1585 6000 1600
rect 5950 1565 5965 1585
rect 5985 1565 6000 1585
rect 5950 1535 6000 1565
rect 5950 1515 5965 1535
rect 5985 1515 6000 1535
rect 5950 1485 6000 1515
rect 5950 1465 5965 1485
rect 5985 1465 6000 1485
rect 5950 1435 6000 1465
rect 5950 1415 5965 1435
rect 5985 1415 6000 1435
rect 5950 1385 6000 1415
rect 5950 1365 5965 1385
rect 5985 1365 6000 1385
rect 5950 1335 6000 1365
rect 5950 1315 5965 1335
rect 5985 1315 6000 1335
rect 5950 1285 6000 1315
rect 5950 1265 5965 1285
rect 5985 1265 6000 1285
rect 5950 1235 6000 1265
rect 5950 1215 5965 1235
rect 5985 1215 6000 1235
rect 5950 1185 6000 1215
rect 5950 1165 5965 1185
rect 5985 1165 6000 1185
rect 5950 1135 6000 1165
rect 5950 1115 5965 1135
rect 5985 1115 6000 1135
rect 5950 1085 6000 1115
rect 5950 1065 5965 1085
rect 5985 1065 6000 1085
rect 5950 1035 6000 1065
rect 5950 1015 5965 1035
rect 5985 1015 6000 1035
rect 5950 985 6000 1015
rect 5950 965 5965 985
rect 5985 965 6000 985
rect 5950 935 6000 965
rect 5950 915 5965 935
rect 5985 915 6000 935
rect 5950 900 6000 915
rect 6100 900 6150 1600
rect 6250 1585 6300 1600
rect 6250 1565 6265 1585
rect 6285 1565 6300 1585
rect 6250 1535 6300 1565
rect 6250 1515 6265 1535
rect 6285 1515 6300 1535
rect 6250 1485 6300 1515
rect 6250 1465 6265 1485
rect 6285 1465 6300 1485
rect 6250 1435 6300 1465
rect 6250 1415 6265 1435
rect 6285 1415 6300 1435
rect 6250 1385 6300 1415
rect 6250 1365 6265 1385
rect 6285 1365 6300 1385
rect 6250 1335 6300 1365
rect 6250 1315 6265 1335
rect 6285 1315 6300 1335
rect 6250 1285 6300 1315
rect 6250 1265 6265 1285
rect 6285 1265 6300 1285
rect 6250 1235 6300 1265
rect 6250 1215 6265 1235
rect 6285 1215 6300 1235
rect 6250 1185 6300 1215
rect 6250 1165 6265 1185
rect 6285 1165 6300 1185
rect 6250 1135 6300 1165
rect 6250 1115 6265 1135
rect 6285 1115 6300 1135
rect 6250 1085 6300 1115
rect 6250 1065 6265 1085
rect 6285 1065 6300 1085
rect 6250 1035 6300 1065
rect 6250 1015 6265 1035
rect 6285 1015 6300 1035
rect 6250 985 6300 1015
rect 6250 965 6265 985
rect 6285 965 6300 985
rect 6250 935 6300 965
rect 6250 915 6265 935
rect 6285 915 6300 935
rect 6250 900 6300 915
rect 6400 900 6450 1600
rect 6550 1585 6600 1600
rect 6550 1565 6565 1585
rect 6585 1565 6600 1585
rect 6550 1535 6600 1565
rect 6550 1515 6565 1535
rect 6585 1515 6600 1535
rect 6550 1485 6600 1515
rect 6550 1465 6565 1485
rect 6585 1465 6600 1485
rect 6550 1435 6600 1465
rect 6550 1415 6565 1435
rect 6585 1415 6600 1435
rect 6550 1385 6600 1415
rect 6550 1365 6565 1385
rect 6585 1365 6600 1385
rect 6550 1335 6600 1365
rect 6550 1315 6565 1335
rect 6585 1315 6600 1335
rect 6550 1285 6600 1315
rect 6550 1265 6565 1285
rect 6585 1265 6600 1285
rect 6550 1235 6600 1265
rect 6550 1215 6565 1235
rect 6585 1215 6600 1235
rect 6550 1185 6600 1215
rect 6550 1165 6565 1185
rect 6585 1165 6600 1185
rect 6550 1135 6600 1165
rect 6550 1115 6565 1135
rect 6585 1115 6600 1135
rect 6550 1085 6600 1115
rect 6550 1065 6565 1085
rect 6585 1065 6600 1085
rect 6550 1035 6600 1065
rect 6550 1015 6565 1035
rect 6585 1015 6600 1035
rect 6550 985 6600 1015
rect 6550 965 6565 985
rect 6585 965 6600 985
rect 6550 935 6600 965
rect 6550 915 6565 935
rect 6585 915 6600 935
rect 6550 900 6600 915
rect 6700 900 6750 1600
rect 6850 1585 6900 1600
rect 6850 1565 6865 1585
rect 6885 1565 6900 1585
rect 6850 1535 6900 1565
rect 6850 1515 6865 1535
rect 6885 1515 6900 1535
rect 6850 1485 6900 1515
rect 6850 1465 6865 1485
rect 6885 1465 6900 1485
rect 6850 1435 6900 1465
rect 6850 1415 6865 1435
rect 6885 1415 6900 1435
rect 6850 1385 6900 1415
rect 6850 1365 6865 1385
rect 6885 1365 6900 1385
rect 6850 1335 6900 1365
rect 6850 1315 6865 1335
rect 6885 1315 6900 1335
rect 6850 1285 6900 1315
rect 6850 1265 6865 1285
rect 6885 1265 6900 1285
rect 6850 1235 6900 1265
rect 6850 1215 6865 1235
rect 6885 1215 6900 1235
rect 6850 1185 6900 1215
rect 6850 1165 6865 1185
rect 6885 1165 6900 1185
rect 6850 1135 6900 1165
rect 6850 1115 6865 1135
rect 6885 1115 6900 1135
rect 6850 1085 6900 1115
rect 6850 1065 6865 1085
rect 6885 1065 6900 1085
rect 6850 1035 6900 1065
rect 6850 1015 6865 1035
rect 6885 1015 6900 1035
rect 6850 985 6900 1015
rect 6850 965 6865 985
rect 6885 965 6900 985
rect 6850 935 6900 965
rect 6850 915 6865 935
rect 6885 915 6900 935
rect 6850 900 6900 915
rect 7000 900 7050 1600
rect 7150 1585 7200 1600
rect 7150 1565 7165 1585
rect 7185 1565 7200 1585
rect 7150 1535 7200 1565
rect 7150 1515 7165 1535
rect 7185 1515 7200 1535
rect 7150 1485 7200 1515
rect 7150 1465 7165 1485
rect 7185 1465 7200 1485
rect 7150 1435 7200 1465
rect 7150 1415 7165 1435
rect 7185 1415 7200 1435
rect 7150 1385 7200 1415
rect 7150 1365 7165 1385
rect 7185 1365 7200 1385
rect 7150 1335 7200 1365
rect 7150 1315 7165 1335
rect 7185 1315 7200 1335
rect 7150 1285 7200 1315
rect 7150 1265 7165 1285
rect 7185 1265 7200 1285
rect 7150 1235 7200 1265
rect 7150 1215 7165 1235
rect 7185 1215 7200 1235
rect 7150 1185 7200 1215
rect 7150 1165 7165 1185
rect 7185 1165 7200 1185
rect 7150 1135 7200 1165
rect 7150 1115 7165 1135
rect 7185 1115 7200 1135
rect 7150 1085 7200 1115
rect 7150 1065 7165 1085
rect 7185 1065 7200 1085
rect 7150 1035 7200 1065
rect 7150 1015 7165 1035
rect 7185 1015 7200 1035
rect 7150 985 7200 1015
rect 7150 965 7165 985
rect 7185 965 7200 985
rect 7150 935 7200 965
rect 7150 915 7165 935
rect 7185 915 7200 935
rect 7150 900 7200 915
rect 7300 900 7350 1600
rect 7450 900 7500 1600
rect 7600 900 7650 1600
rect 7750 900 7800 1600
rect 7900 900 7950 1600
rect 8050 900 8100 1600
rect 8200 900 8250 1600
rect 8350 1585 8400 1600
rect 8350 1565 8365 1585
rect 8385 1565 8400 1585
rect 8350 1535 8400 1565
rect 8350 1515 8365 1535
rect 8385 1515 8400 1535
rect 8350 1485 8400 1515
rect 8350 1465 8365 1485
rect 8385 1465 8400 1485
rect 8350 1435 8400 1465
rect 8350 1415 8365 1435
rect 8385 1415 8400 1435
rect 8350 1385 8400 1415
rect 8350 1365 8365 1385
rect 8385 1365 8400 1385
rect 8350 1335 8400 1365
rect 8350 1315 8365 1335
rect 8385 1315 8400 1335
rect 8350 1285 8400 1315
rect 8350 1265 8365 1285
rect 8385 1265 8400 1285
rect 8350 1235 8400 1265
rect 8350 1215 8365 1235
rect 8385 1215 8400 1235
rect 8350 1185 8400 1215
rect 8350 1165 8365 1185
rect 8385 1165 8400 1185
rect 8350 1135 8400 1165
rect 8350 1115 8365 1135
rect 8385 1115 8400 1135
rect 8350 1085 8400 1115
rect 8350 1065 8365 1085
rect 8385 1065 8400 1085
rect 8350 1035 8400 1065
rect 8350 1015 8365 1035
rect 8385 1015 8400 1035
rect 8350 985 8400 1015
rect 8350 965 8365 985
rect 8385 965 8400 985
rect 8350 935 8400 965
rect 8350 915 8365 935
rect 8385 915 8400 935
rect 8350 900 8400 915
rect 8500 900 8550 1600
rect 8650 900 8700 1600
rect 8800 900 8850 1600
rect 8950 900 9000 1600
rect 9100 900 9150 1600
rect 9250 900 9300 1600
rect 9400 900 9450 1600
rect 9550 1585 9600 1600
rect 9550 1565 9565 1585
rect 9585 1565 9600 1585
rect 9550 1535 9600 1565
rect 9550 1515 9565 1535
rect 9585 1515 9600 1535
rect 9550 1485 9600 1515
rect 9550 1465 9565 1485
rect 9585 1465 9600 1485
rect 9550 1435 9600 1465
rect 9550 1415 9565 1435
rect 9585 1415 9600 1435
rect 9550 1385 9600 1415
rect 9550 1365 9565 1385
rect 9585 1365 9600 1385
rect 9550 1335 9600 1365
rect 9550 1315 9565 1335
rect 9585 1315 9600 1335
rect 9550 1285 9600 1315
rect 9550 1265 9565 1285
rect 9585 1265 9600 1285
rect 9550 1235 9600 1265
rect 9550 1215 9565 1235
rect 9585 1215 9600 1235
rect 9550 1185 9600 1215
rect 9550 1165 9565 1185
rect 9585 1165 9600 1185
rect 9550 1135 9600 1165
rect 9550 1115 9565 1135
rect 9585 1115 9600 1135
rect 9550 1085 9600 1115
rect 9550 1065 9565 1085
rect 9585 1065 9600 1085
rect 9550 1035 9600 1065
rect 9550 1015 9565 1035
rect 9585 1015 9600 1035
rect 9550 985 9600 1015
rect 9550 965 9565 985
rect 9585 965 9600 985
rect 9550 935 9600 965
rect 9550 915 9565 935
rect 9585 915 9600 935
rect 9550 900 9600 915
rect 9700 900 9750 1600
rect 9850 900 9900 1600
rect 10000 900 10050 1600
rect 10150 900 10200 1600
rect 10300 900 10350 1600
rect 10450 900 10500 1600
rect 10600 900 10650 1600
rect 10750 1585 10800 1600
rect 10750 1565 10765 1585
rect 10785 1565 10800 1585
rect 10750 1535 10800 1565
rect 10750 1515 10765 1535
rect 10785 1515 10800 1535
rect 10750 1485 10800 1515
rect 10750 1465 10765 1485
rect 10785 1465 10800 1485
rect 10750 1435 10800 1465
rect 10750 1415 10765 1435
rect 10785 1415 10800 1435
rect 10750 1385 10800 1415
rect 10750 1365 10765 1385
rect 10785 1365 10800 1385
rect 10750 1335 10800 1365
rect 10750 1315 10765 1335
rect 10785 1315 10800 1335
rect 10750 1285 10800 1315
rect 10750 1265 10765 1285
rect 10785 1265 10800 1285
rect 10750 1235 10800 1265
rect 10750 1215 10765 1235
rect 10785 1215 10800 1235
rect 10750 1185 10800 1215
rect 10750 1165 10765 1185
rect 10785 1165 10800 1185
rect 10750 1135 10800 1165
rect 10750 1115 10765 1135
rect 10785 1115 10800 1135
rect 10750 1085 10800 1115
rect 10750 1065 10765 1085
rect 10785 1065 10800 1085
rect 10750 1035 10800 1065
rect 10750 1015 10765 1035
rect 10785 1015 10800 1035
rect 10750 985 10800 1015
rect 10750 965 10765 985
rect 10785 965 10800 985
rect 10750 935 10800 965
rect 10750 915 10765 935
rect 10785 915 10800 935
rect 10750 900 10800 915
rect 10900 900 10950 1600
rect 11050 900 11100 1600
rect 11200 900 11250 1600
rect 11350 900 11400 1600
rect 11500 900 11550 1600
rect 11650 900 11700 1600
rect 11800 900 11850 1600
rect 11950 1585 12000 1600
rect 11950 1565 11965 1585
rect 11985 1565 12000 1585
rect 11950 1535 12000 1565
rect 11950 1515 11965 1535
rect 11985 1515 12000 1535
rect 11950 1485 12000 1515
rect 11950 1465 11965 1485
rect 11985 1465 12000 1485
rect 11950 1435 12000 1465
rect 11950 1415 11965 1435
rect 11985 1415 12000 1435
rect 11950 1385 12000 1415
rect 11950 1365 11965 1385
rect 11985 1365 12000 1385
rect 11950 1335 12000 1365
rect 11950 1315 11965 1335
rect 11985 1315 12000 1335
rect 11950 1285 12000 1315
rect 11950 1265 11965 1285
rect 11985 1265 12000 1285
rect 11950 1235 12000 1265
rect 11950 1215 11965 1235
rect 11985 1215 12000 1235
rect 11950 1185 12000 1215
rect 11950 1165 11965 1185
rect 11985 1165 12000 1185
rect 11950 1135 12000 1165
rect 11950 1115 11965 1135
rect 11985 1115 12000 1135
rect 11950 1085 12000 1115
rect 11950 1065 11965 1085
rect 11985 1065 12000 1085
rect 11950 1035 12000 1065
rect 11950 1015 11965 1035
rect 11985 1015 12000 1035
rect 11950 985 12000 1015
rect 11950 965 11965 985
rect 11985 965 12000 985
rect 11950 935 12000 965
rect 11950 915 11965 935
rect 11985 915 12000 935
rect 11950 900 12000 915
rect 12100 900 12150 1600
rect 12250 1585 12300 1600
rect 12250 1565 12265 1585
rect 12285 1565 12300 1585
rect 12250 1535 12300 1565
rect 12250 1515 12265 1535
rect 12285 1515 12300 1535
rect 12250 1485 12300 1515
rect 12250 1465 12265 1485
rect 12285 1465 12300 1485
rect 12250 1435 12300 1465
rect 12250 1415 12265 1435
rect 12285 1415 12300 1435
rect 12250 1385 12300 1415
rect 12250 1365 12265 1385
rect 12285 1365 12300 1385
rect 12250 1335 12300 1365
rect 12250 1315 12265 1335
rect 12285 1315 12300 1335
rect 12250 1285 12300 1315
rect 12250 1265 12265 1285
rect 12285 1265 12300 1285
rect 12250 1235 12300 1265
rect 12250 1215 12265 1235
rect 12285 1215 12300 1235
rect 12250 1185 12300 1215
rect 12250 1165 12265 1185
rect 12285 1165 12300 1185
rect 12250 1135 12300 1165
rect 12250 1115 12265 1135
rect 12285 1115 12300 1135
rect 12250 1085 12300 1115
rect 12250 1065 12265 1085
rect 12285 1065 12300 1085
rect 12250 1035 12300 1065
rect 12250 1015 12265 1035
rect 12285 1015 12300 1035
rect 12250 985 12300 1015
rect 12250 965 12265 985
rect 12285 965 12300 985
rect 12250 935 12300 965
rect 12250 915 12265 935
rect 12285 915 12300 935
rect 12250 900 12300 915
rect 12400 900 12450 1600
rect 12550 1585 12600 1600
rect 12550 1565 12565 1585
rect 12585 1565 12600 1585
rect 12550 1535 12600 1565
rect 12550 1515 12565 1535
rect 12585 1515 12600 1535
rect 12550 1485 12600 1515
rect 12550 1465 12565 1485
rect 12585 1465 12600 1485
rect 12550 1435 12600 1465
rect 12550 1415 12565 1435
rect 12585 1415 12600 1435
rect 12550 1385 12600 1415
rect 12550 1365 12565 1385
rect 12585 1365 12600 1385
rect 12550 1335 12600 1365
rect 12550 1315 12565 1335
rect 12585 1315 12600 1335
rect 12550 1285 12600 1315
rect 12550 1265 12565 1285
rect 12585 1265 12600 1285
rect 12550 1235 12600 1265
rect 12550 1215 12565 1235
rect 12585 1215 12600 1235
rect 12550 1185 12600 1215
rect 12550 1165 12565 1185
rect 12585 1165 12600 1185
rect 12550 1135 12600 1165
rect 12550 1115 12565 1135
rect 12585 1115 12600 1135
rect 12550 1085 12600 1115
rect 12550 1065 12565 1085
rect 12585 1065 12600 1085
rect 12550 1035 12600 1065
rect 12550 1015 12565 1035
rect 12585 1015 12600 1035
rect 12550 985 12600 1015
rect 12550 965 12565 985
rect 12585 965 12600 985
rect 12550 935 12600 965
rect 12550 915 12565 935
rect 12585 915 12600 935
rect 12550 900 12600 915
rect 12700 900 12750 1600
rect 12850 1585 12900 1600
rect 12850 1565 12865 1585
rect 12885 1565 12900 1585
rect 12850 1535 12900 1565
rect 12850 1515 12865 1535
rect 12885 1515 12900 1535
rect 12850 1485 12900 1515
rect 12850 1465 12865 1485
rect 12885 1465 12900 1485
rect 12850 1435 12900 1465
rect 12850 1415 12865 1435
rect 12885 1415 12900 1435
rect 12850 1385 12900 1415
rect 12850 1365 12865 1385
rect 12885 1365 12900 1385
rect 12850 1335 12900 1365
rect 12850 1315 12865 1335
rect 12885 1315 12900 1335
rect 12850 1285 12900 1315
rect 12850 1265 12865 1285
rect 12885 1265 12900 1285
rect 12850 1235 12900 1265
rect 12850 1215 12865 1235
rect 12885 1215 12900 1235
rect 12850 1185 12900 1215
rect 12850 1165 12865 1185
rect 12885 1165 12900 1185
rect 12850 1135 12900 1165
rect 12850 1115 12865 1135
rect 12885 1115 12900 1135
rect 12850 1085 12900 1115
rect 12850 1065 12865 1085
rect 12885 1065 12900 1085
rect 12850 1035 12900 1065
rect 12850 1015 12865 1035
rect 12885 1015 12900 1035
rect 12850 985 12900 1015
rect 12850 965 12865 985
rect 12885 965 12900 985
rect 12850 935 12900 965
rect 12850 915 12865 935
rect 12885 915 12900 935
rect 12850 900 12900 915
rect 13000 900 13050 1600
rect 13150 1585 13200 1600
rect 13150 1565 13165 1585
rect 13185 1565 13200 1585
rect 13150 1535 13200 1565
rect 13150 1515 13165 1535
rect 13185 1515 13200 1535
rect 13150 1485 13200 1515
rect 13150 1465 13165 1485
rect 13185 1465 13200 1485
rect 13150 1435 13200 1465
rect 13150 1415 13165 1435
rect 13185 1415 13200 1435
rect 13150 1385 13200 1415
rect 13150 1365 13165 1385
rect 13185 1365 13200 1385
rect 13150 1335 13200 1365
rect 13150 1315 13165 1335
rect 13185 1315 13200 1335
rect 13150 1285 13200 1315
rect 13150 1265 13165 1285
rect 13185 1265 13200 1285
rect 13150 1235 13200 1265
rect 13150 1215 13165 1235
rect 13185 1215 13200 1235
rect 13150 1185 13200 1215
rect 13150 1165 13165 1185
rect 13185 1165 13200 1185
rect 13150 1135 13200 1165
rect 13150 1115 13165 1135
rect 13185 1115 13200 1135
rect 13150 1085 13200 1115
rect 13150 1065 13165 1085
rect 13185 1065 13200 1085
rect 13150 1035 13200 1065
rect 13150 1015 13165 1035
rect 13185 1015 13200 1035
rect 13150 985 13200 1015
rect 13150 965 13165 985
rect 13185 965 13200 985
rect 13150 935 13200 965
rect 13150 915 13165 935
rect 13185 915 13200 935
rect 13150 900 13200 915
rect 13300 900 13350 1600
rect 13450 1585 13500 1600
rect 13450 1565 13465 1585
rect 13485 1565 13500 1585
rect 13450 1535 13500 1565
rect 13450 1515 13465 1535
rect 13485 1515 13500 1535
rect 13450 1485 13500 1515
rect 13450 1465 13465 1485
rect 13485 1465 13500 1485
rect 13450 1435 13500 1465
rect 13450 1415 13465 1435
rect 13485 1415 13500 1435
rect 13450 1385 13500 1415
rect 13450 1365 13465 1385
rect 13485 1365 13500 1385
rect 13450 1335 13500 1365
rect 13450 1315 13465 1335
rect 13485 1315 13500 1335
rect 13450 1285 13500 1315
rect 13450 1265 13465 1285
rect 13485 1265 13500 1285
rect 13450 1235 13500 1265
rect 13450 1215 13465 1235
rect 13485 1215 13500 1235
rect 13450 1185 13500 1215
rect 13450 1165 13465 1185
rect 13485 1165 13500 1185
rect 13450 1135 13500 1165
rect 13450 1115 13465 1135
rect 13485 1115 13500 1135
rect 13450 1085 13500 1115
rect 13450 1065 13465 1085
rect 13485 1065 13500 1085
rect 13450 1035 13500 1065
rect 13450 1015 13465 1035
rect 13485 1015 13500 1035
rect 13450 985 13500 1015
rect 13450 965 13465 985
rect 13485 965 13500 985
rect 13450 935 13500 965
rect 13450 915 13465 935
rect 13485 915 13500 935
rect 13450 900 13500 915
rect 13600 900 13650 1600
rect 13750 1585 13800 1600
rect 13750 1565 13765 1585
rect 13785 1565 13800 1585
rect 13750 1535 13800 1565
rect 13750 1515 13765 1535
rect 13785 1515 13800 1535
rect 13750 1485 13800 1515
rect 13750 1465 13765 1485
rect 13785 1465 13800 1485
rect 13750 1435 13800 1465
rect 13750 1415 13765 1435
rect 13785 1415 13800 1435
rect 13750 1385 13800 1415
rect 13750 1365 13765 1385
rect 13785 1365 13800 1385
rect 13750 1335 13800 1365
rect 13750 1315 13765 1335
rect 13785 1315 13800 1335
rect 13750 1285 13800 1315
rect 13750 1265 13765 1285
rect 13785 1265 13800 1285
rect 13750 1235 13800 1265
rect 13750 1215 13765 1235
rect 13785 1215 13800 1235
rect 13750 1185 13800 1215
rect 13750 1165 13765 1185
rect 13785 1165 13800 1185
rect 13750 1135 13800 1165
rect 13750 1115 13765 1135
rect 13785 1115 13800 1135
rect 13750 1085 13800 1115
rect 13750 1065 13765 1085
rect 13785 1065 13800 1085
rect 13750 1035 13800 1065
rect 13750 1015 13765 1035
rect 13785 1015 13800 1035
rect 13750 985 13800 1015
rect 13750 965 13765 985
rect 13785 965 13800 985
rect 13750 935 13800 965
rect 13750 915 13765 935
rect 13785 915 13800 935
rect 13750 900 13800 915
rect 13900 900 13950 1600
rect 14050 1585 14100 1600
rect 14050 1565 14065 1585
rect 14085 1565 14100 1585
rect 14050 1535 14100 1565
rect 14050 1515 14065 1535
rect 14085 1515 14100 1535
rect 14050 1485 14100 1515
rect 14050 1465 14065 1485
rect 14085 1465 14100 1485
rect 14050 1435 14100 1465
rect 14050 1415 14065 1435
rect 14085 1415 14100 1435
rect 14050 1385 14100 1415
rect 14050 1365 14065 1385
rect 14085 1365 14100 1385
rect 14050 1335 14100 1365
rect 14050 1315 14065 1335
rect 14085 1315 14100 1335
rect 14050 1285 14100 1315
rect 14050 1265 14065 1285
rect 14085 1265 14100 1285
rect 14050 1235 14100 1265
rect 14050 1215 14065 1235
rect 14085 1215 14100 1235
rect 14050 1185 14100 1215
rect 14050 1165 14065 1185
rect 14085 1165 14100 1185
rect 14050 1135 14100 1165
rect 14050 1115 14065 1135
rect 14085 1115 14100 1135
rect 14050 1085 14100 1115
rect 14050 1065 14065 1085
rect 14085 1065 14100 1085
rect 14050 1035 14100 1065
rect 14050 1015 14065 1035
rect 14085 1015 14100 1035
rect 14050 985 14100 1015
rect 14050 965 14065 985
rect 14085 965 14100 985
rect 14050 935 14100 965
rect 14050 915 14065 935
rect 14085 915 14100 935
rect 14050 900 14100 915
rect 14200 900 14250 1600
rect 14350 1585 14400 1600
rect 14350 1565 14365 1585
rect 14385 1565 14400 1585
rect 14350 1535 14400 1565
rect 14350 1515 14365 1535
rect 14385 1515 14400 1535
rect 14350 1485 14400 1515
rect 14350 1465 14365 1485
rect 14385 1465 14400 1485
rect 14350 1435 14400 1465
rect 14350 1415 14365 1435
rect 14385 1415 14400 1435
rect 14350 1385 14400 1415
rect 14350 1365 14365 1385
rect 14385 1365 14400 1385
rect 14350 1335 14400 1365
rect 14350 1315 14365 1335
rect 14385 1315 14400 1335
rect 14350 1285 14400 1315
rect 14350 1265 14365 1285
rect 14385 1265 14400 1285
rect 14350 1235 14400 1265
rect 14350 1215 14365 1235
rect 14385 1215 14400 1235
rect 14350 1185 14400 1215
rect 14350 1165 14365 1185
rect 14385 1165 14400 1185
rect 14350 1135 14400 1165
rect 14350 1115 14365 1135
rect 14385 1115 14400 1135
rect 14350 1085 14400 1115
rect 14350 1065 14365 1085
rect 14385 1065 14400 1085
rect 14350 1035 14400 1065
rect 14350 1015 14365 1035
rect 14385 1015 14400 1035
rect 14350 985 14400 1015
rect 14350 965 14365 985
rect 14385 965 14400 985
rect 14350 935 14400 965
rect 14350 915 14365 935
rect 14385 915 14400 935
rect 14350 900 14400 915
rect 14500 900 14550 1600
rect 14650 900 14700 1600
rect 14800 900 14850 1600
rect 14950 900 15000 1600
rect 15100 900 15150 1600
rect 15250 900 15300 1600
rect 15400 900 15450 1600
rect 15550 1585 15600 1600
rect 15550 1565 15565 1585
rect 15585 1565 15600 1585
rect 15550 1535 15600 1565
rect 15550 1515 15565 1535
rect 15585 1515 15600 1535
rect 15550 1485 15600 1515
rect 15550 1465 15565 1485
rect 15585 1465 15600 1485
rect 15550 1435 15600 1465
rect 15550 1415 15565 1435
rect 15585 1415 15600 1435
rect 15550 1385 15600 1415
rect 15550 1365 15565 1385
rect 15585 1365 15600 1385
rect 15550 1335 15600 1365
rect 15550 1315 15565 1335
rect 15585 1315 15600 1335
rect 15550 1285 15600 1315
rect 15550 1265 15565 1285
rect 15585 1265 15600 1285
rect 15550 1235 15600 1265
rect 15550 1215 15565 1235
rect 15585 1215 15600 1235
rect 15550 1185 15600 1215
rect 15550 1165 15565 1185
rect 15585 1165 15600 1185
rect 15550 1135 15600 1165
rect 15550 1115 15565 1135
rect 15585 1115 15600 1135
rect 15550 1085 15600 1115
rect 15550 1065 15565 1085
rect 15585 1065 15600 1085
rect 15550 1035 15600 1065
rect 15550 1015 15565 1035
rect 15585 1015 15600 1035
rect 15550 985 15600 1015
rect 15550 965 15565 985
rect 15585 965 15600 985
rect 15550 935 15600 965
rect 15550 915 15565 935
rect 15585 915 15600 935
rect 15550 900 15600 915
rect 15700 900 15750 1600
rect 15850 900 15900 1600
rect 16000 900 16050 1600
rect 16150 900 16200 1600
rect 16300 900 16350 1600
rect 16450 900 16500 1600
rect 16600 900 16650 1600
rect 16750 1585 16800 1600
rect 16750 1565 16765 1585
rect 16785 1565 16800 1585
rect 16750 1535 16800 1565
rect 16750 1515 16765 1535
rect 16785 1515 16800 1535
rect 16750 1485 16800 1515
rect 16750 1465 16765 1485
rect 16785 1465 16800 1485
rect 16750 1435 16800 1465
rect 16750 1415 16765 1435
rect 16785 1415 16800 1435
rect 16750 1385 16800 1415
rect 16750 1365 16765 1385
rect 16785 1365 16800 1385
rect 16750 1335 16800 1365
rect 16750 1315 16765 1335
rect 16785 1315 16800 1335
rect 16750 1285 16800 1315
rect 16750 1265 16765 1285
rect 16785 1265 16800 1285
rect 16750 1235 16800 1265
rect 16750 1215 16765 1235
rect 16785 1215 16800 1235
rect 16750 1185 16800 1215
rect 16750 1165 16765 1185
rect 16785 1165 16800 1185
rect 16750 1135 16800 1165
rect 16750 1115 16765 1135
rect 16785 1115 16800 1135
rect 16750 1085 16800 1115
rect 16750 1065 16765 1085
rect 16785 1065 16800 1085
rect 16750 1035 16800 1065
rect 16750 1015 16765 1035
rect 16785 1015 16800 1035
rect 16750 985 16800 1015
rect 16750 965 16765 985
rect 16785 965 16800 985
rect 16750 935 16800 965
rect 16750 915 16765 935
rect 16785 915 16800 935
rect 16750 900 16800 915
rect 16900 900 16950 1600
rect 17050 900 17100 1600
rect 17200 900 17250 1600
rect 17350 900 17400 1600
rect 17500 900 17550 1600
rect 17650 900 17700 1600
rect 17800 900 17850 1600
rect 17950 1585 18000 1600
rect 17950 1565 17965 1585
rect 17985 1565 18000 1585
rect 17950 1535 18000 1565
rect 17950 1515 17965 1535
rect 17985 1515 18000 1535
rect 17950 1485 18000 1515
rect 17950 1465 17965 1485
rect 17985 1465 18000 1485
rect 17950 1435 18000 1465
rect 17950 1415 17965 1435
rect 17985 1415 18000 1435
rect 17950 1385 18000 1415
rect 17950 1365 17965 1385
rect 17985 1365 18000 1385
rect 17950 1335 18000 1365
rect 17950 1315 17965 1335
rect 17985 1315 18000 1335
rect 17950 1285 18000 1315
rect 17950 1265 17965 1285
rect 17985 1265 18000 1285
rect 17950 1235 18000 1265
rect 17950 1215 17965 1235
rect 17985 1215 18000 1235
rect 17950 1185 18000 1215
rect 17950 1165 17965 1185
rect 17985 1165 18000 1185
rect 17950 1135 18000 1165
rect 17950 1115 17965 1135
rect 17985 1115 18000 1135
rect 17950 1085 18000 1115
rect 17950 1065 17965 1085
rect 17985 1065 18000 1085
rect 17950 1035 18000 1065
rect 17950 1015 17965 1035
rect 17985 1015 18000 1035
rect 17950 985 18000 1015
rect 17950 965 17965 985
rect 17985 965 18000 985
rect 17950 935 18000 965
rect 17950 915 17965 935
rect 17985 915 18000 935
rect 17950 900 18000 915
rect 18100 900 18150 1600
rect 18250 900 18300 1600
rect 18400 900 18450 1600
rect 18550 900 18600 1600
rect 18700 900 18750 1600
rect 18850 900 18900 1600
rect 19000 900 19050 1600
rect 19150 1585 19200 1600
rect 19150 1565 19165 1585
rect 19185 1565 19200 1585
rect 19150 1535 19200 1565
rect 19150 1515 19165 1535
rect 19185 1515 19200 1535
rect 19150 1485 19200 1515
rect 19150 1465 19165 1485
rect 19185 1465 19200 1485
rect 19150 1435 19200 1465
rect 19150 1415 19165 1435
rect 19185 1415 19200 1435
rect 19150 1385 19200 1415
rect 19150 1365 19165 1385
rect 19185 1365 19200 1385
rect 19150 1335 19200 1365
rect 19150 1315 19165 1335
rect 19185 1315 19200 1335
rect 19150 1285 19200 1315
rect 19150 1265 19165 1285
rect 19185 1265 19200 1285
rect 19150 1235 19200 1265
rect 19150 1215 19165 1235
rect 19185 1215 19200 1235
rect 19150 1185 19200 1215
rect 19150 1165 19165 1185
rect 19185 1165 19200 1185
rect 19150 1135 19200 1165
rect 19150 1115 19165 1135
rect 19185 1115 19200 1135
rect 19150 1085 19200 1115
rect 19150 1065 19165 1085
rect 19185 1065 19200 1085
rect 19150 1035 19200 1065
rect 19150 1015 19165 1035
rect 19185 1015 19200 1035
rect 19150 985 19200 1015
rect 19150 965 19165 985
rect 19185 965 19200 985
rect 19150 935 19200 965
rect 19150 915 19165 935
rect 19185 915 19200 935
rect 19150 900 19200 915
rect 19300 900 19350 1600
rect 19450 900 19500 1600
rect 19600 900 19650 1600
rect 19750 900 19800 1600
rect 19900 900 19950 1600
rect 20050 900 20100 1600
rect 20200 900 20250 1600
rect 20350 1585 20400 1600
rect 20350 1565 20365 1585
rect 20385 1565 20400 1585
rect 20350 1535 20400 1565
rect 20350 1515 20365 1535
rect 20385 1515 20400 1535
rect 20350 1485 20400 1515
rect 20350 1465 20365 1485
rect 20385 1465 20400 1485
rect 20350 1435 20400 1465
rect 20350 1415 20365 1435
rect 20385 1415 20400 1435
rect 20350 1385 20400 1415
rect 20350 1365 20365 1385
rect 20385 1365 20400 1385
rect 20350 1335 20400 1365
rect 20350 1315 20365 1335
rect 20385 1315 20400 1335
rect 20350 1285 20400 1315
rect 20350 1265 20365 1285
rect 20385 1265 20400 1285
rect 20350 1235 20400 1265
rect 20350 1215 20365 1235
rect 20385 1215 20400 1235
rect 20350 1185 20400 1215
rect 20350 1165 20365 1185
rect 20385 1165 20400 1185
rect 20350 1135 20400 1165
rect 20350 1115 20365 1135
rect 20385 1115 20400 1135
rect 20350 1085 20400 1115
rect 20350 1065 20365 1085
rect 20385 1065 20400 1085
rect 20350 1035 20400 1065
rect 20350 1015 20365 1035
rect 20385 1015 20400 1035
rect 20350 985 20400 1015
rect 20350 965 20365 985
rect 20385 965 20400 985
rect 20350 935 20400 965
rect 20350 915 20365 935
rect 20385 915 20400 935
rect 20350 900 20400 915
rect -650 735 -600 750
rect -650 715 -635 735
rect -615 715 -600 735
rect -650 685 -600 715
rect -650 665 -635 685
rect -615 665 -600 685
rect -650 635 -600 665
rect -650 615 -635 635
rect -615 615 -600 635
rect -650 585 -600 615
rect -650 565 -635 585
rect -615 565 -600 585
rect -650 535 -600 565
rect -650 515 -635 535
rect -615 515 -600 535
rect -650 485 -600 515
rect -650 465 -635 485
rect -615 465 -600 485
rect -650 435 -600 465
rect -650 415 -635 435
rect -615 415 -600 435
rect -650 385 -600 415
rect -650 365 -635 385
rect -615 365 -600 385
rect -650 335 -600 365
rect -650 315 -635 335
rect -615 315 -600 335
rect -650 285 -600 315
rect -650 265 -635 285
rect -615 265 -600 285
rect -650 235 -600 265
rect -650 215 -635 235
rect -615 215 -600 235
rect -650 185 -600 215
rect -650 165 -635 185
rect -615 165 -600 185
rect -650 135 -600 165
rect -650 115 -635 135
rect -615 115 -600 135
rect -650 85 -600 115
rect -650 65 -635 85
rect -615 65 -600 85
rect -650 50 -600 65
rect -500 735 -450 750
rect -500 715 -485 735
rect -465 715 -450 735
rect -500 685 -450 715
rect -500 665 -485 685
rect -465 665 -450 685
rect -500 635 -450 665
rect -500 615 -485 635
rect -465 615 -450 635
rect -500 585 -450 615
rect -500 565 -485 585
rect -465 565 -450 585
rect -500 535 -450 565
rect -500 515 -485 535
rect -465 515 -450 535
rect -500 485 -450 515
rect -500 465 -485 485
rect -465 465 -450 485
rect -500 435 -450 465
rect -500 415 -485 435
rect -465 415 -450 435
rect -500 385 -450 415
rect -500 365 -485 385
rect -465 365 -450 385
rect -500 335 -450 365
rect -500 315 -485 335
rect -465 315 -450 335
rect -500 285 -450 315
rect -500 265 -485 285
rect -465 265 -450 285
rect -500 235 -450 265
rect -500 215 -485 235
rect -465 215 -450 235
rect -500 185 -450 215
rect -500 165 -485 185
rect -465 165 -450 185
rect -500 135 -450 165
rect -500 115 -485 135
rect -465 115 -450 135
rect -500 85 -450 115
rect -500 65 -485 85
rect -465 65 -450 85
rect -500 50 -450 65
rect -350 735 -300 750
rect -350 715 -335 735
rect -315 715 -300 735
rect -350 685 -300 715
rect -350 665 -335 685
rect -315 665 -300 685
rect -350 635 -300 665
rect -350 615 -335 635
rect -315 615 -300 635
rect -350 585 -300 615
rect -350 565 -335 585
rect -315 565 -300 585
rect -350 535 -300 565
rect -350 515 -335 535
rect -315 515 -300 535
rect -350 485 -300 515
rect -350 465 -335 485
rect -315 465 -300 485
rect -350 435 -300 465
rect -350 415 -335 435
rect -315 415 -300 435
rect -350 385 -300 415
rect -350 365 -335 385
rect -315 365 -300 385
rect -350 335 -300 365
rect -350 315 -335 335
rect -315 315 -300 335
rect -350 285 -300 315
rect -350 265 -335 285
rect -315 265 -300 285
rect -350 235 -300 265
rect -350 215 -335 235
rect -315 215 -300 235
rect -350 185 -300 215
rect -350 165 -335 185
rect -315 165 -300 185
rect -350 135 -300 165
rect -350 115 -335 135
rect -315 115 -300 135
rect -350 85 -300 115
rect -350 65 -335 85
rect -315 65 -300 85
rect -350 50 -300 65
rect -200 735 -150 750
rect -200 715 -185 735
rect -165 715 -150 735
rect -200 685 -150 715
rect -200 665 -185 685
rect -165 665 -150 685
rect -200 635 -150 665
rect -200 615 -185 635
rect -165 615 -150 635
rect -200 585 -150 615
rect -200 565 -185 585
rect -165 565 -150 585
rect -200 535 -150 565
rect -200 515 -185 535
rect -165 515 -150 535
rect -200 485 -150 515
rect -200 465 -185 485
rect -165 465 -150 485
rect -200 435 -150 465
rect -200 415 -185 435
rect -165 415 -150 435
rect -200 385 -150 415
rect -200 365 -185 385
rect -165 365 -150 385
rect -200 335 -150 365
rect -200 315 -185 335
rect -165 315 -150 335
rect -200 285 -150 315
rect -200 265 -185 285
rect -165 265 -150 285
rect -200 235 -150 265
rect -200 215 -185 235
rect -165 215 -150 235
rect -200 185 -150 215
rect -200 165 -185 185
rect -165 165 -150 185
rect -200 135 -150 165
rect -200 115 -185 135
rect -165 115 -150 135
rect -200 85 -150 115
rect -200 65 -185 85
rect -165 65 -150 85
rect -200 50 -150 65
rect -50 735 0 750
rect -50 715 -35 735
rect -15 715 0 735
rect -50 685 0 715
rect -50 665 -35 685
rect -15 665 0 685
rect -50 635 0 665
rect -50 615 -35 635
rect -15 615 0 635
rect -50 585 0 615
rect -50 565 -35 585
rect -15 565 0 585
rect -50 535 0 565
rect -50 515 -35 535
rect -15 515 0 535
rect -50 485 0 515
rect -50 465 -35 485
rect -15 465 0 485
rect -50 435 0 465
rect -50 415 -35 435
rect -15 415 0 435
rect -50 385 0 415
rect -50 365 -35 385
rect -15 365 0 385
rect -50 335 0 365
rect -50 315 -35 335
rect -15 315 0 335
rect -50 285 0 315
rect -50 265 -35 285
rect -15 265 0 285
rect -50 235 0 265
rect -50 215 -35 235
rect -15 215 0 235
rect -50 185 0 215
rect -50 165 -35 185
rect -15 165 0 185
rect -50 135 0 165
rect -50 115 -35 135
rect -15 115 0 135
rect -50 85 0 115
rect -50 65 -35 85
rect -15 65 0 85
rect -50 50 0 65
rect 100 50 150 750
rect 250 50 300 750
rect 400 50 450 750
rect 550 50 600 750
rect 700 50 750 750
rect 850 50 900 750
rect 1000 50 1050 750
rect 1150 735 1200 750
rect 1150 715 1165 735
rect 1185 715 1200 735
rect 1150 685 1200 715
rect 1150 665 1165 685
rect 1185 665 1200 685
rect 1150 635 1200 665
rect 1150 615 1165 635
rect 1185 615 1200 635
rect 1150 585 1200 615
rect 1150 565 1165 585
rect 1185 565 1200 585
rect 1150 535 1200 565
rect 1150 515 1165 535
rect 1185 515 1200 535
rect 1150 485 1200 515
rect 1150 465 1165 485
rect 1185 465 1200 485
rect 1150 435 1200 465
rect 1150 415 1165 435
rect 1185 415 1200 435
rect 1150 385 1200 415
rect 1150 365 1165 385
rect 1185 365 1200 385
rect 1150 335 1200 365
rect 1150 315 1165 335
rect 1185 315 1200 335
rect 1150 285 1200 315
rect 1150 265 1165 285
rect 1185 265 1200 285
rect 1150 235 1200 265
rect 1150 215 1165 235
rect 1185 215 1200 235
rect 1150 185 1200 215
rect 1150 165 1165 185
rect 1185 165 1200 185
rect 1150 135 1200 165
rect 1150 115 1165 135
rect 1185 115 1200 135
rect 1150 85 1200 115
rect 1150 65 1165 85
rect 1185 65 1200 85
rect 1150 50 1200 65
rect 1300 50 1350 750
rect 1450 735 1500 750
rect 1450 715 1465 735
rect 1485 715 1500 735
rect 1450 685 1500 715
rect 1450 665 1465 685
rect 1485 665 1500 685
rect 1450 635 1500 665
rect 1450 615 1465 635
rect 1485 615 1500 635
rect 1450 585 1500 615
rect 1450 565 1465 585
rect 1485 565 1500 585
rect 1450 535 1500 565
rect 1450 515 1465 535
rect 1485 515 1500 535
rect 1450 485 1500 515
rect 1450 465 1465 485
rect 1485 465 1500 485
rect 1450 435 1500 465
rect 1450 415 1465 435
rect 1485 415 1500 435
rect 1450 385 1500 415
rect 1450 365 1465 385
rect 1485 365 1500 385
rect 1450 335 1500 365
rect 1450 315 1465 335
rect 1485 315 1500 335
rect 1450 285 1500 315
rect 1450 265 1465 285
rect 1485 265 1500 285
rect 1450 235 1500 265
rect 1450 215 1465 235
rect 1485 215 1500 235
rect 1450 185 1500 215
rect 1450 165 1465 185
rect 1485 165 1500 185
rect 1450 135 1500 165
rect 1450 115 1465 135
rect 1485 115 1500 135
rect 1450 85 1500 115
rect 1450 65 1465 85
rect 1485 65 1500 85
rect 1450 50 1500 65
rect 1600 50 1650 750
rect 1750 735 1800 750
rect 1750 715 1765 735
rect 1785 715 1800 735
rect 1750 685 1800 715
rect 1750 665 1765 685
rect 1785 665 1800 685
rect 1750 635 1800 665
rect 1750 615 1765 635
rect 1785 615 1800 635
rect 1750 585 1800 615
rect 1750 565 1765 585
rect 1785 565 1800 585
rect 1750 535 1800 565
rect 1750 515 1765 535
rect 1785 515 1800 535
rect 1750 485 1800 515
rect 1750 465 1765 485
rect 1785 465 1800 485
rect 1750 435 1800 465
rect 1750 415 1765 435
rect 1785 415 1800 435
rect 1750 385 1800 415
rect 1750 365 1765 385
rect 1785 365 1800 385
rect 1750 335 1800 365
rect 1750 315 1765 335
rect 1785 315 1800 335
rect 1750 285 1800 315
rect 1750 265 1765 285
rect 1785 265 1800 285
rect 1750 235 1800 265
rect 1750 215 1765 235
rect 1785 215 1800 235
rect 1750 185 1800 215
rect 1750 165 1765 185
rect 1785 165 1800 185
rect 1750 135 1800 165
rect 1750 115 1765 135
rect 1785 115 1800 135
rect 1750 85 1800 115
rect 1750 65 1765 85
rect 1785 65 1800 85
rect 1750 50 1800 65
rect 1900 50 1950 750
rect 2050 735 2100 750
rect 2050 715 2065 735
rect 2085 715 2100 735
rect 2050 685 2100 715
rect 2050 665 2065 685
rect 2085 665 2100 685
rect 2050 635 2100 665
rect 2050 615 2065 635
rect 2085 615 2100 635
rect 2050 585 2100 615
rect 2050 565 2065 585
rect 2085 565 2100 585
rect 2050 535 2100 565
rect 2050 515 2065 535
rect 2085 515 2100 535
rect 2050 485 2100 515
rect 2050 465 2065 485
rect 2085 465 2100 485
rect 2050 435 2100 465
rect 2050 415 2065 435
rect 2085 415 2100 435
rect 2050 385 2100 415
rect 2050 365 2065 385
rect 2085 365 2100 385
rect 2050 335 2100 365
rect 2050 315 2065 335
rect 2085 315 2100 335
rect 2050 285 2100 315
rect 2050 265 2065 285
rect 2085 265 2100 285
rect 2050 235 2100 265
rect 2050 215 2065 235
rect 2085 215 2100 235
rect 2050 185 2100 215
rect 2050 165 2065 185
rect 2085 165 2100 185
rect 2050 135 2100 165
rect 2050 115 2065 135
rect 2085 115 2100 135
rect 2050 85 2100 115
rect 2050 65 2065 85
rect 2085 65 2100 85
rect 2050 50 2100 65
rect 2200 50 2250 750
rect 2350 735 2400 750
rect 2350 715 2365 735
rect 2385 715 2400 735
rect 2350 685 2400 715
rect 2350 665 2365 685
rect 2385 665 2400 685
rect 2350 635 2400 665
rect 2350 615 2365 635
rect 2385 615 2400 635
rect 2350 585 2400 615
rect 2350 565 2365 585
rect 2385 565 2400 585
rect 2350 535 2400 565
rect 2350 515 2365 535
rect 2385 515 2400 535
rect 2350 485 2400 515
rect 2350 465 2365 485
rect 2385 465 2400 485
rect 2350 435 2400 465
rect 2350 415 2365 435
rect 2385 415 2400 435
rect 2350 385 2400 415
rect 2350 365 2365 385
rect 2385 365 2400 385
rect 2350 335 2400 365
rect 2350 315 2365 335
rect 2385 315 2400 335
rect 2350 285 2400 315
rect 2350 265 2365 285
rect 2385 265 2400 285
rect 2350 235 2400 265
rect 2350 215 2365 235
rect 2385 215 2400 235
rect 2350 185 2400 215
rect 2350 165 2365 185
rect 2385 165 2400 185
rect 2350 135 2400 165
rect 2350 115 2365 135
rect 2385 115 2400 135
rect 2350 85 2400 115
rect 2350 65 2365 85
rect 2385 65 2400 85
rect 2350 50 2400 65
rect 2500 50 2550 750
rect 2650 735 2700 750
rect 2650 715 2665 735
rect 2685 715 2700 735
rect 2650 685 2700 715
rect 2650 665 2665 685
rect 2685 665 2700 685
rect 2650 635 2700 665
rect 2650 615 2665 635
rect 2685 615 2700 635
rect 2650 585 2700 615
rect 2650 565 2665 585
rect 2685 565 2700 585
rect 2650 535 2700 565
rect 2650 515 2665 535
rect 2685 515 2700 535
rect 2650 485 2700 515
rect 2650 465 2665 485
rect 2685 465 2700 485
rect 2650 435 2700 465
rect 2650 415 2665 435
rect 2685 415 2700 435
rect 2650 385 2700 415
rect 2650 365 2665 385
rect 2685 365 2700 385
rect 2650 335 2700 365
rect 2650 315 2665 335
rect 2685 315 2700 335
rect 2650 285 2700 315
rect 2650 265 2665 285
rect 2685 265 2700 285
rect 2650 235 2700 265
rect 2650 215 2665 235
rect 2685 215 2700 235
rect 2650 185 2700 215
rect 2650 165 2665 185
rect 2685 165 2700 185
rect 2650 135 2700 165
rect 2650 115 2665 135
rect 2685 115 2700 135
rect 2650 85 2700 115
rect 2650 65 2665 85
rect 2685 65 2700 85
rect 2650 50 2700 65
rect 2800 50 2850 750
rect 2950 735 3000 750
rect 2950 715 2965 735
rect 2985 715 3000 735
rect 2950 685 3000 715
rect 2950 665 2965 685
rect 2985 665 3000 685
rect 2950 635 3000 665
rect 2950 615 2965 635
rect 2985 615 3000 635
rect 2950 585 3000 615
rect 2950 565 2965 585
rect 2985 565 3000 585
rect 2950 535 3000 565
rect 2950 515 2965 535
rect 2985 515 3000 535
rect 2950 485 3000 515
rect 2950 465 2965 485
rect 2985 465 3000 485
rect 2950 435 3000 465
rect 2950 415 2965 435
rect 2985 415 3000 435
rect 2950 385 3000 415
rect 2950 365 2965 385
rect 2985 365 3000 385
rect 2950 335 3000 365
rect 2950 315 2965 335
rect 2985 315 3000 335
rect 2950 285 3000 315
rect 2950 265 2965 285
rect 2985 265 3000 285
rect 2950 235 3000 265
rect 2950 215 2965 235
rect 2985 215 3000 235
rect 2950 185 3000 215
rect 2950 165 2965 185
rect 2985 165 3000 185
rect 2950 135 3000 165
rect 2950 115 2965 135
rect 2985 115 3000 135
rect 2950 85 3000 115
rect 2950 65 2965 85
rect 2985 65 3000 85
rect 2950 50 3000 65
rect 3100 50 3150 750
rect 3250 735 3300 750
rect 3250 715 3265 735
rect 3285 715 3300 735
rect 3250 685 3300 715
rect 3250 665 3265 685
rect 3285 665 3300 685
rect 3250 635 3300 665
rect 3250 615 3265 635
rect 3285 615 3300 635
rect 3250 585 3300 615
rect 3250 565 3265 585
rect 3285 565 3300 585
rect 3250 535 3300 565
rect 3250 515 3265 535
rect 3285 515 3300 535
rect 3250 485 3300 515
rect 3250 465 3265 485
rect 3285 465 3300 485
rect 3250 435 3300 465
rect 3250 415 3265 435
rect 3285 415 3300 435
rect 3250 385 3300 415
rect 3250 365 3265 385
rect 3285 365 3300 385
rect 3250 335 3300 365
rect 3250 315 3265 335
rect 3285 315 3300 335
rect 3250 285 3300 315
rect 3250 265 3265 285
rect 3285 265 3300 285
rect 3250 235 3300 265
rect 3250 215 3265 235
rect 3285 215 3300 235
rect 3250 185 3300 215
rect 3250 165 3265 185
rect 3285 165 3300 185
rect 3250 135 3300 165
rect 3250 115 3265 135
rect 3285 115 3300 135
rect 3250 85 3300 115
rect 3250 65 3265 85
rect 3285 65 3300 85
rect 3250 50 3300 65
rect 3400 50 3450 750
rect 3550 735 3600 750
rect 3550 715 3565 735
rect 3585 715 3600 735
rect 3550 685 3600 715
rect 3550 665 3565 685
rect 3585 665 3600 685
rect 3550 635 3600 665
rect 3550 615 3565 635
rect 3585 615 3600 635
rect 3550 585 3600 615
rect 3550 565 3565 585
rect 3585 565 3600 585
rect 3550 535 3600 565
rect 3550 515 3565 535
rect 3585 515 3600 535
rect 3550 485 3600 515
rect 3550 465 3565 485
rect 3585 465 3600 485
rect 3550 435 3600 465
rect 3550 415 3565 435
rect 3585 415 3600 435
rect 3550 385 3600 415
rect 3550 365 3565 385
rect 3585 365 3600 385
rect 3550 335 3600 365
rect 3550 315 3565 335
rect 3585 315 3600 335
rect 3550 285 3600 315
rect 3550 265 3565 285
rect 3585 265 3600 285
rect 3550 235 3600 265
rect 3550 215 3565 235
rect 3585 215 3600 235
rect 3550 185 3600 215
rect 3550 165 3565 185
rect 3585 165 3600 185
rect 3550 135 3600 165
rect 3550 115 3565 135
rect 3585 115 3600 135
rect 3550 85 3600 115
rect 3550 65 3565 85
rect 3585 65 3600 85
rect 3550 50 3600 65
rect 3700 735 3750 750
rect 3700 715 3715 735
rect 3735 715 3750 735
rect 3700 685 3750 715
rect 3700 665 3715 685
rect 3735 665 3750 685
rect 3700 635 3750 665
rect 3700 615 3715 635
rect 3735 615 3750 635
rect 3700 585 3750 615
rect 3700 565 3715 585
rect 3735 565 3750 585
rect 3700 535 3750 565
rect 3700 515 3715 535
rect 3735 515 3750 535
rect 3700 485 3750 515
rect 3700 465 3715 485
rect 3735 465 3750 485
rect 3700 435 3750 465
rect 3700 415 3715 435
rect 3735 415 3750 435
rect 3700 385 3750 415
rect 3700 365 3715 385
rect 3735 365 3750 385
rect 3700 335 3750 365
rect 3700 315 3715 335
rect 3735 315 3750 335
rect 3700 285 3750 315
rect 3700 265 3715 285
rect 3735 265 3750 285
rect 3700 235 3750 265
rect 3700 215 3715 235
rect 3735 215 3750 235
rect 3700 185 3750 215
rect 3700 165 3715 185
rect 3735 165 3750 185
rect 3700 135 3750 165
rect 3700 115 3715 135
rect 3735 115 3750 135
rect 3700 85 3750 115
rect 3700 65 3715 85
rect 3735 65 3750 85
rect 3700 50 3750 65
rect 3850 735 3900 750
rect 3850 715 3865 735
rect 3885 715 3900 735
rect 3850 685 3900 715
rect 3850 665 3865 685
rect 3885 665 3900 685
rect 3850 635 3900 665
rect 3850 615 3865 635
rect 3885 615 3900 635
rect 3850 585 3900 615
rect 3850 565 3865 585
rect 3885 565 3900 585
rect 3850 535 3900 565
rect 3850 515 3865 535
rect 3885 515 3900 535
rect 3850 485 3900 515
rect 3850 465 3865 485
rect 3885 465 3900 485
rect 3850 435 3900 465
rect 3850 415 3865 435
rect 3885 415 3900 435
rect 3850 385 3900 415
rect 3850 365 3865 385
rect 3885 365 3900 385
rect 3850 335 3900 365
rect 3850 315 3865 335
rect 3885 315 3900 335
rect 3850 285 3900 315
rect 3850 265 3865 285
rect 3885 265 3900 285
rect 3850 235 3900 265
rect 3850 215 3865 235
rect 3885 215 3900 235
rect 3850 185 3900 215
rect 3850 165 3865 185
rect 3885 165 3900 185
rect 3850 135 3900 165
rect 3850 115 3865 135
rect 3885 115 3900 135
rect 3850 85 3900 115
rect 3850 65 3865 85
rect 3885 65 3900 85
rect 3850 50 3900 65
rect 4000 735 4050 750
rect 4000 715 4015 735
rect 4035 715 4050 735
rect 4000 685 4050 715
rect 4000 665 4015 685
rect 4035 665 4050 685
rect 4000 635 4050 665
rect 4000 615 4015 635
rect 4035 615 4050 635
rect 4000 585 4050 615
rect 4000 565 4015 585
rect 4035 565 4050 585
rect 4000 535 4050 565
rect 4000 515 4015 535
rect 4035 515 4050 535
rect 4000 485 4050 515
rect 4000 465 4015 485
rect 4035 465 4050 485
rect 4000 435 4050 465
rect 4000 415 4015 435
rect 4035 415 4050 435
rect 4000 385 4050 415
rect 4000 365 4015 385
rect 4035 365 4050 385
rect 4000 335 4050 365
rect 4000 315 4015 335
rect 4035 315 4050 335
rect 4000 285 4050 315
rect 4000 265 4015 285
rect 4035 265 4050 285
rect 4000 235 4050 265
rect 4000 215 4015 235
rect 4035 215 4050 235
rect 4000 185 4050 215
rect 4000 165 4015 185
rect 4035 165 4050 185
rect 4000 135 4050 165
rect 4000 115 4015 135
rect 4035 115 4050 135
rect 4000 85 4050 115
rect 4000 65 4015 85
rect 4035 65 4050 85
rect 4000 50 4050 65
rect 4150 735 4200 750
rect 4150 715 4165 735
rect 4185 715 4200 735
rect 4150 685 4200 715
rect 4150 665 4165 685
rect 4185 665 4200 685
rect 4150 635 4200 665
rect 4150 615 4165 635
rect 4185 615 4200 635
rect 4150 585 4200 615
rect 4150 565 4165 585
rect 4185 565 4200 585
rect 4150 535 4200 565
rect 4150 515 4165 535
rect 4185 515 4200 535
rect 4150 485 4200 515
rect 4150 465 4165 485
rect 4185 465 4200 485
rect 4150 435 4200 465
rect 4150 415 4165 435
rect 4185 415 4200 435
rect 4150 385 4200 415
rect 4150 365 4165 385
rect 4185 365 4200 385
rect 4150 335 4200 365
rect 4150 315 4165 335
rect 4185 315 4200 335
rect 4150 285 4200 315
rect 4150 265 4165 285
rect 4185 265 4200 285
rect 4150 235 4200 265
rect 4150 215 4165 235
rect 4185 215 4200 235
rect 4150 185 4200 215
rect 4150 165 4165 185
rect 4185 165 4200 185
rect 4150 135 4200 165
rect 4150 115 4165 135
rect 4185 115 4200 135
rect 4150 85 4200 115
rect 4150 65 4165 85
rect 4185 65 4200 85
rect 4150 50 4200 65
rect 4300 735 4350 750
rect 4300 715 4315 735
rect 4335 715 4350 735
rect 4300 685 4350 715
rect 4300 665 4315 685
rect 4335 665 4350 685
rect 4300 635 4350 665
rect 4300 615 4315 635
rect 4335 615 4350 635
rect 4300 585 4350 615
rect 4300 565 4315 585
rect 4335 565 4350 585
rect 4300 535 4350 565
rect 4300 515 4315 535
rect 4335 515 4350 535
rect 4300 485 4350 515
rect 4300 465 4315 485
rect 4335 465 4350 485
rect 4300 435 4350 465
rect 4300 415 4315 435
rect 4335 415 4350 435
rect 4300 385 4350 415
rect 4300 365 4315 385
rect 4335 365 4350 385
rect 4300 335 4350 365
rect 4300 315 4315 335
rect 4335 315 4350 335
rect 4300 285 4350 315
rect 4300 265 4315 285
rect 4335 265 4350 285
rect 4300 235 4350 265
rect 4300 215 4315 235
rect 4335 215 4350 235
rect 4300 185 4350 215
rect 4300 165 4315 185
rect 4335 165 4350 185
rect 4300 135 4350 165
rect 4300 115 4315 135
rect 4335 115 4350 135
rect 4300 85 4350 115
rect 4300 65 4315 85
rect 4335 65 4350 85
rect 4300 50 4350 65
rect 4450 735 4500 750
rect 4450 715 4465 735
rect 4485 715 4500 735
rect 4450 685 4500 715
rect 4450 665 4465 685
rect 4485 665 4500 685
rect 4450 635 4500 665
rect 4450 615 4465 635
rect 4485 615 4500 635
rect 4450 585 4500 615
rect 4450 565 4465 585
rect 4485 565 4500 585
rect 4450 535 4500 565
rect 4450 515 4465 535
rect 4485 515 4500 535
rect 4450 485 4500 515
rect 4450 465 4465 485
rect 4485 465 4500 485
rect 4450 435 4500 465
rect 4450 415 4465 435
rect 4485 415 4500 435
rect 4450 385 4500 415
rect 4450 365 4465 385
rect 4485 365 4500 385
rect 4450 335 4500 365
rect 4450 315 4465 335
rect 4485 315 4500 335
rect 4450 285 4500 315
rect 4450 265 4465 285
rect 4485 265 4500 285
rect 4450 235 4500 265
rect 4450 215 4465 235
rect 4485 215 4500 235
rect 4450 185 4500 215
rect 4450 165 4465 185
rect 4485 165 4500 185
rect 4450 135 4500 165
rect 4450 115 4465 135
rect 4485 115 4500 135
rect 4450 85 4500 115
rect 4450 65 4465 85
rect 4485 65 4500 85
rect 4450 50 4500 65
rect 4600 735 4650 750
rect 4600 715 4615 735
rect 4635 715 4650 735
rect 4600 685 4650 715
rect 4600 665 4615 685
rect 4635 665 4650 685
rect 4600 635 4650 665
rect 4600 615 4615 635
rect 4635 615 4650 635
rect 4600 585 4650 615
rect 4600 565 4615 585
rect 4635 565 4650 585
rect 4600 535 4650 565
rect 4600 515 4615 535
rect 4635 515 4650 535
rect 4600 485 4650 515
rect 4600 465 4615 485
rect 4635 465 4650 485
rect 4600 435 4650 465
rect 4600 415 4615 435
rect 4635 415 4650 435
rect 4600 385 4650 415
rect 4600 365 4615 385
rect 4635 365 4650 385
rect 4600 335 4650 365
rect 4600 315 4615 335
rect 4635 315 4650 335
rect 4600 285 4650 315
rect 4600 265 4615 285
rect 4635 265 4650 285
rect 4600 235 4650 265
rect 4600 215 4615 235
rect 4635 215 4650 235
rect 4600 185 4650 215
rect 4600 165 4615 185
rect 4635 165 4650 185
rect 4600 135 4650 165
rect 4600 115 4615 135
rect 4635 115 4650 135
rect 4600 85 4650 115
rect 4600 65 4615 85
rect 4635 65 4650 85
rect 4600 50 4650 65
rect 4750 735 4800 750
rect 4750 715 4765 735
rect 4785 715 4800 735
rect 4750 685 4800 715
rect 4750 665 4765 685
rect 4785 665 4800 685
rect 4750 635 4800 665
rect 4750 615 4765 635
rect 4785 615 4800 635
rect 4750 585 4800 615
rect 4750 565 4765 585
rect 4785 565 4800 585
rect 4750 535 4800 565
rect 4750 515 4765 535
rect 4785 515 4800 535
rect 4750 485 4800 515
rect 4750 465 4765 485
rect 4785 465 4800 485
rect 4750 435 4800 465
rect 4750 415 4765 435
rect 4785 415 4800 435
rect 4750 385 4800 415
rect 4750 365 4765 385
rect 4785 365 4800 385
rect 4750 335 4800 365
rect 4750 315 4765 335
rect 4785 315 4800 335
rect 4750 285 4800 315
rect 4750 265 4765 285
rect 4785 265 4800 285
rect 4750 235 4800 265
rect 4750 215 4765 235
rect 4785 215 4800 235
rect 4750 185 4800 215
rect 4750 165 4765 185
rect 4785 165 4800 185
rect 4750 135 4800 165
rect 4750 115 4765 135
rect 4785 115 4800 135
rect 4750 85 4800 115
rect 4750 65 4765 85
rect 4785 65 4800 85
rect 4750 50 4800 65
rect 4900 50 4950 750
rect 5050 735 5100 750
rect 5050 715 5065 735
rect 5085 715 5100 735
rect 5050 685 5100 715
rect 5050 665 5065 685
rect 5085 665 5100 685
rect 5050 635 5100 665
rect 5050 615 5065 635
rect 5085 615 5100 635
rect 5050 585 5100 615
rect 5050 565 5065 585
rect 5085 565 5100 585
rect 5050 535 5100 565
rect 5050 515 5065 535
rect 5085 515 5100 535
rect 5050 485 5100 515
rect 5050 465 5065 485
rect 5085 465 5100 485
rect 5050 435 5100 465
rect 5050 415 5065 435
rect 5085 415 5100 435
rect 5050 385 5100 415
rect 5050 365 5065 385
rect 5085 365 5100 385
rect 5050 335 5100 365
rect 5050 315 5065 335
rect 5085 315 5100 335
rect 5050 285 5100 315
rect 5050 265 5065 285
rect 5085 265 5100 285
rect 5050 235 5100 265
rect 5050 215 5065 235
rect 5085 215 5100 235
rect 5050 185 5100 215
rect 5050 165 5065 185
rect 5085 165 5100 185
rect 5050 135 5100 165
rect 5050 115 5065 135
rect 5085 115 5100 135
rect 5050 85 5100 115
rect 5050 65 5065 85
rect 5085 65 5100 85
rect 5050 50 5100 65
rect 5200 50 5250 750
rect 5350 735 5400 750
rect 5350 715 5365 735
rect 5385 715 5400 735
rect 5350 685 5400 715
rect 5350 665 5365 685
rect 5385 665 5400 685
rect 5350 635 5400 665
rect 5350 615 5365 635
rect 5385 615 5400 635
rect 5350 585 5400 615
rect 5350 565 5365 585
rect 5385 565 5400 585
rect 5350 535 5400 565
rect 5350 515 5365 535
rect 5385 515 5400 535
rect 5350 485 5400 515
rect 5350 465 5365 485
rect 5385 465 5400 485
rect 5350 435 5400 465
rect 5350 415 5365 435
rect 5385 415 5400 435
rect 5350 385 5400 415
rect 5350 365 5365 385
rect 5385 365 5400 385
rect 5350 335 5400 365
rect 5350 315 5365 335
rect 5385 315 5400 335
rect 5350 285 5400 315
rect 5350 265 5365 285
rect 5385 265 5400 285
rect 5350 235 5400 265
rect 5350 215 5365 235
rect 5385 215 5400 235
rect 5350 185 5400 215
rect 5350 165 5365 185
rect 5385 165 5400 185
rect 5350 135 5400 165
rect 5350 115 5365 135
rect 5385 115 5400 135
rect 5350 85 5400 115
rect 5350 65 5365 85
rect 5385 65 5400 85
rect 5350 50 5400 65
rect 5500 50 5550 750
rect 5650 735 5700 750
rect 5650 715 5665 735
rect 5685 715 5700 735
rect 5650 685 5700 715
rect 5650 665 5665 685
rect 5685 665 5700 685
rect 5650 635 5700 665
rect 5650 615 5665 635
rect 5685 615 5700 635
rect 5650 585 5700 615
rect 5650 565 5665 585
rect 5685 565 5700 585
rect 5650 535 5700 565
rect 5650 515 5665 535
rect 5685 515 5700 535
rect 5650 485 5700 515
rect 5650 465 5665 485
rect 5685 465 5700 485
rect 5650 435 5700 465
rect 5650 415 5665 435
rect 5685 415 5700 435
rect 5650 385 5700 415
rect 5650 365 5665 385
rect 5685 365 5700 385
rect 5650 335 5700 365
rect 5650 315 5665 335
rect 5685 315 5700 335
rect 5650 285 5700 315
rect 5650 265 5665 285
rect 5685 265 5700 285
rect 5650 235 5700 265
rect 5650 215 5665 235
rect 5685 215 5700 235
rect 5650 185 5700 215
rect 5650 165 5665 185
rect 5685 165 5700 185
rect 5650 135 5700 165
rect 5650 115 5665 135
rect 5685 115 5700 135
rect 5650 85 5700 115
rect 5650 65 5665 85
rect 5685 65 5700 85
rect 5650 50 5700 65
rect 5800 50 5850 750
rect 5950 735 6000 750
rect 5950 715 5965 735
rect 5985 715 6000 735
rect 5950 685 6000 715
rect 5950 665 5965 685
rect 5985 665 6000 685
rect 5950 635 6000 665
rect 5950 615 5965 635
rect 5985 615 6000 635
rect 5950 585 6000 615
rect 5950 565 5965 585
rect 5985 565 6000 585
rect 5950 535 6000 565
rect 5950 515 5965 535
rect 5985 515 6000 535
rect 5950 485 6000 515
rect 5950 465 5965 485
rect 5985 465 6000 485
rect 5950 435 6000 465
rect 5950 415 5965 435
rect 5985 415 6000 435
rect 5950 385 6000 415
rect 5950 365 5965 385
rect 5985 365 6000 385
rect 5950 335 6000 365
rect 5950 315 5965 335
rect 5985 315 6000 335
rect 5950 285 6000 315
rect 5950 265 5965 285
rect 5985 265 6000 285
rect 5950 235 6000 265
rect 5950 215 5965 235
rect 5985 215 6000 235
rect 5950 185 6000 215
rect 5950 165 5965 185
rect 5985 165 6000 185
rect 5950 135 6000 165
rect 5950 115 5965 135
rect 5985 115 6000 135
rect 5950 85 6000 115
rect 5950 65 5965 85
rect 5985 65 6000 85
rect 5950 50 6000 65
rect 6100 50 6150 750
rect 6250 735 6300 750
rect 6250 715 6265 735
rect 6285 715 6300 735
rect 6250 685 6300 715
rect 6250 665 6265 685
rect 6285 665 6300 685
rect 6250 635 6300 665
rect 6250 615 6265 635
rect 6285 615 6300 635
rect 6250 585 6300 615
rect 6250 565 6265 585
rect 6285 565 6300 585
rect 6250 535 6300 565
rect 6250 515 6265 535
rect 6285 515 6300 535
rect 6250 485 6300 515
rect 6250 465 6265 485
rect 6285 465 6300 485
rect 6250 435 6300 465
rect 6250 415 6265 435
rect 6285 415 6300 435
rect 6250 385 6300 415
rect 6250 365 6265 385
rect 6285 365 6300 385
rect 6250 335 6300 365
rect 6250 315 6265 335
rect 6285 315 6300 335
rect 6250 285 6300 315
rect 6250 265 6265 285
rect 6285 265 6300 285
rect 6250 235 6300 265
rect 6250 215 6265 235
rect 6285 215 6300 235
rect 6250 185 6300 215
rect 6250 165 6265 185
rect 6285 165 6300 185
rect 6250 135 6300 165
rect 6250 115 6265 135
rect 6285 115 6300 135
rect 6250 85 6300 115
rect 6250 65 6265 85
rect 6285 65 6300 85
rect 6250 50 6300 65
rect 6400 50 6450 750
rect 6550 735 6600 750
rect 6550 715 6565 735
rect 6585 715 6600 735
rect 6550 685 6600 715
rect 6550 665 6565 685
rect 6585 665 6600 685
rect 6550 635 6600 665
rect 6550 615 6565 635
rect 6585 615 6600 635
rect 6550 585 6600 615
rect 6550 565 6565 585
rect 6585 565 6600 585
rect 6550 535 6600 565
rect 6550 515 6565 535
rect 6585 515 6600 535
rect 6550 485 6600 515
rect 6550 465 6565 485
rect 6585 465 6600 485
rect 6550 435 6600 465
rect 6550 415 6565 435
rect 6585 415 6600 435
rect 6550 385 6600 415
rect 6550 365 6565 385
rect 6585 365 6600 385
rect 6550 335 6600 365
rect 6550 315 6565 335
rect 6585 315 6600 335
rect 6550 285 6600 315
rect 6550 265 6565 285
rect 6585 265 6600 285
rect 6550 235 6600 265
rect 6550 215 6565 235
rect 6585 215 6600 235
rect 6550 185 6600 215
rect 6550 165 6565 185
rect 6585 165 6600 185
rect 6550 135 6600 165
rect 6550 115 6565 135
rect 6585 115 6600 135
rect 6550 85 6600 115
rect 6550 65 6565 85
rect 6585 65 6600 85
rect 6550 50 6600 65
rect 6700 50 6750 750
rect 6850 735 6900 750
rect 6850 715 6865 735
rect 6885 715 6900 735
rect 6850 685 6900 715
rect 6850 665 6865 685
rect 6885 665 6900 685
rect 6850 635 6900 665
rect 6850 615 6865 635
rect 6885 615 6900 635
rect 6850 585 6900 615
rect 6850 565 6865 585
rect 6885 565 6900 585
rect 6850 535 6900 565
rect 6850 515 6865 535
rect 6885 515 6900 535
rect 6850 485 6900 515
rect 6850 465 6865 485
rect 6885 465 6900 485
rect 6850 435 6900 465
rect 6850 415 6865 435
rect 6885 415 6900 435
rect 6850 385 6900 415
rect 6850 365 6865 385
rect 6885 365 6900 385
rect 6850 335 6900 365
rect 6850 315 6865 335
rect 6885 315 6900 335
rect 6850 285 6900 315
rect 6850 265 6865 285
rect 6885 265 6900 285
rect 6850 235 6900 265
rect 6850 215 6865 235
rect 6885 215 6900 235
rect 6850 185 6900 215
rect 6850 165 6865 185
rect 6885 165 6900 185
rect 6850 135 6900 165
rect 6850 115 6865 135
rect 6885 115 6900 135
rect 6850 85 6900 115
rect 6850 65 6865 85
rect 6885 65 6900 85
rect 6850 50 6900 65
rect 7000 50 7050 750
rect 7150 735 7200 750
rect 7150 715 7165 735
rect 7185 715 7200 735
rect 7150 685 7200 715
rect 7150 665 7165 685
rect 7185 665 7200 685
rect 7150 635 7200 665
rect 7150 615 7165 635
rect 7185 615 7200 635
rect 7150 585 7200 615
rect 7150 565 7165 585
rect 7185 565 7200 585
rect 7150 535 7200 565
rect 7150 515 7165 535
rect 7185 515 7200 535
rect 7150 485 7200 515
rect 7150 465 7165 485
rect 7185 465 7200 485
rect 7150 435 7200 465
rect 7150 415 7165 435
rect 7185 415 7200 435
rect 7150 385 7200 415
rect 7150 365 7165 385
rect 7185 365 7200 385
rect 7150 335 7200 365
rect 7150 315 7165 335
rect 7185 315 7200 335
rect 7150 285 7200 315
rect 7150 265 7165 285
rect 7185 265 7200 285
rect 7150 235 7200 265
rect 7150 215 7165 235
rect 7185 215 7200 235
rect 7150 185 7200 215
rect 7150 165 7165 185
rect 7185 165 7200 185
rect 7150 135 7200 165
rect 7150 115 7165 135
rect 7185 115 7200 135
rect 7150 85 7200 115
rect 7150 65 7165 85
rect 7185 65 7200 85
rect 7150 50 7200 65
rect 7300 50 7350 750
rect 7450 50 7500 750
rect 7600 50 7650 750
rect 7750 50 7800 750
rect 7900 50 7950 750
rect 8050 50 8100 750
rect 8200 50 8250 750
rect 8350 735 8400 750
rect 8350 715 8365 735
rect 8385 715 8400 735
rect 8350 685 8400 715
rect 8350 665 8365 685
rect 8385 665 8400 685
rect 8350 635 8400 665
rect 8350 615 8365 635
rect 8385 615 8400 635
rect 8350 585 8400 615
rect 8350 565 8365 585
rect 8385 565 8400 585
rect 8350 535 8400 565
rect 8350 515 8365 535
rect 8385 515 8400 535
rect 8350 485 8400 515
rect 8350 465 8365 485
rect 8385 465 8400 485
rect 8350 435 8400 465
rect 8350 415 8365 435
rect 8385 415 8400 435
rect 8350 385 8400 415
rect 8350 365 8365 385
rect 8385 365 8400 385
rect 8350 335 8400 365
rect 8350 315 8365 335
rect 8385 315 8400 335
rect 8350 285 8400 315
rect 8350 265 8365 285
rect 8385 265 8400 285
rect 8350 235 8400 265
rect 8350 215 8365 235
rect 8385 215 8400 235
rect 8350 185 8400 215
rect 8350 165 8365 185
rect 8385 165 8400 185
rect 8350 135 8400 165
rect 8350 115 8365 135
rect 8385 115 8400 135
rect 8350 85 8400 115
rect 8350 65 8365 85
rect 8385 65 8400 85
rect 8350 50 8400 65
rect 8500 50 8550 750
rect 8650 50 8700 750
rect 8800 50 8850 750
rect 8950 50 9000 750
rect 9100 50 9150 750
rect 9250 50 9300 750
rect 9400 50 9450 750
rect 9550 735 9600 750
rect 9550 715 9565 735
rect 9585 715 9600 735
rect 9550 685 9600 715
rect 9550 665 9565 685
rect 9585 665 9600 685
rect 9550 635 9600 665
rect 9550 615 9565 635
rect 9585 615 9600 635
rect 9550 585 9600 615
rect 9550 565 9565 585
rect 9585 565 9600 585
rect 9550 535 9600 565
rect 9550 515 9565 535
rect 9585 515 9600 535
rect 9550 485 9600 515
rect 9550 465 9565 485
rect 9585 465 9600 485
rect 9550 435 9600 465
rect 9550 415 9565 435
rect 9585 415 9600 435
rect 9550 385 9600 415
rect 9550 365 9565 385
rect 9585 365 9600 385
rect 9550 335 9600 365
rect 9550 315 9565 335
rect 9585 315 9600 335
rect 9550 285 9600 315
rect 9550 265 9565 285
rect 9585 265 9600 285
rect 9550 235 9600 265
rect 9550 215 9565 235
rect 9585 215 9600 235
rect 9550 185 9600 215
rect 9550 165 9565 185
rect 9585 165 9600 185
rect 9550 135 9600 165
rect 9550 115 9565 135
rect 9585 115 9600 135
rect 9550 85 9600 115
rect 9550 65 9565 85
rect 9585 65 9600 85
rect 9550 50 9600 65
rect 9700 50 9750 750
rect 9850 50 9900 750
rect 10000 50 10050 750
rect 10150 50 10200 750
rect 10300 50 10350 750
rect 10450 50 10500 750
rect 10600 50 10650 750
rect 10750 735 10800 750
rect 10750 715 10765 735
rect 10785 715 10800 735
rect 10750 685 10800 715
rect 10750 665 10765 685
rect 10785 665 10800 685
rect 10750 635 10800 665
rect 10750 615 10765 635
rect 10785 615 10800 635
rect 10750 585 10800 615
rect 10750 565 10765 585
rect 10785 565 10800 585
rect 10750 535 10800 565
rect 10750 515 10765 535
rect 10785 515 10800 535
rect 10750 485 10800 515
rect 10750 465 10765 485
rect 10785 465 10800 485
rect 10750 435 10800 465
rect 10750 415 10765 435
rect 10785 415 10800 435
rect 10750 385 10800 415
rect 10750 365 10765 385
rect 10785 365 10800 385
rect 10750 335 10800 365
rect 10750 315 10765 335
rect 10785 315 10800 335
rect 10750 285 10800 315
rect 10750 265 10765 285
rect 10785 265 10800 285
rect 10750 235 10800 265
rect 10750 215 10765 235
rect 10785 215 10800 235
rect 10750 185 10800 215
rect 10750 165 10765 185
rect 10785 165 10800 185
rect 10750 135 10800 165
rect 10750 115 10765 135
rect 10785 115 10800 135
rect 10750 85 10800 115
rect 10750 65 10765 85
rect 10785 65 10800 85
rect 10750 50 10800 65
rect 10900 50 10950 750
rect 11050 50 11100 750
rect 11200 50 11250 750
rect 11350 50 11400 750
rect 11500 50 11550 750
rect 11650 50 11700 750
rect 11800 50 11850 750
rect 11950 735 12000 750
rect 11950 715 11965 735
rect 11985 715 12000 735
rect 11950 685 12000 715
rect 11950 665 11965 685
rect 11985 665 12000 685
rect 11950 635 12000 665
rect 11950 615 11965 635
rect 11985 615 12000 635
rect 11950 585 12000 615
rect 11950 565 11965 585
rect 11985 565 12000 585
rect 11950 535 12000 565
rect 11950 515 11965 535
rect 11985 515 12000 535
rect 11950 485 12000 515
rect 11950 465 11965 485
rect 11985 465 12000 485
rect 11950 435 12000 465
rect 11950 415 11965 435
rect 11985 415 12000 435
rect 11950 385 12000 415
rect 11950 365 11965 385
rect 11985 365 12000 385
rect 11950 335 12000 365
rect 11950 315 11965 335
rect 11985 315 12000 335
rect 11950 285 12000 315
rect 11950 265 11965 285
rect 11985 265 12000 285
rect 11950 235 12000 265
rect 11950 215 11965 235
rect 11985 215 12000 235
rect 11950 185 12000 215
rect 11950 165 11965 185
rect 11985 165 12000 185
rect 11950 135 12000 165
rect 11950 115 11965 135
rect 11985 115 12000 135
rect 11950 85 12000 115
rect 11950 65 11965 85
rect 11985 65 12000 85
rect 11950 50 12000 65
rect 12100 50 12150 750
rect 12250 735 12300 750
rect 12250 715 12265 735
rect 12285 715 12300 735
rect 12250 685 12300 715
rect 12250 665 12265 685
rect 12285 665 12300 685
rect 12250 635 12300 665
rect 12250 615 12265 635
rect 12285 615 12300 635
rect 12250 585 12300 615
rect 12250 565 12265 585
rect 12285 565 12300 585
rect 12250 535 12300 565
rect 12250 515 12265 535
rect 12285 515 12300 535
rect 12250 485 12300 515
rect 12250 465 12265 485
rect 12285 465 12300 485
rect 12250 435 12300 465
rect 12250 415 12265 435
rect 12285 415 12300 435
rect 12250 385 12300 415
rect 12250 365 12265 385
rect 12285 365 12300 385
rect 12250 335 12300 365
rect 12250 315 12265 335
rect 12285 315 12300 335
rect 12250 285 12300 315
rect 12250 265 12265 285
rect 12285 265 12300 285
rect 12250 235 12300 265
rect 12250 215 12265 235
rect 12285 215 12300 235
rect 12250 185 12300 215
rect 12250 165 12265 185
rect 12285 165 12300 185
rect 12250 135 12300 165
rect 12250 115 12265 135
rect 12285 115 12300 135
rect 12250 85 12300 115
rect 12250 65 12265 85
rect 12285 65 12300 85
rect 12250 50 12300 65
rect 12400 50 12450 750
rect 12550 735 12600 750
rect 12550 715 12565 735
rect 12585 715 12600 735
rect 12550 685 12600 715
rect 12550 665 12565 685
rect 12585 665 12600 685
rect 12550 635 12600 665
rect 12550 615 12565 635
rect 12585 615 12600 635
rect 12550 585 12600 615
rect 12550 565 12565 585
rect 12585 565 12600 585
rect 12550 535 12600 565
rect 12550 515 12565 535
rect 12585 515 12600 535
rect 12550 485 12600 515
rect 12550 465 12565 485
rect 12585 465 12600 485
rect 12550 435 12600 465
rect 12550 415 12565 435
rect 12585 415 12600 435
rect 12550 385 12600 415
rect 12550 365 12565 385
rect 12585 365 12600 385
rect 12550 335 12600 365
rect 12550 315 12565 335
rect 12585 315 12600 335
rect 12550 285 12600 315
rect 12550 265 12565 285
rect 12585 265 12600 285
rect 12550 235 12600 265
rect 12550 215 12565 235
rect 12585 215 12600 235
rect 12550 185 12600 215
rect 12550 165 12565 185
rect 12585 165 12600 185
rect 12550 135 12600 165
rect 12550 115 12565 135
rect 12585 115 12600 135
rect 12550 85 12600 115
rect 12550 65 12565 85
rect 12585 65 12600 85
rect 12550 50 12600 65
rect 12700 50 12750 750
rect 12850 735 12900 750
rect 12850 715 12865 735
rect 12885 715 12900 735
rect 12850 685 12900 715
rect 12850 665 12865 685
rect 12885 665 12900 685
rect 12850 635 12900 665
rect 12850 615 12865 635
rect 12885 615 12900 635
rect 12850 585 12900 615
rect 12850 565 12865 585
rect 12885 565 12900 585
rect 12850 535 12900 565
rect 12850 515 12865 535
rect 12885 515 12900 535
rect 12850 485 12900 515
rect 12850 465 12865 485
rect 12885 465 12900 485
rect 12850 435 12900 465
rect 12850 415 12865 435
rect 12885 415 12900 435
rect 12850 385 12900 415
rect 12850 365 12865 385
rect 12885 365 12900 385
rect 12850 335 12900 365
rect 12850 315 12865 335
rect 12885 315 12900 335
rect 12850 285 12900 315
rect 12850 265 12865 285
rect 12885 265 12900 285
rect 12850 235 12900 265
rect 12850 215 12865 235
rect 12885 215 12900 235
rect 12850 185 12900 215
rect 12850 165 12865 185
rect 12885 165 12900 185
rect 12850 135 12900 165
rect 12850 115 12865 135
rect 12885 115 12900 135
rect 12850 85 12900 115
rect 12850 65 12865 85
rect 12885 65 12900 85
rect 12850 50 12900 65
rect 13000 50 13050 750
rect 13150 735 13200 750
rect 13150 715 13165 735
rect 13185 715 13200 735
rect 13150 685 13200 715
rect 13150 665 13165 685
rect 13185 665 13200 685
rect 13150 635 13200 665
rect 13150 615 13165 635
rect 13185 615 13200 635
rect 13150 585 13200 615
rect 13150 565 13165 585
rect 13185 565 13200 585
rect 13150 535 13200 565
rect 13150 515 13165 535
rect 13185 515 13200 535
rect 13150 485 13200 515
rect 13150 465 13165 485
rect 13185 465 13200 485
rect 13150 435 13200 465
rect 13150 415 13165 435
rect 13185 415 13200 435
rect 13150 385 13200 415
rect 13150 365 13165 385
rect 13185 365 13200 385
rect 13150 335 13200 365
rect 13150 315 13165 335
rect 13185 315 13200 335
rect 13150 285 13200 315
rect 13150 265 13165 285
rect 13185 265 13200 285
rect 13150 235 13200 265
rect 13150 215 13165 235
rect 13185 215 13200 235
rect 13150 185 13200 215
rect 13150 165 13165 185
rect 13185 165 13200 185
rect 13150 135 13200 165
rect 13150 115 13165 135
rect 13185 115 13200 135
rect 13150 85 13200 115
rect 13150 65 13165 85
rect 13185 65 13200 85
rect 13150 50 13200 65
rect 13300 50 13350 750
rect 13450 735 13500 750
rect 13450 715 13465 735
rect 13485 715 13500 735
rect 13450 685 13500 715
rect 13450 665 13465 685
rect 13485 665 13500 685
rect 13450 635 13500 665
rect 13450 615 13465 635
rect 13485 615 13500 635
rect 13450 585 13500 615
rect 13450 565 13465 585
rect 13485 565 13500 585
rect 13450 535 13500 565
rect 13450 515 13465 535
rect 13485 515 13500 535
rect 13450 485 13500 515
rect 13450 465 13465 485
rect 13485 465 13500 485
rect 13450 435 13500 465
rect 13450 415 13465 435
rect 13485 415 13500 435
rect 13450 385 13500 415
rect 13450 365 13465 385
rect 13485 365 13500 385
rect 13450 335 13500 365
rect 13450 315 13465 335
rect 13485 315 13500 335
rect 13450 285 13500 315
rect 13450 265 13465 285
rect 13485 265 13500 285
rect 13450 235 13500 265
rect 13450 215 13465 235
rect 13485 215 13500 235
rect 13450 185 13500 215
rect 13450 165 13465 185
rect 13485 165 13500 185
rect 13450 135 13500 165
rect 13450 115 13465 135
rect 13485 115 13500 135
rect 13450 85 13500 115
rect 13450 65 13465 85
rect 13485 65 13500 85
rect 13450 50 13500 65
rect 13600 50 13650 750
rect 13750 735 13800 750
rect 13750 715 13765 735
rect 13785 715 13800 735
rect 13750 685 13800 715
rect 13750 665 13765 685
rect 13785 665 13800 685
rect 13750 635 13800 665
rect 13750 615 13765 635
rect 13785 615 13800 635
rect 13750 585 13800 615
rect 13750 565 13765 585
rect 13785 565 13800 585
rect 13750 535 13800 565
rect 13750 515 13765 535
rect 13785 515 13800 535
rect 13750 485 13800 515
rect 13750 465 13765 485
rect 13785 465 13800 485
rect 13750 435 13800 465
rect 13750 415 13765 435
rect 13785 415 13800 435
rect 13750 385 13800 415
rect 13750 365 13765 385
rect 13785 365 13800 385
rect 13750 335 13800 365
rect 13750 315 13765 335
rect 13785 315 13800 335
rect 13750 285 13800 315
rect 13750 265 13765 285
rect 13785 265 13800 285
rect 13750 235 13800 265
rect 13750 215 13765 235
rect 13785 215 13800 235
rect 13750 185 13800 215
rect 13750 165 13765 185
rect 13785 165 13800 185
rect 13750 135 13800 165
rect 13750 115 13765 135
rect 13785 115 13800 135
rect 13750 85 13800 115
rect 13750 65 13765 85
rect 13785 65 13800 85
rect 13750 50 13800 65
rect 13900 50 13950 750
rect 14050 735 14100 750
rect 14050 715 14065 735
rect 14085 715 14100 735
rect 14050 685 14100 715
rect 14050 665 14065 685
rect 14085 665 14100 685
rect 14050 635 14100 665
rect 14050 615 14065 635
rect 14085 615 14100 635
rect 14050 585 14100 615
rect 14050 565 14065 585
rect 14085 565 14100 585
rect 14050 535 14100 565
rect 14050 515 14065 535
rect 14085 515 14100 535
rect 14050 485 14100 515
rect 14050 465 14065 485
rect 14085 465 14100 485
rect 14050 435 14100 465
rect 14050 415 14065 435
rect 14085 415 14100 435
rect 14050 385 14100 415
rect 14050 365 14065 385
rect 14085 365 14100 385
rect 14050 335 14100 365
rect 14050 315 14065 335
rect 14085 315 14100 335
rect 14050 285 14100 315
rect 14050 265 14065 285
rect 14085 265 14100 285
rect 14050 235 14100 265
rect 14050 215 14065 235
rect 14085 215 14100 235
rect 14050 185 14100 215
rect 14050 165 14065 185
rect 14085 165 14100 185
rect 14050 135 14100 165
rect 14050 115 14065 135
rect 14085 115 14100 135
rect 14050 85 14100 115
rect 14050 65 14065 85
rect 14085 65 14100 85
rect 14050 50 14100 65
rect 14200 50 14250 750
rect 14350 735 14400 750
rect 14350 715 14365 735
rect 14385 715 14400 735
rect 14350 685 14400 715
rect 14350 665 14365 685
rect 14385 665 14400 685
rect 14350 635 14400 665
rect 14350 615 14365 635
rect 14385 615 14400 635
rect 14350 585 14400 615
rect 14350 565 14365 585
rect 14385 565 14400 585
rect 14350 535 14400 565
rect 14350 515 14365 535
rect 14385 515 14400 535
rect 14350 485 14400 515
rect 14350 465 14365 485
rect 14385 465 14400 485
rect 14350 435 14400 465
rect 14350 415 14365 435
rect 14385 415 14400 435
rect 14350 385 14400 415
rect 14350 365 14365 385
rect 14385 365 14400 385
rect 14350 335 14400 365
rect 14350 315 14365 335
rect 14385 315 14400 335
rect 14350 285 14400 315
rect 14350 265 14365 285
rect 14385 265 14400 285
rect 14350 235 14400 265
rect 14350 215 14365 235
rect 14385 215 14400 235
rect 14350 185 14400 215
rect 14350 165 14365 185
rect 14385 165 14400 185
rect 14350 135 14400 165
rect 14350 115 14365 135
rect 14385 115 14400 135
rect 14350 85 14400 115
rect 14350 65 14365 85
rect 14385 65 14400 85
rect 14350 50 14400 65
rect 14500 50 14550 750
rect 14650 50 14700 750
rect 14800 50 14850 750
rect 14950 50 15000 750
rect 15100 50 15150 750
rect 15250 50 15300 750
rect 15400 50 15450 750
rect 15550 735 15600 750
rect 15550 715 15565 735
rect 15585 715 15600 735
rect 15550 685 15600 715
rect 15550 665 15565 685
rect 15585 665 15600 685
rect 15550 635 15600 665
rect 15550 615 15565 635
rect 15585 615 15600 635
rect 15550 585 15600 615
rect 15550 565 15565 585
rect 15585 565 15600 585
rect 15550 535 15600 565
rect 15550 515 15565 535
rect 15585 515 15600 535
rect 15550 485 15600 515
rect 15550 465 15565 485
rect 15585 465 15600 485
rect 15550 435 15600 465
rect 15550 415 15565 435
rect 15585 415 15600 435
rect 15550 385 15600 415
rect 15550 365 15565 385
rect 15585 365 15600 385
rect 15550 335 15600 365
rect 15550 315 15565 335
rect 15585 315 15600 335
rect 15550 285 15600 315
rect 15550 265 15565 285
rect 15585 265 15600 285
rect 15550 235 15600 265
rect 15550 215 15565 235
rect 15585 215 15600 235
rect 15550 185 15600 215
rect 15550 165 15565 185
rect 15585 165 15600 185
rect 15550 135 15600 165
rect 15550 115 15565 135
rect 15585 115 15600 135
rect 15550 85 15600 115
rect 15550 65 15565 85
rect 15585 65 15600 85
rect 15550 50 15600 65
rect 15700 50 15750 750
rect 15850 50 15900 750
rect 16000 50 16050 750
rect 16150 50 16200 750
rect 16300 50 16350 750
rect 16450 50 16500 750
rect 16600 50 16650 750
rect 16750 735 16800 750
rect 16750 715 16765 735
rect 16785 715 16800 735
rect 16750 685 16800 715
rect 16750 665 16765 685
rect 16785 665 16800 685
rect 16750 635 16800 665
rect 16750 615 16765 635
rect 16785 615 16800 635
rect 16750 585 16800 615
rect 16750 565 16765 585
rect 16785 565 16800 585
rect 16750 535 16800 565
rect 16750 515 16765 535
rect 16785 515 16800 535
rect 16750 485 16800 515
rect 16750 465 16765 485
rect 16785 465 16800 485
rect 16750 435 16800 465
rect 16750 415 16765 435
rect 16785 415 16800 435
rect 16750 385 16800 415
rect 16750 365 16765 385
rect 16785 365 16800 385
rect 16750 335 16800 365
rect 16750 315 16765 335
rect 16785 315 16800 335
rect 16750 285 16800 315
rect 16750 265 16765 285
rect 16785 265 16800 285
rect 16750 235 16800 265
rect 16750 215 16765 235
rect 16785 215 16800 235
rect 16750 185 16800 215
rect 16750 165 16765 185
rect 16785 165 16800 185
rect 16750 135 16800 165
rect 16750 115 16765 135
rect 16785 115 16800 135
rect 16750 85 16800 115
rect 16750 65 16765 85
rect 16785 65 16800 85
rect 16750 50 16800 65
rect 16900 50 16950 750
rect 17050 50 17100 750
rect 17200 50 17250 750
rect 17350 50 17400 750
rect 17500 50 17550 750
rect 17650 50 17700 750
rect 17800 50 17850 750
rect 17950 735 18000 750
rect 17950 715 17965 735
rect 17985 715 18000 735
rect 17950 685 18000 715
rect 17950 665 17965 685
rect 17985 665 18000 685
rect 17950 635 18000 665
rect 17950 615 17965 635
rect 17985 615 18000 635
rect 17950 585 18000 615
rect 17950 565 17965 585
rect 17985 565 18000 585
rect 17950 535 18000 565
rect 17950 515 17965 535
rect 17985 515 18000 535
rect 17950 485 18000 515
rect 17950 465 17965 485
rect 17985 465 18000 485
rect 17950 435 18000 465
rect 17950 415 17965 435
rect 17985 415 18000 435
rect 17950 385 18000 415
rect 17950 365 17965 385
rect 17985 365 18000 385
rect 17950 335 18000 365
rect 17950 315 17965 335
rect 17985 315 18000 335
rect 17950 285 18000 315
rect 17950 265 17965 285
rect 17985 265 18000 285
rect 17950 235 18000 265
rect 17950 215 17965 235
rect 17985 215 18000 235
rect 17950 185 18000 215
rect 17950 165 17965 185
rect 17985 165 18000 185
rect 17950 135 18000 165
rect 17950 115 17965 135
rect 17985 115 18000 135
rect 17950 85 18000 115
rect 17950 65 17965 85
rect 17985 65 18000 85
rect 17950 50 18000 65
rect 18100 50 18150 750
rect 18250 50 18300 750
rect 18400 50 18450 750
rect 18550 50 18600 750
rect 18700 50 18750 750
rect 18850 50 18900 750
rect 19000 50 19050 750
rect 19150 735 19200 750
rect 19150 715 19165 735
rect 19185 715 19200 735
rect 19150 685 19200 715
rect 19150 665 19165 685
rect 19185 665 19200 685
rect 19150 635 19200 665
rect 19150 615 19165 635
rect 19185 615 19200 635
rect 19150 585 19200 615
rect 19150 565 19165 585
rect 19185 565 19200 585
rect 19150 535 19200 565
rect 19150 515 19165 535
rect 19185 515 19200 535
rect 19150 485 19200 515
rect 19150 465 19165 485
rect 19185 465 19200 485
rect 19150 435 19200 465
rect 19150 415 19165 435
rect 19185 415 19200 435
rect 19150 385 19200 415
rect 19150 365 19165 385
rect 19185 365 19200 385
rect 19150 335 19200 365
rect 19150 315 19165 335
rect 19185 315 19200 335
rect 19150 285 19200 315
rect 19150 265 19165 285
rect 19185 265 19200 285
rect 19150 235 19200 265
rect 19150 215 19165 235
rect 19185 215 19200 235
rect 19150 185 19200 215
rect 19150 165 19165 185
rect 19185 165 19200 185
rect 19150 135 19200 165
rect 19150 115 19165 135
rect 19185 115 19200 135
rect 19150 85 19200 115
rect 19150 65 19165 85
rect 19185 65 19200 85
rect 19150 50 19200 65
rect 19300 50 19350 750
rect 19450 50 19500 750
rect 19600 50 19650 750
rect 19750 50 19800 750
rect 19900 50 19950 750
rect 20050 50 20100 750
rect 20200 50 20250 750
rect 20350 735 20400 750
rect 20350 715 20365 735
rect 20385 715 20400 735
rect 20350 685 20400 715
rect 20350 665 20365 685
rect 20385 665 20400 685
rect 20350 635 20400 665
rect 20350 615 20365 635
rect 20385 615 20400 635
rect 20350 585 20400 615
rect 20350 565 20365 585
rect 20385 565 20400 585
rect 20350 535 20400 565
rect 20350 515 20365 535
rect 20385 515 20400 535
rect 20350 485 20400 515
rect 20350 465 20365 485
rect 20385 465 20400 485
rect 20350 435 20400 465
rect 20350 415 20365 435
rect 20385 415 20400 435
rect 20350 385 20400 415
rect 20350 365 20365 385
rect 20385 365 20400 385
rect 20350 335 20400 365
rect 20350 315 20365 335
rect 20385 315 20400 335
rect 20350 285 20400 315
rect 20350 265 20365 285
rect 20385 265 20400 285
rect 20350 235 20400 265
rect 20350 215 20365 235
rect 20385 215 20400 235
rect 20350 185 20400 215
rect 20350 165 20365 185
rect 20385 165 20400 185
rect 20350 135 20400 165
rect 20350 115 20365 135
rect 20385 115 20400 135
rect 20350 85 20400 115
rect 20350 65 20365 85
rect 20385 65 20400 85
rect 20350 50 20400 65
rect -650 -115 -600 -100
rect -650 -135 -635 -115
rect -615 -135 -600 -115
rect -650 -165 -600 -135
rect -650 -185 -635 -165
rect -615 -185 -600 -165
rect -650 -215 -600 -185
rect -650 -235 -635 -215
rect -615 -235 -600 -215
rect -650 -265 -600 -235
rect -650 -285 -635 -265
rect -615 -285 -600 -265
rect -650 -315 -600 -285
rect -650 -335 -635 -315
rect -615 -335 -600 -315
rect -650 -365 -600 -335
rect -650 -385 -635 -365
rect -615 -385 -600 -365
rect -650 -415 -600 -385
rect -650 -435 -635 -415
rect -615 -435 -600 -415
rect -650 -465 -600 -435
rect -650 -485 -635 -465
rect -615 -485 -600 -465
rect -650 -515 -600 -485
rect -650 -535 -635 -515
rect -615 -535 -600 -515
rect -650 -565 -600 -535
rect -650 -585 -635 -565
rect -615 -585 -600 -565
rect -650 -615 -600 -585
rect -650 -635 -635 -615
rect -615 -635 -600 -615
rect -650 -665 -600 -635
rect -650 -685 -635 -665
rect -615 -685 -600 -665
rect -650 -715 -600 -685
rect -650 -735 -635 -715
rect -615 -735 -600 -715
rect -650 -765 -600 -735
rect -650 -785 -635 -765
rect -615 -785 -600 -765
rect -650 -800 -600 -785
rect -500 -115 -450 -100
rect -500 -135 -485 -115
rect -465 -135 -450 -115
rect -500 -165 -450 -135
rect -500 -185 -485 -165
rect -465 -185 -450 -165
rect -500 -215 -450 -185
rect -500 -235 -485 -215
rect -465 -235 -450 -215
rect -500 -265 -450 -235
rect -500 -285 -485 -265
rect -465 -285 -450 -265
rect -500 -315 -450 -285
rect -500 -335 -485 -315
rect -465 -335 -450 -315
rect -500 -365 -450 -335
rect -500 -385 -485 -365
rect -465 -385 -450 -365
rect -500 -415 -450 -385
rect -500 -435 -485 -415
rect -465 -435 -450 -415
rect -500 -465 -450 -435
rect -500 -485 -485 -465
rect -465 -485 -450 -465
rect -500 -515 -450 -485
rect -500 -535 -485 -515
rect -465 -535 -450 -515
rect -500 -565 -450 -535
rect -500 -585 -485 -565
rect -465 -585 -450 -565
rect -500 -615 -450 -585
rect -500 -635 -485 -615
rect -465 -635 -450 -615
rect -500 -665 -450 -635
rect -500 -685 -485 -665
rect -465 -685 -450 -665
rect -500 -715 -450 -685
rect -500 -735 -485 -715
rect -465 -735 -450 -715
rect -500 -765 -450 -735
rect -500 -785 -485 -765
rect -465 -785 -450 -765
rect -500 -800 -450 -785
rect -350 -115 -300 -100
rect -350 -135 -335 -115
rect -315 -135 -300 -115
rect -350 -165 -300 -135
rect -350 -185 -335 -165
rect -315 -185 -300 -165
rect -350 -215 -300 -185
rect -350 -235 -335 -215
rect -315 -235 -300 -215
rect -350 -265 -300 -235
rect -350 -285 -335 -265
rect -315 -285 -300 -265
rect -350 -315 -300 -285
rect -350 -335 -335 -315
rect -315 -335 -300 -315
rect -350 -365 -300 -335
rect -350 -385 -335 -365
rect -315 -385 -300 -365
rect -350 -415 -300 -385
rect -350 -435 -335 -415
rect -315 -435 -300 -415
rect -350 -465 -300 -435
rect -350 -485 -335 -465
rect -315 -485 -300 -465
rect -350 -515 -300 -485
rect -350 -535 -335 -515
rect -315 -535 -300 -515
rect -350 -565 -300 -535
rect -350 -585 -335 -565
rect -315 -585 -300 -565
rect -350 -615 -300 -585
rect -350 -635 -335 -615
rect -315 -635 -300 -615
rect -350 -665 -300 -635
rect -350 -685 -335 -665
rect -315 -685 -300 -665
rect -350 -715 -300 -685
rect -350 -735 -335 -715
rect -315 -735 -300 -715
rect -350 -765 -300 -735
rect -350 -785 -335 -765
rect -315 -785 -300 -765
rect -350 -800 -300 -785
rect -200 -115 -150 -100
rect -200 -135 -185 -115
rect -165 -135 -150 -115
rect -200 -165 -150 -135
rect -200 -185 -185 -165
rect -165 -185 -150 -165
rect -200 -215 -150 -185
rect -200 -235 -185 -215
rect -165 -235 -150 -215
rect -200 -265 -150 -235
rect -200 -285 -185 -265
rect -165 -285 -150 -265
rect -200 -315 -150 -285
rect -200 -335 -185 -315
rect -165 -335 -150 -315
rect -200 -365 -150 -335
rect -200 -385 -185 -365
rect -165 -385 -150 -365
rect -200 -415 -150 -385
rect -200 -435 -185 -415
rect -165 -435 -150 -415
rect -200 -465 -150 -435
rect -200 -485 -185 -465
rect -165 -485 -150 -465
rect -200 -515 -150 -485
rect -200 -535 -185 -515
rect -165 -535 -150 -515
rect -200 -565 -150 -535
rect -200 -585 -185 -565
rect -165 -585 -150 -565
rect -200 -615 -150 -585
rect -200 -635 -185 -615
rect -165 -635 -150 -615
rect -200 -665 -150 -635
rect -200 -685 -185 -665
rect -165 -685 -150 -665
rect -200 -715 -150 -685
rect -200 -735 -185 -715
rect -165 -735 -150 -715
rect -200 -765 -150 -735
rect -200 -785 -185 -765
rect -165 -785 -150 -765
rect -200 -800 -150 -785
rect -50 -115 0 -100
rect -50 -135 -35 -115
rect -15 -135 0 -115
rect -50 -165 0 -135
rect -50 -185 -35 -165
rect -15 -185 0 -165
rect -50 -215 0 -185
rect -50 -235 -35 -215
rect -15 -235 0 -215
rect -50 -265 0 -235
rect -50 -285 -35 -265
rect -15 -285 0 -265
rect -50 -315 0 -285
rect -50 -335 -35 -315
rect -15 -335 0 -315
rect -50 -365 0 -335
rect -50 -385 -35 -365
rect -15 -385 0 -365
rect -50 -415 0 -385
rect -50 -435 -35 -415
rect -15 -435 0 -415
rect -50 -465 0 -435
rect -50 -485 -35 -465
rect -15 -485 0 -465
rect -50 -515 0 -485
rect -50 -535 -35 -515
rect -15 -535 0 -515
rect -50 -565 0 -535
rect -50 -585 -35 -565
rect -15 -585 0 -565
rect -50 -615 0 -585
rect -50 -635 -35 -615
rect -15 -635 0 -615
rect -50 -665 0 -635
rect -50 -685 -35 -665
rect -15 -685 0 -665
rect -50 -715 0 -685
rect -50 -735 -35 -715
rect -15 -735 0 -715
rect -50 -765 0 -735
rect -50 -785 -35 -765
rect -15 -785 0 -765
rect -50 -800 0 -785
rect 100 -800 150 -100
rect 250 -800 300 -100
rect 400 -800 450 -100
rect 550 -800 600 -100
rect 700 -800 750 -100
rect 850 -800 900 -100
rect 1000 -800 1050 -100
rect 1150 -115 1200 -100
rect 1150 -135 1165 -115
rect 1185 -135 1200 -115
rect 1150 -165 1200 -135
rect 1150 -185 1165 -165
rect 1185 -185 1200 -165
rect 1150 -215 1200 -185
rect 1150 -235 1165 -215
rect 1185 -235 1200 -215
rect 1150 -265 1200 -235
rect 1150 -285 1165 -265
rect 1185 -285 1200 -265
rect 1150 -315 1200 -285
rect 1150 -335 1165 -315
rect 1185 -335 1200 -315
rect 1150 -365 1200 -335
rect 1150 -385 1165 -365
rect 1185 -385 1200 -365
rect 1150 -415 1200 -385
rect 1150 -435 1165 -415
rect 1185 -435 1200 -415
rect 1150 -465 1200 -435
rect 1150 -485 1165 -465
rect 1185 -485 1200 -465
rect 1150 -515 1200 -485
rect 1150 -535 1165 -515
rect 1185 -535 1200 -515
rect 1150 -565 1200 -535
rect 1150 -585 1165 -565
rect 1185 -585 1200 -565
rect 1150 -615 1200 -585
rect 1150 -635 1165 -615
rect 1185 -635 1200 -615
rect 1150 -665 1200 -635
rect 1150 -685 1165 -665
rect 1185 -685 1200 -665
rect 1150 -715 1200 -685
rect 1150 -735 1165 -715
rect 1185 -735 1200 -715
rect 1150 -765 1200 -735
rect 1150 -785 1165 -765
rect 1185 -785 1200 -765
rect 1150 -800 1200 -785
rect 1300 -800 1350 -100
rect 1450 -115 1500 -100
rect 1450 -135 1465 -115
rect 1485 -135 1500 -115
rect 1450 -165 1500 -135
rect 1450 -185 1465 -165
rect 1485 -185 1500 -165
rect 1450 -215 1500 -185
rect 1450 -235 1465 -215
rect 1485 -235 1500 -215
rect 1450 -265 1500 -235
rect 1450 -285 1465 -265
rect 1485 -285 1500 -265
rect 1450 -315 1500 -285
rect 1450 -335 1465 -315
rect 1485 -335 1500 -315
rect 1450 -365 1500 -335
rect 1450 -385 1465 -365
rect 1485 -385 1500 -365
rect 1450 -415 1500 -385
rect 1450 -435 1465 -415
rect 1485 -435 1500 -415
rect 1450 -465 1500 -435
rect 1450 -485 1465 -465
rect 1485 -485 1500 -465
rect 1450 -515 1500 -485
rect 1450 -535 1465 -515
rect 1485 -535 1500 -515
rect 1450 -565 1500 -535
rect 1450 -585 1465 -565
rect 1485 -585 1500 -565
rect 1450 -615 1500 -585
rect 1450 -635 1465 -615
rect 1485 -635 1500 -615
rect 1450 -665 1500 -635
rect 1450 -685 1465 -665
rect 1485 -685 1500 -665
rect 1450 -715 1500 -685
rect 1450 -735 1465 -715
rect 1485 -735 1500 -715
rect 1450 -765 1500 -735
rect 1450 -785 1465 -765
rect 1485 -785 1500 -765
rect 1450 -800 1500 -785
rect 1600 -800 1650 -100
rect 1750 -115 1800 -100
rect 1750 -135 1765 -115
rect 1785 -135 1800 -115
rect 1750 -165 1800 -135
rect 1750 -185 1765 -165
rect 1785 -185 1800 -165
rect 1750 -215 1800 -185
rect 1750 -235 1765 -215
rect 1785 -235 1800 -215
rect 1750 -265 1800 -235
rect 1750 -285 1765 -265
rect 1785 -285 1800 -265
rect 1750 -315 1800 -285
rect 1750 -335 1765 -315
rect 1785 -335 1800 -315
rect 1750 -365 1800 -335
rect 1750 -385 1765 -365
rect 1785 -385 1800 -365
rect 1750 -415 1800 -385
rect 1750 -435 1765 -415
rect 1785 -435 1800 -415
rect 1750 -465 1800 -435
rect 1750 -485 1765 -465
rect 1785 -485 1800 -465
rect 1750 -515 1800 -485
rect 1750 -535 1765 -515
rect 1785 -535 1800 -515
rect 1750 -565 1800 -535
rect 1750 -585 1765 -565
rect 1785 -585 1800 -565
rect 1750 -615 1800 -585
rect 1750 -635 1765 -615
rect 1785 -635 1800 -615
rect 1750 -665 1800 -635
rect 1750 -685 1765 -665
rect 1785 -685 1800 -665
rect 1750 -715 1800 -685
rect 1750 -735 1765 -715
rect 1785 -735 1800 -715
rect 1750 -765 1800 -735
rect 1750 -785 1765 -765
rect 1785 -785 1800 -765
rect 1750 -800 1800 -785
rect 1900 -800 1950 -100
rect 2050 -115 2100 -100
rect 2050 -135 2065 -115
rect 2085 -135 2100 -115
rect 2050 -165 2100 -135
rect 2050 -185 2065 -165
rect 2085 -185 2100 -165
rect 2050 -215 2100 -185
rect 2050 -235 2065 -215
rect 2085 -235 2100 -215
rect 2050 -265 2100 -235
rect 2050 -285 2065 -265
rect 2085 -285 2100 -265
rect 2050 -315 2100 -285
rect 2050 -335 2065 -315
rect 2085 -335 2100 -315
rect 2050 -365 2100 -335
rect 2050 -385 2065 -365
rect 2085 -385 2100 -365
rect 2050 -415 2100 -385
rect 2050 -435 2065 -415
rect 2085 -435 2100 -415
rect 2050 -465 2100 -435
rect 2050 -485 2065 -465
rect 2085 -485 2100 -465
rect 2050 -515 2100 -485
rect 2050 -535 2065 -515
rect 2085 -535 2100 -515
rect 2050 -565 2100 -535
rect 2050 -585 2065 -565
rect 2085 -585 2100 -565
rect 2050 -615 2100 -585
rect 2050 -635 2065 -615
rect 2085 -635 2100 -615
rect 2050 -665 2100 -635
rect 2050 -685 2065 -665
rect 2085 -685 2100 -665
rect 2050 -715 2100 -685
rect 2050 -735 2065 -715
rect 2085 -735 2100 -715
rect 2050 -765 2100 -735
rect 2050 -785 2065 -765
rect 2085 -785 2100 -765
rect 2050 -800 2100 -785
rect 2200 -800 2250 -100
rect 2350 -115 2400 -100
rect 2350 -135 2365 -115
rect 2385 -135 2400 -115
rect 2350 -165 2400 -135
rect 2350 -185 2365 -165
rect 2385 -185 2400 -165
rect 2350 -215 2400 -185
rect 2350 -235 2365 -215
rect 2385 -235 2400 -215
rect 2350 -265 2400 -235
rect 2350 -285 2365 -265
rect 2385 -285 2400 -265
rect 2350 -315 2400 -285
rect 2350 -335 2365 -315
rect 2385 -335 2400 -315
rect 2350 -365 2400 -335
rect 2350 -385 2365 -365
rect 2385 -385 2400 -365
rect 2350 -415 2400 -385
rect 2350 -435 2365 -415
rect 2385 -435 2400 -415
rect 2350 -465 2400 -435
rect 2350 -485 2365 -465
rect 2385 -485 2400 -465
rect 2350 -515 2400 -485
rect 2350 -535 2365 -515
rect 2385 -535 2400 -515
rect 2350 -565 2400 -535
rect 2350 -585 2365 -565
rect 2385 -585 2400 -565
rect 2350 -615 2400 -585
rect 2350 -635 2365 -615
rect 2385 -635 2400 -615
rect 2350 -665 2400 -635
rect 2350 -685 2365 -665
rect 2385 -685 2400 -665
rect 2350 -715 2400 -685
rect 2350 -735 2365 -715
rect 2385 -735 2400 -715
rect 2350 -765 2400 -735
rect 2350 -785 2365 -765
rect 2385 -785 2400 -765
rect 2350 -800 2400 -785
rect 2500 -800 2550 -100
rect 2650 -115 2700 -100
rect 2650 -135 2665 -115
rect 2685 -135 2700 -115
rect 2650 -165 2700 -135
rect 2650 -185 2665 -165
rect 2685 -185 2700 -165
rect 2650 -215 2700 -185
rect 2650 -235 2665 -215
rect 2685 -235 2700 -215
rect 2650 -265 2700 -235
rect 2650 -285 2665 -265
rect 2685 -285 2700 -265
rect 2650 -315 2700 -285
rect 2650 -335 2665 -315
rect 2685 -335 2700 -315
rect 2650 -365 2700 -335
rect 2650 -385 2665 -365
rect 2685 -385 2700 -365
rect 2650 -415 2700 -385
rect 2650 -435 2665 -415
rect 2685 -435 2700 -415
rect 2650 -465 2700 -435
rect 2650 -485 2665 -465
rect 2685 -485 2700 -465
rect 2650 -515 2700 -485
rect 2650 -535 2665 -515
rect 2685 -535 2700 -515
rect 2650 -565 2700 -535
rect 2650 -585 2665 -565
rect 2685 -585 2700 -565
rect 2650 -615 2700 -585
rect 2650 -635 2665 -615
rect 2685 -635 2700 -615
rect 2650 -665 2700 -635
rect 2650 -685 2665 -665
rect 2685 -685 2700 -665
rect 2650 -715 2700 -685
rect 2650 -735 2665 -715
rect 2685 -735 2700 -715
rect 2650 -765 2700 -735
rect 2650 -785 2665 -765
rect 2685 -785 2700 -765
rect 2650 -800 2700 -785
rect 2800 -800 2850 -100
rect 2950 -115 3000 -100
rect 2950 -135 2965 -115
rect 2985 -135 3000 -115
rect 2950 -165 3000 -135
rect 2950 -185 2965 -165
rect 2985 -185 3000 -165
rect 2950 -215 3000 -185
rect 2950 -235 2965 -215
rect 2985 -235 3000 -215
rect 2950 -265 3000 -235
rect 2950 -285 2965 -265
rect 2985 -285 3000 -265
rect 2950 -315 3000 -285
rect 2950 -335 2965 -315
rect 2985 -335 3000 -315
rect 2950 -365 3000 -335
rect 2950 -385 2965 -365
rect 2985 -385 3000 -365
rect 2950 -415 3000 -385
rect 2950 -435 2965 -415
rect 2985 -435 3000 -415
rect 2950 -465 3000 -435
rect 2950 -485 2965 -465
rect 2985 -485 3000 -465
rect 2950 -515 3000 -485
rect 2950 -535 2965 -515
rect 2985 -535 3000 -515
rect 2950 -565 3000 -535
rect 2950 -585 2965 -565
rect 2985 -585 3000 -565
rect 2950 -615 3000 -585
rect 2950 -635 2965 -615
rect 2985 -635 3000 -615
rect 2950 -665 3000 -635
rect 2950 -685 2965 -665
rect 2985 -685 3000 -665
rect 2950 -715 3000 -685
rect 2950 -735 2965 -715
rect 2985 -735 3000 -715
rect 2950 -765 3000 -735
rect 2950 -785 2965 -765
rect 2985 -785 3000 -765
rect 2950 -800 3000 -785
rect 3100 -800 3150 -100
rect 3250 -115 3300 -100
rect 3250 -135 3265 -115
rect 3285 -135 3300 -115
rect 3250 -165 3300 -135
rect 3250 -185 3265 -165
rect 3285 -185 3300 -165
rect 3250 -215 3300 -185
rect 3250 -235 3265 -215
rect 3285 -235 3300 -215
rect 3250 -265 3300 -235
rect 3250 -285 3265 -265
rect 3285 -285 3300 -265
rect 3250 -315 3300 -285
rect 3250 -335 3265 -315
rect 3285 -335 3300 -315
rect 3250 -365 3300 -335
rect 3250 -385 3265 -365
rect 3285 -385 3300 -365
rect 3250 -415 3300 -385
rect 3250 -435 3265 -415
rect 3285 -435 3300 -415
rect 3250 -465 3300 -435
rect 3250 -485 3265 -465
rect 3285 -485 3300 -465
rect 3250 -515 3300 -485
rect 3250 -535 3265 -515
rect 3285 -535 3300 -515
rect 3250 -565 3300 -535
rect 3250 -585 3265 -565
rect 3285 -585 3300 -565
rect 3250 -615 3300 -585
rect 3250 -635 3265 -615
rect 3285 -635 3300 -615
rect 3250 -665 3300 -635
rect 3250 -685 3265 -665
rect 3285 -685 3300 -665
rect 3250 -715 3300 -685
rect 3250 -735 3265 -715
rect 3285 -735 3300 -715
rect 3250 -765 3300 -735
rect 3250 -785 3265 -765
rect 3285 -785 3300 -765
rect 3250 -800 3300 -785
rect 3400 -800 3450 -100
rect 3550 -115 3600 -100
rect 3550 -135 3565 -115
rect 3585 -135 3600 -115
rect 3550 -165 3600 -135
rect 3550 -185 3565 -165
rect 3585 -185 3600 -165
rect 3550 -215 3600 -185
rect 3550 -235 3565 -215
rect 3585 -235 3600 -215
rect 3550 -265 3600 -235
rect 3550 -285 3565 -265
rect 3585 -285 3600 -265
rect 3550 -315 3600 -285
rect 3550 -335 3565 -315
rect 3585 -335 3600 -315
rect 3550 -365 3600 -335
rect 3550 -385 3565 -365
rect 3585 -385 3600 -365
rect 3550 -415 3600 -385
rect 3550 -435 3565 -415
rect 3585 -435 3600 -415
rect 3550 -465 3600 -435
rect 3550 -485 3565 -465
rect 3585 -485 3600 -465
rect 3550 -515 3600 -485
rect 3550 -535 3565 -515
rect 3585 -535 3600 -515
rect 3550 -565 3600 -535
rect 3550 -585 3565 -565
rect 3585 -585 3600 -565
rect 3550 -615 3600 -585
rect 3550 -635 3565 -615
rect 3585 -635 3600 -615
rect 3550 -665 3600 -635
rect 3550 -685 3565 -665
rect 3585 -685 3600 -665
rect 3550 -715 3600 -685
rect 3550 -735 3565 -715
rect 3585 -735 3600 -715
rect 3550 -765 3600 -735
rect 3550 -785 3565 -765
rect 3585 -785 3600 -765
rect 3550 -800 3600 -785
rect 3700 -115 3750 -100
rect 3700 -135 3715 -115
rect 3735 -135 3750 -115
rect 3700 -165 3750 -135
rect 3700 -185 3715 -165
rect 3735 -185 3750 -165
rect 3700 -215 3750 -185
rect 3700 -235 3715 -215
rect 3735 -235 3750 -215
rect 3700 -265 3750 -235
rect 3700 -285 3715 -265
rect 3735 -285 3750 -265
rect 3700 -315 3750 -285
rect 3700 -335 3715 -315
rect 3735 -335 3750 -315
rect 3700 -365 3750 -335
rect 3700 -385 3715 -365
rect 3735 -385 3750 -365
rect 3700 -415 3750 -385
rect 3700 -435 3715 -415
rect 3735 -435 3750 -415
rect 3700 -465 3750 -435
rect 3700 -485 3715 -465
rect 3735 -485 3750 -465
rect 3700 -515 3750 -485
rect 3700 -535 3715 -515
rect 3735 -535 3750 -515
rect 3700 -565 3750 -535
rect 3700 -585 3715 -565
rect 3735 -585 3750 -565
rect 3700 -615 3750 -585
rect 3700 -635 3715 -615
rect 3735 -635 3750 -615
rect 3700 -665 3750 -635
rect 3700 -685 3715 -665
rect 3735 -685 3750 -665
rect 3700 -715 3750 -685
rect 3700 -735 3715 -715
rect 3735 -735 3750 -715
rect 3700 -765 3750 -735
rect 3700 -785 3715 -765
rect 3735 -785 3750 -765
rect 3700 -800 3750 -785
rect 3850 -115 3900 -100
rect 3850 -135 3865 -115
rect 3885 -135 3900 -115
rect 3850 -165 3900 -135
rect 3850 -185 3865 -165
rect 3885 -185 3900 -165
rect 3850 -215 3900 -185
rect 3850 -235 3865 -215
rect 3885 -235 3900 -215
rect 3850 -265 3900 -235
rect 3850 -285 3865 -265
rect 3885 -285 3900 -265
rect 3850 -315 3900 -285
rect 3850 -335 3865 -315
rect 3885 -335 3900 -315
rect 3850 -365 3900 -335
rect 3850 -385 3865 -365
rect 3885 -385 3900 -365
rect 3850 -415 3900 -385
rect 3850 -435 3865 -415
rect 3885 -435 3900 -415
rect 3850 -465 3900 -435
rect 3850 -485 3865 -465
rect 3885 -485 3900 -465
rect 3850 -515 3900 -485
rect 3850 -535 3865 -515
rect 3885 -535 3900 -515
rect 3850 -565 3900 -535
rect 3850 -585 3865 -565
rect 3885 -585 3900 -565
rect 3850 -615 3900 -585
rect 3850 -635 3865 -615
rect 3885 -635 3900 -615
rect 3850 -665 3900 -635
rect 3850 -685 3865 -665
rect 3885 -685 3900 -665
rect 3850 -715 3900 -685
rect 3850 -735 3865 -715
rect 3885 -735 3900 -715
rect 3850 -765 3900 -735
rect 3850 -785 3865 -765
rect 3885 -785 3900 -765
rect 3850 -800 3900 -785
rect 4000 -115 4050 -100
rect 4000 -135 4015 -115
rect 4035 -135 4050 -115
rect 4000 -165 4050 -135
rect 4000 -185 4015 -165
rect 4035 -185 4050 -165
rect 4000 -215 4050 -185
rect 4000 -235 4015 -215
rect 4035 -235 4050 -215
rect 4000 -265 4050 -235
rect 4000 -285 4015 -265
rect 4035 -285 4050 -265
rect 4000 -315 4050 -285
rect 4000 -335 4015 -315
rect 4035 -335 4050 -315
rect 4000 -365 4050 -335
rect 4000 -385 4015 -365
rect 4035 -385 4050 -365
rect 4000 -415 4050 -385
rect 4000 -435 4015 -415
rect 4035 -435 4050 -415
rect 4000 -465 4050 -435
rect 4000 -485 4015 -465
rect 4035 -485 4050 -465
rect 4000 -515 4050 -485
rect 4000 -535 4015 -515
rect 4035 -535 4050 -515
rect 4000 -565 4050 -535
rect 4000 -585 4015 -565
rect 4035 -585 4050 -565
rect 4000 -615 4050 -585
rect 4000 -635 4015 -615
rect 4035 -635 4050 -615
rect 4000 -665 4050 -635
rect 4000 -685 4015 -665
rect 4035 -685 4050 -665
rect 4000 -715 4050 -685
rect 4000 -735 4015 -715
rect 4035 -735 4050 -715
rect 4000 -765 4050 -735
rect 4000 -785 4015 -765
rect 4035 -785 4050 -765
rect 4000 -800 4050 -785
rect 4150 -115 4200 -100
rect 4150 -135 4165 -115
rect 4185 -135 4200 -115
rect 4150 -165 4200 -135
rect 4150 -185 4165 -165
rect 4185 -185 4200 -165
rect 4150 -215 4200 -185
rect 4150 -235 4165 -215
rect 4185 -235 4200 -215
rect 4150 -265 4200 -235
rect 4150 -285 4165 -265
rect 4185 -285 4200 -265
rect 4150 -315 4200 -285
rect 4150 -335 4165 -315
rect 4185 -335 4200 -315
rect 4150 -365 4200 -335
rect 4150 -385 4165 -365
rect 4185 -385 4200 -365
rect 4150 -415 4200 -385
rect 4150 -435 4165 -415
rect 4185 -435 4200 -415
rect 4150 -465 4200 -435
rect 4150 -485 4165 -465
rect 4185 -485 4200 -465
rect 4150 -515 4200 -485
rect 4150 -535 4165 -515
rect 4185 -535 4200 -515
rect 4150 -565 4200 -535
rect 4150 -585 4165 -565
rect 4185 -585 4200 -565
rect 4150 -615 4200 -585
rect 4150 -635 4165 -615
rect 4185 -635 4200 -615
rect 4150 -665 4200 -635
rect 4150 -685 4165 -665
rect 4185 -685 4200 -665
rect 4150 -715 4200 -685
rect 4150 -735 4165 -715
rect 4185 -735 4200 -715
rect 4150 -765 4200 -735
rect 4150 -785 4165 -765
rect 4185 -785 4200 -765
rect 4150 -800 4200 -785
rect 4300 -115 4350 -100
rect 4300 -135 4315 -115
rect 4335 -135 4350 -115
rect 4300 -165 4350 -135
rect 4300 -185 4315 -165
rect 4335 -185 4350 -165
rect 4300 -215 4350 -185
rect 4300 -235 4315 -215
rect 4335 -235 4350 -215
rect 4300 -265 4350 -235
rect 4300 -285 4315 -265
rect 4335 -285 4350 -265
rect 4300 -315 4350 -285
rect 4300 -335 4315 -315
rect 4335 -335 4350 -315
rect 4300 -365 4350 -335
rect 4300 -385 4315 -365
rect 4335 -385 4350 -365
rect 4300 -415 4350 -385
rect 4300 -435 4315 -415
rect 4335 -435 4350 -415
rect 4300 -465 4350 -435
rect 4300 -485 4315 -465
rect 4335 -485 4350 -465
rect 4300 -515 4350 -485
rect 4300 -535 4315 -515
rect 4335 -535 4350 -515
rect 4300 -565 4350 -535
rect 4300 -585 4315 -565
rect 4335 -585 4350 -565
rect 4300 -615 4350 -585
rect 4300 -635 4315 -615
rect 4335 -635 4350 -615
rect 4300 -665 4350 -635
rect 4300 -685 4315 -665
rect 4335 -685 4350 -665
rect 4300 -715 4350 -685
rect 4300 -735 4315 -715
rect 4335 -735 4350 -715
rect 4300 -765 4350 -735
rect 4300 -785 4315 -765
rect 4335 -785 4350 -765
rect 4300 -800 4350 -785
rect 4450 -115 4500 -100
rect 4450 -135 4465 -115
rect 4485 -135 4500 -115
rect 4450 -165 4500 -135
rect 4450 -185 4465 -165
rect 4485 -185 4500 -165
rect 4450 -215 4500 -185
rect 4450 -235 4465 -215
rect 4485 -235 4500 -215
rect 4450 -265 4500 -235
rect 4450 -285 4465 -265
rect 4485 -285 4500 -265
rect 4450 -315 4500 -285
rect 4450 -335 4465 -315
rect 4485 -335 4500 -315
rect 4450 -365 4500 -335
rect 4450 -385 4465 -365
rect 4485 -385 4500 -365
rect 4450 -415 4500 -385
rect 4450 -435 4465 -415
rect 4485 -435 4500 -415
rect 4450 -465 4500 -435
rect 4450 -485 4465 -465
rect 4485 -485 4500 -465
rect 4450 -515 4500 -485
rect 4450 -535 4465 -515
rect 4485 -535 4500 -515
rect 4450 -565 4500 -535
rect 4450 -585 4465 -565
rect 4485 -585 4500 -565
rect 4450 -615 4500 -585
rect 4450 -635 4465 -615
rect 4485 -635 4500 -615
rect 4450 -665 4500 -635
rect 4450 -685 4465 -665
rect 4485 -685 4500 -665
rect 4450 -715 4500 -685
rect 4450 -735 4465 -715
rect 4485 -735 4500 -715
rect 4450 -765 4500 -735
rect 4450 -785 4465 -765
rect 4485 -785 4500 -765
rect 4450 -800 4500 -785
rect 4600 -115 4650 -100
rect 4600 -135 4615 -115
rect 4635 -135 4650 -115
rect 4600 -165 4650 -135
rect 4600 -185 4615 -165
rect 4635 -185 4650 -165
rect 4600 -215 4650 -185
rect 4600 -235 4615 -215
rect 4635 -235 4650 -215
rect 4600 -265 4650 -235
rect 4600 -285 4615 -265
rect 4635 -285 4650 -265
rect 4600 -315 4650 -285
rect 4600 -335 4615 -315
rect 4635 -335 4650 -315
rect 4600 -365 4650 -335
rect 4600 -385 4615 -365
rect 4635 -385 4650 -365
rect 4600 -415 4650 -385
rect 4600 -435 4615 -415
rect 4635 -435 4650 -415
rect 4600 -465 4650 -435
rect 4600 -485 4615 -465
rect 4635 -485 4650 -465
rect 4600 -515 4650 -485
rect 4600 -535 4615 -515
rect 4635 -535 4650 -515
rect 4600 -565 4650 -535
rect 4600 -585 4615 -565
rect 4635 -585 4650 -565
rect 4600 -615 4650 -585
rect 4600 -635 4615 -615
rect 4635 -635 4650 -615
rect 4600 -665 4650 -635
rect 4600 -685 4615 -665
rect 4635 -685 4650 -665
rect 4600 -715 4650 -685
rect 4600 -735 4615 -715
rect 4635 -735 4650 -715
rect 4600 -765 4650 -735
rect 4600 -785 4615 -765
rect 4635 -785 4650 -765
rect 4600 -800 4650 -785
rect 4750 -115 4800 -100
rect 4750 -135 4765 -115
rect 4785 -135 4800 -115
rect 4750 -165 4800 -135
rect 4750 -185 4765 -165
rect 4785 -185 4800 -165
rect 4750 -215 4800 -185
rect 4750 -235 4765 -215
rect 4785 -235 4800 -215
rect 4750 -265 4800 -235
rect 4750 -285 4765 -265
rect 4785 -285 4800 -265
rect 4750 -315 4800 -285
rect 4750 -335 4765 -315
rect 4785 -335 4800 -315
rect 4750 -365 4800 -335
rect 4750 -385 4765 -365
rect 4785 -385 4800 -365
rect 4750 -415 4800 -385
rect 4750 -435 4765 -415
rect 4785 -435 4800 -415
rect 4750 -465 4800 -435
rect 4750 -485 4765 -465
rect 4785 -485 4800 -465
rect 4750 -515 4800 -485
rect 4750 -535 4765 -515
rect 4785 -535 4800 -515
rect 4750 -565 4800 -535
rect 4750 -585 4765 -565
rect 4785 -585 4800 -565
rect 4750 -615 4800 -585
rect 4750 -635 4765 -615
rect 4785 -635 4800 -615
rect 4750 -665 4800 -635
rect 4750 -685 4765 -665
rect 4785 -685 4800 -665
rect 4750 -715 4800 -685
rect 4750 -735 4765 -715
rect 4785 -735 4800 -715
rect 4750 -765 4800 -735
rect 4750 -785 4765 -765
rect 4785 -785 4800 -765
rect 4750 -800 4800 -785
rect 4900 -800 4950 -100
rect 5050 -115 5100 -100
rect 5050 -135 5065 -115
rect 5085 -135 5100 -115
rect 5050 -165 5100 -135
rect 5050 -185 5065 -165
rect 5085 -185 5100 -165
rect 5050 -215 5100 -185
rect 5050 -235 5065 -215
rect 5085 -235 5100 -215
rect 5050 -265 5100 -235
rect 5050 -285 5065 -265
rect 5085 -285 5100 -265
rect 5050 -315 5100 -285
rect 5050 -335 5065 -315
rect 5085 -335 5100 -315
rect 5050 -365 5100 -335
rect 5050 -385 5065 -365
rect 5085 -385 5100 -365
rect 5050 -415 5100 -385
rect 5050 -435 5065 -415
rect 5085 -435 5100 -415
rect 5050 -465 5100 -435
rect 5050 -485 5065 -465
rect 5085 -485 5100 -465
rect 5050 -515 5100 -485
rect 5050 -535 5065 -515
rect 5085 -535 5100 -515
rect 5050 -565 5100 -535
rect 5050 -585 5065 -565
rect 5085 -585 5100 -565
rect 5050 -615 5100 -585
rect 5050 -635 5065 -615
rect 5085 -635 5100 -615
rect 5050 -665 5100 -635
rect 5050 -685 5065 -665
rect 5085 -685 5100 -665
rect 5050 -715 5100 -685
rect 5050 -735 5065 -715
rect 5085 -735 5100 -715
rect 5050 -765 5100 -735
rect 5050 -785 5065 -765
rect 5085 -785 5100 -765
rect 5050 -800 5100 -785
rect 5200 -800 5250 -100
rect 5350 -115 5400 -100
rect 5350 -135 5365 -115
rect 5385 -135 5400 -115
rect 5350 -165 5400 -135
rect 5350 -185 5365 -165
rect 5385 -185 5400 -165
rect 5350 -215 5400 -185
rect 5350 -235 5365 -215
rect 5385 -235 5400 -215
rect 5350 -265 5400 -235
rect 5350 -285 5365 -265
rect 5385 -285 5400 -265
rect 5350 -315 5400 -285
rect 5350 -335 5365 -315
rect 5385 -335 5400 -315
rect 5350 -365 5400 -335
rect 5350 -385 5365 -365
rect 5385 -385 5400 -365
rect 5350 -415 5400 -385
rect 5350 -435 5365 -415
rect 5385 -435 5400 -415
rect 5350 -465 5400 -435
rect 5350 -485 5365 -465
rect 5385 -485 5400 -465
rect 5350 -515 5400 -485
rect 5350 -535 5365 -515
rect 5385 -535 5400 -515
rect 5350 -565 5400 -535
rect 5350 -585 5365 -565
rect 5385 -585 5400 -565
rect 5350 -615 5400 -585
rect 5350 -635 5365 -615
rect 5385 -635 5400 -615
rect 5350 -665 5400 -635
rect 5350 -685 5365 -665
rect 5385 -685 5400 -665
rect 5350 -715 5400 -685
rect 5350 -735 5365 -715
rect 5385 -735 5400 -715
rect 5350 -765 5400 -735
rect 5350 -785 5365 -765
rect 5385 -785 5400 -765
rect 5350 -800 5400 -785
rect 5500 -800 5550 -100
rect 5650 -115 5700 -100
rect 5650 -135 5665 -115
rect 5685 -135 5700 -115
rect 5650 -165 5700 -135
rect 5650 -185 5665 -165
rect 5685 -185 5700 -165
rect 5650 -215 5700 -185
rect 5650 -235 5665 -215
rect 5685 -235 5700 -215
rect 5650 -265 5700 -235
rect 5650 -285 5665 -265
rect 5685 -285 5700 -265
rect 5650 -315 5700 -285
rect 5650 -335 5665 -315
rect 5685 -335 5700 -315
rect 5650 -365 5700 -335
rect 5650 -385 5665 -365
rect 5685 -385 5700 -365
rect 5650 -415 5700 -385
rect 5650 -435 5665 -415
rect 5685 -435 5700 -415
rect 5650 -465 5700 -435
rect 5650 -485 5665 -465
rect 5685 -485 5700 -465
rect 5650 -515 5700 -485
rect 5650 -535 5665 -515
rect 5685 -535 5700 -515
rect 5650 -565 5700 -535
rect 5650 -585 5665 -565
rect 5685 -585 5700 -565
rect 5650 -615 5700 -585
rect 5650 -635 5665 -615
rect 5685 -635 5700 -615
rect 5650 -665 5700 -635
rect 5650 -685 5665 -665
rect 5685 -685 5700 -665
rect 5650 -715 5700 -685
rect 5650 -735 5665 -715
rect 5685 -735 5700 -715
rect 5650 -765 5700 -735
rect 5650 -785 5665 -765
rect 5685 -785 5700 -765
rect 5650 -800 5700 -785
rect 5800 -800 5850 -100
rect 5950 -115 6000 -100
rect 5950 -135 5965 -115
rect 5985 -135 6000 -115
rect 5950 -165 6000 -135
rect 5950 -185 5965 -165
rect 5985 -185 6000 -165
rect 5950 -215 6000 -185
rect 5950 -235 5965 -215
rect 5985 -235 6000 -215
rect 5950 -265 6000 -235
rect 5950 -285 5965 -265
rect 5985 -285 6000 -265
rect 5950 -315 6000 -285
rect 5950 -335 5965 -315
rect 5985 -335 6000 -315
rect 5950 -365 6000 -335
rect 5950 -385 5965 -365
rect 5985 -385 6000 -365
rect 5950 -415 6000 -385
rect 5950 -435 5965 -415
rect 5985 -435 6000 -415
rect 5950 -465 6000 -435
rect 5950 -485 5965 -465
rect 5985 -485 6000 -465
rect 5950 -515 6000 -485
rect 5950 -535 5965 -515
rect 5985 -535 6000 -515
rect 5950 -565 6000 -535
rect 5950 -585 5965 -565
rect 5985 -585 6000 -565
rect 5950 -615 6000 -585
rect 5950 -635 5965 -615
rect 5985 -635 6000 -615
rect 5950 -665 6000 -635
rect 5950 -685 5965 -665
rect 5985 -685 6000 -665
rect 5950 -715 6000 -685
rect 5950 -735 5965 -715
rect 5985 -735 6000 -715
rect 5950 -765 6000 -735
rect 5950 -785 5965 -765
rect 5985 -785 6000 -765
rect 5950 -800 6000 -785
rect 6100 -800 6150 -100
rect 6250 -115 6300 -100
rect 6250 -135 6265 -115
rect 6285 -135 6300 -115
rect 6250 -165 6300 -135
rect 6250 -185 6265 -165
rect 6285 -185 6300 -165
rect 6250 -215 6300 -185
rect 6250 -235 6265 -215
rect 6285 -235 6300 -215
rect 6250 -265 6300 -235
rect 6250 -285 6265 -265
rect 6285 -285 6300 -265
rect 6250 -315 6300 -285
rect 6250 -335 6265 -315
rect 6285 -335 6300 -315
rect 6250 -365 6300 -335
rect 6250 -385 6265 -365
rect 6285 -385 6300 -365
rect 6250 -415 6300 -385
rect 6250 -435 6265 -415
rect 6285 -435 6300 -415
rect 6250 -465 6300 -435
rect 6250 -485 6265 -465
rect 6285 -485 6300 -465
rect 6250 -515 6300 -485
rect 6250 -535 6265 -515
rect 6285 -535 6300 -515
rect 6250 -565 6300 -535
rect 6250 -585 6265 -565
rect 6285 -585 6300 -565
rect 6250 -615 6300 -585
rect 6250 -635 6265 -615
rect 6285 -635 6300 -615
rect 6250 -665 6300 -635
rect 6250 -685 6265 -665
rect 6285 -685 6300 -665
rect 6250 -715 6300 -685
rect 6250 -735 6265 -715
rect 6285 -735 6300 -715
rect 6250 -765 6300 -735
rect 6250 -785 6265 -765
rect 6285 -785 6300 -765
rect 6250 -800 6300 -785
rect 6400 -800 6450 -100
rect 6550 -115 6600 -100
rect 6550 -135 6565 -115
rect 6585 -135 6600 -115
rect 6550 -165 6600 -135
rect 6550 -185 6565 -165
rect 6585 -185 6600 -165
rect 6550 -215 6600 -185
rect 6550 -235 6565 -215
rect 6585 -235 6600 -215
rect 6550 -265 6600 -235
rect 6550 -285 6565 -265
rect 6585 -285 6600 -265
rect 6550 -315 6600 -285
rect 6550 -335 6565 -315
rect 6585 -335 6600 -315
rect 6550 -365 6600 -335
rect 6550 -385 6565 -365
rect 6585 -385 6600 -365
rect 6550 -415 6600 -385
rect 6550 -435 6565 -415
rect 6585 -435 6600 -415
rect 6550 -465 6600 -435
rect 6550 -485 6565 -465
rect 6585 -485 6600 -465
rect 6550 -515 6600 -485
rect 6550 -535 6565 -515
rect 6585 -535 6600 -515
rect 6550 -565 6600 -535
rect 6550 -585 6565 -565
rect 6585 -585 6600 -565
rect 6550 -615 6600 -585
rect 6550 -635 6565 -615
rect 6585 -635 6600 -615
rect 6550 -665 6600 -635
rect 6550 -685 6565 -665
rect 6585 -685 6600 -665
rect 6550 -715 6600 -685
rect 6550 -735 6565 -715
rect 6585 -735 6600 -715
rect 6550 -765 6600 -735
rect 6550 -785 6565 -765
rect 6585 -785 6600 -765
rect 6550 -800 6600 -785
rect 6700 -800 6750 -100
rect 6850 -115 6900 -100
rect 6850 -135 6865 -115
rect 6885 -135 6900 -115
rect 6850 -165 6900 -135
rect 6850 -185 6865 -165
rect 6885 -185 6900 -165
rect 6850 -215 6900 -185
rect 6850 -235 6865 -215
rect 6885 -235 6900 -215
rect 6850 -265 6900 -235
rect 6850 -285 6865 -265
rect 6885 -285 6900 -265
rect 6850 -315 6900 -285
rect 6850 -335 6865 -315
rect 6885 -335 6900 -315
rect 6850 -365 6900 -335
rect 6850 -385 6865 -365
rect 6885 -385 6900 -365
rect 6850 -415 6900 -385
rect 6850 -435 6865 -415
rect 6885 -435 6900 -415
rect 6850 -465 6900 -435
rect 6850 -485 6865 -465
rect 6885 -485 6900 -465
rect 6850 -515 6900 -485
rect 6850 -535 6865 -515
rect 6885 -535 6900 -515
rect 6850 -565 6900 -535
rect 6850 -585 6865 -565
rect 6885 -585 6900 -565
rect 6850 -615 6900 -585
rect 6850 -635 6865 -615
rect 6885 -635 6900 -615
rect 6850 -665 6900 -635
rect 6850 -685 6865 -665
rect 6885 -685 6900 -665
rect 6850 -715 6900 -685
rect 6850 -735 6865 -715
rect 6885 -735 6900 -715
rect 6850 -765 6900 -735
rect 6850 -785 6865 -765
rect 6885 -785 6900 -765
rect 6850 -800 6900 -785
rect 7000 -800 7050 -100
rect 7150 -115 7200 -100
rect 7150 -135 7165 -115
rect 7185 -135 7200 -115
rect 7150 -165 7200 -135
rect 7150 -185 7165 -165
rect 7185 -185 7200 -165
rect 7150 -215 7200 -185
rect 7150 -235 7165 -215
rect 7185 -235 7200 -215
rect 7150 -265 7200 -235
rect 7150 -285 7165 -265
rect 7185 -285 7200 -265
rect 7150 -315 7200 -285
rect 7150 -335 7165 -315
rect 7185 -335 7200 -315
rect 7150 -365 7200 -335
rect 7150 -385 7165 -365
rect 7185 -385 7200 -365
rect 7150 -415 7200 -385
rect 7150 -435 7165 -415
rect 7185 -435 7200 -415
rect 7150 -465 7200 -435
rect 7150 -485 7165 -465
rect 7185 -485 7200 -465
rect 7150 -515 7200 -485
rect 7150 -535 7165 -515
rect 7185 -535 7200 -515
rect 7150 -565 7200 -535
rect 7150 -585 7165 -565
rect 7185 -585 7200 -565
rect 7150 -615 7200 -585
rect 7150 -635 7165 -615
rect 7185 -635 7200 -615
rect 7150 -665 7200 -635
rect 7150 -685 7165 -665
rect 7185 -685 7200 -665
rect 7150 -715 7200 -685
rect 7150 -735 7165 -715
rect 7185 -735 7200 -715
rect 7150 -765 7200 -735
rect 7150 -785 7165 -765
rect 7185 -785 7200 -765
rect 7150 -800 7200 -785
rect 7300 -800 7350 -100
rect 7450 -800 7500 -100
rect 7600 -800 7650 -100
rect 7750 -800 7800 -100
rect 7900 -800 7950 -100
rect 8050 -800 8100 -100
rect 8200 -800 8250 -100
rect 8350 -115 8400 -100
rect 8350 -135 8365 -115
rect 8385 -135 8400 -115
rect 8350 -165 8400 -135
rect 8350 -185 8365 -165
rect 8385 -185 8400 -165
rect 8350 -215 8400 -185
rect 8350 -235 8365 -215
rect 8385 -235 8400 -215
rect 8350 -265 8400 -235
rect 8350 -285 8365 -265
rect 8385 -285 8400 -265
rect 8350 -315 8400 -285
rect 8350 -335 8365 -315
rect 8385 -335 8400 -315
rect 8350 -365 8400 -335
rect 8350 -385 8365 -365
rect 8385 -385 8400 -365
rect 8350 -415 8400 -385
rect 8350 -435 8365 -415
rect 8385 -435 8400 -415
rect 8350 -465 8400 -435
rect 8350 -485 8365 -465
rect 8385 -485 8400 -465
rect 8350 -515 8400 -485
rect 8350 -535 8365 -515
rect 8385 -535 8400 -515
rect 8350 -565 8400 -535
rect 8350 -585 8365 -565
rect 8385 -585 8400 -565
rect 8350 -615 8400 -585
rect 8350 -635 8365 -615
rect 8385 -635 8400 -615
rect 8350 -665 8400 -635
rect 8350 -685 8365 -665
rect 8385 -685 8400 -665
rect 8350 -715 8400 -685
rect 8350 -735 8365 -715
rect 8385 -735 8400 -715
rect 8350 -765 8400 -735
rect 8350 -785 8365 -765
rect 8385 -785 8400 -765
rect 8350 -800 8400 -785
rect 8500 -800 8550 -100
rect 8650 -800 8700 -100
rect 8800 -800 8850 -100
rect 8950 -800 9000 -100
rect 9100 -800 9150 -100
rect 9250 -800 9300 -100
rect 9400 -800 9450 -100
rect 9550 -115 9600 -100
rect 9550 -135 9565 -115
rect 9585 -135 9600 -115
rect 9550 -165 9600 -135
rect 9550 -185 9565 -165
rect 9585 -185 9600 -165
rect 9550 -215 9600 -185
rect 9550 -235 9565 -215
rect 9585 -235 9600 -215
rect 9550 -265 9600 -235
rect 9550 -285 9565 -265
rect 9585 -285 9600 -265
rect 9550 -315 9600 -285
rect 9550 -335 9565 -315
rect 9585 -335 9600 -315
rect 9550 -365 9600 -335
rect 9550 -385 9565 -365
rect 9585 -385 9600 -365
rect 9550 -415 9600 -385
rect 9550 -435 9565 -415
rect 9585 -435 9600 -415
rect 9550 -465 9600 -435
rect 9550 -485 9565 -465
rect 9585 -485 9600 -465
rect 9550 -515 9600 -485
rect 9550 -535 9565 -515
rect 9585 -535 9600 -515
rect 9550 -565 9600 -535
rect 9550 -585 9565 -565
rect 9585 -585 9600 -565
rect 9550 -615 9600 -585
rect 9550 -635 9565 -615
rect 9585 -635 9600 -615
rect 9550 -665 9600 -635
rect 9550 -685 9565 -665
rect 9585 -685 9600 -665
rect 9550 -715 9600 -685
rect 9550 -735 9565 -715
rect 9585 -735 9600 -715
rect 9550 -765 9600 -735
rect 9550 -785 9565 -765
rect 9585 -785 9600 -765
rect 9550 -800 9600 -785
rect 9700 -800 9750 -100
rect 9850 -800 9900 -100
rect 10000 -800 10050 -100
rect 10150 -800 10200 -100
rect 10300 -800 10350 -100
rect 10450 -800 10500 -100
rect 10600 -800 10650 -100
rect 10750 -115 10800 -100
rect 10750 -135 10765 -115
rect 10785 -135 10800 -115
rect 10750 -165 10800 -135
rect 10750 -185 10765 -165
rect 10785 -185 10800 -165
rect 10750 -215 10800 -185
rect 10750 -235 10765 -215
rect 10785 -235 10800 -215
rect 10750 -265 10800 -235
rect 10750 -285 10765 -265
rect 10785 -285 10800 -265
rect 10750 -315 10800 -285
rect 10750 -335 10765 -315
rect 10785 -335 10800 -315
rect 10750 -365 10800 -335
rect 10750 -385 10765 -365
rect 10785 -385 10800 -365
rect 10750 -415 10800 -385
rect 10750 -435 10765 -415
rect 10785 -435 10800 -415
rect 10750 -465 10800 -435
rect 10750 -485 10765 -465
rect 10785 -485 10800 -465
rect 10750 -515 10800 -485
rect 10750 -535 10765 -515
rect 10785 -535 10800 -515
rect 10750 -565 10800 -535
rect 10750 -585 10765 -565
rect 10785 -585 10800 -565
rect 10750 -615 10800 -585
rect 10750 -635 10765 -615
rect 10785 -635 10800 -615
rect 10750 -665 10800 -635
rect 10750 -685 10765 -665
rect 10785 -685 10800 -665
rect 10750 -715 10800 -685
rect 10750 -735 10765 -715
rect 10785 -735 10800 -715
rect 10750 -765 10800 -735
rect 10750 -785 10765 -765
rect 10785 -785 10800 -765
rect 10750 -800 10800 -785
rect 10900 -800 10950 -100
rect 11050 -800 11100 -100
rect 11200 -800 11250 -100
rect 11350 -800 11400 -100
rect 11500 -800 11550 -100
rect 11650 -800 11700 -100
rect 11800 -800 11850 -100
rect 11950 -115 12000 -100
rect 11950 -135 11965 -115
rect 11985 -135 12000 -115
rect 11950 -165 12000 -135
rect 11950 -185 11965 -165
rect 11985 -185 12000 -165
rect 11950 -215 12000 -185
rect 11950 -235 11965 -215
rect 11985 -235 12000 -215
rect 11950 -265 12000 -235
rect 11950 -285 11965 -265
rect 11985 -285 12000 -265
rect 11950 -315 12000 -285
rect 11950 -335 11965 -315
rect 11985 -335 12000 -315
rect 11950 -365 12000 -335
rect 11950 -385 11965 -365
rect 11985 -385 12000 -365
rect 11950 -415 12000 -385
rect 11950 -435 11965 -415
rect 11985 -435 12000 -415
rect 11950 -465 12000 -435
rect 11950 -485 11965 -465
rect 11985 -485 12000 -465
rect 11950 -515 12000 -485
rect 11950 -535 11965 -515
rect 11985 -535 12000 -515
rect 11950 -565 12000 -535
rect 11950 -585 11965 -565
rect 11985 -585 12000 -565
rect 11950 -615 12000 -585
rect 11950 -635 11965 -615
rect 11985 -635 12000 -615
rect 11950 -665 12000 -635
rect 11950 -685 11965 -665
rect 11985 -685 12000 -665
rect 11950 -715 12000 -685
rect 11950 -735 11965 -715
rect 11985 -735 12000 -715
rect 11950 -765 12000 -735
rect 11950 -785 11965 -765
rect 11985 -785 12000 -765
rect 11950 -800 12000 -785
rect 12100 -800 12150 -100
rect 12250 -115 12300 -100
rect 12250 -135 12265 -115
rect 12285 -135 12300 -115
rect 12250 -165 12300 -135
rect 12250 -185 12265 -165
rect 12285 -185 12300 -165
rect 12250 -215 12300 -185
rect 12250 -235 12265 -215
rect 12285 -235 12300 -215
rect 12250 -265 12300 -235
rect 12250 -285 12265 -265
rect 12285 -285 12300 -265
rect 12250 -315 12300 -285
rect 12250 -335 12265 -315
rect 12285 -335 12300 -315
rect 12250 -365 12300 -335
rect 12250 -385 12265 -365
rect 12285 -385 12300 -365
rect 12250 -415 12300 -385
rect 12250 -435 12265 -415
rect 12285 -435 12300 -415
rect 12250 -465 12300 -435
rect 12250 -485 12265 -465
rect 12285 -485 12300 -465
rect 12250 -515 12300 -485
rect 12250 -535 12265 -515
rect 12285 -535 12300 -515
rect 12250 -565 12300 -535
rect 12250 -585 12265 -565
rect 12285 -585 12300 -565
rect 12250 -615 12300 -585
rect 12250 -635 12265 -615
rect 12285 -635 12300 -615
rect 12250 -665 12300 -635
rect 12250 -685 12265 -665
rect 12285 -685 12300 -665
rect 12250 -715 12300 -685
rect 12250 -735 12265 -715
rect 12285 -735 12300 -715
rect 12250 -765 12300 -735
rect 12250 -785 12265 -765
rect 12285 -785 12300 -765
rect 12250 -800 12300 -785
rect 12400 -800 12450 -100
rect 12550 -115 12600 -100
rect 12550 -135 12565 -115
rect 12585 -135 12600 -115
rect 12550 -165 12600 -135
rect 12550 -185 12565 -165
rect 12585 -185 12600 -165
rect 12550 -215 12600 -185
rect 12550 -235 12565 -215
rect 12585 -235 12600 -215
rect 12550 -265 12600 -235
rect 12550 -285 12565 -265
rect 12585 -285 12600 -265
rect 12550 -315 12600 -285
rect 12550 -335 12565 -315
rect 12585 -335 12600 -315
rect 12550 -365 12600 -335
rect 12550 -385 12565 -365
rect 12585 -385 12600 -365
rect 12550 -415 12600 -385
rect 12550 -435 12565 -415
rect 12585 -435 12600 -415
rect 12550 -465 12600 -435
rect 12550 -485 12565 -465
rect 12585 -485 12600 -465
rect 12550 -515 12600 -485
rect 12550 -535 12565 -515
rect 12585 -535 12600 -515
rect 12550 -565 12600 -535
rect 12550 -585 12565 -565
rect 12585 -585 12600 -565
rect 12550 -615 12600 -585
rect 12550 -635 12565 -615
rect 12585 -635 12600 -615
rect 12550 -665 12600 -635
rect 12550 -685 12565 -665
rect 12585 -685 12600 -665
rect 12550 -715 12600 -685
rect 12550 -735 12565 -715
rect 12585 -735 12600 -715
rect 12550 -765 12600 -735
rect 12550 -785 12565 -765
rect 12585 -785 12600 -765
rect 12550 -800 12600 -785
rect 12700 -800 12750 -100
rect 12850 -115 12900 -100
rect 12850 -135 12865 -115
rect 12885 -135 12900 -115
rect 12850 -165 12900 -135
rect 12850 -185 12865 -165
rect 12885 -185 12900 -165
rect 12850 -215 12900 -185
rect 12850 -235 12865 -215
rect 12885 -235 12900 -215
rect 12850 -265 12900 -235
rect 12850 -285 12865 -265
rect 12885 -285 12900 -265
rect 12850 -315 12900 -285
rect 12850 -335 12865 -315
rect 12885 -335 12900 -315
rect 12850 -365 12900 -335
rect 12850 -385 12865 -365
rect 12885 -385 12900 -365
rect 12850 -415 12900 -385
rect 12850 -435 12865 -415
rect 12885 -435 12900 -415
rect 12850 -465 12900 -435
rect 12850 -485 12865 -465
rect 12885 -485 12900 -465
rect 12850 -515 12900 -485
rect 12850 -535 12865 -515
rect 12885 -535 12900 -515
rect 12850 -565 12900 -535
rect 12850 -585 12865 -565
rect 12885 -585 12900 -565
rect 12850 -615 12900 -585
rect 12850 -635 12865 -615
rect 12885 -635 12900 -615
rect 12850 -665 12900 -635
rect 12850 -685 12865 -665
rect 12885 -685 12900 -665
rect 12850 -715 12900 -685
rect 12850 -735 12865 -715
rect 12885 -735 12900 -715
rect 12850 -765 12900 -735
rect 12850 -785 12865 -765
rect 12885 -785 12900 -765
rect 12850 -800 12900 -785
rect 13000 -800 13050 -100
rect 13150 -115 13200 -100
rect 13150 -135 13165 -115
rect 13185 -135 13200 -115
rect 13150 -165 13200 -135
rect 13150 -185 13165 -165
rect 13185 -185 13200 -165
rect 13150 -215 13200 -185
rect 13150 -235 13165 -215
rect 13185 -235 13200 -215
rect 13150 -265 13200 -235
rect 13150 -285 13165 -265
rect 13185 -285 13200 -265
rect 13150 -315 13200 -285
rect 13150 -335 13165 -315
rect 13185 -335 13200 -315
rect 13150 -365 13200 -335
rect 13150 -385 13165 -365
rect 13185 -385 13200 -365
rect 13150 -415 13200 -385
rect 13150 -435 13165 -415
rect 13185 -435 13200 -415
rect 13150 -465 13200 -435
rect 13150 -485 13165 -465
rect 13185 -485 13200 -465
rect 13150 -515 13200 -485
rect 13150 -535 13165 -515
rect 13185 -535 13200 -515
rect 13150 -565 13200 -535
rect 13150 -585 13165 -565
rect 13185 -585 13200 -565
rect 13150 -615 13200 -585
rect 13150 -635 13165 -615
rect 13185 -635 13200 -615
rect 13150 -665 13200 -635
rect 13150 -685 13165 -665
rect 13185 -685 13200 -665
rect 13150 -715 13200 -685
rect 13150 -735 13165 -715
rect 13185 -735 13200 -715
rect 13150 -765 13200 -735
rect 13150 -785 13165 -765
rect 13185 -785 13200 -765
rect 13150 -800 13200 -785
rect 13300 -800 13350 -100
rect 13450 -115 13500 -100
rect 13450 -135 13465 -115
rect 13485 -135 13500 -115
rect 13450 -165 13500 -135
rect 13450 -185 13465 -165
rect 13485 -185 13500 -165
rect 13450 -215 13500 -185
rect 13450 -235 13465 -215
rect 13485 -235 13500 -215
rect 13450 -265 13500 -235
rect 13450 -285 13465 -265
rect 13485 -285 13500 -265
rect 13450 -315 13500 -285
rect 13450 -335 13465 -315
rect 13485 -335 13500 -315
rect 13450 -365 13500 -335
rect 13450 -385 13465 -365
rect 13485 -385 13500 -365
rect 13450 -415 13500 -385
rect 13450 -435 13465 -415
rect 13485 -435 13500 -415
rect 13450 -465 13500 -435
rect 13450 -485 13465 -465
rect 13485 -485 13500 -465
rect 13450 -515 13500 -485
rect 13450 -535 13465 -515
rect 13485 -535 13500 -515
rect 13450 -565 13500 -535
rect 13450 -585 13465 -565
rect 13485 -585 13500 -565
rect 13450 -615 13500 -585
rect 13450 -635 13465 -615
rect 13485 -635 13500 -615
rect 13450 -665 13500 -635
rect 13450 -685 13465 -665
rect 13485 -685 13500 -665
rect 13450 -715 13500 -685
rect 13450 -735 13465 -715
rect 13485 -735 13500 -715
rect 13450 -765 13500 -735
rect 13450 -785 13465 -765
rect 13485 -785 13500 -765
rect 13450 -800 13500 -785
rect 13600 -800 13650 -100
rect 13750 -115 13800 -100
rect 13750 -135 13765 -115
rect 13785 -135 13800 -115
rect 13750 -165 13800 -135
rect 13750 -185 13765 -165
rect 13785 -185 13800 -165
rect 13750 -215 13800 -185
rect 13750 -235 13765 -215
rect 13785 -235 13800 -215
rect 13750 -265 13800 -235
rect 13750 -285 13765 -265
rect 13785 -285 13800 -265
rect 13750 -315 13800 -285
rect 13750 -335 13765 -315
rect 13785 -335 13800 -315
rect 13750 -365 13800 -335
rect 13750 -385 13765 -365
rect 13785 -385 13800 -365
rect 13750 -415 13800 -385
rect 13750 -435 13765 -415
rect 13785 -435 13800 -415
rect 13750 -465 13800 -435
rect 13750 -485 13765 -465
rect 13785 -485 13800 -465
rect 13750 -515 13800 -485
rect 13750 -535 13765 -515
rect 13785 -535 13800 -515
rect 13750 -565 13800 -535
rect 13750 -585 13765 -565
rect 13785 -585 13800 -565
rect 13750 -615 13800 -585
rect 13750 -635 13765 -615
rect 13785 -635 13800 -615
rect 13750 -665 13800 -635
rect 13750 -685 13765 -665
rect 13785 -685 13800 -665
rect 13750 -715 13800 -685
rect 13750 -735 13765 -715
rect 13785 -735 13800 -715
rect 13750 -765 13800 -735
rect 13750 -785 13765 -765
rect 13785 -785 13800 -765
rect 13750 -800 13800 -785
rect 13900 -800 13950 -100
rect 14050 -115 14100 -100
rect 14050 -135 14065 -115
rect 14085 -135 14100 -115
rect 14050 -165 14100 -135
rect 14050 -185 14065 -165
rect 14085 -185 14100 -165
rect 14050 -215 14100 -185
rect 14050 -235 14065 -215
rect 14085 -235 14100 -215
rect 14050 -265 14100 -235
rect 14050 -285 14065 -265
rect 14085 -285 14100 -265
rect 14050 -315 14100 -285
rect 14050 -335 14065 -315
rect 14085 -335 14100 -315
rect 14050 -365 14100 -335
rect 14050 -385 14065 -365
rect 14085 -385 14100 -365
rect 14050 -415 14100 -385
rect 14050 -435 14065 -415
rect 14085 -435 14100 -415
rect 14050 -465 14100 -435
rect 14050 -485 14065 -465
rect 14085 -485 14100 -465
rect 14050 -515 14100 -485
rect 14050 -535 14065 -515
rect 14085 -535 14100 -515
rect 14050 -565 14100 -535
rect 14050 -585 14065 -565
rect 14085 -585 14100 -565
rect 14050 -615 14100 -585
rect 14050 -635 14065 -615
rect 14085 -635 14100 -615
rect 14050 -665 14100 -635
rect 14050 -685 14065 -665
rect 14085 -685 14100 -665
rect 14050 -715 14100 -685
rect 14050 -735 14065 -715
rect 14085 -735 14100 -715
rect 14050 -765 14100 -735
rect 14050 -785 14065 -765
rect 14085 -785 14100 -765
rect 14050 -800 14100 -785
rect 14200 -800 14250 -100
rect 14350 -115 14400 -100
rect 14350 -135 14365 -115
rect 14385 -135 14400 -115
rect 14350 -165 14400 -135
rect 14350 -185 14365 -165
rect 14385 -185 14400 -165
rect 14350 -215 14400 -185
rect 14350 -235 14365 -215
rect 14385 -235 14400 -215
rect 14350 -265 14400 -235
rect 14350 -285 14365 -265
rect 14385 -285 14400 -265
rect 14350 -315 14400 -285
rect 14350 -335 14365 -315
rect 14385 -335 14400 -315
rect 14350 -365 14400 -335
rect 14350 -385 14365 -365
rect 14385 -385 14400 -365
rect 14350 -415 14400 -385
rect 14350 -435 14365 -415
rect 14385 -435 14400 -415
rect 14350 -465 14400 -435
rect 14350 -485 14365 -465
rect 14385 -485 14400 -465
rect 14350 -515 14400 -485
rect 14350 -535 14365 -515
rect 14385 -535 14400 -515
rect 14350 -565 14400 -535
rect 14350 -585 14365 -565
rect 14385 -585 14400 -565
rect 14350 -615 14400 -585
rect 14350 -635 14365 -615
rect 14385 -635 14400 -615
rect 14350 -665 14400 -635
rect 14350 -685 14365 -665
rect 14385 -685 14400 -665
rect 14350 -715 14400 -685
rect 14350 -735 14365 -715
rect 14385 -735 14400 -715
rect 14350 -765 14400 -735
rect 14350 -785 14365 -765
rect 14385 -785 14400 -765
rect 14350 -800 14400 -785
rect 14500 -800 14550 -100
rect 14650 -800 14700 -100
rect 14800 -800 14850 -100
rect 14950 -800 15000 -100
rect 15100 -800 15150 -100
rect 15250 -800 15300 -100
rect 15400 -800 15450 -100
rect 15550 -115 15600 -100
rect 15550 -135 15565 -115
rect 15585 -135 15600 -115
rect 15550 -165 15600 -135
rect 15550 -185 15565 -165
rect 15585 -185 15600 -165
rect 15550 -215 15600 -185
rect 15550 -235 15565 -215
rect 15585 -235 15600 -215
rect 15550 -265 15600 -235
rect 15550 -285 15565 -265
rect 15585 -285 15600 -265
rect 15550 -315 15600 -285
rect 15550 -335 15565 -315
rect 15585 -335 15600 -315
rect 15550 -365 15600 -335
rect 15550 -385 15565 -365
rect 15585 -385 15600 -365
rect 15550 -415 15600 -385
rect 15550 -435 15565 -415
rect 15585 -435 15600 -415
rect 15550 -465 15600 -435
rect 15550 -485 15565 -465
rect 15585 -485 15600 -465
rect 15550 -515 15600 -485
rect 15550 -535 15565 -515
rect 15585 -535 15600 -515
rect 15550 -565 15600 -535
rect 15550 -585 15565 -565
rect 15585 -585 15600 -565
rect 15550 -615 15600 -585
rect 15550 -635 15565 -615
rect 15585 -635 15600 -615
rect 15550 -665 15600 -635
rect 15550 -685 15565 -665
rect 15585 -685 15600 -665
rect 15550 -715 15600 -685
rect 15550 -735 15565 -715
rect 15585 -735 15600 -715
rect 15550 -765 15600 -735
rect 15550 -785 15565 -765
rect 15585 -785 15600 -765
rect 15550 -800 15600 -785
rect 15700 -800 15750 -100
rect 15850 -800 15900 -100
rect 16000 -800 16050 -100
rect 16150 -800 16200 -100
rect 16300 -800 16350 -100
rect 16450 -800 16500 -100
rect 16600 -800 16650 -100
rect 16750 -115 16800 -100
rect 16750 -135 16765 -115
rect 16785 -135 16800 -115
rect 16750 -165 16800 -135
rect 16750 -185 16765 -165
rect 16785 -185 16800 -165
rect 16750 -215 16800 -185
rect 16750 -235 16765 -215
rect 16785 -235 16800 -215
rect 16750 -265 16800 -235
rect 16750 -285 16765 -265
rect 16785 -285 16800 -265
rect 16750 -315 16800 -285
rect 16750 -335 16765 -315
rect 16785 -335 16800 -315
rect 16750 -365 16800 -335
rect 16750 -385 16765 -365
rect 16785 -385 16800 -365
rect 16750 -415 16800 -385
rect 16750 -435 16765 -415
rect 16785 -435 16800 -415
rect 16750 -465 16800 -435
rect 16750 -485 16765 -465
rect 16785 -485 16800 -465
rect 16750 -515 16800 -485
rect 16750 -535 16765 -515
rect 16785 -535 16800 -515
rect 16750 -565 16800 -535
rect 16750 -585 16765 -565
rect 16785 -585 16800 -565
rect 16750 -615 16800 -585
rect 16750 -635 16765 -615
rect 16785 -635 16800 -615
rect 16750 -665 16800 -635
rect 16750 -685 16765 -665
rect 16785 -685 16800 -665
rect 16750 -715 16800 -685
rect 16750 -735 16765 -715
rect 16785 -735 16800 -715
rect 16750 -765 16800 -735
rect 16750 -785 16765 -765
rect 16785 -785 16800 -765
rect 16750 -800 16800 -785
rect 16900 -800 16950 -100
rect 17050 -800 17100 -100
rect 17200 -800 17250 -100
rect 17350 -800 17400 -100
rect 17500 -800 17550 -100
rect 17650 -800 17700 -100
rect 17800 -800 17850 -100
rect 17950 -115 18000 -100
rect 17950 -135 17965 -115
rect 17985 -135 18000 -115
rect 17950 -165 18000 -135
rect 17950 -185 17965 -165
rect 17985 -185 18000 -165
rect 17950 -215 18000 -185
rect 17950 -235 17965 -215
rect 17985 -235 18000 -215
rect 17950 -265 18000 -235
rect 17950 -285 17965 -265
rect 17985 -285 18000 -265
rect 17950 -315 18000 -285
rect 17950 -335 17965 -315
rect 17985 -335 18000 -315
rect 17950 -365 18000 -335
rect 17950 -385 17965 -365
rect 17985 -385 18000 -365
rect 17950 -415 18000 -385
rect 17950 -435 17965 -415
rect 17985 -435 18000 -415
rect 17950 -465 18000 -435
rect 17950 -485 17965 -465
rect 17985 -485 18000 -465
rect 17950 -515 18000 -485
rect 17950 -535 17965 -515
rect 17985 -535 18000 -515
rect 17950 -565 18000 -535
rect 17950 -585 17965 -565
rect 17985 -585 18000 -565
rect 17950 -615 18000 -585
rect 17950 -635 17965 -615
rect 17985 -635 18000 -615
rect 17950 -665 18000 -635
rect 17950 -685 17965 -665
rect 17985 -685 18000 -665
rect 17950 -715 18000 -685
rect 17950 -735 17965 -715
rect 17985 -735 18000 -715
rect 17950 -765 18000 -735
rect 17950 -785 17965 -765
rect 17985 -785 18000 -765
rect 17950 -800 18000 -785
rect 18100 -800 18150 -100
rect 18250 -800 18300 -100
rect 18400 -800 18450 -100
rect 18550 -800 18600 -100
rect 18700 -800 18750 -100
rect 18850 -800 18900 -100
rect 19000 -800 19050 -100
rect 19150 -115 19200 -100
rect 19150 -135 19165 -115
rect 19185 -135 19200 -115
rect 19150 -165 19200 -135
rect 19150 -185 19165 -165
rect 19185 -185 19200 -165
rect 19150 -215 19200 -185
rect 19150 -235 19165 -215
rect 19185 -235 19200 -215
rect 19150 -265 19200 -235
rect 19150 -285 19165 -265
rect 19185 -285 19200 -265
rect 19150 -315 19200 -285
rect 19150 -335 19165 -315
rect 19185 -335 19200 -315
rect 19150 -365 19200 -335
rect 19150 -385 19165 -365
rect 19185 -385 19200 -365
rect 19150 -415 19200 -385
rect 19150 -435 19165 -415
rect 19185 -435 19200 -415
rect 19150 -465 19200 -435
rect 19150 -485 19165 -465
rect 19185 -485 19200 -465
rect 19150 -515 19200 -485
rect 19150 -535 19165 -515
rect 19185 -535 19200 -515
rect 19150 -565 19200 -535
rect 19150 -585 19165 -565
rect 19185 -585 19200 -565
rect 19150 -615 19200 -585
rect 19150 -635 19165 -615
rect 19185 -635 19200 -615
rect 19150 -665 19200 -635
rect 19150 -685 19165 -665
rect 19185 -685 19200 -665
rect 19150 -715 19200 -685
rect 19150 -735 19165 -715
rect 19185 -735 19200 -715
rect 19150 -765 19200 -735
rect 19150 -785 19165 -765
rect 19185 -785 19200 -765
rect 19150 -800 19200 -785
rect 19300 -800 19350 -100
rect 19450 -800 19500 -100
rect 19600 -800 19650 -100
rect 19750 -800 19800 -100
rect 19900 -800 19950 -100
rect 20050 -800 20100 -100
rect 20200 -800 20250 -100
rect 20350 -115 20400 -100
rect 20350 -135 20365 -115
rect 20385 -135 20400 -115
rect 20350 -165 20400 -135
rect 20350 -185 20365 -165
rect 20385 -185 20400 -165
rect 20350 -215 20400 -185
rect 20350 -235 20365 -215
rect 20385 -235 20400 -215
rect 20350 -265 20400 -235
rect 20350 -285 20365 -265
rect 20385 -285 20400 -265
rect 20350 -315 20400 -285
rect 20350 -335 20365 -315
rect 20385 -335 20400 -315
rect 20350 -365 20400 -335
rect 20350 -385 20365 -365
rect 20385 -385 20400 -365
rect 20350 -415 20400 -385
rect 20350 -435 20365 -415
rect 20385 -435 20400 -415
rect 20350 -465 20400 -435
rect 20350 -485 20365 -465
rect 20385 -485 20400 -465
rect 20350 -515 20400 -485
rect 20350 -535 20365 -515
rect 20385 -535 20400 -515
rect 20350 -565 20400 -535
rect 20350 -585 20365 -565
rect 20385 -585 20400 -565
rect 20350 -615 20400 -585
rect 20350 -635 20365 -615
rect 20385 -635 20400 -615
rect 20350 -665 20400 -635
rect 20350 -685 20365 -665
rect 20385 -685 20400 -665
rect 20350 -715 20400 -685
rect 20350 -735 20365 -715
rect 20385 -735 20400 -715
rect 20350 -765 20400 -735
rect 20350 -785 20365 -765
rect 20385 -785 20400 -765
rect 20350 -800 20400 -785
rect -650 -965 -600 -950
rect -650 -985 -635 -965
rect -615 -985 -600 -965
rect -650 -1015 -600 -985
rect -650 -1035 -635 -1015
rect -615 -1035 -600 -1015
rect -650 -1065 -600 -1035
rect -650 -1085 -635 -1065
rect -615 -1085 -600 -1065
rect -650 -1115 -600 -1085
rect -650 -1135 -635 -1115
rect -615 -1135 -600 -1115
rect -650 -1165 -600 -1135
rect -650 -1185 -635 -1165
rect -615 -1185 -600 -1165
rect -650 -1215 -600 -1185
rect -650 -1235 -635 -1215
rect -615 -1235 -600 -1215
rect -650 -1265 -600 -1235
rect -650 -1285 -635 -1265
rect -615 -1285 -600 -1265
rect -650 -1315 -600 -1285
rect -650 -1335 -635 -1315
rect -615 -1335 -600 -1315
rect -650 -1365 -600 -1335
rect -650 -1385 -635 -1365
rect -615 -1385 -600 -1365
rect -650 -1415 -600 -1385
rect -650 -1435 -635 -1415
rect -615 -1435 -600 -1415
rect -650 -1465 -600 -1435
rect -650 -1485 -635 -1465
rect -615 -1485 -600 -1465
rect -650 -1515 -600 -1485
rect -650 -1535 -635 -1515
rect -615 -1535 -600 -1515
rect -650 -1565 -600 -1535
rect -650 -1585 -635 -1565
rect -615 -1585 -600 -1565
rect -650 -1615 -600 -1585
rect -650 -1635 -635 -1615
rect -615 -1635 -600 -1615
rect -650 -1650 -600 -1635
rect -500 -965 -450 -950
rect -500 -985 -485 -965
rect -465 -985 -450 -965
rect -500 -1015 -450 -985
rect -500 -1035 -485 -1015
rect -465 -1035 -450 -1015
rect -500 -1065 -450 -1035
rect -500 -1085 -485 -1065
rect -465 -1085 -450 -1065
rect -500 -1115 -450 -1085
rect -500 -1135 -485 -1115
rect -465 -1135 -450 -1115
rect -500 -1165 -450 -1135
rect -500 -1185 -485 -1165
rect -465 -1185 -450 -1165
rect -500 -1215 -450 -1185
rect -500 -1235 -485 -1215
rect -465 -1235 -450 -1215
rect -500 -1265 -450 -1235
rect -500 -1285 -485 -1265
rect -465 -1285 -450 -1265
rect -500 -1315 -450 -1285
rect -500 -1335 -485 -1315
rect -465 -1335 -450 -1315
rect -500 -1365 -450 -1335
rect -500 -1385 -485 -1365
rect -465 -1385 -450 -1365
rect -500 -1415 -450 -1385
rect -500 -1435 -485 -1415
rect -465 -1435 -450 -1415
rect -500 -1465 -450 -1435
rect -500 -1485 -485 -1465
rect -465 -1485 -450 -1465
rect -500 -1515 -450 -1485
rect -500 -1535 -485 -1515
rect -465 -1535 -450 -1515
rect -500 -1565 -450 -1535
rect -500 -1585 -485 -1565
rect -465 -1585 -450 -1565
rect -500 -1615 -450 -1585
rect -500 -1635 -485 -1615
rect -465 -1635 -450 -1615
rect -500 -1650 -450 -1635
rect -350 -965 -300 -950
rect -350 -985 -335 -965
rect -315 -985 -300 -965
rect -350 -1015 -300 -985
rect -350 -1035 -335 -1015
rect -315 -1035 -300 -1015
rect -350 -1065 -300 -1035
rect -350 -1085 -335 -1065
rect -315 -1085 -300 -1065
rect -350 -1115 -300 -1085
rect -350 -1135 -335 -1115
rect -315 -1135 -300 -1115
rect -350 -1165 -300 -1135
rect -350 -1185 -335 -1165
rect -315 -1185 -300 -1165
rect -350 -1215 -300 -1185
rect -350 -1235 -335 -1215
rect -315 -1235 -300 -1215
rect -350 -1265 -300 -1235
rect -350 -1285 -335 -1265
rect -315 -1285 -300 -1265
rect -350 -1315 -300 -1285
rect -350 -1335 -335 -1315
rect -315 -1335 -300 -1315
rect -350 -1365 -300 -1335
rect -350 -1385 -335 -1365
rect -315 -1385 -300 -1365
rect -350 -1415 -300 -1385
rect -350 -1435 -335 -1415
rect -315 -1435 -300 -1415
rect -350 -1465 -300 -1435
rect -350 -1485 -335 -1465
rect -315 -1485 -300 -1465
rect -350 -1515 -300 -1485
rect -350 -1535 -335 -1515
rect -315 -1535 -300 -1515
rect -350 -1565 -300 -1535
rect -350 -1585 -335 -1565
rect -315 -1585 -300 -1565
rect -350 -1615 -300 -1585
rect -350 -1635 -335 -1615
rect -315 -1635 -300 -1615
rect -350 -1650 -300 -1635
rect -200 -965 -150 -950
rect -200 -985 -185 -965
rect -165 -985 -150 -965
rect -200 -1015 -150 -985
rect -200 -1035 -185 -1015
rect -165 -1035 -150 -1015
rect -200 -1065 -150 -1035
rect -200 -1085 -185 -1065
rect -165 -1085 -150 -1065
rect -200 -1115 -150 -1085
rect -200 -1135 -185 -1115
rect -165 -1135 -150 -1115
rect -200 -1165 -150 -1135
rect -200 -1185 -185 -1165
rect -165 -1185 -150 -1165
rect -200 -1215 -150 -1185
rect -200 -1235 -185 -1215
rect -165 -1235 -150 -1215
rect -200 -1265 -150 -1235
rect -200 -1285 -185 -1265
rect -165 -1285 -150 -1265
rect -200 -1315 -150 -1285
rect -200 -1335 -185 -1315
rect -165 -1335 -150 -1315
rect -200 -1365 -150 -1335
rect -200 -1385 -185 -1365
rect -165 -1385 -150 -1365
rect -200 -1415 -150 -1385
rect -200 -1435 -185 -1415
rect -165 -1435 -150 -1415
rect -200 -1465 -150 -1435
rect -200 -1485 -185 -1465
rect -165 -1485 -150 -1465
rect -200 -1515 -150 -1485
rect -200 -1535 -185 -1515
rect -165 -1535 -150 -1515
rect -200 -1565 -150 -1535
rect -200 -1585 -185 -1565
rect -165 -1585 -150 -1565
rect -200 -1615 -150 -1585
rect -200 -1635 -185 -1615
rect -165 -1635 -150 -1615
rect -200 -1650 -150 -1635
rect -50 -965 0 -950
rect -50 -985 -35 -965
rect -15 -985 0 -965
rect -50 -1015 0 -985
rect -50 -1035 -35 -1015
rect -15 -1035 0 -1015
rect -50 -1065 0 -1035
rect -50 -1085 -35 -1065
rect -15 -1085 0 -1065
rect -50 -1115 0 -1085
rect -50 -1135 -35 -1115
rect -15 -1135 0 -1115
rect -50 -1165 0 -1135
rect -50 -1185 -35 -1165
rect -15 -1185 0 -1165
rect -50 -1215 0 -1185
rect -50 -1235 -35 -1215
rect -15 -1235 0 -1215
rect -50 -1265 0 -1235
rect -50 -1285 -35 -1265
rect -15 -1285 0 -1265
rect -50 -1315 0 -1285
rect -50 -1335 -35 -1315
rect -15 -1335 0 -1315
rect -50 -1365 0 -1335
rect -50 -1385 -35 -1365
rect -15 -1385 0 -1365
rect -50 -1415 0 -1385
rect -50 -1435 -35 -1415
rect -15 -1435 0 -1415
rect -50 -1465 0 -1435
rect -50 -1485 -35 -1465
rect -15 -1485 0 -1465
rect -50 -1515 0 -1485
rect -50 -1535 -35 -1515
rect -15 -1535 0 -1515
rect -50 -1565 0 -1535
rect -50 -1585 -35 -1565
rect -15 -1585 0 -1565
rect -50 -1615 0 -1585
rect -50 -1635 -35 -1615
rect -15 -1635 0 -1615
rect -50 -1650 0 -1635
rect 100 -1650 150 -950
rect 250 -1650 300 -950
rect 400 -1650 450 -950
rect 550 -1650 600 -950
rect 700 -1650 750 -950
rect 850 -1650 900 -950
rect 1000 -1650 1050 -950
rect 1150 -965 1200 -950
rect 1150 -985 1165 -965
rect 1185 -985 1200 -965
rect 1150 -1015 1200 -985
rect 1150 -1035 1165 -1015
rect 1185 -1035 1200 -1015
rect 1150 -1065 1200 -1035
rect 1150 -1085 1165 -1065
rect 1185 -1085 1200 -1065
rect 1150 -1115 1200 -1085
rect 1150 -1135 1165 -1115
rect 1185 -1135 1200 -1115
rect 1150 -1165 1200 -1135
rect 1150 -1185 1165 -1165
rect 1185 -1185 1200 -1165
rect 1150 -1215 1200 -1185
rect 1150 -1235 1165 -1215
rect 1185 -1235 1200 -1215
rect 1150 -1265 1200 -1235
rect 1150 -1285 1165 -1265
rect 1185 -1285 1200 -1265
rect 1150 -1315 1200 -1285
rect 1150 -1335 1165 -1315
rect 1185 -1335 1200 -1315
rect 1150 -1365 1200 -1335
rect 1150 -1385 1165 -1365
rect 1185 -1385 1200 -1365
rect 1150 -1415 1200 -1385
rect 1150 -1435 1165 -1415
rect 1185 -1435 1200 -1415
rect 1150 -1465 1200 -1435
rect 1150 -1485 1165 -1465
rect 1185 -1485 1200 -1465
rect 1150 -1515 1200 -1485
rect 1150 -1535 1165 -1515
rect 1185 -1535 1200 -1515
rect 1150 -1565 1200 -1535
rect 1150 -1585 1165 -1565
rect 1185 -1585 1200 -1565
rect 1150 -1615 1200 -1585
rect 1150 -1635 1165 -1615
rect 1185 -1635 1200 -1615
rect 1150 -1650 1200 -1635
rect 1300 -1650 1350 -950
rect 1450 -965 1500 -950
rect 1450 -985 1465 -965
rect 1485 -985 1500 -965
rect 1450 -1015 1500 -985
rect 1450 -1035 1465 -1015
rect 1485 -1035 1500 -1015
rect 1450 -1065 1500 -1035
rect 1450 -1085 1465 -1065
rect 1485 -1085 1500 -1065
rect 1450 -1115 1500 -1085
rect 1450 -1135 1465 -1115
rect 1485 -1135 1500 -1115
rect 1450 -1165 1500 -1135
rect 1450 -1185 1465 -1165
rect 1485 -1185 1500 -1165
rect 1450 -1215 1500 -1185
rect 1450 -1235 1465 -1215
rect 1485 -1235 1500 -1215
rect 1450 -1265 1500 -1235
rect 1450 -1285 1465 -1265
rect 1485 -1285 1500 -1265
rect 1450 -1315 1500 -1285
rect 1450 -1335 1465 -1315
rect 1485 -1335 1500 -1315
rect 1450 -1365 1500 -1335
rect 1450 -1385 1465 -1365
rect 1485 -1385 1500 -1365
rect 1450 -1415 1500 -1385
rect 1450 -1435 1465 -1415
rect 1485 -1435 1500 -1415
rect 1450 -1465 1500 -1435
rect 1450 -1485 1465 -1465
rect 1485 -1485 1500 -1465
rect 1450 -1515 1500 -1485
rect 1450 -1535 1465 -1515
rect 1485 -1535 1500 -1515
rect 1450 -1565 1500 -1535
rect 1450 -1585 1465 -1565
rect 1485 -1585 1500 -1565
rect 1450 -1615 1500 -1585
rect 1450 -1635 1465 -1615
rect 1485 -1635 1500 -1615
rect 1450 -1650 1500 -1635
rect 1600 -1650 1650 -950
rect 1750 -965 1800 -950
rect 1750 -985 1765 -965
rect 1785 -985 1800 -965
rect 1750 -1015 1800 -985
rect 1750 -1035 1765 -1015
rect 1785 -1035 1800 -1015
rect 1750 -1065 1800 -1035
rect 1750 -1085 1765 -1065
rect 1785 -1085 1800 -1065
rect 1750 -1115 1800 -1085
rect 1750 -1135 1765 -1115
rect 1785 -1135 1800 -1115
rect 1750 -1165 1800 -1135
rect 1750 -1185 1765 -1165
rect 1785 -1185 1800 -1165
rect 1750 -1215 1800 -1185
rect 1750 -1235 1765 -1215
rect 1785 -1235 1800 -1215
rect 1750 -1265 1800 -1235
rect 1750 -1285 1765 -1265
rect 1785 -1285 1800 -1265
rect 1750 -1315 1800 -1285
rect 1750 -1335 1765 -1315
rect 1785 -1335 1800 -1315
rect 1750 -1365 1800 -1335
rect 1750 -1385 1765 -1365
rect 1785 -1385 1800 -1365
rect 1750 -1415 1800 -1385
rect 1750 -1435 1765 -1415
rect 1785 -1435 1800 -1415
rect 1750 -1465 1800 -1435
rect 1750 -1485 1765 -1465
rect 1785 -1485 1800 -1465
rect 1750 -1515 1800 -1485
rect 1750 -1535 1765 -1515
rect 1785 -1535 1800 -1515
rect 1750 -1565 1800 -1535
rect 1750 -1585 1765 -1565
rect 1785 -1585 1800 -1565
rect 1750 -1615 1800 -1585
rect 1750 -1635 1765 -1615
rect 1785 -1635 1800 -1615
rect 1750 -1650 1800 -1635
rect 1900 -1650 1950 -950
rect 2050 -965 2100 -950
rect 2050 -985 2065 -965
rect 2085 -985 2100 -965
rect 2050 -1015 2100 -985
rect 2050 -1035 2065 -1015
rect 2085 -1035 2100 -1015
rect 2050 -1065 2100 -1035
rect 2050 -1085 2065 -1065
rect 2085 -1085 2100 -1065
rect 2050 -1115 2100 -1085
rect 2050 -1135 2065 -1115
rect 2085 -1135 2100 -1115
rect 2050 -1165 2100 -1135
rect 2050 -1185 2065 -1165
rect 2085 -1185 2100 -1165
rect 2050 -1215 2100 -1185
rect 2050 -1235 2065 -1215
rect 2085 -1235 2100 -1215
rect 2050 -1265 2100 -1235
rect 2050 -1285 2065 -1265
rect 2085 -1285 2100 -1265
rect 2050 -1315 2100 -1285
rect 2050 -1335 2065 -1315
rect 2085 -1335 2100 -1315
rect 2050 -1365 2100 -1335
rect 2050 -1385 2065 -1365
rect 2085 -1385 2100 -1365
rect 2050 -1415 2100 -1385
rect 2050 -1435 2065 -1415
rect 2085 -1435 2100 -1415
rect 2050 -1465 2100 -1435
rect 2050 -1485 2065 -1465
rect 2085 -1485 2100 -1465
rect 2050 -1515 2100 -1485
rect 2050 -1535 2065 -1515
rect 2085 -1535 2100 -1515
rect 2050 -1565 2100 -1535
rect 2050 -1585 2065 -1565
rect 2085 -1585 2100 -1565
rect 2050 -1615 2100 -1585
rect 2050 -1635 2065 -1615
rect 2085 -1635 2100 -1615
rect 2050 -1650 2100 -1635
rect 2200 -1650 2250 -950
rect 2350 -965 2400 -950
rect 2350 -985 2365 -965
rect 2385 -985 2400 -965
rect 2350 -1015 2400 -985
rect 2350 -1035 2365 -1015
rect 2385 -1035 2400 -1015
rect 2350 -1065 2400 -1035
rect 2350 -1085 2365 -1065
rect 2385 -1085 2400 -1065
rect 2350 -1115 2400 -1085
rect 2350 -1135 2365 -1115
rect 2385 -1135 2400 -1115
rect 2350 -1165 2400 -1135
rect 2350 -1185 2365 -1165
rect 2385 -1185 2400 -1165
rect 2350 -1215 2400 -1185
rect 2350 -1235 2365 -1215
rect 2385 -1235 2400 -1215
rect 2350 -1265 2400 -1235
rect 2350 -1285 2365 -1265
rect 2385 -1285 2400 -1265
rect 2350 -1315 2400 -1285
rect 2350 -1335 2365 -1315
rect 2385 -1335 2400 -1315
rect 2350 -1365 2400 -1335
rect 2350 -1385 2365 -1365
rect 2385 -1385 2400 -1365
rect 2350 -1415 2400 -1385
rect 2350 -1435 2365 -1415
rect 2385 -1435 2400 -1415
rect 2350 -1465 2400 -1435
rect 2350 -1485 2365 -1465
rect 2385 -1485 2400 -1465
rect 2350 -1515 2400 -1485
rect 2350 -1535 2365 -1515
rect 2385 -1535 2400 -1515
rect 2350 -1565 2400 -1535
rect 2350 -1585 2365 -1565
rect 2385 -1585 2400 -1565
rect 2350 -1615 2400 -1585
rect 2350 -1635 2365 -1615
rect 2385 -1635 2400 -1615
rect 2350 -1650 2400 -1635
rect 2500 -1650 2550 -950
rect 2650 -965 2700 -950
rect 2650 -985 2665 -965
rect 2685 -985 2700 -965
rect 2650 -1015 2700 -985
rect 2650 -1035 2665 -1015
rect 2685 -1035 2700 -1015
rect 2650 -1065 2700 -1035
rect 2650 -1085 2665 -1065
rect 2685 -1085 2700 -1065
rect 2650 -1115 2700 -1085
rect 2650 -1135 2665 -1115
rect 2685 -1135 2700 -1115
rect 2650 -1165 2700 -1135
rect 2650 -1185 2665 -1165
rect 2685 -1185 2700 -1165
rect 2650 -1215 2700 -1185
rect 2650 -1235 2665 -1215
rect 2685 -1235 2700 -1215
rect 2650 -1265 2700 -1235
rect 2650 -1285 2665 -1265
rect 2685 -1285 2700 -1265
rect 2650 -1315 2700 -1285
rect 2650 -1335 2665 -1315
rect 2685 -1335 2700 -1315
rect 2650 -1365 2700 -1335
rect 2650 -1385 2665 -1365
rect 2685 -1385 2700 -1365
rect 2650 -1415 2700 -1385
rect 2650 -1435 2665 -1415
rect 2685 -1435 2700 -1415
rect 2650 -1465 2700 -1435
rect 2650 -1485 2665 -1465
rect 2685 -1485 2700 -1465
rect 2650 -1515 2700 -1485
rect 2650 -1535 2665 -1515
rect 2685 -1535 2700 -1515
rect 2650 -1565 2700 -1535
rect 2650 -1585 2665 -1565
rect 2685 -1585 2700 -1565
rect 2650 -1615 2700 -1585
rect 2650 -1635 2665 -1615
rect 2685 -1635 2700 -1615
rect 2650 -1650 2700 -1635
rect 2800 -1650 2850 -950
rect 2950 -965 3000 -950
rect 2950 -985 2965 -965
rect 2985 -985 3000 -965
rect 2950 -1015 3000 -985
rect 2950 -1035 2965 -1015
rect 2985 -1035 3000 -1015
rect 2950 -1065 3000 -1035
rect 2950 -1085 2965 -1065
rect 2985 -1085 3000 -1065
rect 2950 -1115 3000 -1085
rect 2950 -1135 2965 -1115
rect 2985 -1135 3000 -1115
rect 2950 -1165 3000 -1135
rect 2950 -1185 2965 -1165
rect 2985 -1185 3000 -1165
rect 2950 -1215 3000 -1185
rect 2950 -1235 2965 -1215
rect 2985 -1235 3000 -1215
rect 2950 -1265 3000 -1235
rect 2950 -1285 2965 -1265
rect 2985 -1285 3000 -1265
rect 2950 -1315 3000 -1285
rect 2950 -1335 2965 -1315
rect 2985 -1335 3000 -1315
rect 2950 -1365 3000 -1335
rect 2950 -1385 2965 -1365
rect 2985 -1385 3000 -1365
rect 2950 -1415 3000 -1385
rect 2950 -1435 2965 -1415
rect 2985 -1435 3000 -1415
rect 2950 -1465 3000 -1435
rect 2950 -1485 2965 -1465
rect 2985 -1485 3000 -1465
rect 2950 -1515 3000 -1485
rect 2950 -1535 2965 -1515
rect 2985 -1535 3000 -1515
rect 2950 -1565 3000 -1535
rect 2950 -1585 2965 -1565
rect 2985 -1585 3000 -1565
rect 2950 -1615 3000 -1585
rect 2950 -1635 2965 -1615
rect 2985 -1635 3000 -1615
rect 2950 -1650 3000 -1635
rect 3100 -1650 3150 -950
rect 3250 -965 3300 -950
rect 3250 -985 3265 -965
rect 3285 -985 3300 -965
rect 3250 -1015 3300 -985
rect 3250 -1035 3265 -1015
rect 3285 -1035 3300 -1015
rect 3250 -1065 3300 -1035
rect 3250 -1085 3265 -1065
rect 3285 -1085 3300 -1065
rect 3250 -1115 3300 -1085
rect 3250 -1135 3265 -1115
rect 3285 -1135 3300 -1115
rect 3250 -1165 3300 -1135
rect 3250 -1185 3265 -1165
rect 3285 -1185 3300 -1165
rect 3250 -1215 3300 -1185
rect 3250 -1235 3265 -1215
rect 3285 -1235 3300 -1215
rect 3250 -1265 3300 -1235
rect 3250 -1285 3265 -1265
rect 3285 -1285 3300 -1265
rect 3250 -1315 3300 -1285
rect 3250 -1335 3265 -1315
rect 3285 -1335 3300 -1315
rect 3250 -1365 3300 -1335
rect 3250 -1385 3265 -1365
rect 3285 -1385 3300 -1365
rect 3250 -1415 3300 -1385
rect 3250 -1435 3265 -1415
rect 3285 -1435 3300 -1415
rect 3250 -1465 3300 -1435
rect 3250 -1485 3265 -1465
rect 3285 -1485 3300 -1465
rect 3250 -1515 3300 -1485
rect 3250 -1535 3265 -1515
rect 3285 -1535 3300 -1515
rect 3250 -1565 3300 -1535
rect 3250 -1585 3265 -1565
rect 3285 -1585 3300 -1565
rect 3250 -1615 3300 -1585
rect 3250 -1635 3265 -1615
rect 3285 -1635 3300 -1615
rect 3250 -1650 3300 -1635
rect 3400 -1650 3450 -950
rect 3550 -965 3600 -950
rect 3550 -985 3565 -965
rect 3585 -985 3600 -965
rect 3550 -1015 3600 -985
rect 3550 -1035 3565 -1015
rect 3585 -1035 3600 -1015
rect 3550 -1065 3600 -1035
rect 3550 -1085 3565 -1065
rect 3585 -1085 3600 -1065
rect 3550 -1115 3600 -1085
rect 3550 -1135 3565 -1115
rect 3585 -1135 3600 -1115
rect 3550 -1165 3600 -1135
rect 3550 -1185 3565 -1165
rect 3585 -1185 3600 -1165
rect 3550 -1215 3600 -1185
rect 3550 -1235 3565 -1215
rect 3585 -1235 3600 -1215
rect 3550 -1265 3600 -1235
rect 3550 -1285 3565 -1265
rect 3585 -1285 3600 -1265
rect 3550 -1315 3600 -1285
rect 3550 -1335 3565 -1315
rect 3585 -1335 3600 -1315
rect 3550 -1365 3600 -1335
rect 3550 -1385 3565 -1365
rect 3585 -1385 3600 -1365
rect 3550 -1415 3600 -1385
rect 3550 -1435 3565 -1415
rect 3585 -1435 3600 -1415
rect 3550 -1465 3600 -1435
rect 3550 -1485 3565 -1465
rect 3585 -1485 3600 -1465
rect 3550 -1515 3600 -1485
rect 3550 -1535 3565 -1515
rect 3585 -1535 3600 -1515
rect 3550 -1565 3600 -1535
rect 3550 -1585 3565 -1565
rect 3585 -1585 3600 -1565
rect 3550 -1615 3600 -1585
rect 3550 -1635 3565 -1615
rect 3585 -1635 3600 -1615
rect 3550 -1650 3600 -1635
rect 3700 -965 3750 -950
rect 3700 -985 3715 -965
rect 3735 -985 3750 -965
rect 3700 -1015 3750 -985
rect 3700 -1035 3715 -1015
rect 3735 -1035 3750 -1015
rect 3700 -1065 3750 -1035
rect 3700 -1085 3715 -1065
rect 3735 -1085 3750 -1065
rect 3700 -1115 3750 -1085
rect 3700 -1135 3715 -1115
rect 3735 -1135 3750 -1115
rect 3700 -1165 3750 -1135
rect 3700 -1185 3715 -1165
rect 3735 -1185 3750 -1165
rect 3700 -1215 3750 -1185
rect 3700 -1235 3715 -1215
rect 3735 -1235 3750 -1215
rect 3700 -1265 3750 -1235
rect 3700 -1285 3715 -1265
rect 3735 -1285 3750 -1265
rect 3700 -1315 3750 -1285
rect 3700 -1335 3715 -1315
rect 3735 -1335 3750 -1315
rect 3700 -1365 3750 -1335
rect 3700 -1385 3715 -1365
rect 3735 -1385 3750 -1365
rect 3700 -1415 3750 -1385
rect 3700 -1435 3715 -1415
rect 3735 -1435 3750 -1415
rect 3700 -1465 3750 -1435
rect 3700 -1485 3715 -1465
rect 3735 -1485 3750 -1465
rect 3700 -1515 3750 -1485
rect 3700 -1535 3715 -1515
rect 3735 -1535 3750 -1515
rect 3700 -1565 3750 -1535
rect 3700 -1585 3715 -1565
rect 3735 -1585 3750 -1565
rect 3700 -1615 3750 -1585
rect 3700 -1635 3715 -1615
rect 3735 -1635 3750 -1615
rect 3700 -1650 3750 -1635
rect 3850 -965 3900 -950
rect 3850 -985 3865 -965
rect 3885 -985 3900 -965
rect 3850 -1015 3900 -985
rect 3850 -1035 3865 -1015
rect 3885 -1035 3900 -1015
rect 3850 -1065 3900 -1035
rect 3850 -1085 3865 -1065
rect 3885 -1085 3900 -1065
rect 3850 -1115 3900 -1085
rect 3850 -1135 3865 -1115
rect 3885 -1135 3900 -1115
rect 3850 -1165 3900 -1135
rect 3850 -1185 3865 -1165
rect 3885 -1185 3900 -1165
rect 3850 -1215 3900 -1185
rect 3850 -1235 3865 -1215
rect 3885 -1235 3900 -1215
rect 3850 -1265 3900 -1235
rect 3850 -1285 3865 -1265
rect 3885 -1285 3900 -1265
rect 3850 -1315 3900 -1285
rect 3850 -1335 3865 -1315
rect 3885 -1335 3900 -1315
rect 3850 -1365 3900 -1335
rect 3850 -1385 3865 -1365
rect 3885 -1385 3900 -1365
rect 3850 -1415 3900 -1385
rect 3850 -1435 3865 -1415
rect 3885 -1435 3900 -1415
rect 3850 -1465 3900 -1435
rect 3850 -1485 3865 -1465
rect 3885 -1485 3900 -1465
rect 3850 -1515 3900 -1485
rect 3850 -1535 3865 -1515
rect 3885 -1535 3900 -1515
rect 3850 -1565 3900 -1535
rect 3850 -1585 3865 -1565
rect 3885 -1585 3900 -1565
rect 3850 -1615 3900 -1585
rect 3850 -1635 3865 -1615
rect 3885 -1635 3900 -1615
rect 3850 -1650 3900 -1635
rect 4000 -965 4050 -950
rect 4000 -985 4015 -965
rect 4035 -985 4050 -965
rect 4000 -1015 4050 -985
rect 4000 -1035 4015 -1015
rect 4035 -1035 4050 -1015
rect 4000 -1065 4050 -1035
rect 4000 -1085 4015 -1065
rect 4035 -1085 4050 -1065
rect 4000 -1115 4050 -1085
rect 4000 -1135 4015 -1115
rect 4035 -1135 4050 -1115
rect 4000 -1165 4050 -1135
rect 4000 -1185 4015 -1165
rect 4035 -1185 4050 -1165
rect 4000 -1215 4050 -1185
rect 4000 -1235 4015 -1215
rect 4035 -1235 4050 -1215
rect 4000 -1265 4050 -1235
rect 4000 -1285 4015 -1265
rect 4035 -1285 4050 -1265
rect 4000 -1315 4050 -1285
rect 4000 -1335 4015 -1315
rect 4035 -1335 4050 -1315
rect 4000 -1365 4050 -1335
rect 4000 -1385 4015 -1365
rect 4035 -1385 4050 -1365
rect 4000 -1415 4050 -1385
rect 4000 -1435 4015 -1415
rect 4035 -1435 4050 -1415
rect 4000 -1465 4050 -1435
rect 4000 -1485 4015 -1465
rect 4035 -1485 4050 -1465
rect 4000 -1515 4050 -1485
rect 4000 -1535 4015 -1515
rect 4035 -1535 4050 -1515
rect 4000 -1565 4050 -1535
rect 4000 -1585 4015 -1565
rect 4035 -1585 4050 -1565
rect 4000 -1615 4050 -1585
rect 4000 -1635 4015 -1615
rect 4035 -1635 4050 -1615
rect 4000 -1650 4050 -1635
rect 4150 -965 4200 -950
rect 4150 -985 4165 -965
rect 4185 -985 4200 -965
rect 4150 -1015 4200 -985
rect 4150 -1035 4165 -1015
rect 4185 -1035 4200 -1015
rect 4150 -1065 4200 -1035
rect 4150 -1085 4165 -1065
rect 4185 -1085 4200 -1065
rect 4150 -1115 4200 -1085
rect 4150 -1135 4165 -1115
rect 4185 -1135 4200 -1115
rect 4150 -1165 4200 -1135
rect 4150 -1185 4165 -1165
rect 4185 -1185 4200 -1165
rect 4150 -1215 4200 -1185
rect 4150 -1235 4165 -1215
rect 4185 -1235 4200 -1215
rect 4150 -1265 4200 -1235
rect 4150 -1285 4165 -1265
rect 4185 -1285 4200 -1265
rect 4150 -1315 4200 -1285
rect 4150 -1335 4165 -1315
rect 4185 -1335 4200 -1315
rect 4150 -1365 4200 -1335
rect 4150 -1385 4165 -1365
rect 4185 -1385 4200 -1365
rect 4150 -1415 4200 -1385
rect 4150 -1435 4165 -1415
rect 4185 -1435 4200 -1415
rect 4150 -1465 4200 -1435
rect 4150 -1485 4165 -1465
rect 4185 -1485 4200 -1465
rect 4150 -1515 4200 -1485
rect 4150 -1535 4165 -1515
rect 4185 -1535 4200 -1515
rect 4150 -1565 4200 -1535
rect 4150 -1585 4165 -1565
rect 4185 -1585 4200 -1565
rect 4150 -1615 4200 -1585
rect 4150 -1635 4165 -1615
rect 4185 -1635 4200 -1615
rect 4150 -1650 4200 -1635
rect 4300 -965 4350 -950
rect 4300 -985 4315 -965
rect 4335 -985 4350 -965
rect 4300 -1015 4350 -985
rect 4300 -1035 4315 -1015
rect 4335 -1035 4350 -1015
rect 4300 -1065 4350 -1035
rect 4300 -1085 4315 -1065
rect 4335 -1085 4350 -1065
rect 4300 -1115 4350 -1085
rect 4300 -1135 4315 -1115
rect 4335 -1135 4350 -1115
rect 4300 -1165 4350 -1135
rect 4300 -1185 4315 -1165
rect 4335 -1185 4350 -1165
rect 4300 -1215 4350 -1185
rect 4300 -1235 4315 -1215
rect 4335 -1235 4350 -1215
rect 4300 -1265 4350 -1235
rect 4300 -1285 4315 -1265
rect 4335 -1285 4350 -1265
rect 4300 -1315 4350 -1285
rect 4300 -1335 4315 -1315
rect 4335 -1335 4350 -1315
rect 4300 -1365 4350 -1335
rect 4300 -1385 4315 -1365
rect 4335 -1385 4350 -1365
rect 4300 -1415 4350 -1385
rect 4300 -1435 4315 -1415
rect 4335 -1435 4350 -1415
rect 4300 -1465 4350 -1435
rect 4300 -1485 4315 -1465
rect 4335 -1485 4350 -1465
rect 4300 -1515 4350 -1485
rect 4300 -1535 4315 -1515
rect 4335 -1535 4350 -1515
rect 4300 -1565 4350 -1535
rect 4300 -1585 4315 -1565
rect 4335 -1585 4350 -1565
rect 4300 -1615 4350 -1585
rect 4300 -1635 4315 -1615
rect 4335 -1635 4350 -1615
rect 4300 -1650 4350 -1635
rect 4450 -965 4500 -950
rect 4450 -985 4465 -965
rect 4485 -985 4500 -965
rect 4450 -1015 4500 -985
rect 4450 -1035 4465 -1015
rect 4485 -1035 4500 -1015
rect 4450 -1065 4500 -1035
rect 4450 -1085 4465 -1065
rect 4485 -1085 4500 -1065
rect 4450 -1115 4500 -1085
rect 4450 -1135 4465 -1115
rect 4485 -1135 4500 -1115
rect 4450 -1165 4500 -1135
rect 4450 -1185 4465 -1165
rect 4485 -1185 4500 -1165
rect 4450 -1215 4500 -1185
rect 4450 -1235 4465 -1215
rect 4485 -1235 4500 -1215
rect 4450 -1265 4500 -1235
rect 4450 -1285 4465 -1265
rect 4485 -1285 4500 -1265
rect 4450 -1315 4500 -1285
rect 4450 -1335 4465 -1315
rect 4485 -1335 4500 -1315
rect 4450 -1365 4500 -1335
rect 4450 -1385 4465 -1365
rect 4485 -1385 4500 -1365
rect 4450 -1415 4500 -1385
rect 4450 -1435 4465 -1415
rect 4485 -1435 4500 -1415
rect 4450 -1465 4500 -1435
rect 4450 -1485 4465 -1465
rect 4485 -1485 4500 -1465
rect 4450 -1515 4500 -1485
rect 4450 -1535 4465 -1515
rect 4485 -1535 4500 -1515
rect 4450 -1565 4500 -1535
rect 4450 -1585 4465 -1565
rect 4485 -1585 4500 -1565
rect 4450 -1615 4500 -1585
rect 4450 -1635 4465 -1615
rect 4485 -1635 4500 -1615
rect 4450 -1650 4500 -1635
rect 4600 -965 4650 -950
rect 4600 -985 4615 -965
rect 4635 -985 4650 -965
rect 4600 -1015 4650 -985
rect 4600 -1035 4615 -1015
rect 4635 -1035 4650 -1015
rect 4600 -1065 4650 -1035
rect 4600 -1085 4615 -1065
rect 4635 -1085 4650 -1065
rect 4600 -1115 4650 -1085
rect 4600 -1135 4615 -1115
rect 4635 -1135 4650 -1115
rect 4600 -1165 4650 -1135
rect 4600 -1185 4615 -1165
rect 4635 -1185 4650 -1165
rect 4600 -1215 4650 -1185
rect 4600 -1235 4615 -1215
rect 4635 -1235 4650 -1215
rect 4600 -1265 4650 -1235
rect 4600 -1285 4615 -1265
rect 4635 -1285 4650 -1265
rect 4600 -1315 4650 -1285
rect 4600 -1335 4615 -1315
rect 4635 -1335 4650 -1315
rect 4600 -1365 4650 -1335
rect 4600 -1385 4615 -1365
rect 4635 -1385 4650 -1365
rect 4600 -1415 4650 -1385
rect 4600 -1435 4615 -1415
rect 4635 -1435 4650 -1415
rect 4600 -1465 4650 -1435
rect 4600 -1485 4615 -1465
rect 4635 -1485 4650 -1465
rect 4600 -1515 4650 -1485
rect 4600 -1535 4615 -1515
rect 4635 -1535 4650 -1515
rect 4600 -1565 4650 -1535
rect 4600 -1585 4615 -1565
rect 4635 -1585 4650 -1565
rect 4600 -1615 4650 -1585
rect 4600 -1635 4615 -1615
rect 4635 -1635 4650 -1615
rect 4600 -1650 4650 -1635
rect 4750 -965 4800 -950
rect 4750 -985 4765 -965
rect 4785 -985 4800 -965
rect 4750 -1015 4800 -985
rect 4750 -1035 4765 -1015
rect 4785 -1035 4800 -1015
rect 4750 -1065 4800 -1035
rect 4750 -1085 4765 -1065
rect 4785 -1085 4800 -1065
rect 4750 -1115 4800 -1085
rect 4750 -1135 4765 -1115
rect 4785 -1135 4800 -1115
rect 4750 -1165 4800 -1135
rect 4750 -1185 4765 -1165
rect 4785 -1185 4800 -1165
rect 4750 -1215 4800 -1185
rect 4750 -1235 4765 -1215
rect 4785 -1235 4800 -1215
rect 4750 -1265 4800 -1235
rect 4750 -1285 4765 -1265
rect 4785 -1285 4800 -1265
rect 4750 -1315 4800 -1285
rect 4750 -1335 4765 -1315
rect 4785 -1335 4800 -1315
rect 4750 -1365 4800 -1335
rect 4750 -1385 4765 -1365
rect 4785 -1385 4800 -1365
rect 4750 -1415 4800 -1385
rect 4750 -1435 4765 -1415
rect 4785 -1435 4800 -1415
rect 4750 -1465 4800 -1435
rect 4750 -1485 4765 -1465
rect 4785 -1485 4800 -1465
rect 4750 -1515 4800 -1485
rect 4750 -1535 4765 -1515
rect 4785 -1535 4800 -1515
rect 4750 -1565 4800 -1535
rect 4750 -1585 4765 -1565
rect 4785 -1585 4800 -1565
rect 4750 -1615 4800 -1585
rect 4750 -1635 4765 -1615
rect 4785 -1635 4800 -1615
rect 4750 -1650 4800 -1635
rect 4900 -1650 4950 -950
rect 5050 -965 5100 -950
rect 5050 -985 5065 -965
rect 5085 -985 5100 -965
rect 5050 -1015 5100 -985
rect 5050 -1035 5065 -1015
rect 5085 -1035 5100 -1015
rect 5050 -1065 5100 -1035
rect 5050 -1085 5065 -1065
rect 5085 -1085 5100 -1065
rect 5050 -1115 5100 -1085
rect 5050 -1135 5065 -1115
rect 5085 -1135 5100 -1115
rect 5050 -1165 5100 -1135
rect 5050 -1185 5065 -1165
rect 5085 -1185 5100 -1165
rect 5050 -1215 5100 -1185
rect 5050 -1235 5065 -1215
rect 5085 -1235 5100 -1215
rect 5050 -1265 5100 -1235
rect 5050 -1285 5065 -1265
rect 5085 -1285 5100 -1265
rect 5050 -1315 5100 -1285
rect 5050 -1335 5065 -1315
rect 5085 -1335 5100 -1315
rect 5050 -1365 5100 -1335
rect 5050 -1385 5065 -1365
rect 5085 -1385 5100 -1365
rect 5050 -1415 5100 -1385
rect 5050 -1435 5065 -1415
rect 5085 -1435 5100 -1415
rect 5050 -1465 5100 -1435
rect 5050 -1485 5065 -1465
rect 5085 -1485 5100 -1465
rect 5050 -1515 5100 -1485
rect 5050 -1535 5065 -1515
rect 5085 -1535 5100 -1515
rect 5050 -1565 5100 -1535
rect 5050 -1585 5065 -1565
rect 5085 -1585 5100 -1565
rect 5050 -1615 5100 -1585
rect 5050 -1635 5065 -1615
rect 5085 -1635 5100 -1615
rect 5050 -1650 5100 -1635
rect 5200 -1650 5250 -950
rect 5350 -965 5400 -950
rect 5350 -985 5365 -965
rect 5385 -985 5400 -965
rect 5350 -1015 5400 -985
rect 5350 -1035 5365 -1015
rect 5385 -1035 5400 -1015
rect 5350 -1065 5400 -1035
rect 5350 -1085 5365 -1065
rect 5385 -1085 5400 -1065
rect 5350 -1115 5400 -1085
rect 5350 -1135 5365 -1115
rect 5385 -1135 5400 -1115
rect 5350 -1165 5400 -1135
rect 5350 -1185 5365 -1165
rect 5385 -1185 5400 -1165
rect 5350 -1215 5400 -1185
rect 5350 -1235 5365 -1215
rect 5385 -1235 5400 -1215
rect 5350 -1265 5400 -1235
rect 5350 -1285 5365 -1265
rect 5385 -1285 5400 -1265
rect 5350 -1315 5400 -1285
rect 5350 -1335 5365 -1315
rect 5385 -1335 5400 -1315
rect 5350 -1365 5400 -1335
rect 5350 -1385 5365 -1365
rect 5385 -1385 5400 -1365
rect 5350 -1415 5400 -1385
rect 5350 -1435 5365 -1415
rect 5385 -1435 5400 -1415
rect 5350 -1465 5400 -1435
rect 5350 -1485 5365 -1465
rect 5385 -1485 5400 -1465
rect 5350 -1515 5400 -1485
rect 5350 -1535 5365 -1515
rect 5385 -1535 5400 -1515
rect 5350 -1565 5400 -1535
rect 5350 -1585 5365 -1565
rect 5385 -1585 5400 -1565
rect 5350 -1615 5400 -1585
rect 5350 -1635 5365 -1615
rect 5385 -1635 5400 -1615
rect 5350 -1650 5400 -1635
rect 5500 -1650 5550 -950
rect 5650 -965 5700 -950
rect 5650 -985 5665 -965
rect 5685 -985 5700 -965
rect 5650 -1015 5700 -985
rect 5650 -1035 5665 -1015
rect 5685 -1035 5700 -1015
rect 5650 -1065 5700 -1035
rect 5650 -1085 5665 -1065
rect 5685 -1085 5700 -1065
rect 5650 -1115 5700 -1085
rect 5650 -1135 5665 -1115
rect 5685 -1135 5700 -1115
rect 5650 -1165 5700 -1135
rect 5650 -1185 5665 -1165
rect 5685 -1185 5700 -1165
rect 5650 -1215 5700 -1185
rect 5650 -1235 5665 -1215
rect 5685 -1235 5700 -1215
rect 5650 -1265 5700 -1235
rect 5650 -1285 5665 -1265
rect 5685 -1285 5700 -1265
rect 5650 -1315 5700 -1285
rect 5650 -1335 5665 -1315
rect 5685 -1335 5700 -1315
rect 5650 -1365 5700 -1335
rect 5650 -1385 5665 -1365
rect 5685 -1385 5700 -1365
rect 5650 -1415 5700 -1385
rect 5650 -1435 5665 -1415
rect 5685 -1435 5700 -1415
rect 5650 -1465 5700 -1435
rect 5650 -1485 5665 -1465
rect 5685 -1485 5700 -1465
rect 5650 -1515 5700 -1485
rect 5650 -1535 5665 -1515
rect 5685 -1535 5700 -1515
rect 5650 -1565 5700 -1535
rect 5650 -1585 5665 -1565
rect 5685 -1585 5700 -1565
rect 5650 -1615 5700 -1585
rect 5650 -1635 5665 -1615
rect 5685 -1635 5700 -1615
rect 5650 -1650 5700 -1635
rect 5800 -1650 5850 -950
rect 5950 -965 6000 -950
rect 5950 -985 5965 -965
rect 5985 -985 6000 -965
rect 5950 -1015 6000 -985
rect 5950 -1035 5965 -1015
rect 5985 -1035 6000 -1015
rect 5950 -1065 6000 -1035
rect 5950 -1085 5965 -1065
rect 5985 -1085 6000 -1065
rect 5950 -1115 6000 -1085
rect 5950 -1135 5965 -1115
rect 5985 -1135 6000 -1115
rect 5950 -1165 6000 -1135
rect 5950 -1185 5965 -1165
rect 5985 -1185 6000 -1165
rect 5950 -1215 6000 -1185
rect 5950 -1235 5965 -1215
rect 5985 -1235 6000 -1215
rect 5950 -1265 6000 -1235
rect 5950 -1285 5965 -1265
rect 5985 -1285 6000 -1265
rect 5950 -1315 6000 -1285
rect 5950 -1335 5965 -1315
rect 5985 -1335 6000 -1315
rect 5950 -1365 6000 -1335
rect 5950 -1385 5965 -1365
rect 5985 -1385 6000 -1365
rect 5950 -1415 6000 -1385
rect 5950 -1435 5965 -1415
rect 5985 -1435 6000 -1415
rect 5950 -1465 6000 -1435
rect 5950 -1485 5965 -1465
rect 5985 -1485 6000 -1465
rect 5950 -1515 6000 -1485
rect 5950 -1535 5965 -1515
rect 5985 -1535 6000 -1515
rect 5950 -1565 6000 -1535
rect 5950 -1585 5965 -1565
rect 5985 -1585 6000 -1565
rect 5950 -1615 6000 -1585
rect 5950 -1635 5965 -1615
rect 5985 -1635 6000 -1615
rect 5950 -1650 6000 -1635
rect 6100 -1650 6150 -950
rect 6250 -965 6300 -950
rect 6250 -985 6265 -965
rect 6285 -985 6300 -965
rect 6250 -1015 6300 -985
rect 6250 -1035 6265 -1015
rect 6285 -1035 6300 -1015
rect 6250 -1065 6300 -1035
rect 6250 -1085 6265 -1065
rect 6285 -1085 6300 -1065
rect 6250 -1115 6300 -1085
rect 6250 -1135 6265 -1115
rect 6285 -1135 6300 -1115
rect 6250 -1165 6300 -1135
rect 6250 -1185 6265 -1165
rect 6285 -1185 6300 -1165
rect 6250 -1215 6300 -1185
rect 6250 -1235 6265 -1215
rect 6285 -1235 6300 -1215
rect 6250 -1265 6300 -1235
rect 6250 -1285 6265 -1265
rect 6285 -1285 6300 -1265
rect 6250 -1315 6300 -1285
rect 6250 -1335 6265 -1315
rect 6285 -1335 6300 -1315
rect 6250 -1365 6300 -1335
rect 6250 -1385 6265 -1365
rect 6285 -1385 6300 -1365
rect 6250 -1415 6300 -1385
rect 6250 -1435 6265 -1415
rect 6285 -1435 6300 -1415
rect 6250 -1465 6300 -1435
rect 6250 -1485 6265 -1465
rect 6285 -1485 6300 -1465
rect 6250 -1515 6300 -1485
rect 6250 -1535 6265 -1515
rect 6285 -1535 6300 -1515
rect 6250 -1565 6300 -1535
rect 6250 -1585 6265 -1565
rect 6285 -1585 6300 -1565
rect 6250 -1615 6300 -1585
rect 6250 -1635 6265 -1615
rect 6285 -1635 6300 -1615
rect 6250 -1650 6300 -1635
rect 6400 -1650 6450 -950
rect 6550 -965 6600 -950
rect 6550 -985 6565 -965
rect 6585 -985 6600 -965
rect 6550 -1015 6600 -985
rect 6550 -1035 6565 -1015
rect 6585 -1035 6600 -1015
rect 6550 -1065 6600 -1035
rect 6550 -1085 6565 -1065
rect 6585 -1085 6600 -1065
rect 6550 -1115 6600 -1085
rect 6550 -1135 6565 -1115
rect 6585 -1135 6600 -1115
rect 6550 -1165 6600 -1135
rect 6550 -1185 6565 -1165
rect 6585 -1185 6600 -1165
rect 6550 -1215 6600 -1185
rect 6550 -1235 6565 -1215
rect 6585 -1235 6600 -1215
rect 6550 -1265 6600 -1235
rect 6550 -1285 6565 -1265
rect 6585 -1285 6600 -1265
rect 6550 -1315 6600 -1285
rect 6550 -1335 6565 -1315
rect 6585 -1335 6600 -1315
rect 6550 -1365 6600 -1335
rect 6550 -1385 6565 -1365
rect 6585 -1385 6600 -1365
rect 6550 -1415 6600 -1385
rect 6550 -1435 6565 -1415
rect 6585 -1435 6600 -1415
rect 6550 -1465 6600 -1435
rect 6550 -1485 6565 -1465
rect 6585 -1485 6600 -1465
rect 6550 -1515 6600 -1485
rect 6550 -1535 6565 -1515
rect 6585 -1535 6600 -1515
rect 6550 -1565 6600 -1535
rect 6550 -1585 6565 -1565
rect 6585 -1585 6600 -1565
rect 6550 -1615 6600 -1585
rect 6550 -1635 6565 -1615
rect 6585 -1635 6600 -1615
rect 6550 -1650 6600 -1635
rect 6700 -1650 6750 -950
rect 6850 -965 6900 -950
rect 6850 -985 6865 -965
rect 6885 -985 6900 -965
rect 6850 -1015 6900 -985
rect 6850 -1035 6865 -1015
rect 6885 -1035 6900 -1015
rect 6850 -1065 6900 -1035
rect 6850 -1085 6865 -1065
rect 6885 -1085 6900 -1065
rect 6850 -1115 6900 -1085
rect 6850 -1135 6865 -1115
rect 6885 -1135 6900 -1115
rect 6850 -1165 6900 -1135
rect 6850 -1185 6865 -1165
rect 6885 -1185 6900 -1165
rect 6850 -1215 6900 -1185
rect 6850 -1235 6865 -1215
rect 6885 -1235 6900 -1215
rect 6850 -1265 6900 -1235
rect 6850 -1285 6865 -1265
rect 6885 -1285 6900 -1265
rect 6850 -1315 6900 -1285
rect 6850 -1335 6865 -1315
rect 6885 -1335 6900 -1315
rect 6850 -1365 6900 -1335
rect 6850 -1385 6865 -1365
rect 6885 -1385 6900 -1365
rect 6850 -1415 6900 -1385
rect 6850 -1435 6865 -1415
rect 6885 -1435 6900 -1415
rect 6850 -1465 6900 -1435
rect 6850 -1485 6865 -1465
rect 6885 -1485 6900 -1465
rect 6850 -1515 6900 -1485
rect 6850 -1535 6865 -1515
rect 6885 -1535 6900 -1515
rect 6850 -1565 6900 -1535
rect 6850 -1585 6865 -1565
rect 6885 -1585 6900 -1565
rect 6850 -1615 6900 -1585
rect 6850 -1635 6865 -1615
rect 6885 -1635 6900 -1615
rect 6850 -1650 6900 -1635
rect 7000 -1650 7050 -950
rect 7150 -965 7200 -950
rect 7150 -985 7165 -965
rect 7185 -985 7200 -965
rect 7150 -1015 7200 -985
rect 7150 -1035 7165 -1015
rect 7185 -1035 7200 -1015
rect 7150 -1065 7200 -1035
rect 7150 -1085 7165 -1065
rect 7185 -1085 7200 -1065
rect 7150 -1115 7200 -1085
rect 7150 -1135 7165 -1115
rect 7185 -1135 7200 -1115
rect 7150 -1165 7200 -1135
rect 7150 -1185 7165 -1165
rect 7185 -1185 7200 -1165
rect 7150 -1215 7200 -1185
rect 7150 -1235 7165 -1215
rect 7185 -1235 7200 -1215
rect 7150 -1265 7200 -1235
rect 7150 -1285 7165 -1265
rect 7185 -1285 7200 -1265
rect 7150 -1315 7200 -1285
rect 7150 -1335 7165 -1315
rect 7185 -1335 7200 -1315
rect 7150 -1365 7200 -1335
rect 7150 -1385 7165 -1365
rect 7185 -1385 7200 -1365
rect 7150 -1415 7200 -1385
rect 7150 -1435 7165 -1415
rect 7185 -1435 7200 -1415
rect 7150 -1465 7200 -1435
rect 7150 -1485 7165 -1465
rect 7185 -1485 7200 -1465
rect 7150 -1515 7200 -1485
rect 7150 -1535 7165 -1515
rect 7185 -1535 7200 -1515
rect 7150 -1565 7200 -1535
rect 7150 -1585 7165 -1565
rect 7185 -1585 7200 -1565
rect 7150 -1615 7200 -1585
rect 7150 -1635 7165 -1615
rect 7185 -1635 7200 -1615
rect 7150 -1650 7200 -1635
rect 7300 -1650 7350 -950
rect 7450 -1650 7500 -950
rect 7600 -1650 7650 -950
rect 7750 -1650 7800 -950
rect 7900 -1650 7950 -950
rect 8050 -1650 8100 -950
rect 8200 -1650 8250 -950
rect 8350 -965 8400 -950
rect 8350 -985 8365 -965
rect 8385 -985 8400 -965
rect 8350 -1015 8400 -985
rect 8350 -1035 8365 -1015
rect 8385 -1035 8400 -1015
rect 8350 -1065 8400 -1035
rect 8350 -1085 8365 -1065
rect 8385 -1085 8400 -1065
rect 8350 -1115 8400 -1085
rect 8350 -1135 8365 -1115
rect 8385 -1135 8400 -1115
rect 8350 -1165 8400 -1135
rect 8350 -1185 8365 -1165
rect 8385 -1185 8400 -1165
rect 8350 -1215 8400 -1185
rect 8350 -1235 8365 -1215
rect 8385 -1235 8400 -1215
rect 8350 -1265 8400 -1235
rect 8350 -1285 8365 -1265
rect 8385 -1285 8400 -1265
rect 8350 -1315 8400 -1285
rect 8350 -1335 8365 -1315
rect 8385 -1335 8400 -1315
rect 8350 -1365 8400 -1335
rect 8350 -1385 8365 -1365
rect 8385 -1385 8400 -1365
rect 8350 -1415 8400 -1385
rect 8350 -1435 8365 -1415
rect 8385 -1435 8400 -1415
rect 8350 -1465 8400 -1435
rect 8350 -1485 8365 -1465
rect 8385 -1485 8400 -1465
rect 8350 -1515 8400 -1485
rect 8350 -1535 8365 -1515
rect 8385 -1535 8400 -1515
rect 8350 -1565 8400 -1535
rect 8350 -1585 8365 -1565
rect 8385 -1585 8400 -1565
rect 8350 -1615 8400 -1585
rect 8350 -1635 8365 -1615
rect 8385 -1635 8400 -1615
rect 8350 -1650 8400 -1635
rect 8500 -1650 8550 -950
rect 8650 -1650 8700 -950
rect 8800 -1650 8850 -950
rect 8950 -1650 9000 -950
rect 9100 -1650 9150 -950
rect 9250 -1650 9300 -950
rect 9400 -1650 9450 -950
rect 9550 -965 9600 -950
rect 9550 -985 9565 -965
rect 9585 -985 9600 -965
rect 9550 -1015 9600 -985
rect 9550 -1035 9565 -1015
rect 9585 -1035 9600 -1015
rect 9550 -1065 9600 -1035
rect 9550 -1085 9565 -1065
rect 9585 -1085 9600 -1065
rect 9550 -1115 9600 -1085
rect 9550 -1135 9565 -1115
rect 9585 -1135 9600 -1115
rect 9550 -1165 9600 -1135
rect 9550 -1185 9565 -1165
rect 9585 -1185 9600 -1165
rect 9550 -1215 9600 -1185
rect 9550 -1235 9565 -1215
rect 9585 -1235 9600 -1215
rect 9550 -1265 9600 -1235
rect 9550 -1285 9565 -1265
rect 9585 -1285 9600 -1265
rect 9550 -1315 9600 -1285
rect 9550 -1335 9565 -1315
rect 9585 -1335 9600 -1315
rect 9550 -1365 9600 -1335
rect 9550 -1385 9565 -1365
rect 9585 -1385 9600 -1365
rect 9550 -1415 9600 -1385
rect 9550 -1435 9565 -1415
rect 9585 -1435 9600 -1415
rect 9550 -1465 9600 -1435
rect 9550 -1485 9565 -1465
rect 9585 -1485 9600 -1465
rect 9550 -1515 9600 -1485
rect 9550 -1535 9565 -1515
rect 9585 -1535 9600 -1515
rect 9550 -1565 9600 -1535
rect 9550 -1585 9565 -1565
rect 9585 -1585 9600 -1565
rect 9550 -1615 9600 -1585
rect 9550 -1635 9565 -1615
rect 9585 -1635 9600 -1615
rect 9550 -1650 9600 -1635
rect 9700 -1650 9750 -950
rect 9850 -1650 9900 -950
rect 10000 -1650 10050 -950
rect 10150 -1650 10200 -950
rect 10300 -1650 10350 -950
rect 10450 -1650 10500 -950
rect 10600 -1650 10650 -950
rect 10750 -965 10800 -950
rect 10750 -985 10765 -965
rect 10785 -985 10800 -965
rect 10750 -1015 10800 -985
rect 10750 -1035 10765 -1015
rect 10785 -1035 10800 -1015
rect 10750 -1065 10800 -1035
rect 10750 -1085 10765 -1065
rect 10785 -1085 10800 -1065
rect 10750 -1115 10800 -1085
rect 10750 -1135 10765 -1115
rect 10785 -1135 10800 -1115
rect 10750 -1165 10800 -1135
rect 10750 -1185 10765 -1165
rect 10785 -1185 10800 -1165
rect 10750 -1215 10800 -1185
rect 10750 -1235 10765 -1215
rect 10785 -1235 10800 -1215
rect 10750 -1265 10800 -1235
rect 10750 -1285 10765 -1265
rect 10785 -1285 10800 -1265
rect 10750 -1315 10800 -1285
rect 10750 -1335 10765 -1315
rect 10785 -1335 10800 -1315
rect 10750 -1365 10800 -1335
rect 10750 -1385 10765 -1365
rect 10785 -1385 10800 -1365
rect 10750 -1415 10800 -1385
rect 10750 -1435 10765 -1415
rect 10785 -1435 10800 -1415
rect 10750 -1465 10800 -1435
rect 10750 -1485 10765 -1465
rect 10785 -1485 10800 -1465
rect 10750 -1515 10800 -1485
rect 10750 -1535 10765 -1515
rect 10785 -1535 10800 -1515
rect 10750 -1565 10800 -1535
rect 10750 -1585 10765 -1565
rect 10785 -1585 10800 -1565
rect 10750 -1615 10800 -1585
rect 10750 -1635 10765 -1615
rect 10785 -1635 10800 -1615
rect 10750 -1650 10800 -1635
rect 10900 -1650 10950 -950
rect 11050 -1650 11100 -950
rect 11200 -1650 11250 -950
rect 11350 -1650 11400 -950
rect 11500 -1650 11550 -950
rect 11650 -1650 11700 -950
rect 11800 -1650 11850 -950
rect 11950 -965 12000 -950
rect 11950 -985 11965 -965
rect 11985 -985 12000 -965
rect 11950 -1015 12000 -985
rect 11950 -1035 11965 -1015
rect 11985 -1035 12000 -1015
rect 11950 -1065 12000 -1035
rect 11950 -1085 11965 -1065
rect 11985 -1085 12000 -1065
rect 11950 -1115 12000 -1085
rect 11950 -1135 11965 -1115
rect 11985 -1135 12000 -1115
rect 11950 -1165 12000 -1135
rect 11950 -1185 11965 -1165
rect 11985 -1185 12000 -1165
rect 11950 -1215 12000 -1185
rect 11950 -1235 11965 -1215
rect 11985 -1235 12000 -1215
rect 11950 -1265 12000 -1235
rect 11950 -1285 11965 -1265
rect 11985 -1285 12000 -1265
rect 11950 -1315 12000 -1285
rect 11950 -1335 11965 -1315
rect 11985 -1335 12000 -1315
rect 11950 -1365 12000 -1335
rect 11950 -1385 11965 -1365
rect 11985 -1385 12000 -1365
rect 11950 -1415 12000 -1385
rect 11950 -1435 11965 -1415
rect 11985 -1435 12000 -1415
rect 11950 -1465 12000 -1435
rect 11950 -1485 11965 -1465
rect 11985 -1485 12000 -1465
rect 11950 -1515 12000 -1485
rect 11950 -1535 11965 -1515
rect 11985 -1535 12000 -1515
rect 11950 -1565 12000 -1535
rect 11950 -1585 11965 -1565
rect 11985 -1585 12000 -1565
rect 11950 -1615 12000 -1585
rect 11950 -1635 11965 -1615
rect 11985 -1635 12000 -1615
rect 11950 -1650 12000 -1635
rect 12100 -1650 12150 -950
rect 12250 -965 12300 -950
rect 12250 -985 12265 -965
rect 12285 -985 12300 -965
rect 12250 -1015 12300 -985
rect 12250 -1035 12265 -1015
rect 12285 -1035 12300 -1015
rect 12250 -1065 12300 -1035
rect 12250 -1085 12265 -1065
rect 12285 -1085 12300 -1065
rect 12250 -1115 12300 -1085
rect 12250 -1135 12265 -1115
rect 12285 -1135 12300 -1115
rect 12250 -1165 12300 -1135
rect 12250 -1185 12265 -1165
rect 12285 -1185 12300 -1165
rect 12250 -1215 12300 -1185
rect 12250 -1235 12265 -1215
rect 12285 -1235 12300 -1215
rect 12250 -1265 12300 -1235
rect 12250 -1285 12265 -1265
rect 12285 -1285 12300 -1265
rect 12250 -1315 12300 -1285
rect 12250 -1335 12265 -1315
rect 12285 -1335 12300 -1315
rect 12250 -1365 12300 -1335
rect 12250 -1385 12265 -1365
rect 12285 -1385 12300 -1365
rect 12250 -1415 12300 -1385
rect 12250 -1435 12265 -1415
rect 12285 -1435 12300 -1415
rect 12250 -1465 12300 -1435
rect 12250 -1485 12265 -1465
rect 12285 -1485 12300 -1465
rect 12250 -1515 12300 -1485
rect 12250 -1535 12265 -1515
rect 12285 -1535 12300 -1515
rect 12250 -1565 12300 -1535
rect 12250 -1585 12265 -1565
rect 12285 -1585 12300 -1565
rect 12250 -1615 12300 -1585
rect 12250 -1635 12265 -1615
rect 12285 -1635 12300 -1615
rect 12250 -1650 12300 -1635
rect 12400 -1650 12450 -950
rect 12550 -965 12600 -950
rect 12550 -985 12565 -965
rect 12585 -985 12600 -965
rect 12550 -1015 12600 -985
rect 12550 -1035 12565 -1015
rect 12585 -1035 12600 -1015
rect 12550 -1065 12600 -1035
rect 12550 -1085 12565 -1065
rect 12585 -1085 12600 -1065
rect 12550 -1115 12600 -1085
rect 12550 -1135 12565 -1115
rect 12585 -1135 12600 -1115
rect 12550 -1165 12600 -1135
rect 12550 -1185 12565 -1165
rect 12585 -1185 12600 -1165
rect 12550 -1215 12600 -1185
rect 12550 -1235 12565 -1215
rect 12585 -1235 12600 -1215
rect 12550 -1265 12600 -1235
rect 12550 -1285 12565 -1265
rect 12585 -1285 12600 -1265
rect 12550 -1315 12600 -1285
rect 12550 -1335 12565 -1315
rect 12585 -1335 12600 -1315
rect 12550 -1365 12600 -1335
rect 12550 -1385 12565 -1365
rect 12585 -1385 12600 -1365
rect 12550 -1415 12600 -1385
rect 12550 -1435 12565 -1415
rect 12585 -1435 12600 -1415
rect 12550 -1465 12600 -1435
rect 12550 -1485 12565 -1465
rect 12585 -1485 12600 -1465
rect 12550 -1515 12600 -1485
rect 12550 -1535 12565 -1515
rect 12585 -1535 12600 -1515
rect 12550 -1565 12600 -1535
rect 12550 -1585 12565 -1565
rect 12585 -1585 12600 -1565
rect 12550 -1615 12600 -1585
rect 12550 -1635 12565 -1615
rect 12585 -1635 12600 -1615
rect 12550 -1650 12600 -1635
rect 12700 -1650 12750 -950
rect 12850 -965 12900 -950
rect 12850 -985 12865 -965
rect 12885 -985 12900 -965
rect 12850 -1015 12900 -985
rect 12850 -1035 12865 -1015
rect 12885 -1035 12900 -1015
rect 12850 -1065 12900 -1035
rect 12850 -1085 12865 -1065
rect 12885 -1085 12900 -1065
rect 12850 -1115 12900 -1085
rect 12850 -1135 12865 -1115
rect 12885 -1135 12900 -1115
rect 12850 -1165 12900 -1135
rect 12850 -1185 12865 -1165
rect 12885 -1185 12900 -1165
rect 12850 -1215 12900 -1185
rect 12850 -1235 12865 -1215
rect 12885 -1235 12900 -1215
rect 12850 -1265 12900 -1235
rect 12850 -1285 12865 -1265
rect 12885 -1285 12900 -1265
rect 12850 -1315 12900 -1285
rect 12850 -1335 12865 -1315
rect 12885 -1335 12900 -1315
rect 12850 -1365 12900 -1335
rect 12850 -1385 12865 -1365
rect 12885 -1385 12900 -1365
rect 12850 -1415 12900 -1385
rect 12850 -1435 12865 -1415
rect 12885 -1435 12900 -1415
rect 12850 -1465 12900 -1435
rect 12850 -1485 12865 -1465
rect 12885 -1485 12900 -1465
rect 12850 -1515 12900 -1485
rect 12850 -1535 12865 -1515
rect 12885 -1535 12900 -1515
rect 12850 -1565 12900 -1535
rect 12850 -1585 12865 -1565
rect 12885 -1585 12900 -1565
rect 12850 -1615 12900 -1585
rect 12850 -1635 12865 -1615
rect 12885 -1635 12900 -1615
rect 12850 -1650 12900 -1635
rect 13000 -1650 13050 -950
rect 13150 -965 13200 -950
rect 13150 -985 13165 -965
rect 13185 -985 13200 -965
rect 13150 -1015 13200 -985
rect 13150 -1035 13165 -1015
rect 13185 -1035 13200 -1015
rect 13150 -1065 13200 -1035
rect 13150 -1085 13165 -1065
rect 13185 -1085 13200 -1065
rect 13150 -1115 13200 -1085
rect 13150 -1135 13165 -1115
rect 13185 -1135 13200 -1115
rect 13150 -1165 13200 -1135
rect 13150 -1185 13165 -1165
rect 13185 -1185 13200 -1165
rect 13150 -1215 13200 -1185
rect 13150 -1235 13165 -1215
rect 13185 -1235 13200 -1215
rect 13150 -1265 13200 -1235
rect 13150 -1285 13165 -1265
rect 13185 -1285 13200 -1265
rect 13150 -1315 13200 -1285
rect 13150 -1335 13165 -1315
rect 13185 -1335 13200 -1315
rect 13150 -1365 13200 -1335
rect 13150 -1385 13165 -1365
rect 13185 -1385 13200 -1365
rect 13150 -1415 13200 -1385
rect 13150 -1435 13165 -1415
rect 13185 -1435 13200 -1415
rect 13150 -1465 13200 -1435
rect 13150 -1485 13165 -1465
rect 13185 -1485 13200 -1465
rect 13150 -1515 13200 -1485
rect 13150 -1535 13165 -1515
rect 13185 -1535 13200 -1515
rect 13150 -1565 13200 -1535
rect 13150 -1585 13165 -1565
rect 13185 -1585 13200 -1565
rect 13150 -1615 13200 -1585
rect 13150 -1635 13165 -1615
rect 13185 -1635 13200 -1615
rect 13150 -1650 13200 -1635
rect 13300 -1650 13350 -950
rect 13450 -965 13500 -950
rect 13450 -985 13465 -965
rect 13485 -985 13500 -965
rect 13450 -1015 13500 -985
rect 13450 -1035 13465 -1015
rect 13485 -1035 13500 -1015
rect 13450 -1065 13500 -1035
rect 13450 -1085 13465 -1065
rect 13485 -1085 13500 -1065
rect 13450 -1115 13500 -1085
rect 13450 -1135 13465 -1115
rect 13485 -1135 13500 -1115
rect 13450 -1165 13500 -1135
rect 13450 -1185 13465 -1165
rect 13485 -1185 13500 -1165
rect 13450 -1215 13500 -1185
rect 13450 -1235 13465 -1215
rect 13485 -1235 13500 -1215
rect 13450 -1265 13500 -1235
rect 13450 -1285 13465 -1265
rect 13485 -1285 13500 -1265
rect 13450 -1315 13500 -1285
rect 13450 -1335 13465 -1315
rect 13485 -1335 13500 -1315
rect 13450 -1365 13500 -1335
rect 13450 -1385 13465 -1365
rect 13485 -1385 13500 -1365
rect 13450 -1415 13500 -1385
rect 13450 -1435 13465 -1415
rect 13485 -1435 13500 -1415
rect 13450 -1465 13500 -1435
rect 13450 -1485 13465 -1465
rect 13485 -1485 13500 -1465
rect 13450 -1515 13500 -1485
rect 13450 -1535 13465 -1515
rect 13485 -1535 13500 -1515
rect 13450 -1565 13500 -1535
rect 13450 -1585 13465 -1565
rect 13485 -1585 13500 -1565
rect 13450 -1615 13500 -1585
rect 13450 -1635 13465 -1615
rect 13485 -1635 13500 -1615
rect 13450 -1650 13500 -1635
rect 13600 -1650 13650 -950
rect 13750 -965 13800 -950
rect 13750 -985 13765 -965
rect 13785 -985 13800 -965
rect 13750 -1015 13800 -985
rect 13750 -1035 13765 -1015
rect 13785 -1035 13800 -1015
rect 13750 -1065 13800 -1035
rect 13750 -1085 13765 -1065
rect 13785 -1085 13800 -1065
rect 13750 -1115 13800 -1085
rect 13750 -1135 13765 -1115
rect 13785 -1135 13800 -1115
rect 13750 -1165 13800 -1135
rect 13750 -1185 13765 -1165
rect 13785 -1185 13800 -1165
rect 13750 -1215 13800 -1185
rect 13750 -1235 13765 -1215
rect 13785 -1235 13800 -1215
rect 13750 -1265 13800 -1235
rect 13750 -1285 13765 -1265
rect 13785 -1285 13800 -1265
rect 13750 -1315 13800 -1285
rect 13750 -1335 13765 -1315
rect 13785 -1335 13800 -1315
rect 13750 -1365 13800 -1335
rect 13750 -1385 13765 -1365
rect 13785 -1385 13800 -1365
rect 13750 -1415 13800 -1385
rect 13750 -1435 13765 -1415
rect 13785 -1435 13800 -1415
rect 13750 -1465 13800 -1435
rect 13750 -1485 13765 -1465
rect 13785 -1485 13800 -1465
rect 13750 -1515 13800 -1485
rect 13750 -1535 13765 -1515
rect 13785 -1535 13800 -1515
rect 13750 -1565 13800 -1535
rect 13750 -1585 13765 -1565
rect 13785 -1585 13800 -1565
rect 13750 -1615 13800 -1585
rect 13750 -1635 13765 -1615
rect 13785 -1635 13800 -1615
rect 13750 -1650 13800 -1635
rect 13900 -1650 13950 -950
rect 14050 -965 14100 -950
rect 14050 -985 14065 -965
rect 14085 -985 14100 -965
rect 14050 -1015 14100 -985
rect 14050 -1035 14065 -1015
rect 14085 -1035 14100 -1015
rect 14050 -1065 14100 -1035
rect 14050 -1085 14065 -1065
rect 14085 -1085 14100 -1065
rect 14050 -1115 14100 -1085
rect 14050 -1135 14065 -1115
rect 14085 -1135 14100 -1115
rect 14050 -1165 14100 -1135
rect 14050 -1185 14065 -1165
rect 14085 -1185 14100 -1165
rect 14050 -1215 14100 -1185
rect 14050 -1235 14065 -1215
rect 14085 -1235 14100 -1215
rect 14050 -1265 14100 -1235
rect 14050 -1285 14065 -1265
rect 14085 -1285 14100 -1265
rect 14050 -1315 14100 -1285
rect 14050 -1335 14065 -1315
rect 14085 -1335 14100 -1315
rect 14050 -1365 14100 -1335
rect 14050 -1385 14065 -1365
rect 14085 -1385 14100 -1365
rect 14050 -1415 14100 -1385
rect 14050 -1435 14065 -1415
rect 14085 -1435 14100 -1415
rect 14050 -1465 14100 -1435
rect 14050 -1485 14065 -1465
rect 14085 -1485 14100 -1465
rect 14050 -1515 14100 -1485
rect 14050 -1535 14065 -1515
rect 14085 -1535 14100 -1515
rect 14050 -1565 14100 -1535
rect 14050 -1585 14065 -1565
rect 14085 -1585 14100 -1565
rect 14050 -1615 14100 -1585
rect 14050 -1635 14065 -1615
rect 14085 -1635 14100 -1615
rect 14050 -1650 14100 -1635
rect 14200 -1650 14250 -950
rect 14350 -965 14400 -950
rect 14350 -985 14365 -965
rect 14385 -985 14400 -965
rect 14350 -1015 14400 -985
rect 14350 -1035 14365 -1015
rect 14385 -1035 14400 -1015
rect 14350 -1065 14400 -1035
rect 14350 -1085 14365 -1065
rect 14385 -1085 14400 -1065
rect 14350 -1115 14400 -1085
rect 14350 -1135 14365 -1115
rect 14385 -1135 14400 -1115
rect 14350 -1165 14400 -1135
rect 14350 -1185 14365 -1165
rect 14385 -1185 14400 -1165
rect 14350 -1215 14400 -1185
rect 14350 -1235 14365 -1215
rect 14385 -1235 14400 -1215
rect 14350 -1265 14400 -1235
rect 14350 -1285 14365 -1265
rect 14385 -1285 14400 -1265
rect 14350 -1315 14400 -1285
rect 14350 -1335 14365 -1315
rect 14385 -1335 14400 -1315
rect 14350 -1365 14400 -1335
rect 14350 -1385 14365 -1365
rect 14385 -1385 14400 -1365
rect 14350 -1415 14400 -1385
rect 14350 -1435 14365 -1415
rect 14385 -1435 14400 -1415
rect 14350 -1465 14400 -1435
rect 14350 -1485 14365 -1465
rect 14385 -1485 14400 -1465
rect 14350 -1515 14400 -1485
rect 14350 -1535 14365 -1515
rect 14385 -1535 14400 -1515
rect 14350 -1565 14400 -1535
rect 14350 -1585 14365 -1565
rect 14385 -1585 14400 -1565
rect 14350 -1615 14400 -1585
rect 14350 -1635 14365 -1615
rect 14385 -1635 14400 -1615
rect 14350 -1650 14400 -1635
rect 14500 -1650 14550 -950
rect 14650 -1650 14700 -950
rect 14800 -1650 14850 -950
rect 14950 -1650 15000 -950
rect 15100 -1650 15150 -950
rect 15250 -1650 15300 -950
rect 15400 -1650 15450 -950
rect 15550 -965 15600 -950
rect 15550 -985 15565 -965
rect 15585 -985 15600 -965
rect 15550 -1015 15600 -985
rect 15550 -1035 15565 -1015
rect 15585 -1035 15600 -1015
rect 15550 -1065 15600 -1035
rect 15550 -1085 15565 -1065
rect 15585 -1085 15600 -1065
rect 15550 -1115 15600 -1085
rect 15550 -1135 15565 -1115
rect 15585 -1135 15600 -1115
rect 15550 -1165 15600 -1135
rect 15550 -1185 15565 -1165
rect 15585 -1185 15600 -1165
rect 15550 -1215 15600 -1185
rect 15550 -1235 15565 -1215
rect 15585 -1235 15600 -1215
rect 15550 -1265 15600 -1235
rect 15550 -1285 15565 -1265
rect 15585 -1285 15600 -1265
rect 15550 -1315 15600 -1285
rect 15550 -1335 15565 -1315
rect 15585 -1335 15600 -1315
rect 15550 -1365 15600 -1335
rect 15550 -1385 15565 -1365
rect 15585 -1385 15600 -1365
rect 15550 -1415 15600 -1385
rect 15550 -1435 15565 -1415
rect 15585 -1435 15600 -1415
rect 15550 -1465 15600 -1435
rect 15550 -1485 15565 -1465
rect 15585 -1485 15600 -1465
rect 15550 -1515 15600 -1485
rect 15550 -1535 15565 -1515
rect 15585 -1535 15600 -1515
rect 15550 -1565 15600 -1535
rect 15550 -1585 15565 -1565
rect 15585 -1585 15600 -1565
rect 15550 -1615 15600 -1585
rect 15550 -1635 15565 -1615
rect 15585 -1635 15600 -1615
rect 15550 -1650 15600 -1635
rect 15700 -1650 15750 -950
rect 15850 -1650 15900 -950
rect 16000 -1650 16050 -950
rect 16150 -1650 16200 -950
rect 16300 -1650 16350 -950
rect 16450 -1650 16500 -950
rect 16600 -1650 16650 -950
rect 16750 -965 16800 -950
rect 16750 -985 16765 -965
rect 16785 -985 16800 -965
rect 16750 -1015 16800 -985
rect 16750 -1035 16765 -1015
rect 16785 -1035 16800 -1015
rect 16750 -1065 16800 -1035
rect 16750 -1085 16765 -1065
rect 16785 -1085 16800 -1065
rect 16750 -1115 16800 -1085
rect 16750 -1135 16765 -1115
rect 16785 -1135 16800 -1115
rect 16750 -1165 16800 -1135
rect 16750 -1185 16765 -1165
rect 16785 -1185 16800 -1165
rect 16750 -1215 16800 -1185
rect 16750 -1235 16765 -1215
rect 16785 -1235 16800 -1215
rect 16750 -1265 16800 -1235
rect 16750 -1285 16765 -1265
rect 16785 -1285 16800 -1265
rect 16750 -1315 16800 -1285
rect 16750 -1335 16765 -1315
rect 16785 -1335 16800 -1315
rect 16750 -1365 16800 -1335
rect 16750 -1385 16765 -1365
rect 16785 -1385 16800 -1365
rect 16750 -1415 16800 -1385
rect 16750 -1435 16765 -1415
rect 16785 -1435 16800 -1415
rect 16750 -1465 16800 -1435
rect 16750 -1485 16765 -1465
rect 16785 -1485 16800 -1465
rect 16750 -1515 16800 -1485
rect 16750 -1535 16765 -1515
rect 16785 -1535 16800 -1515
rect 16750 -1565 16800 -1535
rect 16750 -1585 16765 -1565
rect 16785 -1585 16800 -1565
rect 16750 -1615 16800 -1585
rect 16750 -1635 16765 -1615
rect 16785 -1635 16800 -1615
rect 16750 -1650 16800 -1635
rect 16900 -1650 16950 -950
rect 17050 -1650 17100 -950
rect 17200 -1650 17250 -950
rect 17350 -1650 17400 -950
rect 17500 -1650 17550 -950
rect 17650 -1650 17700 -950
rect 17800 -1650 17850 -950
rect 17950 -965 18000 -950
rect 17950 -985 17965 -965
rect 17985 -985 18000 -965
rect 17950 -1015 18000 -985
rect 17950 -1035 17965 -1015
rect 17985 -1035 18000 -1015
rect 17950 -1065 18000 -1035
rect 17950 -1085 17965 -1065
rect 17985 -1085 18000 -1065
rect 17950 -1115 18000 -1085
rect 17950 -1135 17965 -1115
rect 17985 -1135 18000 -1115
rect 17950 -1165 18000 -1135
rect 17950 -1185 17965 -1165
rect 17985 -1185 18000 -1165
rect 17950 -1215 18000 -1185
rect 17950 -1235 17965 -1215
rect 17985 -1235 18000 -1215
rect 17950 -1265 18000 -1235
rect 17950 -1285 17965 -1265
rect 17985 -1285 18000 -1265
rect 17950 -1315 18000 -1285
rect 17950 -1335 17965 -1315
rect 17985 -1335 18000 -1315
rect 17950 -1365 18000 -1335
rect 17950 -1385 17965 -1365
rect 17985 -1385 18000 -1365
rect 17950 -1415 18000 -1385
rect 17950 -1435 17965 -1415
rect 17985 -1435 18000 -1415
rect 17950 -1465 18000 -1435
rect 17950 -1485 17965 -1465
rect 17985 -1485 18000 -1465
rect 17950 -1515 18000 -1485
rect 17950 -1535 17965 -1515
rect 17985 -1535 18000 -1515
rect 17950 -1565 18000 -1535
rect 17950 -1585 17965 -1565
rect 17985 -1585 18000 -1565
rect 17950 -1615 18000 -1585
rect 17950 -1635 17965 -1615
rect 17985 -1635 18000 -1615
rect 17950 -1650 18000 -1635
rect 18100 -1650 18150 -950
rect 18250 -1650 18300 -950
rect 18400 -1650 18450 -950
rect 18550 -1650 18600 -950
rect 18700 -1650 18750 -950
rect 18850 -1650 18900 -950
rect 19000 -1650 19050 -950
rect 19150 -965 19200 -950
rect 19150 -985 19165 -965
rect 19185 -985 19200 -965
rect 19150 -1015 19200 -985
rect 19150 -1035 19165 -1015
rect 19185 -1035 19200 -1015
rect 19150 -1065 19200 -1035
rect 19150 -1085 19165 -1065
rect 19185 -1085 19200 -1065
rect 19150 -1115 19200 -1085
rect 19150 -1135 19165 -1115
rect 19185 -1135 19200 -1115
rect 19150 -1165 19200 -1135
rect 19150 -1185 19165 -1165
rect 19185 -1185 19200 -1165
rect 19150 -1215 19200 -1185
rect 19150 -1235 19165 -1215
rect 19185 -1235 19200 -1215
rect 19150 -1265 19200 -1235
rect 19150 -1285 19165 -1265
rect 19185 -1285 19200 -1265
rect 19150 -1315 19200 -1285
rect 19150 -1335 19165 -1315
rect 19185 -1335 19200 -1315
rect 19150 -1365 19200 -1335
rect 19150 -1385 19165 -1365
rect 19185 -1385 19200 -1365
rect 19150 -1415 19200 -1385
rect 19150 -1435 19165 -1415
rect 19185 -1435 19200 -1415
rect 19150 -1465 19200 -1435
rect 19150 -1485 19165 -1465
rect 19185 -1485 19200 -1465
rect 19150 -1515 19200 -1485
rect 19150 -1535 19165 -1515
rect 19185 -1535 19200 -1515
rect 19150 -1565 19200 -1535
rect 19150 -1585 19165 -1565
rect 19185 -1585 19200 -1565
rect 19150 -1615 19200 -1585
rect 19150 -1635 19165 -1615
rect 19185 -1635 19200 -1615
rect 19150 -1650 19200 -1635
rect 19300 -1650 19350 -950
rect 19450 -1650 19500 -950
rect 19600 -1650 19650 -950
rect 19750 -1650 19800 -950
rect 19900 -1650 19950 -950
rect 20050 -1650 20100 -950
rect 20200 -1650 20250 -950
rect 20350 -965 20400 -950
rect 20350 -985 20365 -965
rect 20385 -985 20400 -965
rect 20350 -1015 20400 -985
rect 20350 -1035 20365 -1015
rect 20385 -1035 20400 -1015
rect 20350 -1065 20400 -1035
rect 20350 -1085 20365 -1065
rect 20385 -1085 20400 -1065
rect 20350 -1115 20400 -1085
rect 20350 -1135 20365 -1115
rect 20385 -1135 20400 -1115
rect 20350 -1165 20400 -1135
rect 20350 -1185 20365 -1165
rect 20385 -1185 20400 -1165
rect 20350 -1215 20400 -1185
rect 20350 -1235 20365 -1215
rect 20385 -1235 20400 -1215
rect 20350 -1265 20400 -1235
rect 20350 -1285 20365 -1265
rect 20385 -1285 20400 -1265
rect 20350 -1315 20400 -1285
rect 20350 -1335 20365 -1315
rect 20385 -1335 20400 -1315
rect 20350 -1365 20400 -1335
rect 20350 -1385 20365 -1365
rect 20385 -1385 20400 -1365
rect 20350 -1415 20400 -1385
rect 20350 -1435 20365 -1415
rect 20385 -1435 20400 -1415
rect 20350 -1465 20400 -1435
rect 20350 -1485 20365 -1465
rect 20385 -1485 20400 -1465
rect 20350 -1515 20400 -1485
rect 20350 -1535 20365 -1515
rect 20385 -1535 20400 -1515
rect 20350 -1565 20400 -1535
rect 20350 -1585 20365 -1565
rect 20385 -1585 20400 -1565
rect 20350 -1615 20400 -1585
rect 20350 -1635 20365 -1615
rect 20385 -1635 20400 -1615
rect 20350 -1650 20400 -1635
<< mvpdiff >>
rect -650 5085 -600 5100
rect -650 5065 -635 5085
rect -615 5065 -600 5085
rect -650 5035 -600 5065
rect -650 5015 -635 5035
rect -615 5015 -600 5035
rect -650 4985 -600 5015
rect -650 4965 -635 4985
rect -615 4965 -600 4985
rect -650 4935 -600 4965
rect -650 4915 -635 4935
rect -615 4915 -600 4935
rect -650 4885 -600 4915
rect -650 4865 -635 4885
rect -615 4865 -600 4885
rect -650 4835 -600 4865
rect -650 4815 -635 4835
rect -615 4815 -600 4835
rect -650 4785 -600 4815
rect -650 4765 -635 4785
rect -615 4765 -600 4785
rect -650 4735 -600 4765
rect -650 4715 -635 4735
rect -615 4715 -600 4735
rect -650 4685 -600 4715
rect -650 4665 -635 4685
rect -615 4665 -600 4685
rect -650 4635 -600 4665
rect -650 4615 -635 4635
rect -615 4615 -600 4635
rect -650 4600 -600 4615
rect -500 5085 -450 5100
rect -500 5065 -485 5085
rect -465 5065 -450 5085
rect -500 5035 -450 5065
rect -500 5015 -485 5035
rect -465 5015 -450 5035
rect -500 4985 -450 5015
rect -500 4965 -485 4985
rect -465 4965 -450 4985
rect -500 4935 -450 4965
rect -500 4915 -485 4935
rect -465 4915 -450 4935
rect -500 4885 -450 4915
rect -500 4865 -485 4885
rect -465 4865 -450 4885
rect -500 4835 -450 4865
rect -500 4815 -485 4835
rect -465 4815 -450 4835
rect -500 4785 -450 4815
rect -500 4765 -485 4785
rect -465 4765 -450 4785
rect -500 4735 -450 4765
rect -500 4715 -485 4735
rect -465 4715 -450 4735
rect -500 4685 -450 4715
rect -500 4665 -485 4685
rect -465 4665 -450 4685
rect -500 4635 -450 4665
rect -500 4615 -485 4635
rect -465 4615 -450 4635
rect -500 4600 -450 4615
rect -350 5085 -300 5100
rect -350 5065 -335 5085
rect -315 5065 -300 5085
rect -350 5035 -300 5065
rect -350 5015 -335 5035
rect -315 5015 -300 5035
rect -350 4985 -300 5015
rect -350 4965 -335 4985
rect -315 4965 -300 4985
rect -350 4935 -300 4965
rect -350 4915 -335 4935
rect -315 4915 -300 4935
rect -350 4885 -300 4915
rect -350 4865 -335 4885
rect -315 4865 -300 4885
rect -350 4835 -300 4865
rect -350 4815 -335 4835
rect -315 4815 -300 4835
rect -350 4785 -300 4815
rect -350 4765 -335 4785
rect -315 4765 -300 4785
rect -350 4735 -300 4765
rect -350 4715 -335 4735
rect -315 4715 -300 4735
rect -350 4685 -300 4715
rect -350 4665 -335 4685
rect -315 4665 -300 4685
rect -350 4635 -300 4665
rect -350 4615 -335 4635
rect -315 4615 -300 4635
rect -350 4600 -300 4615
rect -200 5085 -150 5100
rect -200 5065 -185 5085
rect -165 5065 -150 5085
rect -200 5035 -150 5065
rect -200 5015 -185 5035
rect -165 5015 -150 5035
rect -200 4985 -150 5015
rect -200 4965 -185 4985
rect -165 4965 -150 4985
rect -200 4935 -150 4965
rect -200 4915 -185 4935
rect -165 4915 -150 4935
rect -200 4885 -150 4915
rect -200 4865 -185 4885
rect -165 4865 -150 4885
rect -200 4835 -150 4865
rect -200 4815 -185 4835
rect -165 4815 -150 4835
rect -200 4785 -150 4815
rect -200 4765 -185 4785
rect -165 4765 -150 4785
rect -200 4735 -150 4765
rect -200 4715 -185 4735
rect -165 4715 -150 4735
rect -200 4685 -150 4715
rect -200 4665 -185 4685
rect -165 4665 -150 4685
rect -200 4635 -150 4665
rect -200 4615 -185 4635
rect -165 4615 -150 4635
rect -200 4600 -150 4615
rect -50 5085 0 5100
rect -50 5065 -35 5085
rect -15 5065 0 5085
rect -50 5035 0 5065
rect -50 5015 -35 5035
rect -15 5015 0 5035
rect -50 4985 0 5015
rect -50 4965 -35 4985
rect -15 4965 0 4985
rect -50 4935 0 4965
rect -50 4915 -35 4935
rect -15 4915 0 4935
rect -50 4885 0 4915
rect -50 4865 -35 4885
rect -15 4865 0 4885
rect -50 4835 0 4865
rect -50 4815 -35 4835
rect -15 4815 0 4835
rect -50 4785 0 4815
rect -50 4765 -35 4785
rect -15 4765 0 4785
rect -50 4735 0 4765
rect -50 4715 -35 4735
rect -15 4715 0 4735
rect -50 4685 0 4715
rect -50 4665 -35 4685
rect -15 4665 0 4685
rect -50 4635 0 4665
rect -50 4615 -35 4635
rect -15 4615 0 4635
rect -50 4600 0 4615
rect 100 4600 150 5100
rect 250 4600 300 5100
rect 400 4600 450 5100
rect 550 5085 600 5100
rect 550 5065 565 5085
rect 585 5065 600 5085
rect 550 5035 600 5065
rect 550 5015 565 5035
rect 585 5015 600 5035
rect 550 4985 600 5015
rect 550 4965 565 4985
rect 585 4965 600 4985
rect 550 4935 600 4965
rect 550 4915 565 4935
rect 585 4915 600 4935
rect 550 4885 600 4915
rect 550 4865 565 4885
rect 585 4865 600 4885
rect 550 4835 600 4865
rect 550 4815 565 4835
rect 585 4815 600 4835
rect 550 4785 600 4815
rect 550 4765 565 4785
rect 585 4765 600 4785
rect 550 4735 600 4765
rect 550 4715 565 4735
rect 585 4715 600 4735
rect 550 4685 600 4715
rect 550 4665 565 4685
rect 585 4665 600 4685
rect 550 4635 600 4665
rect 550 4615 565 4635
rect 585 4615 600 4635
rect 550 4600 600 4615
rect 700 5085 750 5100
rect 700 5065 715 5085
rect 735 5065 750 5085
rect 700 5035 750 5065
rect 700 5015 715 5035
rect 735 5015 750 5035
rect 700 4985 750 5015
rect 700 4965 715 4985
rect 735 4965 750 4985
rect 700 4935 750 4965
rect 700 4915 715 4935
rect 735 4915 750 4935
rect 700 4885 750 4915
rect 700 4865 715 4885
rect 735 4865 750 4885
rect 700 4835 750 4865
rect 700 4815 715 4835
rect 735 4815 750 4835
rect 700 4785 750 4815
rect 700 4765 715 4785
rect 735 4765 750 4785
rect 700 4735 750 4765
rect 700 4715 715 4735
rect 735 4715 750 4735
rect 700 4685 750 4715
rect 700 4665 715 4685
rect 735 4665 750 4685
rect 700 4635 750 4665
rect 700 4615 715 4635
rect 735 4615 750 4635
rect 700 4600 750 4615
rect 850 5085 900 5100
rect 850 5065 865 5085
rect 885 5065 900 5085
rect 850 5035 900 5065
rect 850 5015 865 5035
rect 885 5015 900 5035
rect 850 4985 900 5015
rect 850 4965 865 4985
rect 885 4965 900 4985
rect 850 4935 900 4965
rect 850 4915 865 4935
rect 885 4915 900 4935
rect 850 4885 900 4915
rect 850 4865 865 4885
rect 885 4865 900 4885
rect 850 4835 900 4865
rect 850 4815 865 4835
rect 885 4815 900 4835
rect 850 4785 900 4815
rect 850 4765 865 4785
rect 885 4765 900 4785
rect 850 4735 900 4765
rect 850 4715 865 4735
rect 885 4715 900 4735
rect 850 4685 900 4715
rect 850 4665 865 4685
rect 885 4665 900 4685
rect 850 4635 900 4665
rect 850 4615 865 4635
rect 885 4615 900 4635
rect 850 4600 900 4615
rect 1000 5085 1050 5100
rect 1000 5065 1015 5085
rect 1035 5065 1050 5085
rect 1000 5035 1050 5065
rect 1000 5015 1015 5035
rect 1035 5015 1050 5035
rect 1000 4985 1050 5015
rect 1000 4965 1015 4985
rect 1035 4965 1050 4985
rect 1000 4935 1050 4965
rect 1000 4915 1015 4935
rect 1035 4915 1050 4935
rect 1000 4885 1050 4915
rect 1000 4865 1015 4885
rect 1035 4865 1050 4885
rect 1000 4835 1050 4865
rect 1000 4815 1015 4835
rect 1035 4815 1050 4835
rect 1000 4785 1050 4815
rect 1000 4765 1015 4785
rect 1035 4765 1050 4785
rect 1000 4735 1050 4765
rect 1000 4715 1015 4735
rect 1035 4715 1050 4735
rect 1000 4685 1050 4715
rect 1000 4665 1015 4685
rect 1035 4665 1050 4685
rect 1000 4635 1050 4665
rect 1000 4615 1015 4635
rect 1035 4615 1050 4635
rect 1000 4600 1050 4615
rect 1150 5085 1200 5100
rect 1150 5065 1165 5085
rect 1185 5065 1200 5085
rect 1150 5035 1200 5065
rect 1150 5015 1165 5035
rect 1185 5015 1200 5035
rect 1150 4985 1200 5015
rect 1150 4965 1165 4985
rect 1185 4965 1200 4985
rect 1150 4935 1200 4965
rect 1150 4915 1165 4935
rect 1185 4915 1200 4935
rect 1150 4885 1200 4915
rect 1150 4865 1165 4885
rect 1185 4865 1200 4885
rect 1150 4835 1200 4865
rect 1150 4815 1165 4835
rect 1185 4815 1200 4835
rect 1150 4785 1200 4815
rect 1150 4765 1165 4785
rect 1185 4765 1200 4785
rect 1150 4735 1200 4765
rect 1150 4715 1165 4735
rect 1185 4715 1200 4735
rect 1150 4685 1200 4715
rect 1150 4665 1165 4685
rect 1185 4665 1200 4685
rect 1150 4635 1200 4665
rect 1150 4615 1165 4635
rect 1185 4615 1200 4635
rect 1150 4600 1200 4615
rect 1300 5085 1350 5100
rect 1300 5065 1315 5085
rect 1335 5065 1350 5085
rect 1300 5035 1350 5065
rect 1300 5015 1315 5035
rect 1335 5015 1350 5035
rect 1300 4985 1350 5015
rect 1300 4965 1315 4985
rect 1335 4965 1350 4985
rect 1300 4935 1350 4965
rect 1300 4915 1315 4935
rect 1335 4915 1350 4935
rect 1300 4885 1350 4915
rect 1300 4865 1315 4885
rect 1335 4865 1350 4885
rect 1300 4835 1350 4865
rect 1300 4815 1315 4835
rect 1335 4815 1350 4835
rect 1300 4785 1350 4815
rect 1300 4765 1315 4785
rect 1335 4765 1350 4785
rect 1300 4735 1350 4765
rect 1300 4715 1315 4735
rect 1335 4715 1350 4735
rect 1300 4685 1350 4715
rect 1300 4665 1315 4685
rect 1335 4665 1350 4685
rect 1300 4635 1350 4665
rect 1300 4615 1315 4635
rect 1335 4615 1350 4635
rect 1300 4600 1350 4615
rect 1450 5085 1500 5100
rect 1450 5065 1465 5085
rect 1485 5065 1500 5085
rect 1450 5035 1500 5065
rect 1450 5015 1465 5035
rect 1485 5015 1500 5035
rect 1450 4985 1500 5015
rect 1450 4965 1465 4985
rect 1485 4965 1500 4985
rect 1450 4935 1500 4965
rect 1450 4915 1465 4935
rect 1485 4915 1500 4935
rect 1450 4885 1500 4915
rect 1450 4865 1465 4885
rect 1485 4865 1500 4885
rect 1450 4835 1500 4865
rect 1450 4815 1465 4835
rect 1485 4815 1500 4835
rect 1450 4785 1500 4815
rect 1450 4765 1465 4785
rect 1485 4765 1500 4785
rect 1450 4735 1500 4765
rect 1450 4715 1465 4735
rect 1485 4715 1500 4735
rect 1450 4685 1500 4715
rect 1450 4665 1465 4685
rect 1485 4665 1500 4685
rect 1450 4635 1500 4665
rect 1450 4615 1465 4635
rect 1485 4615 1500 4635
rect 1450 4600 1500 4615
rect 1600 5085 1650 5100
rect 1600 5065 1615 5085
rect 1635 5065 1650 5085
rect 1600 5035 1650 5065
rect 1600 5015 1615 5035
rect 1635 5015 1650 5035
rect 1600 4985 1650 5015
rect 1600 4965 1615 4985
rect 1635 4965 1650 4985
rect 1600 4935 1650 4965
rect 1600 4915 1615 4935
rect 1635 4915 1650 4935
rect 1600 4885 1650 4915
rect 1600 4865 1615 4885
rect 1635 4865 1650 4885
rect 1600 4835 1650 4865
rect 1600 4815 1615 4835
rect 1635 4815 1650 4835
rect 1600 4785 1650 4815
rect 1600 4765 1615 4785
rect 1635 4765 1650 4785
rect 1600 4735 1650 4765
rect 1600 4715 1615 4735
rect 1635 4715 1650 4735
rect 1600 4685 1650 4715
rect 1600 4665 1615 4685
rect 1635 4665 1650 4685
rect 1600 4635 1650 4665
rect 1600 4615 1615 4635
rect 1635 4615 1650 4635
rect 1600 4600 1650 4615
rect 1750 5085 1800 5100
rect 1750 5065 1765 5085
rect 1785 5065 1800 5085
rect 1750 5035 1800 5065
rect 1750 5015 1765 5035
rect 1785 5015 1800 5035
rect 1750 4985 1800 5015
rect 1750 4965 1765 4985
rect 1785 4965 1800 4985
rect 1750 4935 1800 4965
rect 1750 4915 1765 4935
rect 1785 4915 1800 4935
rect 1750 4885 1800 4915
rect 1750 4865 1765 4885
rect 1785 4865 1800 4885
rect 1750 4835 1800 4865
rect 1750 4815 1765 4835
rect 1785 4815 1800 4835
rect 1750 4785 1800 4815
rect 1750 4765 1765 4785
rect 1785 4765 1800 4785
rect 1750 4735 1800 4765
rect 1750 4715 1765 4735
rect 1785 4715 1800 4735
rect 1750 4685 1800 4715
rect 1750 4665 1765 4685
rect 1785 4665 1800 4685
rect 1750 4635 1800 4665
rect 1750 4615 1765 4635
rect 1785 4615 1800 4635
rect 1750 4600 1800 4615
rect 1900 5085 1950 5100
rect 1900 5065 1915 5085
rect 1935 5065 1950 5085
rect 1900 5035 1950 5065
rect 1900 5015 1915 5035
rect 1935 5015 1950 5035
rect 1900 4985 1950 5015
rect 1900 4965 1915 4985
rect 1935 4965 1950 4985
rect 1900 4935 1950 4965
rect 1900 4915 1915 4935
rect 1935 4915 1950 4935
rect 1900 4885 1950 4915
rect 1900 4865 1915 4885
rect 1935 4865 1950 4885
rect 1900 4835 1950 4865
rect 1900 4815 1915 4835
rect 1935 4815 1950 4835
rect 1900 4785 1950 4815
rect 1900 4765 1915 4785
rect 1935 4765 1950 4785
rect 1900 4735 1950 4765
rect 1900 4715 1915 4735
rect 1935 4715 1950 4735
rect 1900 4685 1950 4715
rect 1900 4665 1915 4685
rect 1935 4665 1950 4685
rect 1900 4635 1950 4665
rect 1900 4615 1915 4635
rect 1935 4615 1950 4635
rect 1900 4600 1950 4615
rect 2050 5085 2100 5100
rect 2050 5065 2065 5085
rect 2085 5065 2100 5085
rect 2050 5035 2100 5065
rect 2050 5015 2065 5035
rect 2085 5015 2100 5035
rect 2050 4985 2100 5015
rect 2050 4965 2065 4985
rect 2085 4965 2100 4985
rect 2050 4935 2100 4965
rect 2050 4915 2065 4935
rect 2085 4915 2100 4935
rect 2050 4885 2100 4915
rect 2050 4865 2065 4885
rect 2085 4865 2100 4885
rect 2050 4835 2100 4865
rect 2050 4815 2065 4835
rect 2085 4815 2100 4835
rect 2050 4785 2100 4815
rect 2050 4765 2065 4785
rect 2085 4765 2100 4785
rect 2050 4735 2100 4765
rect 2050 4715 2065 4735
rect 2085 4715 2100 4735
rect 2050 4685 2100 4715
rect 2050 4665 2065 4685
rect 2085 4665 2100 4685
rect 2050 4635 2100 4665
rect 2050 4615 2065 4635
rect 2085 4615 2100 4635
rect 2050 4600 2100 4615
rect 2200 5085 2250 5100
rect 2200 5065 2215 5085
rect 2235 5065 2250 5085
rect 2200 5035 2250 5065
rect 2200 5015 2215 5035
rect 2235 5015 2250 5035
rect 2200 4985 2250 5015
rect 2200 4965 2215 4985
rect 2235 4965 2250 4985
rect 2200 4935 2250 4965
rect 2200 4915 2215 4935
rect 2235 4915 2250 4935
rect 2200 4885 2250 4915
rect 2200 4865 2215 4885
rect 2235 4865 2250 4885
rect 2200 4835 2250 4865
rect 2200 4815 2215 4835
rect 2235 4815 2250 4835
rect 2200 4785 2250 4815
rect 2200 4765 2215 4785
rect 2235 4765 2250 4785
rect 2200 4735 2250 4765
rect 2200 4715 2215 4735
rect 2235 4715 2250 4735
rect 2200 4685 2250 4715
rect 2200 4665 2215 4685
rect 2235 4665 2250 4685
rect 2200 4635 2250 4665
rect 2200 4615 2215 4635
rect 2235 4615 2250 4635
rect 2200 4600 2250 4615
rect 2350 5085 2400 5100
rect 2350 5065 2365 5085
rect 2385 5065 2400 5085
rect 2350 5035 2400 5065
rect 2350 5015 2365 5035
rect 2385 5015 2400 5035
rect 2350 4985 2400 5015
rect 2350 4965 2365 4985
rect 2385 4965 2400 4985
rect 2350 4935 2400 4965
rect 2350 4915 2365 4935
rect 2385 4915 2400 4935
rect 2350 4885 2400 4915
rect 2350 4865 2365 4885
rect 2385 4865 2400 4885
rect 2350 4835 2400 4865
rect 2350 4815 2365 4835
rect 2385 4815 2400 4835
rect 2350 4785 2400 4815
rect 2350 4765 2365 4785
rect 2385 4765 2400 4785
rect 2350 4735 2400 4765
rect 2350 4715 2365 4735
rect 2385 4715 2400 4735
rect 2350 4685 2400 4715
rect 2350 4665 2365 4685
rect 2385 4665 2400 4685
rect 2350 4635 2400 4665
rect 2350 4615 2365 4635
rect 2385 4615 2400 4635
rect 2350 4600 2400 4615
rect 2500 5085 2550 5100
rect 2500 5065 2515 5085
rect 2535 5065 2550 5085
rect 2500 5035 2550 5065
rect 2500 5015 2515 5035
rect 2535 5015 2550 5035
rect 2500 4985 2550 5015
rect 2500 4965 2515 4985
rect 2535 4965 2550 4985
rect 2500 4935 2550 4965
rect 2500 4915 2515 4935
rect 2535 4915 2550 4935
rect 2500 4885 2550 4915
rect 2500 4865 2515 4885
rect 2535 4865 2550 4885
rect 2500 4835 2550 4865
rect 2500 4815 2515 4835
rect 2535 4815 2550 4835
rect 2500 4785 2550 4815
rect 2500 4765 2515 4785
rect 2535 4765 2550 4785
rect 2500 4735 2550 4765
rect 2500 4715 2515 4735
rect 2535 4715 2550 4735
rect 2500 4685 2550 4715
rect 2500 4665 2515 4685
rect 2535 4665 2550 4685
rect 2500 4635 2550 4665
rect 2500 4615 2515 4635
rect 2535 4615 2550 4635
rect 2500 4600 2550 4615
rect 2650 5085 2700 5100
rect 2650 5065 2665 5085
rect 2685 5065 2700 5085
rect 2650 5035 2700 5065
rect 2650 5015 2665 5035
rect 2685 5015 2700 5035
rect 2650 4985 2700 5015
rect 2650 4965 2665 4985
rect 2685 4965 2700 4985
rect 2650 4935 2700 4965
rect 2650 4915 2665 4935
rect 2685 4915 2700 4935
rect 2650 4885 2700 4915
rect 2650 4865 2665 4885
rect 2685 4865 2700 4885
rect 2650 4835 2700 4865
rect 2650 4815 2665 4835
rect 2685 4815 2700 4835
rect 2650 4785 2700 4815
rect 2650 4765 2665 4785
rect 2685 4765 2700 4785
rect 2650 4735 2700 4765
rect 2650 4715 2665 4735
rect 2685 4715 2700 4735
rect 2650 4685 2700 4715
rect 2650 4665 2665 4685
rect 2685 4665 2700 4685
rect 2650 4635 2700 4665
rect 2650 4615 2665 4635
rect 2685 4615 2700 4635
rect 2650 4600 2700 4615
rect 2800 5085 2850 5100
rect 2800 5065 2815 5085
rect 2835 5065 2850 5085
rect 2800 5035 2850 5065
rect 2800 5015 2815 5035
rect 2835 5015 2850 5035
rect 2800 4985 2850 5015
rect 2800 4965 2815 4985
rect 2835 4965 2850 4985
rect 2800 4935 2850 4965
rect 2800 4915 2815 4935
rect 2835 4915 2850 4935
rect 2800 4885 2850 4915
rect 2800 4865 2815 4885
rect 2835 4865 2850 4885
rect 2800 4835 2850 4865
rect 2800 4815 2815 4835
rect 2835 4815 2850 4835
rect 2800 4785 2850 4815
rect 2800 4765 2815 4785
rect 2835 4765 2850 4785
rect 2800 4735 2850 4765
rect 2800 4715 2815 4735
rect 2835 4715 2850 4735
rect 2800 4685 2850 4715
rect 2800 4665 2815 4685
rect 2835 4665 2850 4685
rect 2800 4635 2850 4665
rect 2800 4615 2815 4635
rect 2835 4615 2850 4635
rect 2800 4600 2850 4615
rect 2950 5085 3000 5100
rect 2950 5065 2965 5085
rect 2985 5065 3000 5085
rect 2950 5035 3000 5065
rect 2950 5015 2965 5035
rect 2985 5015 3000 5035
rect 2950 4985 3000 5015
rect 2950 4965 2965 4985
rect 2985 4965 3000 4985
rect 2950 4935 3000 4965
rect 2950 4915 2965 4935
rect 2985 4915 3000 4935
rect 2950 4885 3000 4915
rect 2950 4865 2965 4885
rect 2985 4865 3000 4885
rect 2950 4835 3000 4865
rect 2950 4815 2965 4835
rect 2985 4815 3000 4835
rect 2950 4785 3000 4815
rect 2950 4765 2965 4785
rect 2985 4765 3000 4785
rect 2950 4735 3000 4765
rect 2950 4715 2965 4735
rect 2985 4715 3000 4735
rect 2950 4685 3000 4715
rect 2950 4665 2965 4685
rect 2985 4665 3000 4685
rect 2950 4635 3000 4665
rect 2950 4615 2965 4635
rect 2985 4615 3000 4635
rect 2950 4600 3000 4615
rect 3100 5085 3150 5100
rect 3100 5065 3115 5085
rect 3135 5065 3150 5085
rect 3100 5035 3150 5065
rect 3100 5015 3115 5035
rect 3135 5015 3150 5035
rect 3100 4985 3150 5015
rect 3100 4965 3115 4985
rect 3135 4965 3150 4985
rect 3100 4935 3150 4965
rect 3100 4915 3115 4935
rect 3135 4915 3150 4935
rect 3100 4885 3150 4915
rect 3100 4865 3115 4885
rect 3135 4865 3150 4885
rect 3100 4835 3150 4865
rect 3100 4815 3115 4835
rect 3135 4815 3150 4835
rect 3100 4785 3150 4815
rect 3100 4765 3115 4785
rect 3135 4765 3150 4785
rect 3100 4735 3150 4765
rect 3100 4715 3115 4735
rect 3135 4715 3150 4735
rect 3100 4685 3150 4715
rect 3100 4665 3115 4685
rect 3135 4665 3150 4685
rect 3100 4635 3150 4665
rect 3100 4615 3115 4635
rect 3135 4615 3150 4635
rect 3100 4600 3150 4615
rect 3250 5085 3300 5100
rect 3250 5065 3265 5085
rect 3285 5065 3300 5085
rect 3250 5035 3300 5065
rect 3250 5015 3265 5035
rect 3285 5015 3300 5035
rect 3250 4985 3300 5015
rect 3250 4965 3265 4985
rect 3285 4965 3300 4985
rect 3250 4935 3300 4965
rect 3250 4915 3265 4935
rect 3285 4915 3300 4935
rect 3250 4885 3300 4915
rect 3250 4865 3265 4885
rect 3285 4865 3300 4885
rect 3250 4835 3300 4865
rect 3250 4815 3265 4835
rect 3285 4815 3300 4835
rect 3250 4785 3300 4815
rect 3250 4765 3265 4785
rect 3285 4765 3300 4785
rect 3250 4735 3300 4765
rect 3250 4715 3265 4735
rect 3285 4715 3300 4735
rect 3250 4685 3300 4715
rect 3250 4665 3265 4685
rect 3285 4665 3300 4685
rect 3250 4635 3300 4665
rect 3250 4615 3265 4635
rect 3285 4615 3300 4635
rect 3250 4600 3300 4615
rect 3400 5085 3450 5100
rect 3400 5065 3415 5085
rect 3435 5065 3450 5085
rect 3400 5035 3450 5065
rect 3400 5015 3415 5035
rect 3435 5015 3450 5035
rect 3400 4985 3450 5015
rect 3400 4965 3415 4985
rect 3435 4965 3450 4985
rect 3400 4935 3450 4965
rect 3400 4915 3415 4935
rect 3435 4915 3450 4935
rect 3400 4885 3450 4915
rect 3400 4865 3415 4885
rect 3435 4865 3450 4885
rect 3400 4835 3450 4865
rect 3400 4815 3415 4835
rect 3435 4815 3450 4835
rect 3400 4785 3450 4815
rect 3400 4765 3415 4785
rect 3435 4765 3450 4785
rect 3400 4735 3450 4765
rect 3400 4715 3415 4735
rect 3435 4715 3450 4735
rect 3400 4685 3450 4715
rect 3400 4665 3415 4685
rect 3435 4665 3450 4685
rect 3400 4635 3450 4665
rect 3400 4615 3415 4635
rect 3435 4615 3450 4635
rect 3400 4600 3450 4615
rect 3550 5085 3600 5100
rect 3550 5065 3565 5085
rect 3585 5065 3600 5085
rect 3550 5035 3600 5065
rect 3550 5015 3565 5035
rect 3585 5015 3600 5035
rect 3550 4985 3600 5015
rect 3550 4965 3565 4985
rect 3585 4965 3600 4985
rect 3550 4935 3600 4965
rect 3550 4915 3565 4935
rect 3585 4915 3600 4935
rect 3550 4885 3600 4915
rect 3550 4865 3565 4885
rect 3585 4865 3600 4885
rect 3550 4835 3600 4865
rect 3550 4815 3565 4835
rect 3585 4815 3600 4835
rect 3550 4785 3600 4815
rect 3550 4765 3565 4785
rect 3585 4765 3600 4785
rect 3550 4735 3600 4765
rect 3550 4715 3565 4735
rect 3585 4715 3600 4735
rect 3550 4685 3600 4715
rect 3550 4665 3565 4685
rect 3585 4665 3600 4685
rect 3550 4635 3600 4665
rect 3550 4615 3565 4635
rect 3585 4615 3600 4635
rect 3550 4600 3600 4615
rect 3700 4600 3750 5100
rect 3850 4600 3900 5100
rect 4000 4600 4050 5100
rect 4150 5085 4200 5100
rect 4150 5065 4165 5085
rect 4185 5065 4200 5085
rect 4150 5035 4200 5065
rect 4150 5015 4165 5035
rect 4185 5015 4200 5035
rect 4150 4985 4200 5015
rect 4150 4965 4165 4985
rect 4185 4965 4200 4985
rect 4150 4935 4200 4965
rect 4150 4915 4165 4935
rect 4185 4915 4200 4935
rect 4150 4885 4200 4915
rect 4150 4865 4165 4885
rect 4185 4865 4200 4885
rect 4150 4835 4200 4865
rect 4150 4815 4165 4835
rect 4185 4815 4200 4835
rect 4150 4785 4200 4815
rect 4150 4765 4165 4785
rect 4185 4765 4200 4785
rect 4150 4735 4200 4765
rect 4150 4715 4165 4735
rect 4185 4715 4200 4735
rect 4150 4685 4200 4715
rect 4150 4665 4165 4685
rect 4185 4665 4200 4685
rect 4150 4635 4200 4665
rect 4150 4615 4165 4635
rect 4185 4615 4200 4635
rect 4150 4600 4200 4615
rect 4300 4600 4350 5100
rect 4450 4600 4500 5100
rect 4600 4600 4650 5100
rect 4750 5085 4800 5100
rect 4750 5065 4765 5085
rect 4785 5065 4800 5085
rect 4750 5035 4800 5065
rect 4750 5015 4765 5035
rect 4785 5015 4800 5035
rect 4750 4985 4800 5015
rect 4750 4965 4765 4985
rect 4785 4965 4800 4985
rect 4750 4935 4800 4965
rect 4750 4915 4765 4935
rect 4785 4915 4800 4935
rect 4750 4885 4800 4915
rect 4750 4865 4765 4885
rect 4785 4865 4800 4885
rect 4750 4835 4800 4865
rect 4750 4815 4765 4835
rect 4785 4815 4800 4835
rect 4750 4785 4800 4815
rect 4750 4765 4765 4785
rect 4785 4765 4800 4785
rect 4750 4735 4800 4765
rect 4750 4715 4765 4735
rect 4785 4715 4800 4735
rect 4750 4685 4800 4715
rect 4750 4665 4765 4685
rect 4785 4665 4800 4685
rect 4750 4635 4800 4665
rect 4750 4615 4765 4635
rect 4785 4615 4800 4635
rect 4750 4600 4800 4615
rect 4900 5085 4950 5100
rect 4900 5065 4915 5085
rect 4935 5065 4950 5085
rect 4900 5035 4950 5065
rect 4900 5015 4915 5035
rect 4935 5015 4950 5035
rect 4900 4985 4950 5015
rect 4900 4965 4915 4985
rect 4935 4965 4950 4985
rect 4900 4935 4950 4965
rect 4900 4915 4915 4935
rect 4935 4915 4950 4935
rect 4900 4885 4950 4915
rect 4900 4865 4915 4885
rect 4935 4865 4950 4885
rect 4900 4835 4950 4865
rect 4900 4815 4915 4835
rect 4935 4815 4950 4835
rect 4900 4785 4950 4815
rect 4900 4765 4915 4785
rect 4935 4765 4950 4785
rect 4900 4735 4950 4765
rect 4900 4715 4915 4735
rect 4935 4715 4950 4735
rect 4900 4685 4950 4715
rect 4900 4665 4915 4685
rect 4935 4665 4950 4685
rect 4900 4635 4950 4665
rect 4900 4615 4915 4635
rect 4935 4615 4950 4635
rect 4900 4600 4950 4615
rect 5050 5085 5100 5100
rect 5050 5065 5065 5085
rect 5085 5065 5100 5085
rect 5050 5035 5100 5065
rect 5050 5015 5065 5035
rect 5085 5015 5100 5035
rect 5050 4985 5100 5015
rect 5050 4965 5065 4985
rect 5085 4965 5100 4985
rect 5050 4935 5100 4965
rect 5050 4915 5065 4935
rect 5085 4915 5100 4935
rect 5050 4885 5100 4915
rect 5050 4865 5065 4885
rect 5085 4865 5100 4885
rect 5050 4835 5100 4865
rect 5050 4815 5065 4835
rect 5085 4815 5100 4835
rect 5050 4785 5100 4815
rect 5050 4765 5065 4785
rect 5085 4765 5100 4785
rect 5050 4735 5100 4765
rect 5050 4715 5065 4735
rect 5085 4715 5100 4735
rect 5050 4685 5100 4715
rect 5050 4665 5065 4685
rect 5085 4665 5100 4685
rect 5050 4635 5100 4665
rect 5050 4615 5065 4635
rect 5085 4615 5100 4635
rect 5050 4600 5100 4615
rect 5200 5085 5250 5100
rect 5200 5065 5215 5085
rect 5235 5065 5250 5085
rect 5200 5035 5250 5065
rect 5200 5015 5215 5035
rect 5235 5015 5250 5035
rect 5200 4985 5250 5015
rect 5200 4965 5215 4985
rect 5235 4965 5250 4985
rect 5200 4935 5250 4965
rect 5200 4915 5215 4935
rect 5235 4915 5250 4935
rect 5200 4885 5250 4915
rect 5200 4865 5215 4885
rect 5235 4865 5250 4885
rect 5200 4835 5250 4865
rect 5200 4815 5215 4835
rect 5235 4815 5250 4835
rect 5200 4785 5250 4815
rect 5200 4765 5215 4785
rect 5235 4765 5250 4785
rect 5200 4735 5250 4765
rect 5200 4715 5215 4735
rect 5235 4715 5250 4735
rect 5200 4685 5250 4715
rect 5200 4665 5215 4685
rect 5235 4665 5250 4685
rect 5200 4635 5250 4665
rect 5200 4615 5215 4635
rect 5235 4615 5250 4635
rect 5200 4600 5250 4615
rect 5350 5085 5400 5100
rect 5350 5065 5365 5085
rect 5385 5065 5400 5085
rect 5350 5035 5400 5065
rect 5350 5015 5365 5035
rect 5385 5015 5400 5035
rect 5350 4985 5400 5015
rect 5350 4965 5365 4985
rect 5385 4965 5400 4985
rect 5350 4935 5400 4965
rect 5350 4915 5365 4935
rect 5385 4915 5400 4935
rect 5350 4885 5400 4915
rect 5350 4865 5365 4885
rect 5385 4865 5400 4885
rect 5350 4835 5400 4865
rect 5350 4815 5365 4835
rect 5385 4815 5400 4835
rect 5350 4785 5400 4815
rect 5350 4765 5365 4785
rect 5385 4765 5400 4785
rect 5350 4735 5400 4765
rect 5350 4715 5365 4735
rect 5385 4715 5400 4735
rect 5350 4685 5400 4715
rect 5350 4665 5365 4685
rect 5385 4665 5400 4685
rect 5350 4635 5400 4665
rect 5350 4615 5365 4635
rect 5385 4615 5400 4635
rect 5350 4600 5400 4615
rect 5500 5085 5550 5100
rect 5500 5065 5515 5085
rect 5535 5065 5550 5085
rect 5500 5035 5550 5065
rect 5500 5015 5515 5035
rect 5535 5015 5550 5035
rect 5500 4985 5550 5015
rect 5500 4965 5515 4985
rect 5535 4965 5550 4985
rect 5500 4935 5550 4965
rect 5500 4915 5515 4935
rect 5535 4915 5550 4935
rect 5500 4885 5550 4915
rect 5500 4865 5515 4885
rect 5535 4865 5550 4885
rect 5500 4835 5550 4865
rect 5500 4815 5515 4835
rect 5535 4815 5550 4835
rect 5500 4785 5550 4815
rect 5500 4765 5515 4785
rect 5535 4765 5550 4785
rect 5500 4735 5550 4765
rect 5500 4715 5515 4735
rect 5535 4715 5550 4735
rect 5500 4685 5550 4715
rect 5500 4665 5515 4685
rect 5535 4665 5550 4685
rect 5500 4635 5550 4665
rect 5500 4615 5515 4635
rect 5535 4615 5550 4635
rect 5500 4600 5550 4615
rect 5650 5085 5700 5100
rect 5650 5065 5665 5085
rect 5685 5065 5700 5085
rect 5650 5035 5700 5065
rect 5650 5015 5665 5035
rect 5685 5015 5700 5035
rect 5650 4985 5700 5015
rect 5650 4965 5665 4985
rect 5685 4965 5700 4985
rect 5650 4935 5700 4965
rect 5650 4915 5665 4935
rect 5685 4915 5700 4935
rect 5650 4885 5700 4915
rect 5650 4865 5665 4885
rect 5685 4865 5700 4885
rect 5650 4835 5700 4865
rect 5650 4815 5665 4835
rect 5685 4815 5700 4835
rect 5650 4785 5700 4815
rect 5650 4765 5665 4785
rect 5685 4765 5700 4785
rect 5650 4735 5700 4765
rect 5650 4715 5665 4735
rect 5685 4715 5700 4735
rect 5650 4685 5700 4715
rect 5650 4665 5665 4685
rect 5685 4665 5700 4685
rect 5650 4635 5700 4665
rect 5650 4615 5665 4635
rect 5685 4615 5700 4635
rect 5650 4600 5700 4615
rect 5800 5085 5850 5100
rect 5800 5065 5815 5085
rect 5835 5065 5850 5085
rect 5800 5035 5850 5065
rect 5800 5015 5815 5035
rect 5835 5015 5850 5035
rect 5800 4985 5850 5015
rect 5800 4965 5815 4985
rect 5835 4965 5850 4985
rect 5800 4935 5850 4965
rect 5800 4915 5815 4935
rect 5835 4915 5850 4935
rect 5800 4885 5850 4915
rect 5800 4865 5815 4885
rect 5835 4865 5850 4885
rect 5800 4835 5850 4865
rect 5800 4815 5815 4835
rect 5835 4815 5850 4835
rect 5800 4785 5850 4815
rect 5800 4765 5815 4785
rect 5835 4765 5850 4785
rect 5800 4735 5850 4765
rect 5800 4715 5815 4735
rect 5835 4715 5850 4735
rect 5800 4685 5850 4715
rect 5800 4665 5815 4685
rect 5835 4665 5850 4685
rect 5800 4635 5850 4665
rect 5800 4615 5815 4635
rect 5835 4615 5850 4635
rect 5800 4600 5850 4615
rect 5950 5085 6000 5100
rect 5950 5065 5965 5085
rect 5985 5065 6000 5085
rect 5950 5035 6000 5065
rect 5950 5015 5965 5035
rect 5985 5015 6000 5035
rect 5950 4985 6000 5015
rect 5950 4965 5965 4985
rect 5985 4965 6000 4985
rect 5950 4935 6000 4965
rect 5950 4915 5965 4935
rect 5985 4915 6000 4935
rect 5950 4885 6000 4915
rect 5950 4865 5965 4885
rect 5985 4865 6000 4885
rect 5950 4835 6000 4865
rect 5950 4815 5965 4835
rect 5985 4815 6000 4835
rect 5950 4785 6000 4815
rect 5950 4765 5965 4785
rect 5985 4765 6000 4785
rect 5950 4735 6000 4765
rect 5950 4715 5965 4735
rect 5985 4715 6000 4735
rect 5950 4685 6000 4715
rect 5950 4665 5965 4685
rect 5985 4665 6000 4685
rect 5950 4635 6000 4665
rect 5950 4615 5965 4635
rect 5985 4615 6000 4635
rect 5950 4600 6000 4615
rect 6100 5085 6150 5100
rect 6100 5065 6115 5085
rect 6135 5065 6150 5085
rect 6100 5035 6150 5065
rect 6100 5015 6115 5035
rect 6135 5015 6150 5035
rect 6100 4985 6150 5015
rect 6100 4965 6115 4985
rect 6135 4965 6150 4985
rect 6100 4935 6150 4965
rect 6100 4915 6115 4935
rect 6135 4915 6150 4935
rect 6100 4885 6150 4915
rect 6100 4865 6115 4885
rect 6135 4865 6150 4885
rect 6100 4835 6150 4865
rect 6100 4815 6115 4835
rect 6135 4815 6150 4835
rect 6100 4785 6150 4815
rect 6100 4765 6115 4785
rect 6135 4765 6150 4785
rect 6100 4735 6150 4765
rect 6100 4715 6115 4735
rect 6135 4715 6150 4735
rect 6100 4685 6150 4715
rect 6100 4665 6115 4685
rect 6135 4665 6150 4685
rect 6100 4635 6150 4665
rect 6100 4615 6115 4635
rect 6135 4615 6150 4635
rect 6100 4600 6150 4615
rect 6250 5085 6300 5100
rect 6250 5065 6265 5085
rect 6285 5065 6300 5085
rect 6250 5035 6300 5065
rect 6250 5015 6265 5035
rect 6285 5015 6300 5035
rect 6250 4985 6300 5015
rect 6250 4965 6265 4985
rect 6285 4965 6300 4985
rect 6250 4935 6300 4965
rect 6250 4915 6265 4935
rect 6285 4915 6300 4935
rect 6250 4885 6300 4915
rect 6250 4865 6265 4885
rect 6285 4865 6300 4885
rect 6250 4835 6300 4865
rect 6250 4815 6265 4835
rect 6285 4815 6300 4835
rect 6250 4785 6300 4815
rect 6250 4765 6265 4785
rect 6285 4765 6300 4785
rect 6250 4735 6300 4765
rect 6250 4715 6265 4735
rect 6285 4715 6300 4735
rect 6250 4685 6300 4715
rect 6250 4665 6265 4685
rect 6285 4665 6300 4685
rect 6250 4635 6300 4665
rect 6250 4615 6265 4635
rect 6285 4615 6300 4635
rect 6250 4600 6300 4615
rect 6400 5085 6450 5100
rect 6400 5065 6415 5085
rect 6435 5065 6450 5085
rect 6400 5035 6450 5065
rect 6400 5015 6415 5035
rect 6435 5015 6450 5035
rect 6400 4985 6450 5015
rect 6400 4965 6415 4985
rect 6435 4965 6450 4985
rect 6400 4935 6450 4965
rect 6400 4915 6415 4935
rect 6435 4915 6450 4935
rect 6400 4885 6450 4915
rect 6400 4865 6415 4885
rect 6435 4865 6450 4885
rect 6400 4835 6450 4865
rect 6400 4815 6415 4835
rect 6435 4815 6450 4835
rect 6400 4785 6450 4815
rect 6400 4765 6415 4785
rect 6435 4765 6450 4785
rect 6400 4735 6450 4765
rect 6400 4715 6415 4735
rect 6435 4715 6450 4735
rect 6400 4685 6450 4715
rect 6400 4665 6415 4685
rect 6435 4665 6450 4685
rect 6400 4635 6450 4665
rect 6400 4615 6415 4635
rect 6435 4615 6450 4635
rect 6400 4600 6450 4615
rect 6550 5085 6600 5100
rect 6550 5065 6565 5085
rect 6585 5065 6600 5085
rect 6550 5035 6600 5065
rect 6550 5015 6565 5035
rect 6585 5015 6600 5035
rect 6550 4985 6600 5015
rect 6550 4965 6565 4985
rect 6585 4965 6600 4985
rect 6550 4935 6600 4965
rect 6550 4915 6565 4935
rect 6585 4915 6600 4935
rect 6550 4885 6600 4915
rect 6550 4865 6565 4885
rect 6585 4865 6600 4885
rect 6550 4835 6600 4865
rect 6550 4815 6565 4835
rect 6585 4815 6600 4835
rect 6550 4785 6600 4815
rect 6550 4765 6565 4785
rect 6585 4765 6600 4785
rect 6550 4735 6600 4765
rect 6550 4715 6565 4735
rect 6585 4715 6600 4735
rect 6550 4685 6600 4715
rect 6550 4665 6565 4685
rect 6585 4665 6600 4685
rect 6550 4635 6600 4665
rect 6550 4615 6565 4635
rect 6585 4615 6600 4635
rect 6550 4600 6600 4615
rect 6700 5085 6750 5100
rect 6700 5065 6715 5085
rect 6735 5065 6750 5085
rect 6700 5035 6750 5065
rect 6700 5015 6715 5035
rect 6735 5015 6750 5035
rect 6700 4985 6750 5015
rect 6700 4965 6715 4985
rect 6735 4965 6750 4985
rect 6700 4935 6750 4965
rect 6700 4915 6715 4935
rect 6735 4915 6750 4935
rect 6700 4885 6750 4915
rect 6700 4865 6715 4885
rect 6735 4865 6750 4885
rect 6700 4835 6750 4865
rect 6700 4815 6715 4835
rect 6735 4815 6750 4835
rect 6700 4785 6750 4815
rect 6700 4765 6715 4785
rect 6735 4765 6750 4785
rect 6700 4735 6750 4765
rect 6700 4715 6715 4735
rect 6735 4715 6750 4735
rect 6700 4685 6750 4715
rect 6700 4665 6715 4685
rect 6735 4665 6750 4685
rect 6700 4635 6750 4665
rect 6700 4615 6715 4635
rect 6735 4615 6750 4635
rect 6700 4600 6750 4615
rect 6850 5085 6900 5100
rect 6850 5065 6865 5085
rect 6885 5065 6900 5085
rect 6850 5035 6900 5065
rect 6850 5015 6865 5035
rect 6885 5015 6900 5035
rect 6850 4985 6900 5015
rect 6850 4965 6865 4985
rect 6885 4965 6900 4985
rect 6850 4935 6900 4965
rect 6850 4915 6865 4935
rect 6885 4915 6900 4935
rect 6850 4885 6900 4915
rect 6850 4865 6865 4885
rect 6885 4865 6900 4885
rect 6850 4835 6900 4865
rect 6850 4815 6865 4835
rect 6885 4815 6900 4835
rect 6850 4785 6900 4815
rect 6850 4765 6865 4785
rect 6885 4765 6900 4785
rect 6850 4735 6900 4765
rect 6850 4715 6865 4735
rect 6885 4715 6900 4735
rect 6850 4685 6900 4715
rect 6850 4665 6865 4685
rect 6885 4665 6900 4685
rect 6850 4635 6900 4665
rect 6850 4615 6865 4635
rect 6885 4615 6900 4635
rect 6850 4600 6900 4615
rect 7000 5085 7050 5100
rect 7000 5065 7015 5085
rect 7035 5065 7050 5085
rect 7000 5035 7050 5065
rect 7000 5015 7015 5035
rect 7035 5015 7050 5035
rect 7000 4985 7050 5015
rect 7000 4965 7015 4985
rect 7035 4965 7050 4985
rect 7000 4935 7050 4965
rect 7000 4915 7015 4935
rect 7035 4915 7050 4935
rect 7000 4885 7050 4915
rect 7000 4865 7015 4885
rect 7035 4865 7050 4885
rect 7000 4835 7050 4865
rect 7000 4815 7015 4835
rect 7035 4815 7050 4835
rect 7000 4785 7050 4815
rect 7000 4765 7015 4785
rect 7035 4765 7050 4785
rect 7000 4735 7050 4765
rect 7000 4715 7015 4735
rect 7035 4715 7050 4735
rect 7000 4685 7050 4715
rect 7000 4665 7015 4685
rect 7035 4665 7050 4685
rect 7000 4635 7050 4665
rect 7000 4615 7015 4635
rect 7035 4615 7050 4635
rect 7000 4600 7050 4615
rect 7150 5085 7200 5100
rect 7150 5065 7165 5085
rect 7185 5065 7200 5085
rect 7150 5035 7200 5065
rect 7150 5015 7165 5035
rect 7185 5015 7200 5035
rect 7150 4985 7200 5015
rect 7150 4965 7165 4985
rect 7185 4965 7200 4985
rect 7150 4935 7200 4965
rect 7150 4915 7165 4935
rect 7185 4915 7200 4935
rect 7150 4885 7200 4915
rect 7150 4865 7165 4885
rect 7185 4865 7200 4885
rect 7150 4835 7200 4865
rect 7150 4815 7165 4835
rect 7185 4815 7200 4835
rect 7150 4785 7200 4815
rect 7150 4765 7165 4785
rect 7185 4765 7200 4785
rect 7150 4735 7200 4765
rect 7150 4715 7165 4735
rect 7185 4715 7200 4735
rect 7150 4685 7200 4715
rect 7150 4665 7165 4685
rect 7185 4665 7200 4685
rect 7150 4635 7200 4665
rect 7150 4615 7165 4635
rect 7185 4615 7200 4635
rect 7150 4600 7200 4615
rect 7300 5085 7350 5100
rect 7300 5065 7315 5085
rect 7335 5065 7350 5085
rect 7300 5035 7350 5065
rect 7300 5015 7315 5035
rect 7335 5015 7350 5035
rect 7300 4985 7350 5015
rect 7300 4965 7315 4985
rect 7335 4965 7350 4985
rect 7300 4935 7350 4965
rect 7300 4915 7315 4935
rect 7335 4915 7350 4935
rect 7300 4885 7350 4915
rect 7300 4865 7315 4885
rect 7335 4865 7350 4885
rect 7300 4835 7350 4865
rect 7300 4815 7315 4835
rect 7335 4815 7350 4835
rect 7300 4785 7350 4815
rect 7300 4765 7315 4785
rect 7335 4765 7350 4785
rect 7300 4735 7350 4765
rect 7300 4715 7315 4735
rect 7335 4715 7350 4735
rect 7300 4685 7350 4715
rect 7300 4665 7315 4685
rect 7335 4665 7350 4685
rect 7300 4635 7350 4665
rect 7300 4615 7315 4635
rect 7335 4615 7350 4635
rect 7300 4600 7350 4615
rect 7450 5085 7500 5100
rect 7450 5065 7465 5085
rect 7485 5065 7500 5085
rect 7450 5035 7500 5065
rect 7450 5015 7465 5035
rect 7485 5015 7500 5035
rect 7450 4985 7500 5015
rect 7450 4965 7465 4985
rect 7485 4965 7500 4985
rect 7450 4935 7500 4965
rect 7450 4915 7465 4935
rect 7485 4915 7500 4935
rect 7450 4885 7500 4915
rect 7450 4865 7465 4885
rect 7485 4865 7500 4885
rect 7450 4835 7500 4865
rect 7450 4815 7465 4835
rect 7485 4815 7500 4835
rect 7450 4785 7500 4815
rect 7450 4765 7465 4785
rect 7485 4765 7500 4785
rect 7450 4735 7500 4765
rect 7450 4715 7465 4735
rect 7485 4715 7500 4735
rect 7450 4685 7500 4715
rect 7450 4665 7465 4685
rect 7485 4665 7500 4685
rect 7450 4635 7500 4665
rect 7450 4615 7465 4635
rect 7485 4615 7500 4635
rect 7450 4600 7500 4615
rect 7600 5085 7650 5100
rect 7600 5065 7615 5085
rect 7635 5065 7650 5085
rect 7600 5035 7650 5065
rect 7600 5015 7615 5035
rect 7635 5015 7650 5035
rect 7600 4985 7650 5015
rect 7600 4965 7615 4985
rect 7635 4965 7650 4985
rect 7600 4935 7650 4965
rect 7600 4915 7615 4935
rect 7635 4915 7650 4935
rect 7600 4885 7650 4915
rect 7600 4865 7615 4885
rect 7635 4865 7650 4885
rect 7600 4835 7650 4865
rect 7600 4815 7615 4835
rect 7635 4815 7650 4835
rect 7600 4785 7650 4815
rect 7600 4765 7615 4785
rect 7635 4765 7650 4785
rect 7600 4735 7650 4765
rect 7600 4715 7615 4735
rect 7635 4715 7650 4735
rect 7600 4685 7650 4715
rect 7600 4665 7615 4685
rect 7635 4665 7650 4685
rect 7600 4635 7650 4665
rect 7600 4615 7615 4635
rect 7635 4615 7650 4635
rect 7600 4600 7650 4615
rect 7750 5085 7800 5100
rect 7750 5065 7765 5085
rect 7785 5065 7800 5085
rect 7750 5035 7800 5065
rect 7750 5015 7765 5035
rect 7785 5015 7800 5035
rect 7750 4985 7800 5015
rect 7750 4965 7765 4985
rect 7785 4965 7800 4985
rect 7750 4935 7800 4965
rect 7750 4915 7765 4935
rect 7785 4915 7800 4935
rect 7750 4885 7800 4915
rect 7750 4865 7765 4885
rect 7785 4865 7800 4885
rect 7750 4835 7800 4865
rect 7750 4815 7765 4835
rect 7785 4815 7800 4835
rect 7750 4785 7800 4815
rect 7750 4765 7765 4785
rect 7785 4765 7800 4785
rect 7750 4735 7800 4765
rect 7750 4715 7765 4735
rect 7785 4715 7800 4735
rect 7750 4685 7800 4715
rect 7750 4665 7765 4685
rect 7785 4665 7800 4685
rect 7750 4635 7800 4665
rect 7750 4615 7765 4635
rect 7785 4615 7800 4635
rect 7750 4600 7800 4615
rect 7900 4600 7950 5100
rect 8050 4600 8100 5100
rect 8200 4600 8250 5100
rect 8350 5085 8400 5100
rect 8350 5065 8365 5085
rect 8385 5065 8400 5085
rect 8350 5035 8400 5065
rect 8350 5015 8365 5035
rect 8385 5015 8400 5035
rect 8350 4985 8400 5015
rect 8350 4965 8365 4985
rect 8385 4965 8400 4985
rect 8350 4935 8400 4965
rect 8350 4915 8365 4935
rect 8385 4915 8400 4935
rect 8350 4885 8400 4915
rect 8350 4865 8365 4885
rect 8385 4865 8400 4885
rect 8350 4835 8400 4865
rect 8350 4815 8365 4835
rect 8385 4815 8400 4835
rect 8350 4785 8400 4815
rect 8350 4765 8365 4785
rect 8385 4765 8400 4785
rect 8350 4735 8400 4765
rect 8350 4715 8365 4735
rect 8385 4715 8400 4735
rect 8350 4685 8400 4715
rect 8350 4665 8365 4685
rect 8385 4665 8400 4685
rect 8350 4635 8400 4665
rect 8350 4615 8365 4635
rect 8385 4615 8400 4635
rect 8350 4600 8400 4615
rect 8500 5085 8550 5100
rect 8500 5065 8515 5085
rect 8535 5065 8550 5085
rect 8500 5035 8550 5065
rect 8500 5015 8515 5035
rect 8535 5015 8550 5035
rect 8500 4985 8550 5015
rect 8500 4965 8515 4985
rect 8535 4965 8550 4985
rect 8500 4935 8550 4965
rect 8500 4915 8515 4935
rect 8535 4915 8550 4935
rect 8500 4885 8550 4915
rect 8500 4865 8515 4885
rect 8535 4865 8550 4885
rect 8500 4835 8550 4865
rect 8500 4815 8515 4835
rect 8535 4815 8550 4835
rect 8500 4785 8550 4815
rect 8500 4765 8515 4785
rect 8535 4765 8550 4785
rect 8500 4735 8550 4765
rect 8500 4715 8515 4735
rect 8535 4715 8550 4735
rect 8500 4685 8550 4715
rect 8500 4665 8515 4685
rect 8535 4665 8550 4685
rect 8500 4635 8550 4665
rect 8500 4615 8515 4635
rect 8535 4615 8550 4635
rect 8500 4600 8550 4615
rect 8650 5085 8700 5100
rect 8650 5065 8665 5085
rect 8685 5065 8700 5085
rect 8650 5035 8700 5065
rect 8650 5015 8665 5035
rect 8685 5015 8700 5035
rect 8650 4985 8700 5015
rect 8650 4965 8665 4985
rect 8685 4965 8700 4985
rect 8650 4935 8700 4965
rect 8650 4915 8665 4935
rect 8685 4915 8700 4935
rect 8650 4885 8700 4915
rect 8650 4865 8665 4885
rect 8685 4865 8700 4885
rect 8650 4835 8700 4865
rect 8650 4815 8665 4835
rect 8685 4815 8700 4835
rect 8650 4785 8700 4815
rect 8650 4765 8665 4785
rect 8685 4765 8700 4785
rect 8650 4735 8700 4765
rect 8650 4715 8665 4735
rect 8685 4715 8700 4735
rect 8650 4685 8700 4715
rect 8650 4665 8665 4685
rect 8685 4665 8700 4685
rect 8650 4635 8700 4665
rect 8650 4615 8665 4635
rect 8685 4615 8700 4635
rect 8650 4600 8700 4615
rect 8800 5085 8850 5100
rect 8800 5065 8815 5085
rect 8835 5065 8850 5085
rect 8800 5035 8850 5065
rect 8800 5015 8815 5035
rect 8835 5015 8850 5035
rect 8800 4985 8850 5015
rect 8800 4965 8815 4985
rect 8835 4965 8850 4985
rect 8800 4935 8850 4965
rect 8800 4915 8815 4935
rect 8835 4915 8850 4935
rect 8800 4885 8850 4915
rect 8800 4865 8815 4885
rect 8835 4865 8850 4885
rect 8800 4835 8850 4865
rect 8800 4815 8815 4835
rect 8835 4815 8850 4835
rect 8800 4785 8850 4815
rect 8800 4765 8815 4785
rect 8835 4765 8850 4785
rect 8800 4735 8850 4765
rect 8800 4715 8815 4735
rect 8835 4715 8850 4735
rect 8800 4685 8850 4715
rect 8800 4665 8815 4685
rect 8835 4665 8850 4685
rect 8800 4635 8850 4665
rect 8800 4615 8815 4635
rect 8835 4615 8850 4635
rect 8800 4600 8850 4615
rect 8950 5085 9000 5100
rect 8950 5065 8965 5085
rect 8985 5065 9000 5085
rect 8950 5035 9000 5065
rect 8950 5015 8965 5035
rect 8985 5015 9000 5035
rect 8950 4985 9000 5015
rect 8950 4965 8965 4985
rect 8985 4965 9000 4985
rect 8950 4935 9000 4965
rect 8950 4915 8965 4935
rect 8985 4915 9000 4935
rect 8950 4885 9000 4915
rect 8950 4865 8965 4885
rect 8985 4865 9000 4885
rect 8950 4835 9000 4865
rect 8950 4815 8965 4835
rect 8985 4815 9000 4835
rect 8950 4785 9000 4815
rect 8950 4765 8965 4785
rect 8985 4765 9000 4785
rect 8950 4735 9000 4765
rect 8950 4715 8965 4735
rect 8985 4715 9000 4735
rect 8950 4685 9000 4715
rect 8950 4665 8965 4685
rect 8985 4665 9000 4685
rect 8950 4635 9000 4665
rect 8950 4615 8965 4635
rect 8985 4615 9000 4635
rect 8950 4600 9000 4615
rect 9100 5085 9150 5100
rect 9100 5065 9115 5085
rect 9135 5065 9150 5085
rect 9100 5035 9150 5065
rect 9100 5015 9115 5035
rect 9135 5015 9150 5035
rect 9100 4985 9150 5015
rect 9100 4965 9115 4985
rect 9135 4965 9150 4985
rect 9100 4935 9150 4965
rect 9100 4915 9115 4935
rect 9135 4915 9150 4935
rect 9100 4885 9150 4915
rect 9100 4865 9115 4885
rect 9135 4865 9150 4885
rect 9100 4835 9150 4865
rect 9100 4815 9115 4835
rect 9135 4815 9150 4835
rect 9100 4785 9150 4815
rect 9100 4765 9115 4785
rect 9135 4765 9150 4785
rect 9100 4735 9150 4765
rect 9100 4715 9115 4735
rect 9135 4715 9150 4735
rect 9100 4685 9150 4715
rect 9100 4665 9115 4685
rect 9135 4665 9150 4685
rect 9100 4635 9150 4665
rect 9100 4615 9115 4635
rect 9135 4615 9150 4635
rect 9100 4600 9150 4615
rect 9250 5085 9300 5100
rect 9250 5065 9265 5085
rect 9285 5065 9300 5085
rect 9250 5035 9300 5065
rect 9250 5015 9265 5035
rect 9285 5015 9300 5035
rect 9250 4985 9300 5015
rect 9250 4965 9265 4985
rect 9285 4965 9300 4985
rect 9250 4935 9300 4965
rect 9250 4915 9265 4935
rect 9285 4915 9300 4935
rect 9250 4885 9300 4915
rect 9250 4865 9265 4885
rect 9285 4865 9300 4885
rect 9250 4835 9300 4865
rect 9250 4815 9265 4835
rect 9285 4815 9300 4835
rect 9250 4785 9300 4815
rect 9250 4765 9265 4785
rect 9285 4765 9300 4785
rect 9250 4735 9300 4765
rect 9250 4715 9265 4735
rect 9285 4715 9300 4735
rect 9250 4685 9300 4715
rect 9250 4665 9265 4685
rect 9285 4665 9300 4685
rect 9250 4635 9300 4665
rect 9250 4615 9265 4635
rect 9285 4615 9300 4635
rect 9250 4600 9300 4615
rect 9400 5085 9450 5100
rect 9400 5065 9415 5085
rect 9435 5065 9450 5085
rect 9400 5035 9450 5065
rect 9400 5015 9415 5035
rect 9435 5015 9450 5035
rect 9400 4985 9450 5015
rect 9400 4965 9415 4985
rect 9435 4965 9450 4985
rect 9400 4935 9450 4965
rect 9400 4915 9415 4935
rect 9435 4915 9450 4935
rect 9400 4885 9450 4915
rect 9400 4865 9415 4885
rect 9435 4865 9450 4885
rect 9400 4835 9450 4865
rect 9400 4815 9415 4835
rect 9435 4815 9450 4835
rect 9400 4785 9450 4815
rect 9400 4765 9415 4785
rect 9435 4765 9450 4785
rect 9400 4735 9450 4765
rect 9400 4715 9415 4735
rect 9435 4715 9450 4735
rect 9400 4685 9450 4715
rect 9400 4665 9415 4685
rect 9435 4665 9450 4685
rect 9400 4635 9450 4665
rect 9400 4615 9415 4635
rect 9435 4615 9450 4635
rect 9400 4600 9450 4615
rect 9550 5085 9600 5100
rect 9550 5065 9565 5085
rect 9585 5065 9600 5085
rect 9550 5035 9600 5065
rect 9550 5015 9565 5035
rect 9585 5015 9600 5035
rect 9550 4985 9600 5015
rect 9550 4965 9565 4985
rect 9585 4965 9600 4985
rect 9550 4935 9600 4965
rect 9550 4915 9565 4935
rect 9585 4915 9600 4935
rect 9550 4885 9600 4915
rect 9550 4865 9565 4885
rect 9585 4865 9600 4885
rect 9550 4835 9600 4865
rect 9550 4815 9565 4835
rect 9585 4815 9600 4835
rect 9550 4785 9600 4815
rect 9550 4765 9565 4785
rect 9585 4765 9600 4785
rect 9550 4735 9600 4765
rect 9550 4715 9565 4735
rect 9585 4715 9600 4735
rect 9550 4685 9600 4715
rect 9550 4665 9565 4685
rect 9585 4665 9600 4685
rect 9550 4635 9600 4665
rect 9550 4615 9565 4635
rect 9585 4615 9600 4635
rect 9550 4600 9600 4615
rect 9700 5085 9750 5100
rect 9700 5065 9715 5085
rect 9735 5065 9750 5085
rect 9700 5035 9750 5065
rect 9700 5015 9715 5035
rect 9735 5015 9750 5035
rect 9700 4985 9750 5015
rect 9700 4965 9715 4985
rect 9735 4965 9750 4985
rect 9700 4935 9750 4965
rect 9700 4915 9715 4935
rect 9735 4915 9750 4935
rect 9700 4885 9750 4915
rect 9700 4865 9715 4885
rect 9735 4865 9750 4885
rect 9700 4835 9750 4865
rect 9700 4815 9715 4835
rect 9735 4815 9750 4835
rect 9700 4785 9750 4815
rect 9700 4765 9715 4785
rect 9735 4765 9750 4785
rect 9700 4735 9750 4765
rect 9700 4715 9715 4735
rect 9735 4715 9750 4735
rect 9700 4685 9750 4715
rect 9700 4665 9715 4685
rect 9735 4665 9750 4685
rect 9700 4635 9750 4665
rect 9700 4615 9715 4635
rect 9735 4615 9750 4635
rect 9700 4600 9750 4615
rect 9850 5085 9900 5100
rect 9850 5065 9865 5085
rect 9885 5065 9900 5085
rect 9850 5035 9900 5065
rect 9850 5015 9865 5035
rect 9885 5015 9900 5035
rect 9850 4985 9900 5015
rect 9850 4965 9865 4985
rect 9885 4965 9900 4985
rect 9850 4935 9900 4965
rect 9850 4915 9865 4935
rect 9885 4915 9900 4935
rect 9850 4885 9900 4915
rect 9850 4865 9865 4885
rect 9885 4865 9900 4885
rect 9850 4835 9900 4865
rect 9850 4815 9865 4835
rect 9885 4815 9900 4835
rect 9850 4785 9900 4815
rect 9850 4765 9865 4785
rect 9885 4765 9900 4785
rect 9850 4735 9900 4765
rect 9850 4715 9865 4735
rect 9885 4715 9900 4735
rect 9850 4685 9900 4715
rect 9850 4665 9865 4685
rect 9885 4665 9900 4685
rect 9850 4635 9900 4665
rect 9850 4615 9865 4635
rect 9885 4615 9900 4635
rect 9850 4600 9900 4615
rect 10000 5085 10050 5100
rect 10000 5065 10015 5085
rect 10035 5065 10050 5085
rect 10000 5035 10050 5065
rect 10000 5015 10015 5035
rect 10035 5015 10050 5035
rect 10000 4985 10050 5015
rect 10000 4965 10015 4985
rect 10035 4965 10050 4985
rect 10000 4935 10050 4965
rect 10000 4915 10015 4935
rect 10035 4915 10050 4935
rect 10000 4885 10050 4915
rect 10000 4865 10015 4885
rect 10035 4865 10050 4885
rect 10000 4835 10050 4865
rect 10000 4815 10015 4835
rect 10035 4815 10050 4835
rect 10000 4785 10050 4815
rect 10000 4765 10015 4785
rect 10035 4765 10050 4785
rect 10000 4735 10050 4765
rect 10000 4715 10015 4735
rect 10035 4715 10050 4735
rect 10000 4685 10050 4715
rect 10000 4665 10015 4685
rect 10035 4665 10050 4685
rect 10000 4635 10050 4665
rect 10000 4615 10015 4635
rect 10035 4615 10050 4635
rect 10000 4600 10050 4615
rect 10150 5085 10200 5100
rect 10150 5065 10165 5085
rect 10185 5065 10200 5085
rect 10150 5035 10200 5065
rect 10150 5015 10165 5035
rect 10185 5015 10200 5035
rect 10150 4985 10200 5015
rect 10150 4965 10165 4985
rect 10185 4965 10200 4985
rect 10150 4935 10200 4965
rect 10150 4915 10165 4935
rect 10185 4915 10200 4935
rect 10150 4885 10200 4915
rect 10150 4865 10165 4885
rect 10185 4865 10200 4885
rect 10150 4835 10200 4865
rect 10150 4815 10165 4835
rect 10185 4815 10200 4835
rect 10150 4785 10200 4815
rect 10150 4765 10165 4785
rect 10185 4765 10200 4785
rect 10150 4735 10200 4765
rect 10150 4715 10165 4735
rect 10185 4715 10200 4735
rect 10150 4685 10200 4715
rect 10150 4665 10165 4685
rect 10185 4665 10200 4685
rect 10150 4635 10200 4665
rect 10150 4615 10165 4635
rect 10185 4615 10200 4635
rect 10150 4600 10200 4615
rect 10300 5085 10350 5100
rect 10300 5065 10315 5085
rect 10335 5065 10350 5085
rect 10300 5035 10350 5065
rect 10300 5015 10315 5035
rect 10335 5015 10350 5035
rect 10300 4985 10350 5015
rect 10300 4965 10315 4985
rect 10335 4965 10350 4985
rect 10300 4935 10350 4965
rect 10300 4915 10315 4935
rect 10335 4915 10350 4935
rect 10300 4885 10350 4915
rect 10300 4865 10315 4885
rect 10335 4865 10350 4885
rect 10300 4835 10350 4865
rect 10300 4815 10315 4835
rect 10335 4815 10350 4835
rect 10300 4785 10350 4815
rect 10300 4765 10315 4785
rect 10335 4765 10350 4785
rect 10300 4735 10350 4765
rect 10300 4715 10315 4735
rect 10335 4715 10350 4735
rect 10300 4685 10350 4715
rect 10300 4665 10315 4685
rect 10335 4665 10350 4685
rect 10300 4635 10350 4665
rect 10300 4615 10315 4635
rect 10335 4615 10350 4635
rect 10300 4600 10350 4615
rect 10450 5085 10500 5100
rect 10450 5065 10465 5085
rect 10485 5065 10500 5085
rect 10450 5035 10500 5065
rect 10450 5015 10465 5035
rect 10485 5015 10500 5035
rect 10450 4985 10500 5015
rect 10450 4965 10465 4985
rect 10485 4965 10500 4985
rect 10450 4935 10500 4965
rect 10450 4915 10465 4935
rect 10485 4915 10500 4935
rect 10450 4885 10500 4915
rect 10450 4865 10465 4885
rect 10485 4865 10500 4885
rect 10450 4835 10500 4865
rect 10450 4815 10465 4835
rect 10485 4815 10500 4835
rect 10450 4785 10500 4815
rect 10450 4765 10465 4785
rect 10485 4765 10500 4785
rect 10450 4735 10500 4765
rect 10450 4715 10465 4735
rect 10485 4715 10500 4735
rect 10450 4685 10500 4715
rect 10450 4665 10465 4685
rect 10485 4665 10500 4685
rect 10450 4635 10500 4665
rect 10450 4615 10465 4635
rect 10485 4615 10500 4635
rect 10450 4600 10500 4615
rect 10600 5085 10650 5100
rect 10600 5065 10615 5085
rect 10635 5065 10650 5085
rect 10600 5035 10650 5065
rect 10600 5015 10615 5035
rect 10635 5015 10650 5035
rect 10600 4985 10650 5015
rect 10600 4965 10615 4985
rect 10635 4965 10650 4985
rect 10600 4935 10650 4965
rect 10600 4915 10615 4935
rect 10635 4915 10650 4935
rect 10600 4885 10650 4915
rect 10600 4865 10615 4885
rect 10635 4865 10650 4885
rect 10600 4835 10650 4865
rect 10600 4815 10615 4835
rect 10635 4815 10650 4835
rect 10600 4785 10650 4815
rect 10600 4765 10615 4785
rect 10635 4765 10650 4785
rect 10600 4735 10650 4765
rect 10600 4715 10615 4735
rect 10635 4715 10650 4735
rect 10600 4685 10650 4715
rect 10600 4665 10615 4685
rect 10635 4665 10650 4685
rect 10600 4635 10650 4665
rect 10600 4615 10615 4635
rect 10635 4615 10650 4635
rect 10600 4600 10650 4615
rect 10750 5085 10800 5100
rect 10750 5065 10765 5085
rect 10785 5065 10800 5085
rect 10750 5035 10800 5065
rect 10750 5015 10765 5035
rect 10785 5015 10800 5035
rect 10750 4985 10800 5015
rect 10750 4965 10765 4985
rect 10785 4965 10800 4985
rect 10750 4935 10800 4965
rect 10750 4915 10765 4935
rect 10785 4915 10800 4935
rect 10750 4885 10800 4915
rect 10750 4865 10765 4885
rect 10785 4865 10800 4885
rect 10750 4835 10800 4865
rect 10750 4815 10765 4835
rect 10785 4815 10800 4835
rect 10750 4785 10800 4815
rect 10750 4765 10765 4785
rect 10785 4765 10800 4785
rect 10750 4735 10800 4765
rect 10750 4715 10765 4735
rect 10785 4715 10800 4735
rect 10750 4685 10800 4715
rect 10750 4665 10765 4685
rect 10785 4665 10800 4685
rect 10750 4635 10800 4665
rect 10750 4615 10765 4635
rect 10785 4615 10800 4635
rect 10750 4600 10800 4615
rect 10900 4600 10950 5100
rect 11050 4600 11100 5100
rect 11200 4600 11250 5100
rect 11350 5085 11400 5100
rect 11350 5065 11365 5085
rect 11385 5065 11400 5085
rect 11350 5035 11400 5065
rect 11350 5015 11365 5035
rect 11385 5015 11400 5035
rect 11350 4985 11400 5015
rect 11350 4965 11365 4985
rect 11385 4965 11400 4985
rect 11350 4935 11400 4965
rect 11350 4915 11365 4935
rect 11385 4915 11400 4935
rect 11350 4885 11400 4915
rect 11350 4865 11365 4885
rect 11385 4865 11400 4885
rect 11350 4835 11400 4865
rect 11350 4815 11365 4835
rect 11385 4815 11400 4835
rect 11350 4785 11400 4815
rect 11350 4765 11365 4785
rect 11385 4765 11400 4785
rect 11350 4735 11400 4765
rect 11350 4715 11365 4735
rect 11385 4715 11400 4735
rect 11350 4685 11400 4715
rect 11350 4665 11365 4685
rect 11385 4665 11400 4685
rect 11350 4635 11400 4665
rect 11350 4615 11365 4635
rect 11385 4615 11400 4635
rect 11350 4600 11400 4615
rect 11500 4600 11550 5100
rect 11650 4600 11700 5100
rect 11800 4600 11850 5100
rect 11950 5085 12000 5100
rect 11950 5065 11965 5085
rect 11985 5065 12000 5085
rect 11950 5035 12000 5065
rect 11950 5015 11965 5035
rect 11985 5015 12000 5035
rect 11950 4985 12000 5015
rect 11950 4965 11965 4985
rect 11985 4965 12000 4985
rect 11950 4935 12000 4965
rect 11950 4915 11965 4935
rect 11985 4915 12000 4935
rect 11950 4885 12000 4915
rect 11950 4865 11965 4885
rect 11985 4865 12000 4885
rect 11950 4835 12000 4865
rect 11950 4815 11965 4835
rect 11985 4815 12000 4835
rect 11950 4785 12000 4815
rect 11950 4765 11965 4785
rect 11985 4765 12000 4785
rect 11950 4735 12000 4765
rect 11950 4715 11965 4735
rect 11985 4715 12000 4735
rect 11950 4685 12000 4715
rect 11950 4665 11965 4685
rect 11985 4665 12000 4685
rect 11950 4635 12000 4665
rect 11950 4615 11965 4635
rect 11985 4615 12000 4635
rect 11950 4600 12000 4615
rect 12100 4600 12150 5100
rect 12250 4600 12300 5100
rect 12400 4600 12450 5100
rect 12550 5085 12600 5100
rect 12550 5065 12565 5085
rect 12585 5065 12600 5085
rect 12550 5035 12600 5065
rect 12550 5015 12565 5035
rect 12585 5015 12600 5035
rect 12550 4985 12600 5015
rect 12550 4965 12565 4985
rect 12585 4965 12600 4985
rect 12550 4935 12600 4965
rect 12550 4915 12565 4935
rect 12585 4915 12600 4935
rect 12550 4885 12600 4915
rect 12550 4865 12565 4885
rect 12585 4865 12600 4885
rect 12550 4835 12600 4865
rect 12550 4815 12565 4835
rect 12585 4815 12600 4835
rect 12550 4785 12600 4815
rect 12550 4765 12565 4785
rect 12585 4765 12600 4785
rect 12550 4735 12600 4765
rect 12550 4715 12565 4735
rect 12585 4715 12600 4735
rect 12550 4685 12600 4715
rect 12550 4665 12565 4685
rect 12585 4665 12600 4685
rect 12550 4635 12600 4665
rect 12550 4615 12565 4635
rect 12585 4615 12600 4635
rect 12550 4600 12600 4615
rect 12700 4600 12750 5100
rect 12850 4600 12900 5100
rect 13000 4600 13050 5100
rect 13150 5085 13200 5100
rect 13150 5065 13165 5085
rect 13185 5065 13200 5085
rect 13150 5035 13200 5065
rect 13150 5015 13165 5035
rect 13185 5015 13200 5035
rect 13150 4985 13200 5015
rect 13150 4965 13165 4985
rect 13185 4965 13200 4985
rect 13150 4935 13200 4965
rect 13150 4915 13165 4935
rect 13185 4915 13200 4935
rect 13150 4885 13200 4915
rect 13150 4865 13165 4885
rect 13185 4865 13200 4885
rect 13150 4835 13200 4865
rect 13150 4815 13165 4835
rect 13185 4815 13200 4835
rect 13150 4785 13200 4815
rect 13150 4765 13165 4785
rect 13185 4765 13200 4785
rect 13150 4735 13200 4765
rect 13150 4715 13165 4735
rect 13185 4715 13200 4735
rect 13150 4685 13200 4715
rect 13150 4665 13165 4685
rect 13185 4665 13200 4685
rect 13150 4635 13200 4665
rect 13150 4615 13165 4635
rect 13185 4615 13200 4635
rect 13150 4600 13200 4615
rect 13300 4600 13350 5100
rect 13450 4600 13500 5100
rect 13600 4600 13650 5100
rect 13750 5085 13800 5100
rect 13750 5065 13765 5085
rect 13785 5065 13800 5085
rect 13750 5035 13800 5065
rect 13750 5015 13765 5035
rect 13785 5015 13800 5035
rect 13750 4985 13800 5015
rect 13750 4965 13765 4985
rect 13785 4965 13800 4985
rect 13750 4935 13800 4965
rect 13750 4915 13765 4935
rect 13785 4915 13800 4935
rect 13750 4885 13800 4915
rect 13750 4865 13765 4885
rect 13785 4865 13800 4885
rect 13750 4835 13800 4865
rect 13750 4815 13765 4835
rect 13785 4815 13800 4835
rect 13750 4785 13800 4815
rect 13750 4765 13765 4785
rect 13785 4765 13800 4785
rect 13750 4735 13800 4765
rect 13750 4715 13765 4735
rect 13785 4715 13800 4735
rect 13750 4685 13800 4715
rect 13750 4665 13765 4685
rect 13785 4665 13800 4685
rect 13750 4635 13800 4665
rect 13750 4615 13765 4635
rect 13785 4615 13800 4635
rect 13750 4600 13800 4615
rect 13900 4600 13950 5100
rect 14050 4600 14100 5100
rect 14200 4600 14250 5100
rect 14350 5085 14400 5100
rect 14350 5065 14365 5085
rect 14385 5065 14400 5085
rect 14350 5035 14400 5065
rect 14350 5015 14365 5035
rect 14385 5015 14400 5035
rect 14350 4985 14400 5015
rect 14350 4965 14365 4985
rect 14385 4965 14400 4985
rect 14350 4935 14400 4965
rect 14350 4915 14365 4935
rect 14385 4915 14400 4935
rect 14350 4885 14400 4915
rect 14350 4865 14365 4885
rect 14385 4865 14400 4885
rect 14350 4835 14400 4865
rect 14350 4815 14365 4835
rect 14385 4815 14400 4835
rect 14350 4785 14400 4815
rect 14350 4765 14365 4785
rect 14385 4765 14400 4785
rect 14350 4735 14400 4765
rect 14350 4715 14365 4735
rect 14385 4715 14400 4735
rect 14350 4685 14400 4715
rect 14350 4665 14365 4685
rect 14385 4665 14400 4685
rect 14350 4635 14400 4665
rect 14350 4615 14365 4635
rect 14385 4615 14400 4635
rect 14350 4600 14400 4615
rect 14500 4600 14550 5100
rect 14650 4600 14700 5100
rect 14800 4600 14850 5100
rect 14950 5085 15000 5100
rect 14950 5065 14965 5085
rect 14985 5065 15000 5085
rect 14950 5035 15000 5065
rect 14950 5015 14965 5035
rect 14985 5015 15000 5035
rect 14950 4985 15000 5015
rect 14950 4965 14965 4985
rect 14985 4965 15000 4985
rect 14950 4935 15000 4965
rect 14950 4915 14965 4935
rect 14985 4915 15000 4935
rect 14950 4885 15000 4915
rect 14950 4865 14965 4885
rect 14985 4865 15000 4885
rect 14950 4835 15000 4865
rect 14950 4815 14965 4835
rect 14985 4815 15000 4835
rect 14950 4785 15000 4815
rect 14950 4765 14965 4785
rect 14985 4765 15000 4785
rect 14950 4735 15000 4765
rect 14950 4715 14965 4735
rect 14985 4715 15000 4735
rect 14950 4685 15000 4715
rect 14950 4665 14965 4685
rect 14985 4665 15000 4685
rect 14950 4635 15000 4665
rect 14950 4615 14965 4635
rect 14985 4615 15000 4635
rect 14950 4600 15000 4615
rect 15100 4600 15150 5100
rect 15250 4600 15300 5100
rect 15400 4600 15450 5100
rect 15550 5085 15600 5100
rect 15550 5065 15565 5085
rect 15585 5065 15600 5085
rect 15550 5035 15600 5065
rect 15550 5015 15565 5035
rect 15585 5015 15600 5035
rect 15550 4985 15600 5015
rect 15550 4965 15565 4985
rect 15585 4965 15600 4985
rect 15550 4935 15600 4965
rect 15550 4915 15565 4935
rect 15585 4915 15600 4935
rect 15550 4885 15600 4915
rect 15550 4865 15565 4885
rect 15585 4865 15600 4885
rect 15550 4835 15600 4865
rect 15550 4815 15565 4835
rect 15585 4815 15600 4835
rect 15550 4785 15600 4815
rect 15550 4765 15565 4785
rect 15585 4765 15600 4785
rect 15550 4735 15600 4765
rect 15550 4715 15565 4735
rect 15585 4715 15600 4735
rect 15550 4685 15600 4715
rect 15550 4665 15565 4685
rect 15585 4665 15600 4685
rect 15550 4635 15600 4665
rect 15550 4615 15565 4635
rect 15585 4615 15600 4635
rect 15550 4600 15600 4615
rect 15700 4600 15750 5100
rect 15850 4600 15900 5100
rect 16000 4600 16050 5100
rect 16150 5085 16200 5100
rect 16150 5065 16165 5085
rect 16185 5065 16200 5085
rect 16150 5035 16200 5065
rect 16150 5015 16165 5035
rect 16185 5015 16200 5035
rect 16150 4985 16200 5015
rect 16150 4965 16165 4985
rect 16185 4965 16200 4985
rect 16150 4935 16200 4965
rect 16150 4915 16165 4935
rect 16185 4915 16200 4935
rect 16150 4885 16200 4915
rect 16150 4865 16165 4885
rect 16185 4865 16200 4885
rect 16150 4835 16200 4865
rect 16150 4815 16165 4835
rect 16185 4815 16200 4835
rect 16150 4785 16200 4815
rect 16150 4765 16165 4785
rect 16185 4765 16200 4785
rect 16150 4735 16200 4765
rect 16150 4715 16165 4735
rect 16185 4715 16200 4735
rect 16150 4685 16200 4715
rect 16150 4665 16165 4685
rect 16185 4665 16200 4685
rect 16150 4635 16200 4665
rect 16150 4615 16165 4635
rect 16185 4615 16200 4635
rect 16150 4600 16200 4615
rect 16300 5085 16350 5100
rect 16300 5065 16315 5085
rect 16335 5065 16350 5085
rect 16300 5035 16350 5065
rect 16300 5015 16315 5035
rect 16335 5015 16350 5035
rect 16300 4985 16350 5015
rect 16300 4965 16315 4985
rect 16335 4965 16350 4985
rect 16300 4935 16350 4965
rect 16300 4915 16315 4935
rect 16335 4915 16350 4935
rect 16300 4885 16350 4915
rect 16300 4865 16315 4885
rect 16335 4865 16350 4885
rect 16300 4835 16350 4865
rect 16300 4815 16315 4835
rect 16335 4815 16350 4835
rect 16300 4785 16350 4815
rect 16300 4765 16315 4785
rect 16335 4765 16350 4785
rect 16300 4735 16350 4765
rect 16300 4715 16315 4735
rect 16335 4715 16350 4735
rect 16300 4685 16350 4715
rect 16300 4665 16315 4685
rect 16335 4665 16350 4685
rect 16300 4635 16350 4665
rect 16300 4615 16315 4635
rect 16335 4615 16350 4635
rect 16300 4600 16350 4615
rect 16450 5085 16500 5100
rect 16450 5065 16465 5085
rect 16485 5065 16500 5085
rect 16450 5035 16500 5065
rect 16450 5015 16465 5035
rect 16485 5015 16500 5035
rect 16450 4985 16500 5015
rect 16450 4965 16465 4985
rect 16485 4965 16500 4985
rect 16450 4935 16500 4965
rect 16450 4915 16465 4935
rect 16485 4915 16500 4935
rect 16450 4885 16500 4915
rect 16450 4865 16465 4885
rect 16485 4865 16500 4885
rect 16450 4835 16500 4865
rect 16450 4815 16465 4835
rect 16485 4815 16500 4835
rect 16450 4785 16500 4815
rect 16450 4765 16465 4785
rect 16485 4765 16500 4785
rect 16450 4735 16500 4765
rect 16450 4715 16465 4735
rect 16485 4715 16500 4735
rect 16450 4685 16500 4715
rect 16450 4665 16465 4685
rect 16485 4665 16500 4685
rect 16450 4635 16500 4665
rect 16450 4615 16465 4635
rect 16485 4615 16500 4635
rect 16450 4600 16500 4615
rect 16600 5085 16650 5100
rect 16600 5065 16615 5085
rect 16635 5065 16650 5085
rect 16600 5035 16650 5065
rect 16600 5015 16615 5035
rect 16635 5015 16650 5035
rect 16600 4985 16650 5015
rect 16600 4965 16615 4985
rect 16635 4965 16650 4985
rect 16600 4935 16650 4965
rect 16600 4915 16615 4935
rect 16635 4915 16650 4935
rect 16600 4885 16650 4915
rect 16600 4865 16615 4885
rect 16635 4865 16650 4885
rect 16600 4835 16650 4865
rect 16600 4815 16615 4835
rect 16635 4815 16650 4835
rect 16600 4785 16650 4815
rect 16600 4765 16615 4785
rect 16635 4765 16650 4785
rect 16600 4735 16650 4765
rect 16600 4715 16615 4735
rect 16635 4715 16650 4735
rect 16600 4685 16650 4715
rect 16600 4665 16615 4685
rect 16635 4665 16650 4685
rect 16600 4635 16650 4665
rect 16600 4615 16615 4635
rect 16635 4615 16650 4635
rect 16600 4600 16650 4615
rect 16750 5085 16800 5100
rect 16750 5065 16765 5085
rect 16785 5065 16800 5085
rect 16750 5035 16800 5065
rect 16750 5015 16765 5035
rect 16785 5015 16800 5035
rect 16750 4985 16800 5015
rect 16750 4965 16765 4985
rect 16785 4965 16800 4985
rect 16750 4935 16800 4965
rect 16750 4915 16765 4935
rect 16785 4915 16800 4935
rect 16750 4885 16800 4915
rect 16750 4865 16765 4885
rect 16785 4865 16800 4885
rect 16750 4835 16800 4865
rect 16750 4815 16765 4835
rect 16785 4815 16800 4835
rect 16750 4785 16800 4815
rect 16750 4765 16765 4785
rect 16785 4765 16800 4785
rect 16750 4735 16800 4765
rect 16750 4715 16765 4735
rect 16785 4715 16800 4735
rect 16750 4685 16800 4715
rect 16750 4665 16765 4685
rect 16785 4665 16800 4685
rect 16750 4635 16800 4665
rect 16750 4615 16765 4635
rect 16785 4615 16800 4635
rect 16750 4600 16800 4615
rect 16900 5085 16950 5100
rect 16900 5065 16915 5085
rect 16935 5065 16950 5085
rect 16900 5035 16950 5065
rect 16900 5015 16915 5035
rect 16935 5015 16950 5035
rect 16900 4985 16950 5015
rect 16900 4965 16915 4985
rect 16935 4965 16950 4985
rect 16900 4935 16950 4965
rect 16900 4915 16915 4935
rect 16935 4915 16950 4935
rect 16900 4885 16950 4915
rect 16900 4865 16915 4885
rect 16935 4865 16950 4885
rect 16900 4835 16950 4865
rect 16900 4815 16915 4835
rect 16935 4815 16950 4835
rect 16900 4785 16950 4815
rect 16900 4765 16915 4785
rect 16935 4765 16950 4785
rect 16900 4735 16950 4765
rect 16900 4715 16915 4735
rect 16935 4715 16950 4735
rect 16900 4685 16950 4715
rect 16900 4665 16915 4685
rect 16935 4665 16950 4685
rect 16900 4635 16950 4665
rect 16900 4615 16915 4635
rect 16935 4615 16950 4635
rect 16900 4600 16950 4615
rect 17050 5085 17100 5100
rect 17050 5065 17065 5085
rect 17085 5065 17100 5085
rect 17050 5035 17100 5065
rect 17050 5015 17065 5035
rect 17085 5015 17100 5035
rect 17050 4985 17100 5015
rect 17050 4965 17065 4985
rect 17085 4965 17100 4985
rect 17050 4935 17100 4965
rect 17050 4915 17065 4935
rect 17085 4915 17100 4935
rect 17050 4885 17100 4915
rect 17050 4865 17065 4885
rect 17085 4865 17100 4885
rect 17050 4835 17100 4865
rect 17050 4815 17065 4835
rect 17085 4815 17100 4835
rect 17050 4785 17100 4815
rect 17050 4765 17065 4785
rect 17085 4765 17100 4785
rect 17050 4735 17100 4765
rect 17050 4715 17065 4735
rect 17085 4715 17100 4735
rect 17050 4685 17100 4715
rect 17050 4665 17065 4685
rect 17085 4665 17100 4685
rect 17050 4635 17100 4665
rect 17050 4615 17065 4635
rect 17085 4615 17100 4635
rect 17050 4600 17100 4615
rect 17200 5085 17250 5100
rect 17200 5065 17215 5085
rect 17235 5065 17250 5085
rect 17200 5035 17250 5065
rect 17200 5015 17215 5035
rect 17235 5015 17250 5035
rect 17200 4985 17250 5015
rect 17200 4965 17215 4985
rect 17235 4965 17250 4985
rect 17200 4935 17250 4965
rect 17200 4915 17215 4935
rect 17235 4915 17250 4935
rect 17200 4885 17250 4915
rect 17200 4865 17215 4885
rect 17235 4865 17250 4885
rect 17200 4835 17250 4865
rect 17200 4815 17215 4835
rect 17235 4815 17250 4835
rect 17200 4785 17250 4815
rect 17200 4765 17215 4785
rect 17235 4765 17250 4785
rect 17200 4735 17250 4765
rect 17200 4715 17215 4735
rect 17235 4715 17250 4735
rect 17200 4685 17250 4715
rect 17200 4665 17215 4685
rect 17235 4665 17250 4685
rect 17200 4635 17250 4665
rect 17200 4615 17215 4635
rect 17235 4615 17250 4635
rect 17200 4600 17250 4615
rect 17350 5085 17400 5100
rect 17350 5065 17365 5085
rect 17385 5065 17400 5085
rect 17350 5035 17400 5065
rect 17350 5015 17365 5035
rect 17385 5015 17400 5035
rect 17350 4985 17400 5015
rect 17350 4965 17365 4985
rect 17385 4965 17400 4985
rect 17350 4935 17400 4965
rect 17350 4915 17365 4935
rect 17385 4915 17400 4935
rect 17350 4885 17400 4915
rect 17350 4865 17365 4885
rect 17385 4865 17400 4885
rect 17350 4835 17400 4865
rect 17350 4815 17365 4835
rect 17385 4815 17400 4835
rect 17350 4785 17400 4815
rect 17350 4765 17365 4785
rect 17385 4765 17400 4785
rect 17350 4735 17400 4765
rect 17350 4715 17365 4735
rect 17385 4715 17400 4735
rect 17350 4685 17400 4715
rect 17350 4665 17365 4685
rect 17385 4665 17400 4685
rect 17350 4635 17400 4665
rect 17350 4615 17365 4635
rect 17385 4615 17400 4635
rect 17350 4600 17400 4615
rect 17500 4600 17550 5100
rect 17650 4600 17700 5100
rect 17800 4600 17850 5100
rect 17950 5085 18000 5100
rect 17950 5065 17965 5085
rect 17985 5065 18000 5085
rect 17950 5035 18000 5065
rect 17950 5015 17965 5035
rect 17985 5015 18000 5035
rect 17950 4985 18000 5015
rect 17950 4965 17965 4985
rect 17985 4965 18000 4985
rect 17950 4935 18000 4965
rect 17950 4915 17965 4935
rect 17985 4915 18000 4935
rect 17950 4885 18000 4915
rect 17950 4865 17965 4885
rect 17985 4865 18000 4885
rect 17950 4835 18000 4865
rect 17950 4815 17965 4835
rect 17985 4815 18000 4835
rect 17950 4785 18000 4815
rect 17950 4765 17965 4785
rect 17985 4765 18000 4785
rect 17950 4735 18000 4765
rect 17950 4715 17965 4735
rect 17985 4715 18000 4735
rect 17950 4685 18000 4715
rect 17950 4665 17965 4685
rect 17985 4665 18000 4685
rect 17950 4635 18000 4665
rect 17950 4615 17965 4635
rect 17985 4615 18000 4635
rect 17950 4600 18000 4615
rect 18100 4600 18150 5100
rect 18250 4600 18300 5100
rect 18400 4600 18450 5100
rect 18550 5085 18600 5100
rect 18550 5065 18565 5085
rect 18585 5065 18600 5085
rect 18550 5035 18600 5065
rect 18550 5015 18565 5035
rect 18585 5015 18600 5035
rect 18550 4985 18600 5015
rect 18550 4965 18565 4985
rect 18585 4965 18600 4985
rect 18550 4935 18600 4965
rect 18550 4915 18565 4935
rect 18585 4915 18600 4935
rect 18550 4885 18600 4915
rect 18550 4865 18565 4885
rect 18585 4865 18600 4885
rect 18550 4835 18600 4865
rect 18550 4815 18565 4835
rect 18585 4815 18600 4835
rect 18550 4785 18600 4815
rect 18550 4765 18565 4785
rect 18585 4765 18600 4785
rect 18550 4735 18600 4765
rect 18550 4715 18565 4735
rect 18585 4715 18600 4735
rect 18550 4685 18600 4715
rect 18550 4665 18565 4685
rect 18585 4665 18600 4685
rect 18550 4635 18600 4665
rect 18550 4615 18565 4635
rect 18585 4615 18600 4635
rect 18550 4600 18600 4615
rect 18700 5085 18750 5100
rect 18700 5065 18715 5085
rect 18735 5065 18750 5085
rect 18700 5035 18750 5065
rect 18700 5015 18715 5035
rect 18735 5015 18750 5035
rect 18700 4985 18750 5015
rect 18700 4965 18715 4985
rect 18735 4965 18750 4985
rect 18700 4935 18750 4965
rect 18700 4915 18715 4935
rect 18735 4915 18750 4935
rect 18700 4885 18750 4915
rect 18700 4865 18715 4885
rect 18735 4865 18750 4885
rect 18700 4835 18750 4865
rect 18700 4815 18715 4835
rect 18735 4815 18750 4835
rect 18700 4785 18750 4815
rect 18700 4765 18715 4785
rect 18735 4765 18750 4785
rect 18700 4735 18750 4765
rect 18700 4715 18715 4735
rect 18735 4715 18750 4735
rect 18700 4685 18750 4715
rect 18700 4665 18715 4685
rect 18735 4665 18750 4685
rect 18700 4635 18750 4665
rect 18700 4615 18715 4635
rect 18735 4615 18750 4635
rect 18700 4600 18750 4615
rect 18850 5085 18900 5100
rect 18850 5065 18865 5085
rect 18885 5065 18900 5085
rect 18850 5035 18900 5065
rect 18850 5015 18865 5035
rect 18885 5015 18900 5035
rect 18850 4985 18900 5015
rect 18850 4965 18865 4985
rect 18885 4965 18900 4985
rect 18850 4935 18900 4965
rect 18850 4915 18865 4935
rect 18885 4915 18900 4935
rect 18850 4885 18900 4915
rect 18850 4865 18865 4885
rect 18885 4865 18900 4885
rect 18850 4835 18900 4865
rect 18850 4815 18865 4835
rect 18885 4815 18900 4835
rect 18850 4785 18900 4815
rect 18850 4765 18865 4785
rect 18885 4765 18900 4785
rect 18850 4735 18900 4765
rect 18850 4715 18865 4735
rect 18885 4715 18900 4735
rect 18850 4685 18900 4715
rect 18850 4665 18865 4685
rect 18885 4665 18900 4685
rect 18850 4635 18900 4665
rect 18850 4615 18865 4635
rect 18885 4615 18900 4635
rect 18850 4600 18900 4615
rect 19000 5085 19050 5100
rect 19000 5065 19015 5085
rect 19035 5065 19050 5085
rect 19000 5035 19050 5065
rect 19000 5015 19015 5035
rect 19035 5015 19050 5035
rect 19000 4985 19050 5015
rect 19000 4965 19015 4985
rect 19035 4965 19050 4985
rect 19000 4935 19050 4965
rect 19000 4915 19015 4935
rect 19035 4915 19050 4935
rect 19000 4885 19050 4915
rect 19000 4865 19015 4885
rect 19035 4865 19050 4885
rect 19000 4835 19050 4865
rect 19000 4815 19015 4835
rect 19035 4815 19050 4835
rect 19000 4785 19050 4815
rect 19000 4765 19015 4785
rect 19035 4765 19050 4785
rect 19000 4735 19050 4765
rect 19000 4715 19015 4735
rect 19035 4715 19050 4735
rect 19000 4685 19050 4715
rect 19000 4665 19015 4685
rect 19035 4665 19050 4685
rect 19000 4635 19050 4665
rect 19000 4615 19015 4635
rect 19035 4615 19050 4635
rect 19000 4600 19050 4615
rect 19150 5085 19200 5100
rect 19150 5065 19165 5085
rect 19185 5065 19200 5085
rect 19150 5035 19200 5065
rect 19150 5015 19165 5035
rect 19185 5015 19200 5035
rect 19150 4985 19200 5015
rect 19150 4965 19165 4985
rect 19185 4965 19200 4985
rect 19150 4935 19200 4965
rect 19150 4915 19165 4935
rect 19185 4915 19200 4935
rect 19150 4885 19200 4915
rect 19150 4865 19165 4885
rect 19185 4865 19200 4885
rect 19150 4835 19200 4865
rect 19150 4815 19165 4835
rect 19185 4815 19200 4835
rect 19150 4785 19200 4815
rect 19150 4765 19165 4785
rect 19185 4765 19200 4785
rect 19150 4735 19200 4765
rect 19150 4715 19165 4735
rect 19185 4715 19200 4735
rect 19150 4685 19200 4715
rect 19150 4665 19165 4685
rect 19185 4665 19200 4685
rect 19150 4635 19200 4665
rect 19150 4615 19165 4635
rect 19185 4615 19200 4635
rect 19150 4600 19200 4615
rect 19300 5085 19350 5100
rect 19300 5065 19315 5085
rect 19335 5065 19350 5085
rect 19300 5035 19350 5065
rect 19300 5015 19315 5035
rect 19335 5015 19350 5035
rect 19300 4985 19350 5015
rect 19300 4965 19315 4985
rect 19335 4965 19350 4985
rect 19300 4935 19350 4965
rect 19300 4915 19315 4935
rect 19335 4915 19350 4935
rect 19300 4885 19350 4915
rect 19300 4865 19315 4885
rect 19335 4865 19350 4885
rect 19300 4835 19350 4865
rect 19300 4815 19315 4835
rect 19335 4815 19350 4835
rect 19300 4785 19350 4815
rect 19300 4765 19315 4785
rect 19335 4765 19350 4785
rect 19300 4735 19350 4765
rect 19300 4715 19315 4735
rect 19335 4715 19350 4735
rect 19300 4685 19350 4715
rect 19300 4665 19315 4685
rect 19335 4665 19350 4685
rect 19300 4635 19350 4665
rect 19300 4615 19315 4635
rect 19335 4615 19350 4635
rect 19300 4600 19350 4615
rect 19450 5085 19500 5100
rect 19450 5065 19465 5085
rect 19485 5065 19500 5085
rect 19450 5035 19500 5065
rect 19450 5015 19465 5035
rect 19485 5015 19500 5035
rect 19450 4985 19500 5015
rect 19450 4965 19465 4985
rect 19485 4965 19500 4985
rect 19450 4935 19500 4965
rect 19450 4915 19465 4935
rect 19485 4915 19500 4935
rect 19450 4885 19500 4915
rect 19450 4865 19465 4885
rect 19485 4865 19500 4885
rect 19450 4835 19500 4865
rect 19450 4815 19465 4835
rect 19485 4815 19500 4835
rect 19450 4785 19500 4815
rect 19450 4765 19465 4785
rect 19485 4765 19500 4785
rect 19450 4735 19500 4765
rect 19450 4715 19465 4735
rect 19485 4715 19500 4735
rect 19450 4685 19500 4715
rect 19450 4665 19465 4685
rect 19485 4665 19500 4685
rect 19450 4635 19500 4665
rect 19450 4615 19465 4635
rect 19485 4615 19500 4635
rect 19450 4600 19500 4615
rect 19600 5085 19650 5100
rect 19600 5065 19615 5085
rect 19635 5065 19650 5085
rect 19600 5035 19650 5065
rect 19600 5015 19615 5035
rect 19635 5015 19650 5035
rect 19600 4985 19650 5015
rect 19600 4965 19615 4985
rect 19635 4965 19650 4985
rect 19600 4935 19650 4965
rect 19600 4915 19615 4935
rect 19635 4915 19650 4935
rect 19600 4885 19650 4915
rect 19600 4865 19615 4885
rect 19635 4865 19650 4885
rect 19600 4835 19650 4865
rect 19600 4815 19615 4835
rect 19635 4815 19650 4835
rect 19600 4785 19650 4815
rect 19600 4765 19615 4785
rect 19635 4765 19650 4785
rect 19600 4735 19650 4765
rect 19600 4715 19615 4735
rect 19635 4715 19650 4735
rect 19600 4685 19650 4715
rect 19600 4665 19615 4685
rect 19635 4665 19650 4685
rect 19600 4635 19650 4665
rect 19600 4615 19615 4635
rect 19635 4615 19650 4635
rect 19600 4600 19650 4615
rect 19750 5085 19800 5100
rect 19750 5065 19765 5085
rect 19785 5065 19800 5085
rect 19750 5035 19800 5065
rect 19750 5015 19765 5035
rect 19785 5015 19800 5035
rect 19750 4985 19800 5015
rect 19750 4965 19765 4985
rect 19785 4965 19800 4985
rect 19750 4935 19800 4965
rect 19750 4915 19765 4935
rect 19785 4915 19800 4935
rect 19750 4885 19800 4915
rect 19750 4865 19765 4885
rect 19785 4865 19800 4885
rect 19750 4835 19800 4865
rect 19750 4815 19765 4835
rect 19785 4815 19800 4835
rect 19750 4785 19800 4815
rect 19750 4765 19765 4785
rect 19785 4765 19800 4785
rect 19750 4735 19800 4765
rect 19750 4715 19765 4735
rect 19785 4715 19800 4735
rect 19750 4685 19800 4715
rect 19750 4665 19765 4685
rect 19785 4665 19800 4685
rect 19750 4635 19800 4665
rect 19750 4615 19765 4635
rect 19785 4615 19800 4635
rect 19750 4600 19800 4615
rect 19900 4600 19950 5100
rect 20050 4600 20100 5100
rect 20200 4600 20250 5100
rect 20350 5085 20400 5100
rect 20350 5065 20365 5085
rect 20385 5065 20400 5085
rect 20350 5035 20400 5065
rect 20350 5015 20365 5035
rect 20385 5015 20400 5035
rect 20350 4985 20400 5015
rect 20350 4965 20365 4985
rect 20385 4965 20400 4985
rect 20350 4935 20400 4965
rect 20350 4915 20365 4935
rect 20385 4915 20400 4935
rect 20350 4885 20400 4915
rect 20350 4865 20365 4885
rect 20385 4865 20400 4885
rect 20350 4835 20400 4865
rect 20350 4815 20365 4835
rect 20385 4815 20400 4835
rect 20350 4785 20400 4815
rect 20350 4765 20365 4785
rect 20385 4765 20400 4785
rect 20350 4735 20400 4765
rect 20350 4715 20365 4735
rect 20385 4715 20400 4735
rect 20350 4685 20400 4715
rect 20350 4665 20365 4685
rect 20385 4665 20400 4685
rect 20350 4635 20400 4665
rect 20350 4615 20365 4635
rect 20385 4615 20400 4635
rect 20350 4600 20400 4615
rect -650 4435 -600 4450
rect -650 4415 -635 4435
rect -615 4415 -600 4435
rect -650 4385 -600 4415
rect -650 4365 -635 4385
rect -615 4365 -600 4385
rect -650 4335 -600 4365
rect -650 4315 -635 4335
rect -615 4315 -600 4335
rect -650 4285 -600 4315
rect -650 4265 -635 4285
rect -615 4265 -600 4285
rect -650 4235 -600 4265
rect -650 4215 -635 4235
rect -615 4215 -600 4235
rect -650 4185 -600 4215
rect -650 4165 -635 4185
rect -615 4165 -600 4185
rect -650 4135 -600 4165
rect -650 4115 -635 4135
rect -615 4115 -600 4135
rect -650 4085 -600 4115
rect -650 4065 -635 4085
rect -615 4065 -600 4085
rect -650 4035 -600 4065
rect -650 4015 -635 4035
rect -615 4015 -600 4035
rect -650 3985 -600 4015
rect -650 3965 -635 3985
rect -615 3965 -600 3985
rect -650 3950 -600 3965
rect -500 4435 -450 4450
rect -500 4415 -485 4435
rect -465 4415 -450 4435
rect -500 4385 -450 4415
rect -500 4365 -485 4385
rect -465 4365 -450 4385
rect -500 4335 -450 4365
rect -500 4315 -485 4335
rect -465 4315 -450 4335
rect -500 4285 -450 4315
rect -500 4265 -485 4285
rect -465 4265 -450 4285
rect -500 4235 -450 4265
rect -500 4215 -485 4235
rect -465 4215 -450 4235
rect -500 4185 -450 4215
rect -500 4165 -485 4185
rect -465 4165 -450 4185
rect -500 4135 -450 4165
rect -500 4115 -485 4135
rect -465 4115 -450 4135
rect -500 4085 -450 4115
rect -500 4065 -485 4085
rect -465 4065 -450 4085
rect -500 4035 -450 4065
rect -500 4015 -485 4035
rect -465 4015 -450 4035
rect -500 3985 -450 4015
rect -500 3965 -485 3985
rect -465 3965 -450 3985
rect -500 3950 -450 3965
rect -350 4435 -300 4450
rect -350 4415 -335 4435
rect -315 4415 -300 4435
rect -350 4385 -300 4415
rect -350 4365 -335 4385
rect -315 4365 -300 4385
rect -350 4335 -300 4365
rect -350 4315 -335 4335
rect -315 4315 -300 4335
rect -350 4285 -300 4315
rect -350 4265 -335 4285
rect -315 4265 -300 4285
rect -350 4235 -300 4265
rect -350 4215 -335 4235
rect -315 4215 -300 4235
rect -350 4185 -300 4215
rect -350 4165 -335 4185
rect -315 4165 -300 4185
rect -350 4135 -300 4165
rect -350 4115 -335 4135
rect -315 4115 -300 4135
rect -350 4085 -300 4115
rect -350 4065 -335 4085
rect -315 4065 -300 4085
rect -350 4035 -300 4065
rect -350 4015 -335 4035
rect -315 4015 -300 4035
rect -350 3985 -300 4015
rect -350 3965 -335 3985
rect -315 3965 -300 3985
rect -350 3950 -300 3965
rect -200 4435 -150 4450
rect -200 4415 -185 4435
rect -165 4415 -150 4435
rect -200 4385 -150 4415
rect -200 4365 -185 4385
rect -165 4365 -150 4385
rect -200 4335 -150 4365
rect -200 4315 -185 4335
rect -165 4315 -150 4335
rect -200 4285 -150 4315
rect -200 4265 -185 4285
rect -165 4265 -150 4285
rect -200 4235 -150 4265
rect -200 4215 -185 4235
rect -165 4215 -150 4235
rect -200 4185 -150 4215
rect -200 4165 -185 4185
rect -165 4165 -150 4185
rect -200 4135 -150 4165
rect -200 4115 -185 4135
rect -165 4115 -150 4135
rect -200 4085 -150 4115
rect -200 4065 -185 4085
rect -165 4065 -150 4085
rect -200 4035 -150 4065
rect -200 4015 -185 4035
rect -165 4015 -150 4035
rect -200 3985 -150 4015
rect -200 3965 -185 3985
rect -165 3965 -150 3985
rect -200 3950 -150 3965
rect -50 4435 0 4450
rect -50 4415 -35 4435
rect -15 4415 0 4435
rect -50 4385 0 4415
rect -50 4365 -35 4385
rect -15 4365 0 4385
rect -50 4335 0 4365
rect -50 4315 -35 4335
rect -15 4315 0 4335
rect -50 4285 0 4315
rect -50 4265 -35 4285
rect -15 4265 0 4285
rect -50 4235 0 4265
rect -50 4215 -35 4235
rect -15 4215 0 4235
rect -50 4185 0 4215
rect -50 4165 -35 4185
rect -15 4165 0 4185
rect -50 4135 0 4165
rect -50 4115 -35 4135
rect -15 4115 0 4135
rect -50 4085 0 4115
rect -50 4065 -35 4085
rect -15 4065 0 4085
rect -50 4035 0 4065
rect -50 4015 -35 4035
rect -15 4015 0 4035
rect -50 3985 0 4015
rect -50 3965 -35 3985
rect -15 3965 0 3985
rect -50 3950 0 3965
rect 100 3950 150 4450
rect 250 3950 300 4450
rect 400 3950 450 4450
rect 550 4435 600 4450
rect 550 4415 565 4435
rect 585 4415 600 4435
rect 550 4385 600 4415
rect 550 4365 565 4385
rect 585 4365 600 4385
rect 550 4335 600 4365
rect 550 4315 565 4335
rect 585 4315 600 4335
rect 550 4285 600 4315
rect 550 4265 565 4285
rect 585 4265 600 4285
rect 550 4235 600 4265
rect 550 4215 565 4235
rect 585 4215 600 4235
rect 550 4185 600 4215
rect 550 4165 565 4185
rect 585 4165 600 4185
rect 550 4135 600 4165
rect 550 4115 565 4135
rect 585 4115 600 4135
rect 550 4085 600 4115
rect 550 4065 565 4085
rect 585 4065 600 4085
rect 550 4035 600 4065
rect 550 4015 565 4035
rect 585 4015 600 4035
rect 550 3985 600 4015
rect 550 3965 565 3985
rect 585 3965 600 3985
rect 550 3950 600 3965
rect 700 4435 750 4450
rect 700 4415 715 4435
rect 735 4415 750 4435
rect 700 4385 750 4415
rect 700 4365 715 4385
rect 735 4365 750 4385
rect 700 4335 750 4365
rect 700 4315 715 4335
rect 735 4315 750 4335
rect 700 4285 750 4315
rect 700 4265 715 4285
rect 735 4265 750 4285
rect 700 4235 750 4265
rect 700 4215 715 4235
rect 735 4215 750 4235
rect 700 4185 750 4215
rect 700 4165 715 4185
rect 735 4165 750 4185
rect 700 4135 750 4165
rect 700 4115 715 4135
rect 735 4115 750 4135
rect 700 4085 750 4115
rect 700 4065 715 4085
rect 735 4065 750 4085
rect 700 4035 750 4065
rect 700 4015 715 4035
rect 735 4015 750 4035
rect 700 3985 750 4015
rect 700 3965 715 3985
rect 735 3965 750 3985
rect 700 3950 750 3965
rect 850 4435 900 4450
rect 850 4415 865 4435
rect 885 4415 900 4435
rect 850 4385 900 4415
rect 850 4365 865 4385
rect 885 4365 900 4385
rect 850 4335 900 4365
rect 850 4315 865 4335
rect 885 4315 900 4335
rect 850 4285 900 4315
rect 850 4265 865 4285
rect 885 4265 900 4285
rect 850 4235 900 4265
rect 850 4215 865 4235
rect 885 4215 900 4235
rect 850 4185 900 4215
rect 850 4165 865 4185
rect 885 4165 900 4185
rect 850 4135 900 4165
rect 850 4115 865 4135
rect 885 4115 900 4135
rect 850 4085 900 4115
rect 850 4065 865 4085
rect 885 4065 900 4085
rect 850 4035 900 4065
rect 850 4015 865 4035
rect 885 4015 900 4035
rect 850 3985 900 4015
rect 850 3965 865 3985
rect 885 3965 900 3985
rect 850 3950 900 3965
rect 1000 4435 1050 4450
rect 1000 4415 1015 4435
rect 1035 4415 1050 4435
rect 1000 4385 1050 4415
rect 1000 4365 1015 4385
rect 1035 4365 1050 4385
rect 1000 4335 1050 4365
rect 1000 4315 1015 4335
rect 1035 4315 1050 4335
rect 1000 4285 1050 4315
rect 1000 4265 1015 4285
rect 1035 4265 1050 4285
rect 1000 4235 1050 4265
rect 1000 4215 1015 4235
rect 1035 4215 1050 4235
rect 1000 4185 1050 4215
rect 1000 4165 1015 4185
rect 1035 4165 1050 4185
rect 1000 4135 1050 4165
rect 1000 4115 1015 4135
rect 1035 4115 1050 4135
rect 1000 4085 1050 4115
rect 1000 4065 1015 4085
rect 1035 4065 1050 4085
rect 1000 4035 1050 4065
rect 1000 4015 1015 4035
rect 1035 4015 1050 4035
rect 1000 3985 1050 4015
rect 1000 3965 1015 3985
rect 1035 3965 1050 3985
rect 1000 3950 1050 3965
rect 1150 4435 1200 4450
rect 1150 4415 1165 4435
rect 1185 4415 1200 4435
rect 1150 4385 1200 4415
rect 1150 4365 1165 4385
rect 1185 4365 1200 4385
rect 1150 4335 1200 4365
rect 1150 4315 1165 4335
rect 1185 4315 1200 4335
rect 1150 4285 1200 4315
rect 1150 4265 1165 4285
rect 1185 4265 1200 4285
rect 1150 4235 1200 4265
rect 1150 4215 1165 4235
rect 1185 4215 1200 4235
rect 1150 4185 1200 4215
rect 1150 4165 1165 4185
rect 1185 4165 1200 4185
rect 1150 4135 1200 4165
rect 1150 4115 1165 4135
rect 1185 4115 1200 4135
rect 1150 4085 1200 4115
rect 1150 4065 1165 4085
rect 1185 4065 1200 4085
rect 1150 4035 1200 4065
rect 1150 4015 1165 4035
rect 1185 4015 1200 4035
rect 1150 3985 1200 4015
rect 1150 3965 1165 3985
rect 1185 3965 1200 3985
rect 1150 3950 1200 3965
rect 1300 4435 1350 4450
rect 1300 4415 1315 4435
rect 1335 4415 1350 4435
rect 1300 4385 1350 4415
rect 1300 4365 1315 4385
rect 1335 4365 1350 4385
rect 1300 4335 1350 4365
rect 1300 4315 1315 4335
rect 1335 4315 1350 4335
rect 1300 4285 1350 4315
rect 1300 4265 1315 4285
rect 1335 4265 1350 4285
rect 1300 4235 1350 4265
rect 1300 4215 1315 4235
rect 1335 4215 1350 4235
rect 1300 4185 1350 4215
rect 1300 4165 1315 4185
rect 1335 4165 1350 4185
rect 1300 4135 1350 4165
rect 1300 4115 1315 4135
rect 1335 4115 1350 4135
rect 1300 4085 1350 4115
rect 1300 4065 1315 4085
rect 1335 4065 1350 4085
rect 1300 4035 1350 4065
rect 1300 4015 1315 4035
rect 1335 4015 1350 4035
rect 1300 3985 1350 4015
rect 1300 3965 1315 3985
rect 1335 3965 1350 3985
rect 1300 3950 1350 3965
rect 1450 4435 1500 4450
rect 1450 4415 1465 4435
rect 1485 4415 1500 4435
rect 1450 4385 1500 4415
rect 1450 4365 1465 4385
rect 1485 4365 1500 4385
rect 1450 4335 1500 4365
rect 1450 4315 1465 4335
rect 1485 4315 1500 4335
rect 1450 4285 1500 4315
rect 1450 4265 1465 4285
rect 1485 4265 1500 4285
rect 1450 4235 1500 4265
rect 1450 4215 1465 4235
rect 1485 4215 1500 4235
rect 1450 4185 1500 4215
rect 1450 4165 1465 4185
rect 1485 4165 1500 4185
rect 1450 4135 1500 4165
rect 1450 4115 1465 4135
rect 1485 4115 1500 4135
rect 1450 4085 1500 4115
rect 1450 4065 1465 4085
rect 1485 4065 1500 4085
rect 1450 4035 1500 4065
rect 1450 4015 1465 4035
rect 1485 4015 1500 4035
rect 1450 3985 1500 4015
rect 1450 3965 1465 3985
rect 1485 3965 1500 3985
rect 1450 3950 1500 3965
rect 1600 4435 1650 4450
rect 1600 4415 1615 4435
rect 1635 4415 1650 4435
rect 1600 4385 1650 4415
rect 1600 4365 1615 4385
rect 1635 4365 1650 4385
rect 1600 4335 1650 4365
rect 1600 4315 1615 4335
rect 1635 4315 1650 4335
rect 1600 4285 1650 4315
rect 1600 4265 1615 4285
rect 1635 4265 1650 4285
rect 1600 4235 1650 4265
rect 1600 4215 1615 4235
rect 1635 4215 1650 4235
rect 1600 4185 1650 4215
rect 1600 4165 1615 4185
rect 1635 4165 1650 4185
rect 1600 4135 1650 4165
rect 1600 4115 1615 4135
rect 1635 4115 1650 4135
rect 1600 4085 1650 4115
rect 1600 4065 1615 4085
rect 1635 4065 1650 4085
rect 1600 4035 1650 4065
rect 1600 4015 1615 4035
rect 1635 4015 1650 4035
rect 1600 3985 1650 4015
rect 1600 3965 1615 3985
rect 1635 3965 1650 3985
rect 1600 3950 1650 3965
rect 1750 4435 1800 4450
rect 1750 4415 1765 4435
rect 1785 4415 1800 4435
rect 1750 4385 1800 4415
rect 1750 4365 1765 4385
rect 1785 4365 1800 4385
rect 1750 4335 1800 4365
rect 1750 4315 1765 4335
rect 1785 4315 1800 4335
rect 1750 4285 1800 4315
rect 1750 4265 1765 4285
rect 1785 4265 1800 4285
rect 1750 4235 1800 4265
rect 1750 4215 1765 4235
rect 1785 4215 1800 4235
rect 1750 4185 1800 4215
rect 1750 4165 1765 4185
rect 1785 4165 1800 4185
rect 1750 4135 1800 4165
rect 1750 4115 1765 4135
rect 1785 4115 1800 4135
rect 1750 4085 1800 4115
rect 1750 4065 1765 4085
rect 1785 4065 1800 4085
rect 1750 4035 1800 4065
rect 1750 4015 1765 4035
rect 1785 4015 1800 4035
rect 1750 3985 1800 4015
rect 1750 3965 1765 3985
rect 1785 3965 1800 3985
rect 1750 3950 1800 3965
rect 1900 4435 1950 4450
rect 1900 4415 1915 4435
rect 1935 4415 1950 4435
rect 1900 4385 1950 4415
rect 1900 4365 1915 4385
rect 1935 4365 1950 4385
rect 1900 4335 1950 4365
rect 1900 4315 1915 4335
rect 1935 4315 1950 4335
rect 1900 4285 1950 4315
rect 1900 4265 1915 4285
rect 1935 4265 1950 4285
rect 1900 4235 1950 4265
rect 1900 4215 1915 4235
rect 1935 4215 1950 4235
rect 1900 4185 1950 4215
rect 1900 4165 1915 4185
rect 1935 4165 1950 4185
rect 1900 4135 1950 4165
rect 1900 4115 1915 4135
rect 1935 4115 1950 4135
rect 1900 4085 1950 4115
rect 1900 4065 1915 4085
rect 1935 4065 1950 4085
rect 1900 4035 1950 4065
rect 1900 4015 1915 4035
rect 1935 4015 1950 4035
rect 1900 3985 1950 4015
rect 1900 3965 1915 3985
rect 1935 3965 1950 3985
rect 1900 3950 1950 3965
rect 2050 4435 2100 4450
rect 2050 4415 2065 4435
rect 2085 4415 2100 4435
rect 2050 4385 2100 4415
rect 2050 4365 2065 4385
rect 2085 4365 2100 4385
rect 2050 4335 2100 4365
rect 2050 4315 2065 4335
rect 2085 4315 2100 4335
rect 2050 4285 2100 4315
rect 2050 4265 2065 4285
rect 2085 4265 2100 4285
rect 2050 4235 2100 4265
rect 2050 4215 2065 4235
rect 2085 4215 2100 4235
rect 2050 4185 2100 4215
rect 2050 4165 2065 4185
rect 2085 4165 2100 4185
rect 2050 4135 2100 4165
rect 2050 4115 2065 4135
rect 2085 4115 2100 4135
rect 2050 4085 2100 4115
rect 2050 4065 2065 4085
rect 2085 4065 2100 4085
rect 2050 4035 2100 4065
rect 2050 4015 2065 4035
rect 2085 4015 2100 4035
rect 2050 3985 2100 4015
rect 2050 3965 2065 3985
rect 2085 3965 2100 3985
rect 2050 3950 2100 3965
rect 2200 4435 2250 4450
rect 2200 4415 2215 4435
rect 2235 4415 2250 4435
rect 2200 4385 2250 4415
rect 2200 4365 2215 4385
rect 2235 4365 2250 4385
rect 2200 4335 2250 4365
rect 2200 4315 2215 4335
rect 2235 4315 2250 4335
rect 2200 4285 2250 4315
rect 2200 4265 2215 4285
rect 2235 4265 2250 4285
rect 2200 4235 2250 4265
rect 2200 4215 2215 4235
rect 2235 4215 2250 4235
rect 2200 4185 2250 4215
rect 2200 4165 2215 4185
rect 2235 4165 2250 4185
rect 2200 4135 2250 4165
rect 2200 4115 2215 4135
rect 2235 4115 2250 4135
rect 2200 4085 2250 4115
rect 2200 4065 2215 4085
rect 2235 4065 2250 4085
rect 2200 4035 2250 4065
rect 2200 4015 2215 4035
rect 2235 4015 2250 4035
rect 2200 3985 2250 4015
rect 2200 3965 2215 3985
rect 2235 3965 2250 3985
rect 2200 3950 2250 3965
rect 2350 4435 2400 4450
rect 2350 4415 2365 4435
rect 2385 4415 2400 4435
rect 2350 4385 2400 4415
rect 2350 4365 2365 4385
rect 2385 4365 2400 4385
rect 2350 4335 2400 4365
rect 2350 4315 2365 4335
rect 2385 4315 2400 4335
rect 2350 4285 2400 4315
rect 2350 4265 2365 4285
rect 2385 4265 2400 4285
rect 2350 4235 2400 4265
rect 2350 4215 2365 4235
rect 2385 4215 2400 4235
rect 2350 4185 2400 4215
rect 2350 4165 2365 4185
rect 2385 4165 2400 4185
rect 2350 4135 2400 4165
rect 2350 4115 2365 4135
rect 2385 4115 2400 4135
rect 2350 4085 2400 4115
rect 2350 4065 2365 4085
rect 2385 4065 2400 4085
rect 2350 4035 2400 4065
rect 2350 4015 2365 4035
rect 2385 4015 2400 4035
rect 2350 3985 2400 4015
rect 2350 3965 2365 3985
rect 2385 3965 2400 3985
rect 2350 3950 2400 3965
rect 2500 4435 2550 4450
rect 2500 4415 2515 4435
rect 2535 4415 2550 4435
rect 2500 4385 2550 4415
rect 2500 4365 2515 4385
rect 2535 4365 2550 4385
rect 2500 4335 2550 4365
rect 2500 4315 2515 4335
rect 2535 4315 2550 4335
rect 2500 4285 2550 4315
rect 2500 4265 2515 4285
rect 2535 4265 2550 4285
rect 2500 4235 2550 4265
rect 2500 4215 2515 4235
rect 2535 4215 2550 4235
rect 2500 4185 2550 4215
rect 2500 4165 2515 4185
rect 2535 4165 2550 4185
rect 2500 4135 2550 4165
rect 2500 4115 2515 4135
rect 2535 4115 2550 4135
rect 2500 4085 2550 4115
rect 2500 4065 2515 4085
rect 2535 4065 2550 4085
rect 2500 4035 2550 4065
rect 2500 4015 2515 4035
rect 2535 4015 2550 4035
rect 2500 3985 2550 4015
rect 2500 3965 2515 3985
rect 2535 3965 2550 3985
rect 2500 3950 2550 3965
rect 2650 4435 2700 4450
rect 2650 4415 2665 4435
rect 2685 4415 2700 4435
rect 2650 4385 2700 4415
rect 2650 4365 2665 4385
rect 2685 4365 2700 4385
rect 2650 4335 2700 4365
rect 2650 4315 2665 4335
rect 2685 4315 2700 4335
rect 2650 4285 2700 4315
rect 2650 4265 2665 4285
rect 2685 4265 2700 4285
rect 2650 4235 2700 4265
rect 2650 4215 2665 4235
rect 2685 4215 2700 4235
rect 2650 4185 2700 4215
rect 2650 4165 2665 4185
rect 2685 4165 2700 4185
rect 2650 4135 2700 4165
rect 2650 4115 2665 4135
rect 2685 4115 2700 4135
rect 2650 4085 2700 4115
rect 2650 4065 2665 4085
rect 2685 4065 2700 4085
rect 2650 4035 2700 4065
rect 2650 4015 2665 4035
rect 2685 4015 2700 4035
rect 2650 3985 2700 4015
rect 2650 3965 2665 3985
rect 2685 3965 2700 3985
rect 2650 3950 2700 3965
rect 2800 4435 2850 4450
rect 2800 4415 2815 4435
rect 2835 4415 2850 4435
rect 2800 4385 2850 4415
rect 2800 4365 2815 4385
rect 2835 4365 2850 4385
rect 2800 4335 2850 4365
rect 2800 4315 2815 4335
rect 2835 4315 2850 4335
rect 2800 4285 2850 4315
rect 2800 4265 2815 4285
rect 2835 4265 2850 4285
rect 2800 4235 2850 4265
rect 2800 4215 2815 4235
rect 2835 4215 2850 4235
rect 2800 4185 2850 4215
rect 2800 4165 2815 4185
rect 2835 4165 2850 4185
rect 2800 4135 2850 4165
rect 2800 4115 2815 4135
rect 2835 4115 2850 4135
rect 2800 4085 2850 4115
rect 2800 4065 2815 4085
rect 2835 4065 2850 4085
rect 2800 4035 2850 4065
rect 2800 4015 2815 4035
rect 2835 4015 2850 4035
rect 2800 3985 2850 4015
rect 2800 3965 2815 3985
rect 2835 3965 2850 3985
rect 2800 3950 2850 3965
rect 2950 4435 3000 4450
rect 2950 4415 2965 4435
rect 2985 4415 3000 4435
rect 2950 4385 3000 4415
rect 2950 4365 2965 4385
rect 2985 4365 3000 4385
rect 2950 4335 3000 4365
rect 2950 4315 2965 4335
rect 2985 4315 3000 4335
rect 2950 4285 3000 4315
rect 2950 4265 2965 4285
rect 2985 4265 3000 4285
rect 2950 4235 3000 4265
rect 2950 4215 2965 4235
rect 2985 4215 3000 4235
rect 2950 4185 3000 4215
rect 2950 4165 2965 4185
rect 2985 4165 3000 4185
rect 2950 4135 3000 4165
rect 2950 4115 2965 4135
rect 2985 4115 3000 4135
rect 2950 4085 3000 4115
rect 2950 4065 2965 4085
rect 2985 4065 3000 4085
rect 2950 4035 3000 4065
rect 2950 4015 2965 4035
rect 2985 4015 3000 4035
rect 2950 3985 3000 4015
rect 2950 3965 2965 3985
rect 2985 3965 3000 3985
rect 2950 3950 3000 3965
rect 3100 4435 3150 4450
rect 3100 4415 3115 4435
rect 3135 4415 3150 4435
rect 3100 4385 3150 4415
rect 3100 4365 3115 4385
rect 3135 4365 3150 4385
rect 3100 4335 3150 4365
rect 3100 4315 3115 4335
rect 3135 4315 3150 4335
rect 3100 4285 3150 4315
rect 3100 4265 3115 4285
rect 3135 4265 3150 4285
rect 3100 4235 3150 4265
rect 3100 4215 3115 4235
rect 3135 4215 3150 4235
rect 3100 4185 3150 4215
rect 3100 4165 3115 4185
rect 3135 4165 3150 4185
rect 3100 4135 3150 4165
rect 3100 4115 3115 4135
rect 3135 4115 3150 4135
rect 3100 4085 3150 4115
rect 3100 4065 3115 4085
rect 3135 4065 3150 4085
rect 3100 4035 3150 4065
rect 3100 4015 3115 4035
rect 3135 4015 3150 4035
rect 3100 3985 3150 4015
rect 3100 3965 3115 3985
rect 3135 3965 3150 3985
rect 3100 3950 3150 3965
rect 3250 4435 3300 4450
rect 3250 4415 3265 4435
rect 3285 4415 3300 4435
rect 3250 4385 3300 4415
rect 3250 4365 3265 4385
rect 3285 4365 3300 4385
rect 3250 4335 3300 4365
rect 3250 4315 3265 4335
rect 3285 4315 3300 4335
rect 3250 4285 3300 4315
rect 3250 4265 3265 4285
rect 3285 4265 3300 4285
rect 3250 4235 3300 4265
rect 3250 4215 3265 4235
rect 3285 4215 3300 4235
rect 3250 4185 3300 4215
rect 3250 4165 3265 4185
rect 3285 4165 3300 4185
rect 3250 4135 3300 4165
rect 3250 4115 3265 4135
rect 3285 4115 3300 4135
rect 3250 4085 3300 4115
rect 3250 4065 3265 4085
rect 3285 4065 3300 4085
rect 3250 4035 3300 4065
rect 3250 4015 3265 4035
rect 3285 4015 3300 4035
rect 3250 3985 3300 4015
rect 3250 3965 3265 3985
rect 3285 3965 3300 3985
rect 3250 3950 3300 3965
rect 3400 4435 3450 4450
rect 3400 4415 3415 4435
rect 3435 4415 3450 4435
rect 3400 4385 3450 4415
rect 3400 4365 3415 4385
rect 3435 4365 3450 4385
rect 3400 4335 3450 4365
rect 3400 4315 3415 4335
rect 3435 4315 3450 4335
rect 3400 4285 3450 4315
rect 3400 4265 3415 4285
rect 3435 4265 3450 4285
rect 3400 4235 3450 4265
rect 3400 4215 3415 4235
rect 3435 4215 3450 4235
rect 3400 4185 3450 4215
rect 3400 4165 3415 4185
rect 3435 4165 3450 4185
rect 3400 4135 3450 4165
rect 3400 4115 3415 4135
rect 3435 4115 3450 4135
rect 3400 4085 3450 4115
rect 3400 4065 3415 4085
rect 3435 4065 3450 4085
rect 3400 4035 3450 4065
rect 3400 4015 3415 4035
rect 3435 4015 3450 4035
rect 3400 3985 3450 4015
rect 3400 3965 3415 3985
rect 3435 3965 3450 3985
rect 3400 3950 3450 3965
rect 3550 4435 3600 4450
rect 3550 4415 3565 4435
rect 3585 4415 3600 4435
rect 3550 4385 3600 4415
rect 3550 4365 3565 4385
rect 3585 4365 3600 4385
rect 3550 4335 3600 4365
rect 3550 4315 3565 4335
rect 3585 4315 3600 4335
rect 3550 4285 3600 4315
rect 3550 4265 3565 4285
rect 3585 4265 3600 4285
rect 3550 4235 3600 4265
rect 3550 4215 3565 4235
rect 3585 4215 3600 4235
rect 3550 4185 3600 4215
rect 3550 4165 3565 4185
rect 3585 4165 3600 4185
rect 3550 4135 3600 4165
rect 3550 4115 3565 4135
rect 3585 4115 3600 4135
rect 3550 4085 3600 4115
rect 3550 4065 3565 4085
rect 3585 4065 3600 4085
rect 3550 4035 3600 4065
rect 3550 4015 3565 4035
rect 3585 4015 3600 4035
rect 3550 3985 3600 4015
rect 3550 3965 3565 3985
rect 3585 3965 3600 3985
rect 3550 3950 3600 3965
rect 3700 3950 3750 4450
rect 3850 3950 3900 4450
rect 4000 3950 4050 4450
rect 4150 4435 4200 4450
rect 4150 4415 4165 4435
rect 4185 4415 4200 4435
rect 4150 4385 4200 4415
rect 4150 4365 4165 4385
rect 4185 4365 4200 4385
rect 4150 4335 4200 4365
rect 4150 4315 4165 4335
rect 4185 4315 4200 4335
rect 4150 4285 4200 4315
rect 4150 4265 4165 4285
rect 4185 4265 4200 4285
rect 4150 4235 4200 4265
rect 4150 4215 4165 4235
rect 4185 4215 4200 4235
rect 4150 4185 4200 4215
rect 4150 4165 4165 4185
rect 4185 4165 4200 4185
rect 4150 4135 4200 4165
rect 4150 4115 4165 4135
rect 4185 4115 4200 4135
rect 4150 4085 4200 4115
rect 4150 4065 4165 4085
rect 4185 4065 4200 4085
rect 4150 4035 4200 4065
rect 4150 4015 4165 4035
rect 4185 4015 4200 4035
rect 4150 3985 4200 4015
rect 4150 3965 4165 3985
rect 4185 3965 4200 3985
rect 4150 3950 4200 3965
rect 4300 3950 4350 4450
rect 4450 3950 4500 4450
rect 4600 3950 4650 4450
rect 4750 4435 4800 4450
rect 4750 4415 4765 4435
rect 4785 4415 4800 4435
rect 4750 4385 4800 4415
rect 4750 4365 4765 4385
rect 4785 4365 4800 4385
rect 4750 4335 4800 4365
rect 4750 4315 4765 4335
rect 4785 4315 4800 4335
rect 4750 4285 4800 4315
rect 4750 4265 4765 4285
rect 4785 4265 4800 4285
rect 4750 4235 4800 4265
rect 4750 4215 4765 4235
rect 4785 4215 4800 4235
rect 4750 4185 4800 4215
rect 4750 4165 4765 4185
rect 4785 4165 4800 4185
rect 4750 4135 4800 4165
rect 4750 4115 4765 4135
rect 4785 4115 4800 4135
rect 4750 4085 4800 4115
rect 4750 4065 4765 4085
rect 4785 4065 4800 4085
rect 4750 4035 4800 4065
rect 4750 4015 4765 4035
rect 4785 4015 4800 4035
rect 4750 3985 4800 4015
rect 4750 3965 4765 3985
rect 4785 3965 4800 3985
rect 4750 3950 4800 3965
rect 4900 4435 4950 4450
rect 4900 4415 4915 4435
rect 4935 4415 4950 4435
rect 4900 4385 4950 4415
rect 4900 4365 4915 4385
rect 4935 4365 4950 4385
rect 4900 4335 4950 4365
rect 4900 4315 4915 4335
rect 4935 4315 4950 4335
rect 4900 4285 4950 4315
rect 4900 4265 4915 4285
rect 4935 4265 4950 4285
rect 4900 4235 4950 4265
rect 4900 4215 4915 4235
rect 4935 4215 4950 4235
rect 4900 4185 4950 4215
rect 4900 4165 4915 4185
rect 4935 4165 4950 4185
rect 4900 4135 4950 4165
rect 4900 4115 4915 4135
rect 4935 4115 4950 4135
rect 4900 4085 4950 4115
rect 4900 4065 4915 4085
rect 4935 4065 4950 4085
rect 4900 4035 4950 4065
rect 4900 4015 4915 4035
rect 4935 4015 4950 4035
rect 4900 3985 4950 4015
rect 4900 3965 4915 3985
rect 4935 3965 4950 3985
rect 4900 3950 4950 3965
rect 5050 4435 5100 4450
rect 5050 4415 5065 4435
rect 5085 4415 5100 4435
rect 5050 4385 5100 4415
rect 5050 4365 5065 4385
rect 5085 4365 5100 4385
rect 5050 4335 5100 4365
rect 5050 4315 5065 4335
rect 5085 4315 5100 4335
rect 5050 4285 5100 4315
rect 5050 4265 5065 4285
rect 5085 4265 5100 4285
rect 5050 4235 5100 4265
rect 5050 4215 5065 4235
rect 5085 4215 5100 4235
rect 5050 4185 5100 4215
rect 5050 4165 5065 4185
rect 5085 4165 5100 4185
rect 5050 4135 5100 4165
rect 5050 4115 5065 4135
rect 5085 4115 5100 4135
rect 5050 4085 5100 4115
rect 5050 4065 5065 4085
rect 5085 4065 5100 4085
rect 5050 4035 5100 4065
rect 5050 4015 5065 4035
rect 5085 4015 5100 4035
rect 5050 3985 5100 4015
rect 5050 3965 5065 3985
rect 5085 3965 5100 3985
rect 5050 3950 5100 3965
rect 5200 4435 5250 4450
rect 5200 4415 5215 4435
rect 5235 4415 5250 4435
rect 5200 4385 5250 4415
rect 5200 4365 5215 4385
rect 5235 4365 5250 4385
rect 5200 4335 5250 4365
rect 5200 4315 5215 4335
rect 5235 4315 5250 4335
rect 5200 4285 5250 4315
rect 5200 4265 5215 4285
rect 5235 4265 5250 4285
rect 5200 4235 5250 4265
rect 5200 4215 5215 4235
rect 5235 4215 5250 4235
rect 5200 4185 5250 4215
rect 5200 4165 5215 4185
rect 5235 4165 5250 4185
rect 5200 4135 5250 4165
rect 5200 4115 5215 4135
rect 5235 4115 5250 4135
rect 5200 4085 5250 4115
rect 5200 4065 5215 4085
rect 5235 4065 5250 4085
rect 5200 4035 5250 4065
rect 5200 4015 5215 4035
rect 5235 4015 5250 4035
rect 5200 3985 5250 4015
rect 5200 3965 5215 3985
rect 5235 3965 5250 3985
rect 5200 3950 5250 3965
rect 5350 4435 5400 4450
rect 5350 4415 5365 4435
rect 5385 4415 5400 4435
rect 5350 4385 5400 4415
rect 5350 4365 5365 4385
rect 5385 4365 5400 4385
rect 5350 4335 5400 4365
rect 5350 4315 5365 4335
rect 5385 4315 5400 4335
rect 5350 4285 5400 4315
rect 5350 4265 5365 4285
rect 5385 4265 5400 4285
rect 5350 4235 5400 4265
rect 5350 4215 5365 4235
rect 5385 4215 5400 4235
rect 5350 4185 5400 4215
rect 5350 4165 5365 4185
rect 5385 4165 5400 4185
rect 5350 4135 5400 4165
rect 5350 4115 5365 4135
rect 5385 4115 5400 4135
rect 5350 4085 5400 4115
rect 5350 4065 5365 4085
rect 5385 4065 5400 4085
rect 5350 4035 5400 4065
rect 5350 4015 5365 4035
rect 5385 4015 5400 4035
rect 5350 3985 5400 4015
rect 5350 3965 5365 3985
rect 5385 3965 5400 3985
rect 5350 3950 5400 3965
rect 5500 4435 5550 4450
rect 5500 4415 5515 4435
rect 5535 4415 5550 4435
rect 5500 4385 5550 4415
rect 5500 4365 5515 4385
rect 5535 4365 5550 4385
rect 5500 4335 5550 4365
rect 5500 4315 5515 4335
rect 5535 4315 5550 4335
rect 5500 4285 5550 4315
rect 5500 4265 5515 4285
rect 5535 4265 5550 4285
rect 5500 4235 5550 4265
rect 5500 4215 5515 4235
rect 5535 4215 5550 4235
rect 5500 4185 5550 4215
rect 5500 4165 5515 4185
rect 5535 4165 5550 4185
rect 5500 4135 5550 4165
rect 5500 4115 5515 4135
rect 5535 4115 5550 4135
rect 5500 4085 5550 4115
rect 5500 4065 5515 4085
rect 5535 4065 5550 4085
rect 5500 4035 5550 4065
rect 5500 4015 5515 4035
rect 5535 4015 5550 4035
rect 5500 3985 5550 4015
rect 5500 3965 5515 3985
rect 5535 3965 5550 3985
rect 5500 3950 5550 3965
rect 5650 4435 5700 4450
rect 5650 4415 5665 4435
rect 5685 4415 5700 4435
rect 5650 4385 5700 4415
rect 5650 4365 5665 4385
rect 5685 4365 5700 4385
rect 5650 4335 5700 4365
rect 5650 4315 5665 4335
rect 5685 4315 5700 4335
rect 5650 4285 5700 4315
rect 5650 4265 5665 4285
rect 5685 4265 5700 4285
rect 5650 4235 5700 4265
rect 5650 4215 5665 4235
rect 5685 4215 5700 4235
rect 5650 4185 5700 4215
rect 5650 4165 5665 4185
rect 5685 4165 5700 4185
rect 5650 4135 5700 4165
rect 5650 4115 5665 4135
rect 5685 4115 5700 4135
rect 5650 4085 5700 4115
rect 5650 4065 5665 4085
rect 5685 4065 5700 4085
rect 5650 4035 5700 4065
rect 5650 4015 5665 4035
rect 5685 4015 5700 4035
rect 5650 3985 5700 4015
rect 5650 3965 5665 3985
rect 5685 3965 5700 3985
rect 5650 3950 5700 3965
rect 5800 4435 5850 4450
rect 5800 4415 5815 4435
rect 5835 4415 5850 4435
rect 5800 4385 5850 4415
rect 5800 4365 5815 4385
rect 5835 4365 5850 4385
rect 5800 4335 5850 4365
rect 5800 4315 5815 4335
rect 5835 4315 5850 4335
rect 5800 4285 5850 4315
rect 5800 4265 5815 4285
rect 5835 4265 5850 4285
rect 5800 4235 5850 4265
rect 5800 4215 5815 4235
rect 5835 4215 5850 4235
rect 5800 4185 5850 4215
rect 5800 4165 5815 4185
rect 5835 4165 5850 4185
rect 5800 4135 5850 4165
rect 5800 4115 5815 4135
rect 5835 4115 5850 4135
rect 5800 4085 5850 4115
rect 5800 4065 5815 4085
rect 5835 4065 5850 4085
rect 5800 4035 5850 4065
rect 5800 4015 5815 4035
rect 5835 4015 5850 4035
rect 5800 3985 5850 4015
rect 5800 3965 5815 3985
rect 5835 3965 5850 3985
rect 5800 3950 5850 3965
rect 5950 4435 6000 4450
rect 5950 4415 5965 4435
rect 5985 4415 6000 4435
rect 5950 4385 6000 4415
rect 5950 4365 5965 4385
rect 5985 4365 6000 4385
rect 5950 4335 6000 4365
rect 5950 4315 5965 4335
rect 5985 4315 6000 4335
rect 5950 4285 6000 4315
rect 5950 4265 5965 4285
rect 5985 4265 6000 4285
rect 5950 4235 6000 4265
rect 5950 4215 5965 4235
rect 5985 4215 6000 4235
rect 5950 4185 6000 4215
rect 5950 4165 5965 4185
rect 5985 4165 6000 4185
rect 5950 4135 6000 4165
rect 5950 4115 5965 4135
rect 5985 4115 6000 4135
rect 5950 4085 6000 4115
rect 5950 4065 5965 4085
rect 5985 4065 6000 4085
rect 5950 4035 6000 4065
rect 5950 4015 5965 4035
rect 5985 4015 6000 4035
rect 5950 3985 6000 4015
rect 5950 3965 5965 3985
rect 5985 3965 6000 3985
rect 5950 3950 6000 3965
rect 6100 4435 6150 4450
rect 6100 4415 6115 4435
rect 6135 4415 6150 4435
rect 6100 4385 6150 4415
rect 6100 4365 6115 4385
rect 6135 4365 6150 4385
rect 6100 4335 6150 4365
rect 6100 4315 6115 4335
rect 6135 4315 6150 4335
rect 6100 4285 6150 4315
rect 6100 4265 6115 4285
rect 6135 4265 6150 4285
rect 6100 4235 6150 4265
rect 6100 4215 6115 4235
rect 6135 4215 6150 4235
rect 6100 4185 6150 4215
rect 6100 4165 6115 4185
rect 6135 4165 6150 4185
rect 6100 4135 6150 4165
rect 6100 4115 6115 4135
rect 6135 4115 6150 4135
rect 6100 4085 6150 4115
rect 6100 4065 6115 4085
rect 6135 4065 6150 4085
rect 6100 4035 6150 4065
rect 6100 4015 6115 4035
rect 6135 4015 6150 4035
rect 6100 3985 6150 4015
rect 6100 3965 6115 3985
rect 6135 3965 6150 3985
rect 6100 3950 6150 3965
rect 6250 4435 6300 4450
rect 6250 4415 6265 4435
rect 6285 4415 6300 4435
rect 6250 4385 6300 4415
rect 6250 4365 6265 4385
rect 6285 4365 6300 4385
rect 6250 4335 6300 4365
rect 6250 4315 6265 4335
rect 6285 4315 6300 4335
rect 6250 4285 6300 4315
rect 6250 4265 6265 4285
rect 6285 4265 6300 4285
rect 6250 4235 6300 4265
rect 6250 4215 6265 4235
rect 6285 4215 6300 4235
rect 6250 4185 6300 4215
rect 6250 4165 6265 4185
rect 6285 4165 6300 4185
rect 6250 4135 6300 4165
rect 6250 4115 6265 4135
rect 6285 4115 6300 4135
rect 6250 4085 6300 4115
rect 6250 4065 6265 4085
rect 6285 4065 6300 4085
rect 6250 4035 6300 4065
rect 6250 4015 6265 4035
rect 6285 4015 6300 4035
rect 6250 3985 6300 4015
rect 6250 3965 6265 3985
rect 6285 3965 6300 3985
rect 6250 3950 6300 3965
rect 6400 4435 6450 4450
rect 6400 4415 6415 4435
rect 6435 4415 6450 4435
rect 6400 4385 6450 4415
rect 6400 4365 6415 4385
rect 6435 4365 6450 4385
rect 6400 4335 6450 4365
rect 6400 4315 6415 4335
rect 6435 4315 6450 4335
rect 6400 4285 6450 4315
rect 6400 4265 6415 4285
rect 6435 4265 6450 4285
rect 6400 4235 6450 4265
rect 6400 4215 6415 4235
rect 6435 4215 6450 4235
rect 6400 4185 6450 4215
rect 6400 4165 6415 4185
rect 6435 4165 6450 4185
rect 6400 4135 6450 4165
rect 6400 4115 6415 4135
rect 6435 4115 6450 4135
rect 6400 4085 6450 4115
rect 6400 4065 6415 4085
rect 6435 4065 6450 4085
rect 6400 4035 6450 4065
rect 6400 4015 6415 4035
rect 6435 4015 6450 4035
rect 6400 3985 6450 4015
rect 6400 3965 6415 3985
rect 6435 3965 6450 3985
rect 6400 3950 6450 3965
rect 6550 4435 6600 4450
rect 6550 4415 6565 4435
rect 6585 4415 6600 4435
rect 6550 4385 6600 4415
rect 6550 4365 6565 4385
rect 6585 4365 6600 4385
rect 6550 4335 6600 4365
rect 6550 4315 6565 4335
rect 6585 4315 6600 4335
rect 6550 4285 6600 4315
rect 6550 4265 6565 4285
rect 6585 4265 6600 4285
rect 6550 4235 6600 4265
rect 6550 4215 6565 4235
rect 6585 4215 6600 4235
rect 6550 4185 6600 4215
rect 6550 4165 6565 4185
rect 6585 4165 6600 4185
rect 6550 4135 6600 4165
rect 6550 4115 6565 4135
rect 6585 4115 6600 4135
rect 6550 4085 6600 4115
rect 6550 4065 6565 4085
rect 6585 4065 6600 4085
rect 6550 4035 6600 4065
rect 6550 4015 6565 4035
rect 6585 4015 6600 4035
rect 6550 3985 6600 4015
rect 6550 3965 6565 3985
rect 6585 3965 6600 3985
rect 6550 3950 6600 3965
rect 6700 4435 6750 4450
rect 6700 4415 6715 4435
rect 6735 4415 6750 4435
rect 6700 4385 6750 4415
rect 6700 4365 6715 4385
rect 6735 4365 6750 4385
rect 6700 4335 6750 4365
rect 6700 4315 6715 4335
rect 6735 4315 6750 4335
rect 6700 4285 6750 4315
rect 6700 4265 6715 4285
rect 6735 4265 6750 4285
rect 6700 4235 6750 4265
rect 6700 4215 6715 4235
rect 6735 4215 6750 4235
rect 6700 4185 6750 4215
rect 6700 4165 6715 4185
rect 6735 4165 6750 4185
rect 6700 4135 6750 4165
rect 6700 4115 6715 4135
rect 6735 4115 6750 4135
rect 6700 4085 6750 4115
rect 6700 4065 6715 4085
rect 6735 4065 6750 4085
rect 6700 4035 6750 4065
rect 6700 4015 6715 4035
rect 6735 4015 6750 4035
rect 6700 3985 6750 4015
rect 6700 3965 6715 3985
rect 6735 3965 6750 3985
rect 6700 3950 6750 3965
rect 6850 4435 6900 4450
rect 6850 4415 6865 4435
rect 6885 4415 6900 4435
rect 6850 4385 6900 4415
rect 6850 4365 6865 4385
rect 6885 4365 6900 4385
rect 6850 4335 6900 4365
rect 6850 4315 6865 4335
rect 6885 4315 6900 4335
rect 6850 4285 6900 4315
rect 6850 4265 6865 4285
rect 6885 4265 6900 4285
rect 6850 4235 6900 4265
rect 6850 4215 6865 4235
rect 6885 4215 6900 4235
rect 6850 4185 6900 4215
rect 6850 4165 6865 4185
rect 6885 4165 6900 4185
rect 6850 4135 6900 4165
rect 6850 4115 6865 4135
rect 6885 4115 6900 4135
rect 6850 4085 6900 4115
rect 6850 4065 6865 4085
rect 6885 4065 6900 4085
rect 6850 4035 6900 4065
rect 6850 4015 6865 4035
rect 6885 4015 6900 4035
rect 6850 3985 6900 4015
rect 6850 3965 6865 3985
rect 6885 3965 6900 3985
rect 6850 3950 6900 3965
rect 7000 4435 7050 4450
rect 7000 4415 7015 4435
rect 7035 4415 7050 4435
rect 7000 4385 7050 4415
rect 7000 4365 7015 4385
rect 7035 4365 7050 4385
rect 7000 4335 7050 4365
rect 7000 4315 7015 4335
rect 7035 4315 7050 4335
rect 7000 4285 7050 4315
rect 7000 4265 7015 4285
rect 7035 4265 7050 4285
rect 7000 4235 7050 4265
rect 7000 4215 7015 4235
rect 7035 4215 7050 4235
rect 7000 4185 7050 4215
rect 7000 4165 7015 4185
rect 7035 4165 7050 4185
rect 7000 4135 7050 4165
rect 7000 4115 7015 4135
rect 7035 4115 7050 4135
rect 7000 4085 7050 4115
rect 7000 4065 7015 4085
rect 7035 4065 7050 4085
rect 7000 4035 7050 4065
rect 7000 4015 7015 4035
rect 7035 4015 7050 4035
rect 7000 3985 7050 4015
rect 7000 3965 7015 3985
rect 7035 3965 7050 3985
rect 7000 3950 7050 3965
rect 7150 4435 7200 4450
rect 7150 4415 7165 4435
rect 7185 4415 7200 4435
rect 7150 4385 7200 4415
rect 7150 4365 7165 4385
rect 7185 4365 7200 4385
rect 7150 4335 7200 4365
rect 7150 4315 7165 4335
rect 7185 4315 7200 4335
rect 7150 4285 7200 4315
rect 7150 4265 7165 4285
rect 7185 4265 7200 4285
rect 7150 4235 7200 4265
rect 7150 4215 7165 4235
rect 7185 4215 7200 4235
rect 7150 4185 7200 4215
rect 7150 4165 7165 4185
rect 7185 4165 7200 4185
rect 7150 4135 7200 4165
rect 7150 4115 7165 4135
rect 7185 4115 7200 4135
rect 7150 4085 7200 4115
rect 7150 4065 7165 4085
rect 7185 4065 7200 4085
rect 7150 4035 7200 4065
rect 7150 4015 7165 4035
rect 7185 4015 7200 4035
rect 7150 3985 7200 4015
rect 7150 3965 7165 3985
rect 7185 3965 7200 3985
rect 7150 3950 7200 3965
rect 7300 4435 7350 4450
rect 7300 4415 7315 4435
rect 7335 4415 7350 4435
rect 7300 4385 7350 4415
rect 7300 4365 7315 4385
rect 7335 4365 7350 4385
rect 7300 4335 7350 4365
rect 7300 4315 7315 4335
rect 7335 4315 7350 4335
rect 7300 4285 7350 4315
rect 7300 4265 7315 4285
rect 7335 4265 7350 4285
rect 7300 4235 7350 4265
rect 7300 4215 7315 4235
rect 7335 4215 7350 4235
rect 7300 4185 7350 4215
rect 7300 4165 7315 4185
rect 7335 4165 7350 4185
rect 7300 4135 7350 4165
rect 7300 4115 7315 4135
rect 7335 4115 7350 4135
rect 7300 4085 7350 4115
rect 7300 4065 7315 4085
rect 7335 4065 7350 4085
rect 7300 4035 7350 4065
rect 7300 4015 7315 4035
rect 7335 4015 7350 4035
rect 7300 3985 7350 4015
rect 7300 3965 7315 3985
rect 7335 3965 7350 3985
rect 7300 3950 7350 3965
rect 7450 4435 7500 4450
rect 7450 4415 7465 4435
rect 7485 4415 7500 4435
rect 7450 4385 7500 4415
rect 7450 4365 7465 4385
rect 7485 4365 7500 4385
rect 7450 4335 7500 4365
rect 7450 4315 7465 4335
rect 7485 4315 7500 4335
rect 7450 4285 7500 4315
rect 7450 4265 7465 4285
rect 7485 4265 7500 4285
rect 7450 4235 7500 4265
rect 7450 4215 7465 4235
rect 7485 4215 7500 4235
rect 7450 4185 7500 4215
rect 7450 4165 7465 4185
rect 7485 4165 7500 4185
rect 7450 4135 7500 4165
rect 7450 4115 7465 4135
rect 7485 4115 7500 4135
rect 7450 4085 7500 4115
rect 7450 4065 7465 4085
rect 7485 4065 7500 4085
rect 7450 4035 7500 4065
rect 7450 4015 7465 4035
rect 7485 4015 7500 4035
rect 7450 3985 7500 4015
rect 7450 3965 7465 3985
rect 7485 3965 7500 3985
rect 7450 3950 7500 3965
rect 7600 4435 7650 4450
rect 7600 4415 7615 4435
rect 7635 4415 7650 4435
rect 7600 4385 7650 4415
rect 7600 4365 7615 4385
rect 7635 4365 7650 4385
rect 7600 4335 7650 4365
rect 7600 4315 7615 4335
rect 7635 4315 7650 4335
rect 7600 4285 7650 4315
rect 7600 4265 7615 4285
rect 7635 4265 7650 4285
rect 7600 4235 7650 4265
rect 7600 4215 7615 4235
rect 7635 4215 7650 4235
rect 7600 4185 7650 4215
rect 7600 4165 7615 4185
rect 7635 4165 7650 4185
rect 7600 4135 7650 4165
rect 7600 4115 7615 4135
rect 7635 4115 7650 4135
rect 7600 4085 7650 4115
rect 7600 4065 7615 4085
rect 7635 4065 7650 4085
rect 7600 4035 7650 4065
rect 7600 4015 7615 4035
rect 7635 4015 7650 4035
rect 7600 3985 7650 4015
rect 7600 3965 7615 3985
rect 7635 3965 7650 3985
rect 7600 3950 7650 3965
rect 7750 4435 7800 4450
rect 7750 4415 7765 4435
rect 7785 4415 7800 4435
rect 7750 4385 7800 4415
rect 7750 4365 7765 4385
rect 7785 4365 7800 4385
rect 7750 4335 7800 4365
rect 7750 4315 7765 4335
rect 7785 4315 7800 4335
rect 7750 4285 7800 4315
rect 7750 4265 7765 4285
rect 7785 4265 7800 4285
rect 7750 4235 7800 4265
rect 7750 4215 7765 4235
rect 7785 4215 7800 4235
rect 7750 4185 7800 4215
rect 7750 4165 7765 4185
rect 7785 4165 7800 4185
rect 7750 4135 7800 4165
rect 7750 4115 7765 4135
rect 7785 4115 7800 4135
rect 7750 4085 7800 4115
rect 7750 4065 7765 4085
rect 7785 4065 7800 4085
rect 7750 4035 7800 4065
rect 7750 4015 7765 4035
rect 7785 4015 7800 4035
rect 7750 3985 7800 4015
rect 7750 3965 7765 3985
rect 7785 3965 7800 3985
rect 7750 3950 7800 3965
rect 7900 3950 7950 4450
rect 8050 3950 8100 4450
rect 8200 3950 8250 4450
rect 8350 4435 8400 4450
rect 8350 4415 8365 4435
rect 8385 4415 8400 4435
rect 8350 4385 8400 4415
rect 8350 4365 8365 4385
rect 8385 4365 8400 4385
rect 8350 4335 8400 4365
rect 8350 4315 8365 4335
rect 8385 4315 8400 4335
rect 8350 4285 8400 4315
rect 8350 4265 8365 4285
rect 8385 4265 8400 4285
rect 8350 4235 8400 4265
rect 8350 4215 8365 4235
rect 8385 4215 8400 4235
rect 8350 4185 8400 4215
rect 8350 4165 8365 4185
rect 8385 4165 8400 4185
rect 8350 4135 8400 4165
rect 8350 4115 8365 4135
rect 8385 4115 8400 4135
rect 8350 4085 8400 4115
rect 8350 4065 8365 4085
rect 8385 4065 8400 4085
rect 8350 4035 8400 4065
rect 8350 4015 8365 4035
rect 8385 4015 8400 4035
rect 8350 3985 8400 4015
rect 8350 3965 8365 3985
rect 8385 3965 8400 3985
rect 8350 3950 8400 3965
rect 8500 4435 8550 4450
rect 8500 4415 8515 4435
rect 8535 4415 8550 4435
rect 8500 4385 8550 4415
rect 8500 4365 8515 4385
rect 8535 4365 8550 4385
rect 8500 4335 8550 4365
rect 8500 4315 8515 4335
rect 8535 4315 8550 4335
rect 8500 4285 8550 4315
rect 8500 4265 8515 4285
rect 8535 4265 8550 4285
rect 8500 4235 8550 4265
rect 8500 4215 8515 4235
rect 8535 4215 8550 4235
rect 8500 4185 8550 4215
rect 8500 4165 8515 4185
rect 8535 4165 8550 4185
rect 8500 4135 8550 4165
rect 8500 4115 8515 4135
rect 8535 4115 8550 4135
rect 8500 4085 8550 4115
rect 8500 4065 8515 4085
rect 8535 4065 8550 4085
rect 8500 4035 8550 4065
rect 8500 4015 8515 4035
rect 8535 4015 8550 4035
rect 8500 3985 8550 4015
rect 8500 3965 8515 3985
rect 8535 3965 8550 3985
rect 8500 3950 8550 3965
rect 8650 4435 8700 4450
rect 8650 4415 8665 4435
rect 8685 4415 8700 4435
rect 8650 4385 8700 4415
rect 8650 4365 8665 4385
rect 8685 4365 8700 4385
rect 8650 4335 8700 4365
rect 8650 4315 8665 4335
rect 8685 4315 8700 4335
rect 8650 4285 8700 4315
rect 8650 4265 8665 4285
rect 8685 4265 8700 4285
rect 8650 4235 8700 4265
rect 8650 4215 8665 4235
rect 8685 4215 8700 4235
rect 8650 4185 8700 4215
rect 8650 4165 8665 4185
rect 8685 4165 8700 4185
rect 8650 4135 8700 4165
rect 8650 4115 8665 4135
rect 8685 4115 8700 4135
rect 8650 4085 8700 4115
rect 8650 4065 8665 4085
rect 8685 4065 8700 4085
rect 8650 4035 8700 4065
rect 8650 4015 8665 4035
rect 8685 4015 8700 4035
rect 8650 3985 8700 4015
rect 8650 3965 8665 3985
rect 8685 3965 8700 3985
rect 8650 3950 8700 3965
rect 8800 4435 8850 4450
rect 8800 4415 8815 4435
rect 8835 4415 8850 4435
rect 8800 4385 8850 4415
rect 8800 4365 8815 4385
rect 8835 4365 8850 4385
rect 8800 4335 8850 4365
rect 8800 4315 8815 4335
rect 8835 4315 8850 4335
rect 8800 4285 8850 4315
rect 8800 4265 8815 4285
rect 8835 4265 8850 4285
rect 8800 4235 8850 4265
rect 8800 4215 8815 4235
rect 8835 4215 8850 4235
rect 8800 4185 8850 4215
rect 8800 4165 8815 4185
rect 8835 4165 8850 4185
rect 8800 4135 8850 4165
rect 8800 4115 8815 4135
rect 8835 4115 8850 4135
rect 8800 4085 8850 4115
rect 8800 4065 8815 4085
rect 8835 4065 8850 4085
rect 8800 4035 8850 4065
rect 8800 4015 8815 4035
rect 8835 4015 8850 4035
rect 8800 3985 8850 4015
rect 8800 3965 8815 3985
rect 8835 3965 8850 3985
rect 8800 3950 8850 3965
rect 8950 4435 9000 4450
rect 8950 4415 8965 4435
rect 8985 4415 9000 4435
rect 8950 4385 9000 4415
rect 8950 4365 8965 4385
rect 8985 4365 9000 4385
rect 8950 4335 9000 4365
rect 8950 4315 8965 4335
rect 8985 4315 9000 4335
rect 8950 4285 9000 4315
rect 8950 4265 8965 4285
rect 8985 4265 9000 4285
rect 8950 4235 9000 4265
rect 8950 4215 8965 4235
rect 8985 4215 9000 4235
rect 8950 4185 9000 4215
rect 8950 4165 8965 4185
rect 8985 4165 9000 4185
rect 8950 4135 9000 4165
rect 8950 4115 8965 4135
rect 8985 4115 9000 4135
rect 8950 4085 9000 4115
rect 8950 4065 8965 4085
rect 8985 4065 9000 4085
rect 8950 4035 9000 4065
rect 8950 4015 8965 4035
rect 8985 4015 9000 4035
rect 8950 3985 9000 4015
rect 8950 3965 8965 3985
rect 8985 3965 9000 3985
rect 8950 3950 9000 3965
rect 9100 4435 9150 4450
rect 9100 4415 9115 4435
rect 9135 4415 9150 4435
rect 9100 4385 9150 4415
rect 9100 4365 9115 4385
rect 9135 4365 9150 4385
rect 9100 4335 9150 4365
rect 9100 4315 9115 4335
rect 9135 4315 9150 4335
rect 9100 4285 9150 4315
rect 9100 4265 9115 4285
rect 9135 4265 9150 4285
rect 9100 4235 9150 4265
rect 9100 4215 9115 4235
rect 9135 4215 9150 4235
rect 9100 4185 9150 4215
rect 9100 4165 9115 4185
rect 9135 4165 9150 4185
rect 9100 4135 9150 4165
rect 9100 4115 9115 4135
rect 9135 4115 9150 4135
rect 9100 4085 9150 4115
rect 9100 4065 9115 4085
rect 9135 4065 9150 4085
rect 9100 4035 9150 4065
rect 9100 4015 9115 4035
rect 9135 4015 9150 4035
rect 9100 3985 9150 4015
rect 9100 3965 9115 3985
rect 9135 3965 9150 3985
rect 9100 3950 9150 3965
rect 9250 4435 9300 4450
rect 9250 4415 9265 4435
rect 9285 4415 9300 4435
rect 9250 4385 9300 4415
rect 9250 4365 9265 4385
rect 9285 4365 9300 4385
rect 9250 4335 9300 4365
rect 9250 4315 9265 4335
rect 9285 4315 9300 4335
rect 9250 4285 9300 4315
rect 9250 4265 9265 4285
rect 9285 4265 9300 4285
rect 9250 4235 9300 4265
rect 9250 4215 9265 4235
rect 9285 4215 9300 4235
rect 9250 4185 9300 4215
rect 9250 4165 9265 4185
rect 9285 4165 9300 4185
rect 9250 4135 9300 4165
rect 9250 4115 9265 4135
rect 9285 4115 9300 4135
rect 9250 4085 9300 4115
rect 9250 4065 9265 4085
rect 9285 4065 9300 4085
rect 9250 4035 9300 4065
rect 9250 4015 9265 4035
rect 9285 4015 9300 4035
rect 9250 3985 9300 4015
rect 9250 3965 9265 3985
rect 9285 3965 9300 3985
rect 9250 3950 9300 3965
rect 9400 4435 9450 4450
rect 9400 4415 9415 4435
rect 9435 4415 9450 4435
rect 9400 4385 9450 4415
rect 9400 4365 9415 4385
rect 9435 4365 9450 4385
rect 9400 4335 9450 4365
rect 9400 4315 9415 4335
rect 9435 4315 9450 4335
rect 9400 4285 9450 4315
rect 9400 4265 9415 4285
rect 9435 4265 9450 4285
rect 9400 4235 9450 4265
rect 9400 4215 9415 4235
rect 9435 4215 9450 4235
rect 9400 4185 9450 4215
rect 9400 4165 9415 4185
rect 9435 4165 9450 4185
rect 9400 4135 9450 4165
rect 9400 4115 9415 4135
rect 9435 4115 9450 4135
rect 9400 4085 9450 4115
rect 9400 4065 9415 4085
rect 9435 4065 9450 4085
rect 9400 4035 9450 4065
rect 9400 4015 9415 4035
rect 9435 4015 9450 4035
rect 9400 3985 9450 4015
rect 9400 3965 9415 3985
rect 9435 3965 9450 3985
rect 9400 3950 9450 3965
rect 9550 4435 9600 4450
rect 9550 4415 9565 4435
rect 9585 4415 9600 4435
rect 9550 4385 9600 4415
rect 9550 4365 9565 4385
rect 9585 4365 9600 4385
rect 9550 4335 9600 4365
rect 9550 4315 9565 4335
rect 9585 4315 9600 4335
rect 9550 4285 9600 4315
rect 9550 4265 9565 4285
rect 9585 4265 9600 4285
rect 9550 4235 9600 4265
rect 9550 4215 9565 4235
rect 9585 4215 9600 4235
rect 9550 4185 9600 4215
rect 9550 4165 9565 4185
rect 9585 4165 9600 4185
rect 9550 4135 9600 4165
rect 9550 4115 9565 4135
rect 9585 4115 9600 4135
rect 9550 4085 9600 4115
rect 9550 4065 9565 4085
rect 9585 4065 9600 4085
rect 9550 4035 9600 4065
rect 9550 4015 9565 4035
rect 9585 4015 9600 4035
rect 9550 3985 9600 4015
rect 9550 3965 9565 3985
rect 9585 3965 9600 3985
rect 9550 3950 9600 3965
rect 9700 4435 9750 4450
rect 9700 4415 9715 4435
rect 9735 4415 9750 4435
rect 9700 4385 9750 4415
rect 9700 4365 9715 4385
rect 9735 4365 9750 4385
rect 9700 4335 9750 4365
rect 9700 4315 9715 4335
rect 9735 4315 9750 4335
rect 9700 4285 9750 4315
rect 9700 4265 9715 4285
rect 9735 4265 9750 4285
rect 9700 4235 9750 4265
rect 9700 4215 9715 4235
rect 9735 4215 9750 4235
rect 9700 4185 9750 4215
rect 9700 4165 9715 4185
rect 9735 4165 9750 4185
rect 9700 4135 9750 4165
rect 9700 4115 9715 4135
rect 9735 4115 9750 4135
rect 9700 4085 9750 4115
rect 9700 4065 9715 4085
rect 9735 4065 9750 4085
rect 9700 4035 9750 4065
rect 9700 4015 9715 4035
rect 9735 4015 9750 4035
rect 9700 3985 9750 4015
rect 9700 3965 9715 3985
rect 9735 3965 9750 3985
rect 9700 3950 9750 3965
rect 9850 4435 9900 4450
rect 9850 4415 9865 4435
rect 9885 4415 9900 4435
rect 9850 4385 9900 4415
rect 9850 4365 9865 4385
rect 9885 4365 9900 4385
rect 9850 4335 9900 4365
rect 9850 4315 9865 4335
rect 9885 4315 9900 4335
rect 9850 4285 9900 4315
rect 9850 4265 9865 4285
rect 9885 4265 9900 4285
rect 9850 4235 9900 4265
rect 9850 4215 9865 4235
rect 9885 4215 9900 4235
rect 9850 4185 9900 4215
rect 9850 4165 9865 4185
rect 9885 4165 9900 4185
rect 9850 4135 9900 4165
rect 9850 4115 9865 4135
rect 9885 4115 9900 4135
rect 9850 4085 9900 4115
rect 9850 4065 9865 4085
rect 9885 4065 9900 4085
rect 9850 4035 9900 4065
rect 9850 4015 9865 4035
rect 9885 4015 9900 4035
rect 9850 3985 9900 4015
rect 9850 3965 9865 3985
rect 9885 3965 9900 3985
rect 9850 3950 9900 3965
rect 10000 4435 10050 4450
rect 10000 4415 10015 4435
rect 10035 4415 10050 4435
rect 10000 4385 10050 4415
rect 10000 4365 10015 4385
rect 10035 4365 10050 4385
rect 10000 4335 10050 4365
rect 10000 4315 10015 4335
rect 10035 4315 10050 4335
rect 10000 4285 10050 4315
rect 10000 4265 10015 4285
rect 10035 4265 10050 4285
rect 10000 4235 10050 4265
rect 10000 4215 10015 4235
rect 10035 4215 10050 4235
rect 10000 4185 10050 4215
rect 10000 4165 10015 4185
rect 10035 4165 10050 4185
rect 10000 4135 10050 4165
rect 10000 4115 10015 4135
rect 10035 4115 10050 4135
rect 10000 4085 10050 4115
rect 10000 4065 10015 4085
rect 10035 4065 10050 4085
rect 10000 4035 10050 4065
rect 10000 4015 10015 4035
rect 10035 4015 10050 4035
rect 10000 3985 10050 4015
rect 10000 3965 10015 3985
rect 10035 3965 10050 3985
rect 10000 3950 10050 3965
rect 10150 4435 10200 4450
rect 10150 4415 10165 4435
rect 10185 4415 10200 4435
rect 10150 4385 10200 4415
rect 10150 4365 10165 4385
rect 10185 4365 10200 4385
rect 10150 4335 10200 4365
rect 10150 4315 10165 4335
rect 10185 4315 10200 4335
rect 10150 4285 10200 4315
rect 10150 4265 10165 4285
rect 10185 4265 10200 4285
rect 10150 4235 10200 4265
rect 10150 4215 10165 4235
rect 10185 4215 10200 4235
rect 10150 4185 10200 4215
rect 10150 4165 10165 4185
rect 10185 4165 10200 4185
rect 10150 4135 10200 4165
rect 10150 4115 10165 4135
rect 10185 4115 10200 4135
rect 10150 4085 10200 4115
rect 10150 4065 10165 4085
rect 10185 4065 10200 4085
rect 10150 4035 10200 4065
rect 10150 4015 10165 4035
rect 10185 4015 10200 4035
rect 10150 3985 10200 4015
rect 10150 3965 10165 3985
rect 10185 3965 10200 3985
rect 10150 3950 10200 3965
rect 10300 4435 10350 4450
rect 10300 4415 10315 4435
rect 10335 4415 10350 4435
rect 10300 4385 10350 4415
rect 10300 4365 10315 4385
rect 10335 4365 10350 4385
rect 10300 4335 10350 4365
rect 10300 4315 10315 4335
rect 10335 4315 10350 4335
rect 10300 4285 10350 4315
rect 10300 4265 10315 4285
rect 10335 4265 10350 4285
rect 10300 4235 10350 4265
rect 10300 4215 10315 4235
rect 10335 4215 10350 4235
rect 10300 4185 10350 4215
rect 10300 4165 10315 4185
rect 10335 4165 10350 4185
rect 10300 4135 10350 4165
rect 10300 4115 10315 4135
rect 10335 4115 10350 4135
rect 10300 4085 10350 4115
rect 10300 4065 10315 4085
rect 10335 4065 10350 4085
rect 10300 4035 10350 4065
rect 10300 4015 10315 4035
rect 10335 4015 10350 4035
rect 10300 3985 10350 4015
rect 10300 3965 10315 3985
rect 10335 3965 10350 3985
rect 10300 3950 10350 3965
rect 10450 4435 10500 4450
rect 10450 4415 10465 4435
rect 10485 4415 10500 4435
rect 10450 4385 10500 4415
rect 10450 4365 10465 4385
rect 10485 4365 10500 4385
rect 10450 4335 10500 4365
rect 10450 4315 10465 4335
rect 10485 4315 10500 4335
rect 10450 4285 10500 4315
rect 10450 4265 10465 4285
rect 10485 4265 10500 4285
rect 10450 4235 10500 4265
rect 10450 4215 10465 4235
rect 10485 4215 10500 4235
rect 10450 4185 10500 4215
rect 10450 4165 10465 4185
rect 10485 4165 10500 4185
rect 10450 4135 10500 4165
rect 10450 4115 10465 4135
rect 10485 4115 10500 4135
rect 10450 4085 10500 4115
rect 10450 4065 10465 4085
rect 10485 4065 10500 4085
rect 10450 4035 10500 4065
rect 10450 4015 10465 4035
rect 10485 4015 10500 4035
rect 10450 3985 10500 4015
rect 10450 3965 10465 3985
rect 10485 3965 10500 3985
rect 10450 3950 10500 3965
rect 10600 4435 10650 4450
rect 10600 4415 10615 4435
rect 10635 4415 10650 4435
rect 10600 4385 10650 4415
rect 10600 4365 10615 4385
rect 10635 4365 10650 4385
rect 10600 4335 10650 4365
rect 10600 4315 10615 4335
rect 10635 4315 10650 4335
rect 10600 4285 10650 4315
rect 10600 4265 10615 4285
rect 10635 4265 10650 4285
rect 10600 4235 10650 4265
rect 10600 4215 10615 4235
rect 10635 4215 10650 4235
rect 10600 4185 10650 4215
rect 10600 4165 10615 4185
rect 10635 4165 10650 4185
rect 10600 4135 10650 4165
rect 10600 4115 10615 4135
rect 10635 4115 10650 4135
rect 10600 4085 10650 4115
rect 10600 4065 10615 4085
rect 10635 4065 10650 4085
rect 10600 4035 10650 4065
rect 10600 4015 10615 4035
rect 10635 4015 10650 4035
rect 10600 3985 10650 4015
rect 10600 3965 10615 3985
rect 10635 3965 10650 3985
rect 10600 3950 10650 3965
rect 10750 4435 10800 4450
rect 10750 4415 10765 4435
rect 10785 4415 10800 4435
rect 10750 4385 10800 4415
rect 10750 4365 10765 4385
rect 10785 4365 10800 4385
rect 10750 4335 10800 4365
rect 10750 4315 10765 4335
rect 10785 4315 10800 4335
rect 10750 4285 10800 4315
rect 10750 4265 10765 4285
rect 10785 4265 10800 4285
rect 10750 4235 10800 4265
rect 10750 4215 10765 4235
rect 10785 4215 10800 4235
rect 10750 4185 10800 4215
rect 10750 4165 10765 4185
rect 10785 4165 10800 4185
rect 10750 4135 10800 4165
rect 10750 4115 10765 4135
rect 10785 4115 10800 4135
rect 10750 4085 10800 4115
rect 10750 4065 10765 4085
rect 10785 4065 10800 4085
rect 10750 4035 10800 4065
rect 10750 4015 10765 4035
rect 10785 4015 10800 4035
rect 10750 3985 10800 4015
rect 10750 3965 10765 3985
rect 10785 3965 10800 3985
rect 10750 3950 10800 3965
rect 10900 3950 10950 4450
rect 11050 3950 11100 4450
rect 11200 3950 11250 4450
rect 11350 4435 11400 4450
rect 11350 4415 11365 4435
rect 11385 4415 11400 4435
rect 11350 4385 11400 4415
rect 11350 4365 11365 4385
rect 11385 4365 11400 4385
rect 11350 4335 11400 4365
rect 11350 4315 11365 4335
rect 11385 4315 11400 4335
rect 11350 4285 11400 4315
rect 11350 4265 11365 4285
rect 11385 4265 11400 4285
rect 11350 4235 11400 4265
rect 11350 4215 11365 4235
rect 11385 4215 11400 4235
rect 11350 4185 11400 4215
rect 11350 4165 11365 4185
rect 11385 4165 11400 4185
rect 11350 4135 11400 4165
rect 11350 4115 11365 4135
rect 11385 4115 11400 4135
rect 11350 4085 11400 4115
rect 11350 4065 11365 4085
rect 11385 4065 11400 4085
rect 11350 4035 11400 4065
rect 11350 4015 11365 4035
rect 11385 4015 11400 4035
rect 11350 3985 11400 4015
rect 11350 3965 11365 3985
rect 11385 3965 11400 3985
rect 11350 3950 11400 3965
rect 11500 3950 11550 4450
rect 11650 3950 11700 4450
rect 11800 3950 11850 4450
rect 11950 4435 12000 4450
rect 11950 4415 11965 4435
rect 11985 4415 12000 4435
rect 11950 4385 12000 4415
rect 11950 4365 11965 4385
rect 11985 4365 12000 4385
rect 11950 4335 12000 4365
rect 11950 4315 11965 4335
rect 11985 4315 12000 4335
rect 11950 4285 12000 4315
rect 11950 4265 11965 4285
rect 11985 4265 12000 4285
rect 11950 4235 12000 4265
rect 11950 4215 11965 4235
rect 11985 4215 12000 4235
rect 11950 4185 12000 4215
rect 11950 4165 11965 4185
rect 11985 4165 12000 4185
rect 11950 4135 12000 4165
rect 11950 4115 11965 4135
rect 11985 4115 12000 4135
rect 11950 4085 12000 4115
rect 11950 4065 11965 4085
rect 11985 4065 12000 4085
rect 11950 4035 12000 4065
rect 11950 4015 11965 4035
rect 11985 4015 12000 4035
rect 11950 3985 12000 4015
rect 11950 3965 11965 3985
rect 11985 3965 12000 3985
rect 11950 3950 12000 3965
rect 12100 3950 12150 4450
rect 12250 3950 12300 4450
rect 12400 3950 12450 4450
rect 12550 4435 12600 4450
rect 12550 4415 12565 4435
rect 12585 4415 12600 4435
rect 12550 4385 12600 4415
rect 12550 4365 12565 4385
rect 12585 4365 12600 4385
rect 12550 4335 12600 4365
rect 12550 4315 12565 4335
rect 12585 4315 12600 4335
rect 12550 4285 12600 4315
rect 12550 4265 12565 4285
rect 12585 4265 12600 4285
rect 12550 4235 12600 4265
rect 12550 4215 12565 4235
rect 12585 4215 12600 4235
rect 12550 4185 12600 4215
rect 12550 4165 12565 4185
rect 12585 4165 12600 4185
rect 12550 4135 12600 4165
rect 12550 4115 12565 4135
rect 12585 4115 12600 4135
rect 12550 4085 12600 4115
rect 12550 4065 12565 4085
rect 12585 4065 12600 4085
rect 12550 4035 12600 4065
rect 12550 4015 12565 4035
rect 12585 4015 12600 4035
rect 12550 3985 12600 4015
rect 12550 3965 12565 3985
rect 12585 3965 12600 3985
rect 12550 3950 12600 3965
rect 12700 3950 12750 4450
rect 12850 3950 12900 4450
rect 13000 3950 13050 4450
rect 13150 4435 13200 4450
rect 13150 4415 13165 4435
rect 13185 4415 13200 4435
rect 13150 4385 13200 4415
rect 13150 4365 13165 4385
rect 13185 4365 13200 4385
rect 13150 4335 13200 4365
rect 13150 4315 13165 4335
rect 13185 4315 13200 4335
rect 13150 4285 13200 4315
rect 13150 4265 13165 4285
rect 13185 4265 13200 4285
rect 13150 4235 13200 4265
rect 13150 4215 13165 4235
rect 13185 4215 13200 4235
rect 13150 4185 13200 4215
rect 13150 4165 13165 4185
rect 13185 4165 13200 4185
rect 13150 4135 13200 4165
rect 13150 4115 13165 4135
rect 13185 4115 13200 4135
rect 13150 4085 13200 4115
rect 13150 4065 13165 4085
rect 13185 4065 13200 4085
rect 13150 4035 13200 4065
rect 13150 4015 13165 4035
rect 13185 4015 13200 4035
rect 13150 3985 13200 4015
rect 13150 3965 13165 3985
rect 13185 3965 13200 3985
rect 13150 3950 13200 3965
rect 13300 3950 13350 4450
rect 13450 3950 13500 4450
rect 13600 3950 13650 4450
rect 13750 4435 13800 4450
rect 13750 4415 13765 4435
rect 13785 4415 13800 4435
rect 13750 4385 13800 4415
rect 13750 4365 13765 4385
rect 13785 4365 13800 4385
rect 13750 4335 13800 4365
rect 13750 4315 13765 4335
rect 13785 4315 13800 4335
rect 13750 4285 13800 4315
rect 13750 4265 13765 4285
rect 13785 4265 13800 4285
rect 13750 4235 13800 4265
rect 13750 4215 13765 4235
rect 13785 4215 13800 4235
rect 13750 4185 13800 4215
rect 13750 4165 13765 4185
rect 13785 4165 13800 4185
rect 13750 4135 13800 4165
rect 13750 4115 13765 4135
rect 13785 4115 13800 4135
rect 13750 4085 13800 4115
rect 13750 4065 13765 4085
rect 13785 4065 13800 4085
rect 13750 4035 13800 4065
rect 13750 4015 13765 4035
rect 13785 4015 13800 4035
rect 13750 3985 13800 4015
rect 13750 3965 13765 3985
rect 13785 3965 13800 3985
rect 13750 3950 13800 3965
rect 13900 3950 13950 4450
rect 14050 3950 14100 4450
rect 14200 3950 14250 4450
rect 14350 4435 14400 4450
rect 14350 4415 14365 4435
rect 14385 4415 14400 4435
rect 14350 4385 14400 4415
rect 14350 4365 14365 4385
rect 14385 4365 14400 4385
rect 14350 4335 14400 4365
rect 14350 4315 14365 4335
rect 14385 4315 14400 4335
rect 14350 4285 14400 4315
rect 14350 4265 14365 4285
rect 14385 4265 14400 4285
rect 14350 4235 14400 4265
rect 14350 4215 14365 4235
rect 14385 4215 14400 4235
rect 14350 4185 14400 4215
rect 14350 4165 14365 4185
rect 14385 4165 14400 4185
rect 14350 4135 14400 4165
rect 14350 4115 14365 4135
rect 14385 4115 14400 4135
rect 14350 4085 14400 4115
rect 14350 4065 14365 4085
rect 14385 4065 14400 4085
rect 14350 4035 14400 4065
rect 14350 4015 14365 4035
rect 14385 4015 14400 4035
rect 14350 3985 14400 4015
rect 14350 3965 14365 3985
rect 14385 3965 14400 3985
rect 14350 3950 14400 3965
rect 14500 3950 14550 4450
rect 14650 3950 14700 4450
rect 14800 3950 14850 4450
rect 14950 4435 15000 4450
rect 14950 4415 14965 4435
rect 14985 4415 15000 4435
rect 14950 4385 15000 4415
rect 14950 4365 14965 4385
rect 14985 4365 15000 4385
rect 14950 4335 15000 4365
rect 14950 4315 14965 4335
rect 14985 4315 15000 4335
rect 14950 4285 15000 4315
rect 14950 4265 14965 4285
rect 14985 4265 15000 4285
rect 14950 4235 15000 4265
rect 14950 4215 14965 4235
rect 14985 4215 15000 4235
rect 14950 4185 15000 4215
rect 14950 4165 14965 4185
rect 14985 4165 15000 4185
rect 14950 4135 15000 4165
rect 14950 4115 14965 4135
rect 14985 4115 15000 4135
rect 14950 4085 15000 4115
rect 14950 4065 14965 4085
rect 14985 4065 15000 4085
rect 14950 4035 15000 4065
rect 14950 4015 14965 4035
rect 14985 4015 15000 4035
rect 14950 3985 15000 4015
rect 14950 3965 14965 3985
rect 14985 3965 15000 3985
rect 14950 3950 15000 3965
rect 15100 3950 15150 4450
rect 15250 3950 15300 4450
rect 15400 3950 15450 4450
rect 15550 4435 15600 4450
rect 15550 4415 15565 4435
rect 15585 4415 15600 4435
rect 15550 4385 15600 4415
rect 15550 4365 15565 4385
rect 15585 4365 15600 4385
rect 15550 4335 15600 4365
rect 15550 4315 15565 4335
rect 15585 4315 15600 4335
rect 15550 4285 15600 4315
rect 15550 4265 15565 4285
rect 15585 4265 15600 4285
rect 15550 4235 15600 4265
rect 15550 4215 15565 4235
rect 15585 4215 15600 4235
rect 15550 4185 15600 4215
rect 15550 4165 15565 4185
rect 15585 4165 15600 4185
rect 15550 4135 15600 4165
rect 15550 4115 15565 4135
rect 15585 4115 15600 4135
rect 15550 4085 15600 4115
rect 15550 4065 15565 4085
rect 15585 4065 15600 4085
rect 15550 4035 15600 4065
rect 15550 4015 15565 4035
rect 15585 4015 15600 4035
rect 15550 3985 15600 4015
rect 15550 3965 15565 3985
rect 15585 3965 15600 3985
rect 15550 3950 15600 3965
rect 15700 3950 15750 4450
rect 15850 3950 15900 4450
rect 16000 3950 16050 4450
rect 16150 4435 16200 4450
rect 16150 4415 16165 4435
rect 16185 4415 16200 4435
rect 16150 4385 16200 4415
rect 16150 4365 16165 4385
rect 16185 4365 16200 4385
rect 16150 4335 16200 4365
rect 16150 4315 16165 4335
rect 16185 4315 16200 4335
rect 16150 4285 16200 4315
rect 16150 4265 16165 4285
rect 16185 4265 16200 4285
rect 16150 4235 16200 4265
rect 16150 4215 16165 4235
rect 16185 4215 16200 4235
rect 16150 4185 16200 4215
rect 16150 4165 16165 4185
rect 16185 4165 16200 4185
rect 16150 4135 16200 4165
rect 16150 4115 16165 4135
rect 16185 4115 16200 4135
rect 16150 4085 16200 4115
rect 16150 4065 16165 4085
rect 16185 4065 16200 4085
rect 16150 4035 16200 4065
rect 16150 4015 16165 4035
rect 16185 4015 16200 4035
rect 16150 3985 16200 4015
rect 16150 3965 16165 3985
rect 16185 3965 16200 3985
rect 16150 3950 16200 3965
rect 16300 4435 16350 4450
rect 16300 4415 16315 4435
rect 16335 4415 16350 4435
rect 16300 4385 16350 4415
rect 16300 4365 16315 4385
rect 16335 4365 16350 4385
rect 16300 4335 16350 4365
rect 16300 4315 16315 4335
rect 16335 4315 16350 4335
rect 16300 4285 16350 4315
rect 16300 4265 16315 4285
rect 16335 4265 16350 4285
rect 16300 4235 16350 4265
rect 16300 4215 16315 4235
rect 16335 4215 16350 4235
rect 16300 4185 16350 4215
rect 16300 4165 16315 4185
rect 16335 4165 16350 4185
rect 16300 4135 16350 4165
rect 16300 4115 16315 4135
rect 16335 4115 16350 4135
rect 16300 4085 16350 4115
rect 16300 4065 16315 4085
rect 16335 4065 16350 4085
rect 16300 4035 16350 4065
rect 16300 4015 16315 4035
rect 16335 4015 16350 4035
rect 16300 3985 16350 4015
rect 16300 3965 16315 3985
rect 16335 3965 16350 3985
rect 16300 3950 16350 3965
rect 16450 4435 16500 4450
rect 16450 4415 16465 4435
rect 16485 4415 16500 4435
rect 16450 4385 16500 4415
rect 16450 4365 16465 4385
rect 16485 4365 16500 4385
rect 16450 4335 16500 4365
rect 16450 4315 16465 4335
rect 16485 4315 16500 4335
rect 16450 4285 16500 4315
rect 16450 4265 16465 4285
rect 16485 4265 16500 4285
rect 16450 4235 16500 4265
rect 16450 4215 16465 4235
rect 16485 4215 16500 4235
rect 16450 4185 16500 4215
rect 16450 4165 16465 4185
rect 16485 4165 16500 4185
rect 16450 4135 16500 4165
rect 16450 4115 16465 4135
rect 16485 4115 16500 4135
rect 16450 4085 16500 4115
rect 16450 4065 16465 4085
rect 16485 4065 16500 4085
rect 16450 4035 16500 4065
rect 16450 4015 16465 4035
rect 16485 4015 16500 4035
rect 16450 3985 16500 4015
rect 16450 3965 16465 3985
rect 16485 3965 16500 3985
rect 16450 3950 16500 3965
rect 16600 4435 16650 4450
rect 16600 4415 16615 4435
rect 16635 4415 16650 4435
rect 16600 4385 16650 4415
rect 16600 4365 16615 4385
rect 16635 4365 16650 4385
rect 16600 4335 16650 4365
rect 16600 4315 16615 4335
rect 16635 4315 16650 4335
rect 16600 4285 16650 4315
rect 16600 4265 16615 4285
rect 16635 4265 16650 4285
rect 16600 4235 16650 4265
rect 16600 4215 16615 4235
rect 16635 4215 16650 4235
rect 16600 4185 16650 4215
rect 16600 4165 16615 4185
rect 16635 4165 16650 4185
rect 16600 4135 16650 4165
rect 16600 4115 16615 4135
rect 16635 4115 16650 4135
rect 16600 4085 16650 4115
rect 16600 4065 16615 4085
rect 16635 4065 16650 4085
rect 16600 4035 16650 4065
rect 16600 4015 16615 4035
rect 16635 4015 16650 4035
rect 16600 3985 16650 4015
rect 16600 3965 16615 3985
rect 16635 3965 16650 3985
rect 16600 3950 16650 3965
rect 16750 4435 16800 4450
rect 16750 4415 16765 4435
rect 16785 4415 16800 4435
rect 16750 4385 16800 4415
rect 16750 4365 16765 4385
rect 16785 4365 16800 4385
rect 16750 4335 16800 4365
rect 16750 4315 16765 4335
rect 16785 4315 16800 4335
rect 16750 4285 16800 4315
rect 16750 4265 16765 4285
rect 16785 4265 16800 4285
rect 16750 4235 16800 4265
rect 16750 4215 16765 4235
rect 16785 4215 16800 4235
rect 16750 4185 16800 4215
rect 16750 4165 16765 4185
rect 16785 4165 16800 4185
rect 16750 4135 16800 4165
rect 16750 4115 16765 4135
rect 16785 4115 16800 4135
rect 16750 4085 16800 4115
rect 16750 4065 16765 4085
rect 16785 4065 16800 4085
rect 16750 4035 16800 4065
rect 16750 4015 16765 4035
rect 16785 4015 16800 4035
rect 16750 3985 16800 4015
rect 16750 3965 16765 3985
rect 16785 3965 16800 3985
rect 16750 3950 16800 3965
rect 16900 4435 16950 4450
rect 16900 4415 16915 4435
rect 16935 4415 16950 4435
rect 16900 4385 16950 4415
rect 16900 4365 16915 4385
rect 16935 4365 16950 4385
rect 16900 4335 16950 4365
rect 16900 4315 16915 4335
rect 16935 4315 16950 4335
rect 16900 4285 16950 4315
rect 16900 4265 16915 4285
rect 16935 4265 16950 4285
rect 16900 4235 16950 4265
rect 16900 4215 16915 4235
rect 16935 4215 16950 4235
rect 16900 4185 16950 4215
rect 16900 4165 16915 4185
rect 16935 4165 16950 4185
rect 16900 4135 16950 4165
rect 16900 4115 16915 4135
rect 16935 4115 16950 4135
rect 16900 4085 16950 4115
rect 16900 4065 16915 4085
rect 16935 4065 16950 4085
rect 16900 4035 16950 4065
rect 16900 4015 16915 4035
rect 16935 4015 16950 4035
rect 16900 3985 16950 4015
rect 16900 3965 16915 3985
rect 16935 3965 16950 3985
rect 16900 3950 16950 3965
rect 17050 4435 17100 4450
rect 17050 4415 17065 4435
rect 17085 4415 17100 4435
rect 17050 4385 17100 4415
rect 17050 4365 17065 4385
rect 17085 4365 17100 4385
rect 17050 4335 17100 4365
rect 17050 4315 17065 4335
rect 17085 4315 17100 4335
rect 17050 4285 17100 4315
rect 17050 4265 17065 4285
rect 17085 4265 17100 4285
rect 17050 4235 17100 4265
rect 17050 4215 17065 4235
rect 17085 4215 17100 4235
rect 17050 4185 17100 4215
rect 17050 4165 17065 4185
rect 17085 4165 17100 4185
rect 17050 4135 17100 4165
rect 17050 4115 17065 4135
rect 17085 4115 17100 4135
rect 17050 4085 17100 4115
rect 17050 4065 17065 4085
rect 17085 4065 17100 4085
rect 17050 4035 17100 4065
rect 17050 4015 17065 4035
rect 17085 4015 17100 4035
rect 17050 3985 17100 4015
rect 17050 3965 17065 3985
rect 17085 3965 17100 3985
rect 17050 3950 17100 3965
rect 17200 4435 17250 4450
rect 17200 4415 17215 4435
rect 17235 4415 17250 4435
rect 17200 4385 17250 4415
rect 17200 4365 17215 4385
rect 17235 4365 17250 4385
rect 17200 4335 17250 4365
rect 17200 4315 17215 4335
rect 17235 4315 17250 4335
rect 17200 4285 17250 4315
rect 17200 4265 17215 4285
rect 17235 4265 17250 4285
rect 17200 4235 17250 4265
rect 17200 4215 17215 4235
rect 17235 4215 17250 4235
rect 17200 4185 17250 4215
rect 17200 4165 17215 4185
rect 17235 4165 17250 4185
rect 17200 4135 17250 4165
rect 17200 4115 17215 4135
rect 17235 4115 17250 4135
rect 17200 4085 17250 4115
rect 17200 4065 17215 4085
rect 17235 4065 17250 4085
rect 17200 4035 17250 4065
rect 17200 4015 17215 4035
rect 17235 4015 17250 4035
rect 17200 3985 17250 4015
rect 17200 3965 17215 3985
rect 17235 3965 17250 3985
rect 17200 3950 17250 3965
rect 17350 4435 17400 4450
rect 17350 4415 17365 4435
rect 17385 4415 17400 4435
rect 17350 4385 17400 4415
rect 17350 4365 17365 4385
rect 17385 4365 17400 4385
rect 17350 4335 17400 4365
rect 17350 4315 17365 4335
rect 17385 4315 17400 4335
rect 17350 4285 17400 4315
rect 17350 4265 17365 4285
rect 17385 4265 17400 4285
rect 17350 4235 17400 4265
rect 17350 4215 17365 4235
rect 17385 4215 17400 4235
rect 17350 4185 17400 4215
rect 17350 4165 17365 4185
rect 17385 4165 17400 4185
rect 17350 4135 17400 4165
rect 17350 4115 17365 4135
rect 17385 4115 17400 4135
rect 17350 4085 17400 4115
rect 17350 4065 17365 4085
rect 17385 4065 17400 4085
rect 17350 4035 17400 4065
rect 17350 4015 17365 4035
rect 17385 4015 17400 4035
rect 17350 3985 17400 4015
rect 17350 3965 17365 3985
rect 17385 3965 17400 3985
rect 17350 3950 17400 3965
rect 17500 3950 17550 4450
rect 17650 3950 17700 4450
rect 17800 3950 17850 4450
rect 17950 4435 18000 4450
rect 17950 4415 17965 4435
rect 17985 4415 18000 4435
rect 17950 4385 18000 4415
rect 17950 4365 17965 4385
rect 17985 4365 18000 4385
rect 17950 4335 18000 4365
rect 17950 4315 17965 4335
rect 17985 4315 18000 4335
rect 17950 4285 18000 4315
rect 17950 4265 17965 4285
rect 17985 4265 18000 4285
rect 17950 4235 18000 4265
rect 17950 4215 17965 4235
rect 17985 4215 18000 4235
rect 17950 4185 18000 4215
rect 17950 4165 17965 4185
rect 17985 4165 18000 4185
rect 17950 4135 18000 4165
rect 17950 4115 17965 4135
rect 17985 4115 18000 4135
rect 17950 4085 18000 4115
rect 17950 4065 17965 4085
rect 17985 4065 18000 4085
rect 17950 4035 18000 4065
rect 17950 4015 17965 4035
rect 17985 4015 18000 4035
rect 17950 3985 18000 4015
rect 17950 3965 17965 3985
rect 17985 3965 18000 3985
rect 17950 3950 18000 3965
rect 18100 3950 18150 4450
rect 18250 3950 18300 4450
rect 18400 3950 18450 4450
rect 18550 4435 18600 4450
rect 18550 4415 18565 4435
rect 18585 4415 18600 4435
rect 18550 4385 18600 4415
rect 18550 4365 18565 4385
rect 18585 4365 18600 4385
rect 18550 4335 18600 4365
rect 18550 4315 18565 4335
rect 18585 4315 18600 4335
rect 18550 4285 18600 4315
rect 18550 4265 18565 4285
rect 18585 4265 18600 4285
rect 18550 4235 18600 4265
rect 18550 4215 18565 4235
rect 18585 4215 18600 4235
rect 18550 4185 18600 4215
rect 18550 4165 18565 4185
rect 18585 4165 18600 4185
rect 18550 4135 18600 4165
rect 18550 4115 18565 4135
rect 18585 4115 18600 4135
rect 18550 4085 18600 4115
rect 18550 4065 18565 4085
rect 18585 4065 18600 4085
rect 18550 4035 18600 4065
rect 18550 4015 18565 4035
rect 18585 4015 18600 4035
rect 18550 3985 18600 4015
rect 18550 3965 18565 3985
rect 18585 3965 18600 3985
rect 18550 3950 18600 3965
rect 18700 4435 18750 4450
rect 18700 4415 18715 4435
rect 18735 4415 18750 4435
rect 18700 4385 18750 4415
rect 18700 4365 18715 4385
rect 18735 4365 18750 4385
rect 18700 4335 18750 4365
rect 18700 4315 18715 4335
rect 18735 4315 18750 4335
rect 18700 4285 18750 4315
rect 18700 4265 18715 4285
rect 18735 4265 18750 4285
rect 18700 4235 18750 4265
rect 18700 4215 18715 4235
rect 18735 4215 18750 4235
rect 18700 4185 18750 4215
rect 18700 4165 18715 4185
rect 18735 4165 18750 4185
rect 18700 4135 18750 4165
rect 18700 4115 18715 4135
rect 18735 4115 18750 4135
rect 18700 4085 18750 4115
rect 18700 4065 18715 4085
rect 18735 4065 18750 4085
rect 18700 4035 18750 4065
rect 18700 4015 18715 4035
rect 18735 4015 18750 4035
rect 18700 3985 18750 4015
rect 18700 3965 18715 3985
rect 18735 3965 18750 3985
rect 18700 3950 18750 3965
rect 18850 4435 18900 4450
rect 18850 4415 18865 4435
rect 18885 4415 18900 4435
rect 18850 4385 18900 4415
rect 18850 4365 18865 4385
rect 18885 4365 18900 4385
rect 18850 4335 18900 4365
rect 18850 4315 18865 4335
rect 18885 4315 18900 4335
rect 18850 4285 18900 4315
rect 18850 4265 18865 4285
rect 18885 4265 18900 4285
rect 18850 4235 18900 4265
rect 18850 4215 18865 4235
rect 18885 4215 18900 4235
rect 18850 4185 18900 4215
rect 18850 4165 18865 4185
rect 18885 4165 18900 4185
rect 18850 4135 18900 4165
rect 18850 4115 18865 4135
rect 18885 4115 18900 4135
rect 18850 4085 18900 4115
rect 18850 4065 18865 4085
rect 18885 4065 18900 4085
rect 18850 4035 18900 4065
rect 18850 4015 18865 4035
rect 18885 4015 18900 4035
rect 18850 3985 18900 4015
rect 18850 3965 18865 3985
rect 18885 3965 18900 3985
rect 18850 3950 18900 3965
rect 19000 4435 19050 4450
rect 19000 4415 19015 4435
rect 19035 4415 19050 4435
rect 19000 4385 19050 4415
rect 19000 4365 19015 4385
rect 19035 4365 19050 4385
rect 19000 4335 19050 4365
rect 19000 4315 19015 4335
rect 19035 4315 19050 4335
rect 19000 4285 19050 4315
rect 19000 4265 19015 4285
rect 19035 4265 19050 4285
rect 19000 4235 19050 4265
rect 19000 4215 19015 4235
rect 19035 4215 19050 4235
rect 19000 4185 19050 4215
rect 19000 4165 19015 4185
rect 19035 4165 19050 4185
rect 19000 4135 19050 4165
rect 19000 4115 19015 4135
rect 19035 4115 19050 4135
rect 19000 4085 19050 4115
rect 19000 4065 19015 4085
rect 19035 4065 19050 4085
rect 19000 4035 19050 4065
rect 19000 4015 19015 4035
rect 19035 4015 19050 4035
rect 19000 3985 19050 4015
rect 19000 3965 19015 3985
rect 19035 3965 19050 3985
rect 19000 3950 19050 3965
rect 19150 4435 19200 4450
rect 19150 4415 19165 4435
rect 19185 4415 19200 4435
rect 19150 4385 19200 4415
rect 19150 4365 19165 4385
rect 19185 4365 19200 4385
rect 19150 4335 19200 4365
rect 19150 4315 19165 4335
rect 19185 4315 19200 4335
rect 19150 4285 19200 4315
rect 19150 4265 19165 4285
rect 19185 4265 19200 4285
rect 19150 4235 19200 4265
rect 19150 4215 19165 4235
rect 19185 4215 19200 4235
rect 19150 4185 19200 4215
rect 19150 4165 19165 4185
rect 19185 4165 19200 4185
rect 19150 4135 19200 4165
rect 19150 4115 19165 4135
rect 19185 4115 19200 4135
rect 19150 4085 19200 4115
rect 19150 4065 19165 4085
rect 19185 4065 19200 4085
rect 19150 4035 19200 4065
rect 19150 4015 19165 4035
rect 19185 4015 19200 4035
rect 19150 3985 19200 4015
rect 19150 3965 19165 3985
rect 19185 3965 19200 3985
rect 19150 3950 19200 3965
rect 19300 4435 19350 4450
rect 19300 4415 19315 4435
rect 19335 4415 19350 4435
rect 19300 4385 19350 4415
rect 19300 4365 19315 4385
rect 19335 4365 19350 4385
rect 19300 4335 19350 4365
rect 19300 4315 19315 4335
rect 19335 4315 19350 4335
rect 19300 4285 19350 4315
rect 19300 4265 19315 4285
rect 19335 4265 19350 4285
rect 19300 4235 19350 4265
rect 19300 4215 19315 4235
rect 19335 4215 19350 4235
rect 19300 4185 19350 4215
rect 19300 4165 19315 4185
rect 19335 4165 19350 4185
rect 19300 4135 19350 4165
rect 19300 4115 19315 4135
rect 19335 4115 19350 4135
rect 19300 4085 19350 4115
rect 19300 4065 19315 4085
rect 19335 4065 19350 4085
rect 19300 4035 19350 4065
rect 19300 4015 19315 4035
rect 19335 4015 19350 4035
rect 19300 3985 19350 4015
rect 19300 3965 19315 3985
rect 19335 3965 19350 3985
rect 19300 3950 19350 3965
rect 19450 4435 19500 4450
rect 19450 4415 19465 4435
rect 19485 4415 19500 4435
rect 19450 4385 19500 4415
rect 19450 4365 19465 4385
rect 19485 4365 19500 4385
rect 19450 4335 19500 4365
rect 19450 4315 19465 4335
rect 19485 4315 19500 4335
rect 19450 4285 19500 4315
rect 19450 4265 19465 4285
rect 19485 4265 19500 4285
rect 19450 4235 19500 4265
rect 19450 4215 19465 4235
rect 19485 4215 19500 4235
rect 19450 4185 19500 4215
rect 19450 4165 19465 4185
rect 19485 4165 19500 4185
rect 19450 4135 19500 4165
rect 19450 4115 19465 4135
rect 19485 4115 19500 4135
rect 19450 4085 19500 4115
rect 19450 4065 19465 4085
rect 19485 4065 19500 4085
rect 19450 4035 19500 4065
rect 19450 4015 19465 4035
rect 19485 4015 19500 4035
rect 19450 3985 19500 4015
rect 19450 3965 19465 3985
rect 19485 3965 19500 3985
rect 19450 3950 19500 3965
rect 19600 4435 19650 4450
rect 19600 4415 19615 4435
rect 19635 4415 19650 4435
rect 19600 4385 19650 4415
rect 19600 4365 19615 4385
rect 19635 4365 19650 4385
rect 19600 4335 19650 4365
rect 19600 4315 19615 4335
rect 19635 4315 19650 4335
rect 19600 4285 19650 4315
rect 19600 4265 19615 4285
rect 19635 4265 19650 4285
rect 19600 4235 19650 4265
rect 19600 4215 19615 4235
rect 19635 4215 19650 4235
rect 19600 4185 19650 4215
rect 19600 4165 19615 4185
rect 19635 4165 19650 4185
rect 19600 4135 19650 4165
rect 19600 4115 19615 4135
rect 19635 4115 19650 4135
rect 19600 4085 19650 4115
rect 19600 4065 19615 4085
rect 19635 4065 19650 4085
rect 19600 4035 19650 4065
rect 19600 4015 19615 4035
rect 19635 4015 19650 4035
rect 19600 3985 19650 4015
rect 19600 3965 19615 3985
rect 19635 3965 19650 3985
rect 19600 3950 19650 3965
rect 19750 4435 19800 4450
rect 19750 4415 19765 4435
rect 19785 4415 19800 4435
rect 19750 4385 19800 4415
rect 19750 4365 19765 4385
rect 19785 4365 19800 4385
rect 19750 4335 19800 4365
rect 19750 4315 19765 4335
rect 19785 4315 19800 4335
rect 19750 4285 19800 4315
rect 19750 4265 19765 4285
rect 19785 4265 19800 4285
rect 19750 4235 19800 4265
rect 19750 4215 19765 4235
rect 19785 4215 19800 4235
rect 19750 4185 19800 4215
rect 19750 4165 19765 4185
rect 19785 4165 19800 4185
rect 19750 4135 19800 4165
rect 19750 4115 19765 4135
rect 19785 4115 19800 4135
rect 19750 4085 19800 4115
rect 19750 4065 19765 4085
rect 19785 4065 19800 4085
rect 19750 4035 19800 4065
rect 19750 4015 19765 4035
rect 19785 4015 19800 4035
rect 19750 3985 19800 4015
rect 19750 3965 19765 3985
rect 19785 3965 19800 3985
rect 19750 3950 19800 3965
rect 19900 3950 19950 4450
rect 20050 3950 20100 4450
rect 20200 3950 20250 4450
rect 20350 4435 20400 4450
rect 20350 4415 20365 4435
rect 20385 4415 20400 4435
rect 20350 4385 20400 4415
rect 20350 4365 20365 4385
rect 20385 4365 20400 4385
rect 20350 4335 20400 4365
rect 20350 4315 20365 4335
rect 20385 4315 20400 4335
rect 20350 4285 20400 4315
rect 20350 4265 20365 4285
rect 20385 4265 20400 4285
rect 20350 4235 20400 4265
rect 20350 4215 20365 4235
rect 20385 4215 20400 4235
rect 20350 4185 20400 4215
rect 20350 4165 20365 4185
rect 20385 4165 20400 4185
rect 20350 4135 20400 4165
rect 20350 4115 20365 4135
rect 20385 4115 20400 4135
rect 20350 4085 20400 4115
rect 20350 4065 20365 4085
rect 20385 4065 20400 4085
rect 20350 4035 20400 4065
rect 20350 4015 20365 4035
rect 20385 4015 20400 4035
rect 20350 3985 20400 4015
rect 20350 3965 20365 3985
rect 20385 3965 20400 3985
rect 20350 3950 20400 3965
rect -650 3785 -600 3800
rect -650 3765 -635 3785
rect -615 3765 -600 3785
rect -650 3735 -600 3765
rect -650 3715 -635 3735
rect -615 3715 -600 3735
rect -650 3685 -600 3715
rect -650 3665 -635 3685
rect -615 3665 -600 3685
rect -650 3635 -600 3665
rect -650 3615 -635 3635
rect -615 3615 -600 3635
rect -650 3585 -600 3615
rect -650 3565 -635 3585
rect -615 3565 -600 3585
rect -650 3535 -600 3565
rect -650 3515 -635 3535
rect -615 3515 -600 3535
rect -650 3485 -600 3515
rect -650 3465 -635 3485
rect -615 3465 -600 3485
rect -650 3435 -600 3465
rect -650 3415 -635 3435
rect -615 3415 -600 3435
rect -650 3385 -600 3415
rect -650 3365 -635 3385
rect -615 3365 -600 3385
rect -650 3335 -600 3365
rect -650 3315 -635 3335
rect -615 3315 -600 3335
rect -650 3300 -600 3315
rect -500 3785 -450 3800
rect -500 3765 -485 3785
rect -465 3765 -450 3785
rect -500 3735 -450 3765
rect -500 3715 -485 3735
rect -465 3715 -450 3735
rect -500 3685 -450 3715
rect -500 3665 -485 3685
rect -465 3665 -450 3685
rect -500 3635 -450 3665
rect -500 3615 -485 3635
rect -465 3615 -450 3635
rect -500 3585 -450 3615
rect -500 3565 -485 3585
rect -465 3565 -450 3585
rect -500 3535 -450 3565
rect -500 3515 -485 3535
rect -465 3515 -450 3535
rect -500 3485 -450 3515
rect -500 3465 -485 3485
rect -465 3465 -450 3485
rect -500 3435 -450 3465
rect -500 3415 -485 3435
rect -465 3415 -450 3435
rect -500 3385 -450 3415
rect -500 3365 -485 3385
rect -465 3365 -450 3385
rect -500 3335 -450 3365
rect -500 3315 -485 3335
rect -465 3315 -450 3335
rect -500 3300 -450 3315
rect -350 3785 -300 3800
rect -350 3765 -335 3785
rect -315 3765 -300 3785
rect -350 3735 -300 3765
rect -350 3715 -335 3735
rect -315 3715 -300 3735
rect -350 3685 -300 3715
rect -350 3665 -335 3685
rect -315 3665 -300 3685
rect -350 3635 -300 3665
rect -350 3615 -335 3635
rect -315 3615 -300 3635
rect -350 3585 -300 3615
rect -350 3565 -335 3585
rect -315 3565 -300 3585
rect -350 3535 -300 3565
rect -350 3515 -335 3535
rect -315 3515 -300 3535
rect -350 3485 -300 3515
rect -350 3465 -335 3485
rect -315 3465 -300 3485
rect -350 3435 -300 3465
rect -350 3415 -335 3435
rect -315 3415 -300 3435
rect -350 3385 -300 3415
rect -350 3365 -335 3385
rect -315 3365 -300 3385
rect -350 3335 -300 3365
rect -350 3315 -335 3335
rect -315 3315 -300 3335
rect -350 3300 -300 3315
rect -200 3785 -150 3800
rect -200 3765 -185 3785
rect -165 3765 -150 3785
rect -200 3735 -150 3765
rect -200 3715 -185 3735
rect -165 3715 -150 3735
rect -200 3685 -150 3715
rect -200 3665 -185 3685
rect -165 3665 -150 3685
rect -200 3635 -150 3665
rect -200 3615 -185 3635
rect -165 3615 -150 3635
rect -200 3585 -150 3615
rect -200 3565 -185 3585
rect -165 3565 -150 3585
rect -200 3535 -150 3565
rect -200 3515 -185 3535
rect -165 3515 -150 3535
rect -200 3485 -150 3515
rect -200 3465 -185 3485
rect -165 3465 -150 3485
rect -200 3435 -150 3465
rect -200 3415 -185 3435
rect -165 3415 -150 3435
rect -200 3385 -150 3415
rect -200 3365 -185 3385
rect -165 3365 -150 3385
rect -200 3335 -150 3365
rect -200 3315 -185 3335
rect -165 3315 -150 3335
rect -200 3300 -150 3315
rect -50 3785 0 3800
rect -50 3765 -35 3785
rect -15 3765 0 3785
rect -50 3735 0 3765
rect -50 3715 -35 3735
rect -15 3715 0 3735
rect -50 3685 0 3715
rect -50 3665 -35 3685
rect -15 3665 0 3685
rect -50 3635 0 3665
rect -50 3615 -35 3635
rect -15 3615 0 3635
rect -50 3585 0 3615
rect -50 3565 -35 3585
rect -15 3565 0 3585
rect -50 3535 0 3565
rect -50 3515 -35 3535
rect -15 3515 0 3535
rect -50 3485 0 3515
rect -50 3465 -35 3485
rect -15 3465 0 3485
rect -50 3435 0 3465
rect -50 3415 -35 3435
rect -15 3415 0 3435
rect -50 3385 0 3415
rect -50 3365 -35 3385
rect -15 3365 0 3385
rect -50 3335 0 3365
rect -50 3315 -35 3335
rect -15 3315 0 3335
rect -50 3300 0 3315
rect 100 3300 150 3800
rect 250 3300 300 3800
rect 400 3300 450 3800
rect 550 3785 600 3800
rect 550 3765 565 3785
rect 585 3765 600 3785
rect 550 3735 600 3765
rect 550 3715 565 3735
rect 585 3715 600 3735
rect 550 3685 600 3715
rect 550 3665 565 3685
rect 585 3665 600 3685
rect 550 3635 600 3665
rect 550 3615 565 3635
rect 585 3615 600 3635
rect 550 3585 600 3615
rect 550 3565 565 3585
rect 585 3565 600 3585
rect 550 3535 600 3565
rect 550 3515 565 3535
rect 585 3515 600 3535
rect 550 3485 600 3515
rect 550 3465 565 3485
rect 585 3465 600 3485
rect 550 3435 600 3465
rect 550 3415 565 3435
rect 585 3415 600 3435
rect 550 3385 600 3415
rect 550 3365 565 3385
rect 585 3365 600 3385
rect 550 3335 600 3365
rect 550 3315 565 3335
rect 585 3315 600 3335
rect 550 3300 600 3315
rect 700 3785 750 3800
rect 700 3765 715 3785
rect 735 3765 750 3785
rect 700 3735 750 3765
rect 700 3715 715 3735
rect 735 3715 750 3735
rect 700 3685 750 3715
rect 700 3665 715 3685
rect 735 3665 750 3685
rect 700 3635 750 3665
rect 700 3615 715 3635
rect 735 3615 750 3635
rect 700 3585 750 3615
rect 700 3565 715 3585
rect 735 3565 750 3585
rect 700 3535 750 3565
rect 700 3515 715 3535
rect 735 3515 750 3535
rect 700 3485 750 3515
rect 700 3465 715 3485
rect 735 3465 750 3485
rect 700 3435 750 3465
rect 700 3415 715 3435
rect 735 3415 750 3435
rect 700 3385 750 3415
rect 700 3365 715 3385
rect 735 3365 750 3385
rect 700 3335 750 3365
rect 700 3315 715 3335
rect 735 3315 750 3335
rect 700 3300 750 3315
rect 850 3785 900 3800
rect 850 3765 865 3785
rect 885 3765 900 3785
rect 850 3735 900 3765
rect 850 3715 865 3735
rect 885 3715 900 3735
rect 850 3685 900 3715
rect 850 3665 865 3685
rect 885 3665 900 3685
rect 850 3635 900 3665
rect 850 3615 865 3635
rect 885 3615 900 3635
rect 850 3585 900 3615
rect 850 3565 865 3585
rect 885 3565 900 3585
rect 850 3535 900 3565
rect 850 3515 865 3535
rect 885 3515 900 3535
rect 850 3485 900 3515
rect 850 3465 865 3485
rect 885 3465 900 3485
rect 850 3435 900 3465
rect 850 3415 865 3435
rect 885 3415 900 3435
rect 850 3385 900 3415
rect 850 3365 865 3385
rect 885 3365 900 3385
rect 850 3335 900 3365
rect 850 3315 865 3335
rect 885 3315 900 3335
rect 850 3300 900 3315
rect 1000 3785 1050 3800
rect 1000 3765 1015 3785
rect 1035 3765 1050 3785
rect 1000 3735 1050 3765
rect 1000 3715 1015 3735
rect 1035 3715 1050 3735
rect 1000 3685 1050 3715
rect 1000 3665 1015 3685
rect 1035 3665 1050 3685
rect 1000 3635 1050 3665
rect 1000 3615 1015 3635
rect 1035 3615 1050 3635
rect 1000 3585 1050 3615
rect 1000 3565 1015 3585
rect 1035 3565 1050 3585
rect 1000 3535 1050 3565
rect 1000 3515 1015 3535
rect 1035 3515 1050 3535
rect 1000 3485 1050 3515
rect 1000 3465 1015 3485
rect 1035 3465 1050 3485
rect 1000 3435 1050 3465
rect 1000 3415 1015 3435
rect 1035 3415 1050 3435
rect 1000 3385 1050 3415
rect 1000 3365 1015 3385
rect 1035 3365 1050 3385
rect 1000 3335 1050 3365
rect 1000 3315 1015 3335
rect 1035 3315 1050 3335
rect 1000 3300 1050 3315
rect 1150 3785 1200 3800
rect 1150 3765 1165 3785
rect 1185 3765 1200 3785
rect 1150 3735 1200 3765
rect 1150 3715 1165 3735
rect 1185 3715 1200 3735
rect 1150 3685 1200 3715
rect 1150 3665 1165 3685
rect 1185 3665 1200 3685
rect 1150 3635 1200 3665
rect 1150 3615 1165 3635
rect 1185 3615 1200 3635
rect 1150 3585 1200 3615
rect 1150 3565 1165 3585
rect 1185 3565 1200 3585
rect 1150 3535 1200 3565
rect 1150 3515 1165 3535
rect 1185 3515 1200 3535
rect 1150 3485 1200 3515
rect 1150 3465 1165 3485
rect 1185 3465 1200 3485
rect 1150 3435 1200 3465
rect 1150 3415 1165 3435
rect 1185 3415 1200 3435
rect 1150 3385 1200 3415
rect 1150 3365 1165 3385
rect 1185 3365 1200 3385
rect 1150 3335 1200 3365
rect 1150 3315 1165 3335
rect 1185 3315 1200 3335
rect 1150 3300 1200 3315
rect 1300 3785 1350 3800
rect 1300 3765 1315 3785
rect 1335 3765 1350 3785
rect 1300 3735 1350 3765
rect 1300 3715 1315 3735
rect 1335 3715 1350 3735
rect 1300 3685 1350 3715
rect 1300 3665 1315 3685
rect 1335 3665 1350 3685
rect 1300 3635 1350 3665
rect 1300 3615 1315 3635
rect 1335 3615 1350 3635
rect 1300 3585 1350 3615
rect 1300 3565 1315 3585
rect 1335 3565 1350 3585
rect 1300 3535 1350 3565
rect 1300 3515 1315 3535
rect 1335 3515 1350 3535
rect 1300 3485 1350 3515
rect 1300 3465 1315 3485
rect 1335 3465 1350 3485
rect 1300 3435 1350 3465
rect 1300 3415 1315 3435
rect 1335 3415 1350 3435
rect 1300 3385 1350 3415
rect 1300 3365 1315 3385
rect 1335 3365 1350 3385
rect 1300 3335 1350 3365
rect 1300 3315 1315 3335
rect 1335 3315 1350 3335
rect 1300 3300 1350 3315
rect 1450 3785 1500 3800
rect 1450 3765 1465 3785
rect 1485 3765 1500 3785
rect 1450 3735 1500 3765
rect 1450 3715 1465 3735
rect 1485 3715 1500 3735
rect 1450 3685 1500 3715
rect 1450 3665 1465 3685
rect 1485 3665 1500 3685
rect 1450 3635 1500 3665
rect 1450 3615 1465 3635
rect 1485 3615 1500 3635
rect 1450 3585 1500 3615
rect 1450 3565 1465 3585
rect 1485 3565 1500 3585
rect 1450 3535 1500 3565
rect 1450 3515 1465 3535
rect 1485 3515 1500 3535
rect 1450 3485 1500 3515
rect 1450 3465 1465 3485
rect 1485 3465 1500 3485
rect 1450 3435 1500 3465
rect 1450 3415 1465 3435
rect 1485 3415 1500 3435
rect 1450 3385 1500 3415
rect 1450 3365 1465 3385
rect 1485 3365 1500 3385
rect 1450 3335 1500 3365
rect 1450 3315 1465 3335
rect 1485 3315 1500 3335
rect 1450 3300 1500 3315
rect 1600 3785 1650 3800
rect 1600 3765 1615 3785
rect 1635 3765 1650 3785
rect 1600 3735 1650 3765
rect 1600 3715 1615 3735
rect 1635 3715 1650 3735
rect 1600 3685 1650 3715
rect 1600 3665 1615 3685
rect 1635 3665 1650 3685
rect 1600 3635 1650 3665
rect 1600 3615 1615 3635
rect 1635 3615 1650 3635
rect 1600 3585 1650 3615
rect 1600 3565 1615 3585
rect 1635 3565 1650 3585
rect 1600 3535 1650 3565
rect 1600 3515 1615 3535
rect 1635 3515 1650 3535
rect 1600 3485 1650 3515
rect 1600 3465 1615 3485
rect 1635 3465 1650 3485
rect 1600 3435 1650 3465
rect 1600 3415 1615 3435
rect 1635 3415 1650 3435
rect 1600 3385 1650 3415
rect 1600 3365 1615 3385
rect 1635 3365 1650 3385
rect 1600 3335 1650 3365
rect 1600 3315 1615 3335
rect 1635 3315 1650 3335
rect 1600 3300 1650 3315
rect 1750 3785 1800 3800
rect 1750 3765 1765 3785
rect 1785 3765 1800 3785
rect 1750 3735 1800 3765
rect 1750 3715 1765 3735
rect 1785 3715 1800 3735
rect 1750 3685 1800 3715
rect 1750 3665 1765 3685
rect 1785 3665 1800 3685
rect 1750 3635 1800 3665
rect 1750 3615 1765 3635
rect 1785 3615 1800 3635
rect 1750 3585 1800 3615
rect 1750 3565 1765 3585
rect 1785 3565 1800 3585
rect 1750 3535 1800 3565
rect 1750 3515 1765 3535
rect 1785 3515 1800 3535
rect 1750 3485 1800 3515
rect 1750 3465 1765 3485
rect 1785 3465 1800 3485
rect 1750 3435 1800 3465
rect 1750 3415 1765 3435
rect 1785 3415 1800 3435
rect 1750 3385 1800 3415
rect 1750 3365 1765 3385
rect 1785 3365 1800 3385
rect 1750 3335 1800 3365
rect 1750 3315 1765 3335
rect 1785 3315 1800 3335
rect 1750 3300 1800 3315
rect 1900 3785 1950 3800
rect 1900 3765 1915 3785
rect 1935 3765 1950 3785
rect 1900 3735 1950 3765
rect 1900 3715 1915 3735
rect 1935 3715 1950 3735
rect 1900 3685 1950 3715
rect 1900 3665 1915 3685
rect 1935 3665 1950 3685
rect 1900 3635 1950 3665
rect 1900 3615 1915 3635
rect 1935 3615 1950 3635
rect 1900 3585 1950 3615
rect 1900 3565 1915 3585
rect 1935 3565 1950 3585
rect 1900 3535 1950 3565
rect 1900 3515 1915 3535
rect 1935 3515 1950 3535
rect 1900 3485 1950 3515
rect 1900 3465 1915 3485
rect 1935 3465 1950 3485
rect 1900 3435 1950 3465
rect 1900 3415 1915 3435
rect 1935 3415 1950 3435
rect 1900 3385 1950 3415
rect 1900 3365 1915 3385
rect 1935 3365 1950 3385
rect 1900 3335 1950 3365
rect 1900 3315 1915 3335
rect 1935 3315 1950 3335
rect 1900 3300 1950 3315
rect 2050 3785 2100 3800
rect 2050 3765 2065 3785
rect 2085 3765 2100 3785
rect 2050 3735 2100 3765
rect 2050 3715 2065 3735
rect 2085 3715 2100 3735
rect 2050 3685 2100 3715
rect 2050 3665 2065 3685
rect 2085 3665 2100 3685
rect 2050 3635 2100 3665
rect 2050 3615 2065 3635
rect 2085 3615 2100 3635
rect 2050 3585 2100 3615
rect 2050 3565 2065 3585
rect 2085 3565 2100 3585
rect 2050 3535 2100 3565
rect 2050 3515 2065 3535
rect 2085 3515 2100 3535
rect 2050 3485 2100 3515
rect 2050 3465 2065 3485
rect 2085 3465 2100 3485
rect 2050 3435 2100 3465
rect 2050 3415 2065 3435
rect 2085 3415 2100 3435
rect 2050 3385 2100 3415
rect 2050 3365 2065 3385
rect 2085 3365 2100 3385
rect 2050 3335 2100 3365
rect 2050 3315 2065 3335
rect 2085 3315 2100 3335
rect 2050 3300 2100 3315
rect 2200 3785 2250 3800
rect 2200 3765 2215 3785
rect 2235 3765 2250 3785
rect 2200 3735 2250 3765
rect 2200 3715 2215 3735
rect 2235 3715 2250 3735
rect 2200 3685 2250 3715
rect 2200 3665 2215 3685
rect 2235 3665 2250 3685
rect 2200 3635 2250 3665
rect 2200 3615 2215 3635
rect 2235 3615 2250 3635
rect 2200 3585 2250 3615
rect 2200 3565 2215 3585
rect 2235 3565 2250 3585
rect 2200 3535 2250 3565
rect 2200 3515 2215 3535
rect 2235 3515 2250 3535
rect 2200 3485 2250 3515
rect 2200 3465 2215 3485
rect 2235 3465 2250 3485
rect 2200 3435 2250 3465
rect 2200 3415 2215 3435
rect 2235 3415 2250 3435
rect 2200 3385 2250 3415
rect 2200 3365 2215 3385
rect 2235 3365 2250 3385
rect 2200 3335 2250 3365
rect 2200 3315 2215 3335
rect 2235 3315 2250 3335
rect 2200 3300 2250 3315
rect 2350 3785 2400 3800
rect 2350 3765 2365 3785
rect 2385 3765 2400 3785
rect 2350 3735 2400 3765
rect 2350 3715 2365 3735
rect 2385 3715 2400 3735
rect 2350 3685 2400 3715
rect 2350 3665 2365 3685
rect 2385 3665 2400 3685
rect 2350 3635 2400 3665
rect 2350 3615 2365 3635
rect 2385 3615 2400 3635
rect 2350 3585 2400 3615
rect 2350 3565 2365 3585
rect 2385 3565 2400 3585
rect 2350 3535 2400 3565
rect 2350 3515 2365 3535
rect 2385 3515 2400 3535
rect 2350 3485 2400 3515
rect 2350 3465 2365 3485
rect 2385 3465 2400 3485
rect 2350 3435 2400 3465
rect 2350 3415 2365 3435
rect 2385 3415 2400 3435
rect 2350 3385 2400 3415
rect 2350 3365 2365 3385
rect 2385 3365 2400 3385
rect 2350 3335 2400 3365
rect 2350 3315 2365 3335
rect 2385 3315 2400 3335
rect 2350 3300 2400 3315
rect 2500 3785 2550 3800
rect 2500 3765 2515 3785
rect 2535 3765 2550 3785
rect 2500 3735 2550 3765
rect 2500 3715 2515 3735
rect 2535 3715 2550 3735
rect 2500 3685 2550 3715
rect 2500 3665 2515 3685
rect 2535 3665 2550 3685
rect 2500 3635 2550 3665
rect 2500 3615 2515 3635
rect 2535 3615 2550 3635
rect 2500 3585 2550 3615
rect 2500 3565 2515 3585
rect 2535 3565 2550 3585
rect 2500 3535 2550 3565
rect 2500 3515 2515 3535
rect 2535 3515 2550 3535
rect 2500 3485 2550 3515
rect 2500 3465 2515 3485
rect 2535 3465 2550 3485
rect 2500 3435 2550 3465
rect 2500 3415 2515 3435
rect 2535 3415 2550 3435
rect 2500 3385 2550 3415
rect 2500 3365 2515 3385
rect 2535 3365 2550 3385
rect 2500 3335 2550 3365
rect 2500 3315 2515 3335
rect 2535 3315 2550 3335
rect 2500 3300 2550 3315
rect 2650 3785 2700 3800
rect 2650 3765 2665 3785
rect 2685 3765 2700 3785
rect 2650 3735 2700 3765
rect 2650 3715 2665 3735
rect 2685 3715 2700 3735
rect 2650 3685 2700 3715
rect 2650 3665 2665 3685
rect 2685 3665 2700 3685
rect 2650 3635 2700 3665
rect 2650 3615 2665 3635
rect 2685 3615 2700 3635
rect 2650 3585 2700 3615
rect 2650 3565 2665 3585
rect 2685 3565 2700 3585
rect 2650 3535 2700 3565
rect 2650 3515 2665 3535
rect 2685 3515 2700 3535
rect 2650 3485 2700 3515
rect 2650 3465 2665 3485
rect 2685 3465 2700 3485
rect 2650 3435 2700 3465
rect 2650 3415 2665 3435
rect 2685 3415 2700 3435
rect 2650 3385 2700 3415
rect 2650 3365 2665 3385
rect 2685 3365 2700 3385
rect 2650 3335 2700 3365
rect 2650 3315 2665 3335
rect 2685 3315 2700 3335
rect 2650 3300 2700 3315
rect 2800 3785 2850 3800
rect 2800 3765 2815 3785
rect 2835 3765 2850 3785
rect 2800 3735 2850 3765
rect 2800 3715 2815 3735
rect 2835 3715 2850 3735
rect 2800 3685 2850 3715
rect 2800 3665 2815 3685
rect 2835 3665 2850 3685
rect 2800 3635 2850 3665
rect 2800 3615 2815 3635
rect 2835 3615 2850 3635
rect 2800 3585 2850 3615
rect 2800 3565 2815 3585
rect 2835 3565 2850 3585
rect 2800 3535 2850 3565
rect 2800 3515 2815 3535
rect 2835 3515 2850 3535
rect 2800 3485 2850 3515
rect 2800 3465 2815 3485
rect 2835 3465 2850 3485
rect 2800 3435 2850 3465
rect 2800 3415 2815 3435
rect 2835 3415 2850 3435
rect 2800 3385 2850 3415
rect 2800 3365 2815 3385
rect 2835 3365 2850 3385
rect 2800 3335 2850 3365
rect 2800 3315 2815 3335
rect 2835 3315 2850 3335
rect 2800 3300 2850 3315
rect 2950 3785 3000 3800
rect 2950 3765 2965 3785
rect 2985 3765 3000 3785
rect 2950 3735 3000 3765
rect 2950 3715 2965 3735
rect 2985 3715 3000 3735
rect 2950 3685 3000 3715
rect 2950 3665 2965 3685
rect 2985 3665 3000 3685
rect 2950 3635 3000 3665
rect 2950 3615 2965 3635
rect 2985 3615 3000 3635
rect 2950 3585 3000 3615
rect 2950 3565 2965 3585
rect 2985 3565 3000 3585
rect 2950 3535 3000 3565
rect 2950 3515 2965 3535
rect 2985 3515 3000 3535
rect 2950 3485 3000 3515
rect 2950 3465 2965 3485
rect 2985 3465 3000 3485
rect 2950 3435 3000 3465
rect 2950 3415 2965 3435
rect 2985 3415 3000 3435
rect 2950 3385 3000 3415
rect 2950 3365 2965 3385
rect 2985 3365 3000 3385
rect 2950 3335 3000 3365
rect 2950 3315 2965 3335
rect 2985 3315 3000 3335
rect 2950 3300 3000 3315
rect 3100 3785 3150 3800
rect 3100 3765 3115 3785
rect 3135 3765 3150 3785
rect 3100 3735 3150 3765
rect 3100 3715 3115 3735
rect 3135 3715 3150 3735
rect 3100 3685 3150 3715
rect 3100 3665 3115 3685
rect 3135 3665 3150 3685
rect 3100 3635 3150 3665
rect 3100 3615 3115 3635
rect 3135 3615 3150 3635
rect 3100 3585 3150 3615
rect 3100 3565 3115 3585
rect 3135 3565 3150 3585
rect 3100 3535 3150 3565
rect 3100 3515 3115 3535
rect 3135 3515 3150 3535
rect 3100 3485 3150 3515
rect 3100 3465 3115 3485
rect 3135 3465 3150 3485
rect 3100 3435 3150 3465
rect 3100 3415 3115 3435
rect 3135 3415 3150 3435
rect 3100 3385 3150 3415
rect 3100 3365 3115 3385
rect 3135 3365 3150 3385
rect 3100 3335 3150 3365
rect 3100 3315 3115 3335
rect 3135 3315 3150 3335
rect 3100 3300 3150 3315
rect 3250 3785 3300 3800
rect 3250 3765 3265 3785
rect 3285 3765 3300 3785
rect 3250 3735 3300 3765
rect 3250 3715 3265 3735
rect 3285 3715 3300 3735
rect 3250 3685 3300 3715
rect 3250 3665 3265 3685
rect 3285 3665 3300 3685
rect 3250 3635 3300 3665
rect 3250 3615 3265 3635
rect 3285 3615 3300 3635
rect 3250 3585 3300 3615
rect 3250 3565 3265 3585
rect 3285 3565 3300 3585
rect 3250 3535 3300 3565
rect 3250 3515 3265 3535
rect 3285 3515 3300 3535
rect 3250 3485 3300 3515
rect 3250 3465 3265 3485
rect 3285 3465 3300 3485
rect 3250 3435 3300 3465
rect 3250 3415 3265 3435
rect 3285 3415 3300 3435
rect 3250 3385 3300 3415
rect 3250 3365 3265 3385
rect 3285 3365 3300 3385
rect 3250 3335 3300 3365
rect 3250 3315 3265 3335
rect 3285 3315 3300 3335
rect 3250 3300 3300 3315
rect 3400 3785 3450 3800
rect 3400 3765 3415 3785
rect 3435 3765 3450 3785
rect 3400 3735 3450 3765
rect 3400 3715 3415 3735
rect 3435 3715 3450 3735
rect 3400 3685 3450 3715
rect 3400 3665 3415 3685
rect 3435 3665 3450 3685
rect 3400 3635 3450 3665
rect 3400 3615 3415 3635
rect 3435 3615 3450 3635
rect 3400 3585 3450 3615
rect 3400 3565 3415 3585
rect 3435 3565 3450 3585
rect 3400 3535 3450 3565
rect 3400 3515 3415 3535
rect 3435 3515 3450 3535
rect 3400 3485 3450 3515
rect 3400 3465 3415 3485
rect 3435 3465 3450 3485
rect 3400 3435 3450 3465
rect 3400 3415 3415 3435
rect 3435 3415 3450 3435
rect 3400 3385 3450 3415
rect 3400 3365 3415 3385
rect 3435 3365 3450 3385
rect 3400 3335 3450 3365
rect 3400 3315 3415 3335
rect 3435 3315 3450 3335
rect 3400 3300 3450 3315
rect 3550 3785 3600 3800
rect 3550 3765 3565 3785
rect 3585 3765 3600 3785
rect 3550 3735 3600 3765
rect 3550 3715 3565 3735
rect 3585 3715 3600 3735
rect 3550 3685 3600 3715
rect 3550 3665 3565 3685
rect 3585 3665 3600 3685
rect 3550 3635 3600 3665
rect 3550 3615 3565 3635
rect 3585 3615 3600 3635
rect 3550 3585 3600 3615
rect 3550 3565 3565 3585
rect 3585 3565 3600 3585
rect 3550 3535 3600 3565
rect 3550 3515 3565 3535
rect 3585 3515 3600 3535
rect 3550 3485 3600 3515
rect 3550 3465 3565 3485
rect 3585 3465 3600 3485
rect 3550 3435 3600 3465
rect 3550 3415 3565 3435
rect 3585 3415 3600 3435
rect 3550 3385 3600 3415
rect 3550 3365 3565 3385
rect 3585 3365 3600 3385
rect 3550 3335 3600 3365
rect 3550 3315 3565 3335
rect 3585 3315 3600 3335
rect 3550 3300 3600 3315
rect 3700 3300 3750 3800
rect 3850 3300 3900 3800
rect 4000 3300 4050 3800
rect 4150 3785 4200 3800
rect 4150 3765 4165 3785
rect 4185 3765 4200 3785
rect 4150 3735 4200 3765
rect 4150 3715 4165 3735
rect 4185 3715 4200 3735
rect 4150 3685 4200 3715
rect 4150 3665 4165 3685
rect 4185 3665 4200 3685
rect 4150 3635 4200 3665
rect 4150 3615 4165 3635
rect 4185 3615 4200 3635
rect 4150 3585 4200 3615
rect 4150 3565 4165 3585
rect 4185 3565 4200 3585
rect 4150 3535 4200 3565
rect 4150 3515 4165 3535
rect 4185 3515 4200 3535
rect 4150 3485 4200 3515
rect 4150 3465 4165 3485
rect 4185 3465 4200 3485
rect 4150 3435 4200 3465
rect 4150 3415 4165 3435
rect 4185 3415 4200 3435
rect 4150 3385 4200 3415
rect 4150 3365 4165 3385
rect 4185 3365 4200 3385
rect 4150 3335 4200 3365
rect 4150 3315 4165 3335
rect 4185 3315 4200 3335
rect 4150 3300 4200 3315
rect 4300 3300 4350 3800
rect 4450 3300 4500 3800
rect 4600 3300 4650 3800
rect 4750 3785 4800 3800
rect 4750 3765 4765 3785
rect 4785 3765 4800 3785
rect 4750 3735 4800 3765
rect 4750 3715 4765 3735
rect 4785 3715 4800 3735
rect 4750 3685 4800 3715
rect 4750 3665 4765 3685
rect 4785 3665 4800 3685
rect 4750 3635 4800 3665
rect 4750 3615 4765 3635
rect 4785 3615 4800 3635
rect 4750 3585 4800 3615
rect 4750 3565 4765 3585
rect 4785 3565 4800 3585
rect 4750 3535 4800 3565
rect 4750 3515 4765 3535
rect 4785 3515 4800 3535
rect 4750 3485 4800 3515
rect 4750 3465 4765 3485
rect 4785 3465 4800 3485
rect 4750 3435 4800 3465
rect 4750 3415 4765 3435
rect 4785 3415 4800 3435
rect 4750 3385 4800 3415
rect 4750 3365 4765 3385
rect 4785 3365 4800 3385
rect 4750 3335 4800 3365
rect 4750 3315 4765 3335
rect 4785 3315 4800 3335
rect 4750 3300 4800 3315
rect 4900 3785 4950 3800
rect 4900 3765 4915 3785
rect 4935 3765 4950 3785
rect 4900 3735 4950 3765
rect 4900 3715 4915 3735
rect 4935 3715 4950 3735
rect 4900 3685 4950 3715
rect 4900 3665 4915 3685
rect 4935 3665 4950 3685
rect 4900 3635 4950 3665
rect 4900 3615 4915 3635
rect 4935 3615 4950 3635
rect 4900 3585 4950 3615
rect 4900 3565 4915 3585
rect 4935 3565 4950 3585
rect 4900 3535 4950 3565
rect 4900 3515 4915 3535
rect 4935 3515 4950 3535
rect 4900 3485 4950 3515
rect 4900 3465 4915 3485
rect 4935 3465 4950 3485
rect 4900 3435 4950 3465
rect 4900 3415 4915 3435
rect 4935 3415 4950 3435
rect 4900 3385 4950 3415
rect 4900 3365 4915 3385
rect 4935 3365 4950 3385
rect 4900 3335 4950 3365
rect 4900 3315 4915 3335
rect 4935 3315 4950 3335
rect 4900 3300 4950 3315
rect 5050 3785 5100 3800
rect 5050 3765 5065 3785
rect 5085 3765 5100 3785
rect 5050 3735 5100 3765
rect 5050 3715 5065 3735
rect 5085 3715 5100 3735
rect 5050 3685 5100 3715
rect 5050 3665 5065 3685
rect 5085 3665 5100 3685
rect 5050 3635 5100 3665
rect 5050 3615 5065 3635
rect 5085 3615 5100 3635
rect 5050 3585 5100 3615
rect 5050 3565 5065 3585
rect 5085 3565 5100 3585
rect 5050 3535 5100 3565
rect 5050 3515 5065 3535
rect 5085 3515 5100 3535
rect 5050 3485 5100 3515
rect 5050 3465 5065 3485
rect 5085 3465 5100 3485
rect 5050 3435 5100 3465
rect 5050 3415 5065 3435
rect 5085 3415 5100 3435
rect 5050 3385 5100 3415
rect 5050 3365 5065 3385
rect 5085 3365 5100 3385
rect 5050 3335 5100 3365
rect 5050 3315 5065 3335
rect 5085 3315 5100 3335
rect 5050 3300 5100 3315
rect 5200 3785 5250 3800
rect 5200 3765 5215 3785
rect 5235 3765 5250 3785
rect 5200 3735 5250 3765
rect 5200 3715 5215 3735
rect 5235 3715 5250 3735
rect 5200 3685 5250 3715
rect 5200 3665 5215 3685
rect 5235 3665 5250 3685
rect 5200 3635 5250 3665
rect 5200 3615 5215 3635
rect 5235 3615 5250 3635
rect 5200 3585 5250 3615
rect 5200 3565 5215 3585
rect 5235 3565 5250 3585
rect 5200 3535 5250 3565
rect 5200 3515 5215 3535
rect 5235 3515 5250 3535
rect 5200 3485 5250 3515
rect 5200 3465 5215 3485
rect 5235 3465 5250 3485
rect 5200 3435 5250 3465
rect 5200 3415 5215 3435
rect 5235 3415 5250 3435
rect 5200 3385 5250 3415
rect 5200 3365 5215 3385
rect 5235 3365 5250 3385
rect 5200 3335 5250 3365
rect 5200 3315 5215 3335
rect 5235 3315 5250 3335
rect 5200 3300 5250 3315
rect 5350 3785 5400 3800
rect 5350 3765 5365 3785
rect 5385 3765 5400 3785
rect 5350 3735 5400 3765
rect 5350 3715 5365 3735
rect 5385 3715 5400 3735
rect 5350 3685 5400 3715
rect 5350 3665 5365 3685
rect 5385 3665 5400 3685
rect 5350 3635 5400 3665
rect 5350 3615 5365 3635
rect 5385 3615 5400 3635
rect 5350 3585 5400 3615
rect 5350 3565 5365 3585
rect 5385 3565 5400 3585
rect 5350 3535 5400 3565
rect 5350 3515 5365 3535
rect 5385 3515 5400 3535
rect 5350 3485 5400 3515
rect 5350 3465 5365 3485
rect 5385 3465 5400 3485
rect 5350 3435 5400 3465
rect 5350 3415 5365 3435
rect 5385 3415 5400 3435
rect 5350 3385 5400 3415
rect 5350 3365 5365 3385
rect 5385 3365 5400 3385
rect 5350 3335 5400 3365
rect 5350 3315 5365 3335
rect 5385 3315 5400 3335
rect 5350 3300 5400 3315
rect 5500 3785 5550 3800
rect 5500 3765 5515 3785
rect 5535 3765 5550 3785
rect 5500 3735 5550 3765
rect 5500 3715 5515 3735
rect 5535 3715 5550 3735
rect 5500 3685 5550 3715
rect 5500 3665 5515 3685
rect 5535 3665 5550 3685
rect 5500 3635 5550 3665
rect 5500 3615 5515 3635
rect 5535 3615 5550 3635
rect 5500 3585 5550 3615
rect 5500 3565 5515 3585
rect 5535 3565 5550 3585
rect 5500 3535 5550 3565
rect 5500 3515 5515 3535
rect 5535 3515 5550 3535
rect 5500 3485 5550 3515
rect 5500 3465 5515 3485
rect 5535 3465 5550 3485
rect 5500 3435 5550 3465
rect 5500 3415 5515 3435
rect 5535 3415 5550 3435
rect 5500 3385 5550 3415
rect 5500 3365 5515 3385
rect 5535 3365 5550 3385
rect 5500 3335 5550 3365
rect 5500 3315 5515 3335
rect 5535 3315 5550 3335
rect 5500 3300 5550 3315
rect 5650 3785 5700 3800
rect 5650 3765 5665 3785
rect 5685 3765 5700 3785
rect 5650 3735 5700 3765
rect 5650 3715 5665 3735
rect 5685 3715 5700 3735
rect 5650 3685 5700 3715
rect 5650 3665 5665 3685
rect 5685 3665 5700 3685
rect 5650 3635 5700 3665
rect 5650 3615 5665 3635
rect 5685 3615 5700 3635
rect 5650 3585 5700 3615
rect 5650 3565 5665 3585
rect 5685 3565 5700 3585
rect 5650 3535 5700 3565
rect 5650 3515 5665 3535
rect 5685 3515 5700 3535
rect 5650 3485 5700 3515
rect 5650 3465 5665 3485
rect 5685 3465 5700 3485
rect 5650 3435 5700 3465
rect 5650 3415 5665 3435
rect 5685 3415 5700 3435
rect 5650 3385 5700 3415
rect 5650 3365 5665 3385
rect 5685 3365 5700 3385
rect 5650 3335 5700 3365
rect 5650 3315 5665 3335
rect 5685 3315 5700 3335
rect 5650 3300 5700 3315
rect 5800 3785 5850 3800
rect 5800 3765 5815 3785
rect 5835 3765 5850 3785
rect 5800 3735 5850 3765
rect 5800 3715 5815 3735
rect 5835 3715 5850 3735
rect 5800 3685 5850 3715
rect 5800 3665 5815 3685
rect 5835 3665 5850 3685
rect 5800 3635 5850 3665
rect 5800 3615 5815 3635
rect 5835 3615 5850 3635
rect 5800 3585 5850 3615
rect 5800 3565 5815 3585
rect 5835 3565 5850 3585
rect 5800 3535 5850 3565
rect 5800 3515 5815 3535
rect 5835 3515 5850 3535
rect 5800 3485 5850 3515
rect 5800 3465 5815 3485
rect 5835 3465 5850 3485
rect 5800 3435 5850 3465
rect 5800 3415 5815 3435
rect 5835 3415 5850 3435
rect 5800 3385 5850 3415
rect 5800 3365 5815 3385
rect 5835 3365 5850 3385
rect 5800 3335 5850 3365
rect 5800 3315 5815 3335
rect 5835 3315 5850 3335
rect 5800 3300 5850 3315
rect 5950 3785 6000 3800
rect 5950 3765 5965 3785
rect 5985 3765 6000 3785
rect 5950 3735 6000 3765
rect 5950 3715 5965 3735
rect 5985 3715 6000 3735
rect 5950 3685 6000 3715
rect 5950 3665 5965 3685
rect 5985 3665 6000 3685
rect 5950 3635 6000 3665
rect 5950 3615 5965 3635
rect 5985 3615 6000 3635
rect 5950 3585 6000 3615
rect 5950 3565 5965 3585
rect 5985 3565 6000 3585
rect 5950 3535 6000 3565
rect 5950 3515 5965 3535
rect 5985 3515 6000 3535
rect 5950 3485 6000 3515
rect 5950 3465 5965 3485
rect 5985 3465 6000 3485
rect 5950 3435 6000 3465
rect 5950 3415 5965 3435
rect 5985 3415 6000 3435
rect 5950 3385 6000 3415
rect 5950 3365 5965 3385
rect 5985 3365 6000 3385
rect 5950 3335 6000 3365
rect 5950 3315 5965 3335
rect 5985 3315 6000 3335
rect 5950 3300 6000 3315
rect 6100 3785 6150 3800
rect 6100 3765 6115 3785
rect 6135 3765 6150 3785
rect 6100 3735 6150 3765
rect 6100 3715 6115 3735
rect 6135 3715 6150 3735
rect 6100 3685 6150 3715
rect 6100 3665 6115 3685
rect 6135 3665 6150 3685
rect 6100 3635 6150 3665
rect 6100 3615 6115 3635
rect 6135 3615 6150 3635
rect 6100 3585 6150 3615
rect 6100 3565 6115 3585
rect 6135 3565 6150 3585
rect 6100 3535 6150 3565
rect 6100 3515 6115 3535
rect 6135 3515 6150 3535
rect 6100 3485 6150 3515
rect 6100 3465 6115 3485
rect 6135 3465 6150 3485
rect 6100 3435 6150 3465
rect 6100 3415 6115 3435
rect 6135 3415 6150 3435
rect 6100 3385 6150 3415
rect 6100 3365 6115 3385
rect 6135 3365 6150 3385
rect 6100 3335 6150 3365
rect 6100 3315 6115 3335
rect 6135 3315 6150 3335
rect 6100 3300 6150 3315
rect 6250 3785 6300 3800
rect 6250 3765 6265 3785
rect 6285 3765 6300 3785
rect 6250 3735 6300 3765
rect 6250 3715 6265 3735
rect 6285 3715 6300 3735
rect 6250 3685 6300 3715
rect 6250 3665 6265 3685
rect 6285 3665 6300 3685
rect 6250 3635 6300 3665
rect 6250 3615 6265 3635
rect 6285 3615 6300 3635
rect 6250 3585 6300 3615
rect 6250 3565 6265 3585
rect 6285 3565 6300 3585
rect 6250 3535 6300 3565
rect 6250 3515 6265 3535
rect 6285 3515 6300 3535
rect 6250 3485 6300 3515
rect 6250 3465 6265 3485
rect 6285 3465 6300 3485
rect 6250 3435 6300 3465
rect 6250 3415 6265 3435
rect 6285 3415 6300 3435
rect 6250 3385 6300 3415
rect 6250 3365 6265 3385
rect 6285 3365 6300 3385
rect 6250 3335 6300 3365
rect 6250 3315 6265 3335
rect 6285 3315 6300 3335
rect 6250 3300 6300 3315
rect 6400 3785 6450 3800
rect 6400 3765 6415 3785
rect 6435 3765 6450 3785
rect 6400 3735 6450 3765
rect 6400 3715 6415 3735
rect 6435 3715 6450 3735
rect 6400 3685 6450 3715
rect 6400 3665 6415 3685
rect 6435 3665 6450 3685
rect 6400 3635 6450 3665
rect 6400 3615 6415 3635
rect 6435 3615 6450 3635
rect 6400 3585 6450 3615
rect 6400 3565 6415 3585
rect 6435 3565 6450 3585
rect 6400 3535 6450 3565
rect 6400 3515 6415 3535
rect 6435 3515 6450 3535
rect 6400 3485 6450 3515
rect 6400 3465 6415 3485
rect 6435 3465 6450 3485
rect 6400 3435 6450 3465
rect 6400 3415 6415 3435
rect 6435 3415 6450 3435
rect 6400 3385 6450 3415
rect 6400 3365 6415 3385
rect 6435 3365 6450 3385
rect 6400 3335 6450 3365
rect 6400 3315 6415 3335
rect 6435 3315 6450 3335
rect 6400 3300 6450 3315
rect 6550 3785 6600 3800
rect 6550 3765 6565 3785
rect 6585 3765 6600 3785
rect 6550 3735 6600 3765
rect 6550 3715 6565 3735
rect 6585 3715 6600 3735
rect 6550 3685 6600 3715
rect 6550 3665 6565 3685
rect 6585 3665 6600 3685
rect 6550 3635 6600 3665
rect 6550 3615 6565 3635
rect 6585 3615 6600 3635
rect 6550 3585 6600 3615
rect 6550 3565 6565 3585
rect 6585 3565 6600 3585
rect 6550 3535 6600 3565
rect 6550 3515 6565 3535
rect 6585 3515 6600 3535
rect 6550 3485 6600 3515
rect 6550 3465 6565 3485
rect 6585 3465 6600 3485
rect 6550 3435 6600 3465
rect 6550 3415 6565 3435
rect 6585 3415 6600 3435
rect 6550 3385 6600 3415
rect 6550 3365 6565 3385
rect 6585 3365 6600 3385
rect 6550 3335 6600 3365
rect 6550 3315 6565 3335
rect 6585 3315 6600 3335
rect 6550 3300 6600 3315
rect 6700 3785 6750 3800
rect 6700 3765 6715 3785
rect 6735 3765 6750 3785
rect 6700 3735 6750 3765
rect 6700 3715 6715 3735
rect 6735 3715 6750 3735
rect 6700 3685 6750 3715
rect 6700 3665 6715 3685
rect 6735 3665 6750 3685
rect 6700 3635 6750 3665
rect 6700 3615 6715 3635
rect 6735 3615 6750 3635
rect 6700 3585 6750 3615
rect 6700 3565 6715 3585
rect 6735 3565 6750 3585
rect 6700 3535 6750 3565
rect 6700 3515 6715 3535
rect 6735 3515 6750 3535
rect 6700 3485 6750 3515
rect 6700 3465 6715 3485
rect 6735 3465 6750 3485
rect 6700 3435 6750 3465
rect 6700 3415 6715 3435
rect 6735 3415 6750 3435
rect 6700 3385 6750 3415
rect 6700 3365 6715 3385
rect 6735 3365 6750 3385
rect 6700 3335 6750 3365
rect 6700 3315 6715 3335
rect 6735 3315 6750 3335
rect 6700 3300 6750 3315
rect 6850 3785 6900 3800
rect 6850 3765 6865 3785
rect 6885 3765 6900 3785
rect 6850 3735 6900 3765
rect 6850 3715 6865 3735
rect 6885 3715 6900 3735
rect 6850 3685 6900 3715
rect 6850 3665 6865 3685
rect 6885 3665 6900 3685
rect 6850 3635 6900 3665
rect 6850 3615 6865 3635
rect 6885 3615 6900 3635
rect 6850 3585 6900 3615
rect 6850 3565 6865 3585
rect 6885 3565 6900 3585
rect 6850 3535 6900 3565
rect 6850 3515 6865 3535
rect 6885 3515 6900 3535
rect 6850 3485 6900 3515
rect 6850 3465 6865 3485
rect 6885 3465 6900 3485
rect 6850 3435 6900 3465
rect 6850 3415 6865 3435
rect 6885 3415 6900 3435
rect 6850 3385 6900 3415
rect 6850 3365 6865 3385
rect 6885 3365 6900 3385
rect 6850 3335 6900 3365
rect 6850 3315 6865 3335
rect 6885 3315 6900 3335
rect 6850 3300 6900 3315
rect 7000 3785 7050 3800
rect 7000 3765 7015 3785
rect 7035 3765 7050 3785
rect 7000 3735 7050 3765
rect 7000 3715 7015 3735
rect 7035 3715 7050 3735
rect 7000 3685 7050 3715
rect 7000 3665 7015 3685
rect 7035 3665 7050 3685
rect 7000 3635 7050 3665
rect 7000 3615 7015 3635
rect 7035 3615 7050 3635
rect 7000 3585 7050 3615
rect 7000 3565 7015 3585
rect 7035 3565 7050 3585
rect 7000 3535 7050 3565
rect 7000 3515 7015 3535
rect 7035 3515 7050 3535
rect 7000 3485 7050 3515
rect 7000 3465 7015 3485
rect 7035 3465 7050 3485
rect 7000 3435 7050 3465
rect 7000 3415 7015 3435
rect 7035 3415 7050 3435
rect 7000 3385 7050 3415
rect 7000 3365 7015 3385
rect 7035 3365 7050 3385
rect 7000 3335 7050 3365
rect 7000 3315 7015 3335
rect 7035 3315 7050 3335
rect 7000 3300 7050 3315
rect 7150 3785 7200 3800
rect 7150 3765 7165 3785
rect 7185 3765 7200 3785
rect 7150 3735 7200 3765
rect 7150 3715 7165 3735
rect 7185 3715 7200 3735
rect 7150 3685 7200 3715
rect 7150 3665 7165 3685
rect 7185 3665 7200 3685
rect 7150 3635 7200 3665
rect 7150 3615 7165 3635
rect 7185 3615 7200 3635
rect 7150 3585 7200 3615
rect 7150 3565 7165 3585
rect 7185 3565 7200 3585
rect 7150 3535 7200 3565
rect 7150 3515 7165 3535
rect 7185 3515 7200 3535
rect 7150 3485 7200 3515
rect 7150 3465 7165 3485
rect 7185 3465 7200 3485
rect 7150 3435 7200 3465
rect 7150 3415 7165 3435
rect 7185 3415 7200 3435
rect 7150 3385 7200 3415
rect 7150 3365 7165 3385
rect 7185 3365 7200 3385
rect 7150 3335 7200 3365
rect 7150 3315 7165 3335
rect 7185 3315 7200 3335
rect 7150 3300 7200 3315
rect 7300 3785 7350 3800
rect 7300 3765 7315 3785
rect 7335 3765 7350 3785
rect 7300 3735 7350 3765
rect 7300 3715 7315 3735
rect 7335 3715 7350 3735
rect 7300 3685 7350 3715
rect 7300 3665 7315 3685
rect 7335 3665 7350 3685
rect 7300 3635 7350 3665
rect 7300 3615 7315 3635
rect 7335 3615 7350 3635
rect 7300 3585 7350 3615
rect 7300 3565 7315 3585
rect 7335 3565 7350 3585
rect 7300 3535 7350 3565
rect 7300 3515 7315 3535
rect 7335 3515 7350 3535
rect 7300 3485 7350 3515
rect 7300 3465 7315 3485
rect 7335 3465 7350 3485
rect 7300 3435 7350 3465
rect 7300 3415 7315 3435
rect 7335 3415 7350 3435
rect 7300 3385 7350 3415
rect 7300 3365 7315 3385
rect 7335 3365 7350 3385
rect 7300 3335 7350 3365
rect 7300 3315 7315 3335
rect 7335 3315 7350 3335
rect 7300 3300 7350 3315
rect 7450 3785 7500 3800
rect 7450 3765 7465 3785
rect 7485 3765 7500 3785
rect 7450 3735 7500 3765
rect 7450 3715 7465 3735
rect 7485 3715 7500 3735
rect 7450 3685 7500 3715
rect 7450 3665 7465 3685
rect 7485 3665 7500 3685
rect 7450 3635 7500 3665
rect 7450 3615 7465 3635
rect 7485 3615 7500 3635
rect 7450 3585 7500 3615
rect 7450 3565 7465 3585
rect 7485 3565 7500 3585
rect 7450 3535 7500 3565
rect 7450 3515 7465 3535
rect 7485 3515 7500 3535
rect 7450 3485 7500 3515
rect 7450 3465 7465 3485
rect 7485 3465 7500 3485
rect 7450 3435 7500 3465
rect 7450 3415 7465 3435
rect 7485 3415 7500 3435
rect 7450 3385 7500 3415
rect 7450 3365 7465 3385
rect 7485 3365 7500 3385
rect 7450 3335 7500 3365
rect 7450 3315 7465 3335
rect 7485 3315 7500 3335
rect 7450 3300 7500 3315
rect 7600 3785 7650 3800
rect 7600 3765 7615 3785
rect 7635 3765 7650 3785
rect 7600 3735 7650 3765
rect 7600 3715 7615 3735
rect 7635 3715 7650 3735
rect 7600 3685 7650 3715
rect 7600 3665 7615 3685
rect 7635 3665 7650 3685
rect 7600 3635 7650 3665
rect 7600 3615 7615 3635
rect 7635 3615 7650 3635
rect 7600 3585 7650 3615
rect 7600 3565 7615 3585
rect 7635 3565 7650 3585
rect 7600 3535 7650 3565
rect 7600 3515 7615 3535
rect 7635 3515 7650 3535
rect 7600 3485 7650 3515
rect 7600 3465 7615 3485
rect 7635 3465 7650 3485
rect 7600 3435 7650 3465
rect 7600 3415 7615 3435
rect 7635 3415 7650 3435
rect 7600 3385 7650 3415
rect 7600 3365 7615 3385
rect 7635 3365 7650 3385
rect 7600 3335 7650 3365
rect 7600 3315 7615 3335
rect 7635 3315 7650 3335
rect 7600 3300 7650 3315
rect 7750 3785 7800 3800
rect 7750 3765 7765 3785
rect 7785 3765 7800 3785
rect 7750 3735 7800 3765
rect 7750 3715 7765 3735
rect 7785 3715 7800 3735
rect 7750 3685 7800 3715
rect 7750 3665 7765 3685
rect 7785 3665 7800 3685
rect 7750 3635 7800 3665
rect 7750 3615 7765 3635
rect 7785 3615 7800 3635
rect 7750 3585 7800 3615
rect 7750 3565 7765 3585
rect 7785 3565 7800 3585
rect 7750 3535 7800 3565
rect 7750 3515 7765 3535
rect 7785 3515 7800 3535
rect 7750 3485 7800 3515
rect 7750 3465 7765 3485
rect 7785 3465 7800 3485
rect 7750 3435 7800 3465
rect 7750 3415 7765 3435
rect 7785 3415 7800 3435
rect 7750 3385 7800 3415
rect 7750 3365 7765 3385
rect 7785 3365 7800 3385
rect 7750 3335 7800 3365
rect 7750 3315 7765 3335
rect 7785 3315 7800 3335
rect 7750 3300 7800 3315
rect 7900 3300 7950 3800
rect 8050 3300 8100 3800
rect 8200 3300 8250 3800
rect 8350 3785 8400 3800
rect 8350 3765 8365 3785
rect 8385 3765 8400 3785
rect 8350 3735 8400 3765
rect 8350 3715 8365 3735
rect 8385 3715 8400 3735
rect 8350 3685 8400 3715
rect 8350 3665 8365 3685
rect 8385 3665 8400 3685
rect 8350 3635 8400 3665
rect 8350 3615 8365 3635
rect 8385 3615 8400 3635
rect 8350 3585 8400 3615
rect 8350 3565 8365 3585
rect 8385 3565 8400 3585
rect 8350 3535 8400 3565
rect 8350 3515 8365 3535
rect 8385 3515 8400 3535
rect 8350 3485 8400 3515
rect 8350 3465 8365 3485
rect 8385 3465 8400 3485
rect 8350 3435 8400 3465
rect 8350 3415 8365 3435
rect 8385 3415 8400 3435
rect 8350 3385 8400 3415
rect 8350 3365 8365 3385
rect 8385 3365 8400 3385
rect 8350 3335 8400 3365
rect 8350 3315 8365 3335
rect 8385 3315 8400 3335
rect 8350 3300 8400 3315
rect 8500 3785 8550 3800
rect 8500 3765 8515 3785
rect 8535 3765 8550 3785
rect 8500 3735 8550 3765
rect 8500 3715 8515 3735
rect 8535 3715 8550 3735
rect 8500 3685 8550 3715
rect 8500 3665 8515 3685
rect 8535 3665 8550 3685
rect 8500 3635 8550 3665
rect 8500 3615 8515 3635
rect 8535 3615 8550 3635
rect 8500 3585 8550 3615
rect 8500 3565 8515 3585
rect 8535 3565 8550 3585
rect 8500 3535 8550 3565
rect 8500 3515 8515 3535
rect 8535 3515 8550 3535
rect 8500 3485 8550 3515
rect 8500 3465 8515 3485
rect 8535 3465 8550 3485
rect 8500 3435 8550 3465
rect 8500 3415 8515 3435
rect 8535 3415 8550 3435
rect 8500 3385 8550 3415
rect 8500 3365 8515 3385
rect 8535 3365 8550 3385
rect 8500 3335 8550 3365
rect 8500 3315 8515 3335
rect 8535 3315 8550 3335
rect 8500 3300 8550 3315
rect 8650 3785 8700 3800
rect 8650 3765 8665 3785
rect 8685 3765 8700 3785
rect 8650 3735 8700 3765
rect 8650 3715 8665 3735
rect 8685 3715 8700 3735
rect 8650 3685 8700 3715
rect 8650 3665 8665 3685
rect 8685 3665 8700 3685
rect 8650 3635 8700 3665
rect 8650 3615 8665 3635
rect 8685 3615 8700 3635
rect 8650 3585 8700 3615
rect 8650 3565 8665 3585
rect 8685 3565 8700 3585
rect 8650 3535 8700 3565
rect 8650 3515 8665 3535
rect 8685 3515 8700 3535
rect 8650 3485 8700 3515
rect 8650 3465 8665 3485
rect 8685 3465 8700 3485
rect 8650 3435 8700 3465
rect 8650 3415 8665 3435
rect 8685 3415 8700 3435
rect 8650 3385 8700 3415
rect 8650 3365 8665 3385
rect 8685 3365 8700 3385
rect 8650 3335 8700 3365
rect 8650 3315 8665 3335
rect 8685 3315 8700 3335
rect 8650 3300 8700 3315
rect 8800 3785 8850 3800
rect 8800 3765 8815 3785
rect 8835 3765 8850 3785
rect 8800 3735 8850 3765
rect 8800 3715 8815 3735
rect 8835 3715 8850 3735
rect 8800 3685 8850 3715
rect 8800 3665 8815 3685
rect 8835 3665 8850 3685
rect 8800 3635 8850 3665
rect 8800 3615 8815 3635
rect 8835 3615 8850 3635
rect 8800 3585 8850 3615
rect 8800 3565 8815 3585
rect 8835 3565 8850 3585
rect 8800 3535 8850 3565
rect 8800 3515 8815 3535
rect 8835 3515 8850 3535
rect 8800 3485 8850 3515
rect 8800 3465 8815 3485
rect 8835 3465 8850 3485
rect 8800 3435 8850 3465
rect 8800 3415 8815 3435
rect 8835 3415 8850 3435
rect 8800 3385 8850 3415
rect 8800 3365 8815 3385
rect 8835 3365 8850 3385
rect 8800 3335 8850 3365
rect 8800 3315 8815 3335
rect 8835 3315 8850 3335
rect 8800 3300 8850 3315
rect 8950 3785 9000 3800
rect 8950 3765 8965 3785
rect 8985 3765 9000 3785
rect 8950 3735 9000 3765
rect 8950 3715 8965 3735
rect 8985 3715 9000 3735
rect 8950 3685 9000 3715
rect 8950 3665 8965 3685
rect 8985 3665 9000 3685
rect 8950 3635 9000 3665
rect 8950 3615 8965 3635
rect 8985 3615 9000 3635
rect 8950 3585 9000 3615
rect 8950 3565 8965 3585
rect 8985 3565 9000 3585
rect 8950 3535 9000 3565
rect 8950 3515 8965 3535
rect 8985 3515 9000 3535
rect 8950 3485 9000 3515
rect 8950 3465 8965 3485
rect 8985 3465 9000 3485
rect 8950 3435 9000 3465
rect 8950 3415 8965 3435
rect 8985 3415 9000 3435
rect 8950 3385 9000 3415
rect 8950 3365 8965 3385
rect 8985 3365 9000 3385
rect 8950 3335 9000 3365
rect 8950 3315 8965 3335
rect 8985 3315 9000 3335
rect 8950 3300 9000 3315
rect 9100 3785 9150 3800
rect 9100 3765 9115 3785
rect 9135 3765 9150 3785
rect 9100 3735 9150 3765
rect 9100 3715 9115 3735
rect 9135 3715 9150 3735
rect 9100 3685 9150 3715
rect 9100 3665 9115 3685
rect 9135 3665 9150 3685
rect 9100 3635 9150 3665
rect 9100 3615 9115 3635
rect 9135 3615 9150 3635
rect 9100 3585 9150 3615
rect 9100 3565 9115 3585
rect 9135 3565 9150 3585
rect 9100 3535 9150 3565
rect 9100 3515 9115 3535
rect 9135 3515 9150 3535
rect 9100 3485 9150 3515
rect 9100 3465 9115 3485
rect 9135 3465 9150 3485
rect 9100 3435 9150 3465
rect 9100 3415 9115 3435
rect 9135 3415 9150 3435
rect 9100 3385 9150 3415
rect 9100 3365 9115 3385
rect 9135 3365 9150 3385
rect 9100 3335 9150 3365
rect 9100 3315 9115 3335
rect 9135 3315 9150 3335
rect 9100 3300 9150 3315
rect 9250 3785 9300 3800
rect 9250 3765 9265 3785
rect 9285 3765 9300 3785
rect 9250 3735 9300 3765
rect 9250 3715 9265 3735
rect 9285 3715 9300 3735
rect 9250 3685 9300 3715
rect 9250 3665 9265 3685
rect 9285 3665 9300 3685
rect 9250 3635 9300 3665
rect 9250 3615 9265 3635
rect 9285 3615 9300 3635
rect 9250 3585 9300 3615
rect 9250 3565 9265 3585
rect 9285 3565 9300 3585
rect 9250 3535 9300 3565
rect 9250 3515 9265 3535
rect 9285 3515 9300 3535
rect 9250 3485 9300 3515
rect 9250 3465 9265 3485
rect 9285 3465 9300 3485
rect 9250 3435 9300 3465
rect 9250 3415 9265 3435
rect 9285 3415 9300 3435
rect 9250 3385 9300 3415
rect 9250 3365 9265 3385
rect 9285 3365 9300 3385
rect 9250 3335 9300 3365
rect 9250 3315 9265 3335
rect 9285 3315 9300 3335
rect 9250 3300 9300 3315
rect 9400 3785 9450 3800
rect 9400 3765 9415 3785
rect 9435 3765 9450 3785
rect 9400 3735 9450 3765
rect 9400 3715 9415 3735
rect 9435 3715 9450 3735
rect 9400 3685 9450 3715
rect 9400 3665 9415 3685
rect 9435 3665 9450 3685
rect 9400 3635 9450 3665
rect 9400 3615 9415 3635
rect 9435 3615 9450 3635
rect 9400 3585 9450 3615
rect 9400 3565 9415 3585
rect 9435 3565 9450 3585
rect 9400 3535 9450 3565
rect 9400 3515 9415 3535
rect 9435 3515 9450 3535
rect 9400 3485 9450 3515
rect 9400 3465 9415 3485
rect 9435 3465 9450 3485
rect 9400 3435 9450 3465
rect 9400 3415 9415 3435
rect 9435 3415 9450 3435
rect 9400 3385 9450 3415
rect 9400 3365 9415 3385
rect 9435 3365 9450 3385
rect 9400 3335 9450 3365
rect 9400 3315 9415 3335
rect 9435 3315 9450 3335
rect 9400 3300 9450 3315
rect 9550 3785 9600 3800
rect 9550 3765 9565 3785
rect 9585 3765 9600 3785
rect 9550 3735 9600 3765
rect 9550 3715 9565 3735
rect 9585 3715 9600 3735
rect 9550 3685 9600 3715
rect 9550 3665 9565 3685
rect 9585 3665 9600 3685
rect 9550 3635 9600 3665
rect 9550 3615 9565 3635
rect 9585 3615 9600 3635
rect 9550 3585 9600 3615
rect 9550 3565 9565 3585
rect 9585 3565 9600 3585
rect 9550 3535 9600 3565
rect 9550 3515 9565 3535
rect 9585 3515 9600 3535
rect 9550 3485 9600 3515
rect 9550 3465 9565 3485
rect 9585 3465 9600 3485
rect 9550 3435 9600 3465
rect 9550 3415 9565 3435
rect 9585 3415 9600 3435
rect 9550 3385 9600 3415
rect 9550 3365 9565 3385
rect 9585 3365 9600 3385
rect 9550 3335 9600 3365
rect 9550 3315 9565 3335
rect 9585 3315 9600 3335
rect 9550 3300 9600 3315
rect 9700 3785 9750 3800
rect 9700 3765 9715 3785
rect 9735 3765 9750 3785
rect 9700 3735 9750 3765
rect 9700 3715 9715 3735
rect 9735 3715 9750 3735
rect 9700 3685 9750 3715
rect 9700 3665 9715 3685
rect 9735 3665 9750 3685
rect 9700 3635 9750 3665
rect 9700 3615 9715 3635
rect 9735 3615 9750 3635
rect 9700 3585 9750 3615
rect 9700 3565 9715 3585
rect 9735 3565 9750 3585
rect 9700 3535 9750 3565
rect 9700 3515 9715 3535
rect 9735 3515 9750 3535
rect 9700 3485 9750 3515
rect 9700 3465 9715 3485
rect 9735 3465 9750 3485
rect 9700 3435 9750 3465
rect 9700 3415 9715 3435
rect 9735 3415 9750 3435
rect 9700 3385 9750 3415
rect 9700 3365 9715 3385
rect 9735 3365 9750 3385
rect 9700 3335 9750 3365
rect 9700 3315 9715 3335
rect 9735 3315 9750 3335
rect 9700 3300 9750 3315
rect 9850 3785 9900 3800
rect 9850 3765 9865 3785
rect 9885 3765 9900 3785
rect 9850 3735 9900 3765
rect 9850 3715 9865 3735
rect 9885 3715 9900 3735
rect 9850 3685 9900 3715
rect 9850 3665 9865 3685
rect 9885 3665 9900 3685
rect 9850 3635 9900 3665
rect 9850 3615 9865 3635
rect 9885 3615 9900 3635
rect 9850 3585 9900 3615
rect 9850 3565 9865 3585
rect 9885 3565 9900 3585
rect 9850 3535 9900 3565
rect 9850 3515 9865 3535
rect 9885 3515 9900 3535
rect 9850 3485 9900 3515
rect 9850 3465 9865 3485
rect 9885 3465 9900 3485
rect 9850 3435 9900 3465
rect 9850 3415 9865 3435
rect 9885 3415 9900 3435
rect 9850 3385 9900 3415
rect 9850 3365 9865 3385
rect 9885 3365 9900 3385
rect 9850 3335 9900 3365
rect 9850 3315 9865 3335
rect 9885 3315 9900 3335
rect 9850 3300 9900 3315
rect 10000 3785 10050 3800
rect 10000 3765 10015 3785
rect 10035 3765 10050 3785
rect 10000 3735 10050 3765
rect 10000 3715 10015 3735
rect 10035 3715 10050 3735
rect 10000 3685 10050 3715
rect 10000 3665 10015 3685
rect 10035 3665 10050 3685
rect 10000 3635 10050 3665
rect 10000 3615 10015 3635
rect 10035 3615 10050 3635
rect 10000 3585 10050 3615
rect 10000 3565 10015 3585
rect 10035 3565 10050 3585
rect 10000 3535 10050 3565
rect 10000 3515 10015 3535
rect 10035 3515 10050 3535
rect 10000 3485 10050 3515
rect 10000 3465 10015 3485
rect 10035 3465 10050 3485
rect 10000 3435 10050 3465
rect 10000 3415 10015 3435
rect 10035 3415 10050 3435
rect 10000 3385 10050 3415
rect 10000 3365 10015 3385
rect 10035 3365 10050 3385
rect 10000 3335 10050 3365
rect 10000 3315 10015 3335
rect 10035 3315 10050 3335
rect 10000 3300 10050 3315
rect 10150 3785 10200 3800
rect 10150 3765 10165 3785
rect 10185 3765 10200 3785
rect 10150 3735 10200 3765
rect 10150 3715 10165 3735
rect 10185 3715 10200 3735
rect 10150 3685 10200 3715
rect 10150 3665 10165 3685
rect 10185 3665 10200 3685
rect 10150 3635 10200 3665
rect 10150 3615 10165 3635
rect 10185 3615 10200 3635
rect 10150 3585 10200 3615
rect 10150 3565 10165 3585
rect 10185 3565 10200 3585
rect 10150 3535 10200 3565
rect 10150 3515 10165 3535
rect 10185 3515 10200 3535
rect 10150 3485 10200 3515
rect 10150 3465 10165 3485
rect 10185 3465 10200 3485
rect 10150 3435 10200 3465
rect 10150 3415 10165 3435
rect 10185 3415 10200 3435
rect 10150 3385 10200 3415
rect 10150 3365 10165 3385
rect 10185 3365 10200 3385
rect 10150 3335 10200 3365
rect 10150 3315 10165 3335
rect 10185 3315 10200 3335
rect 10150 3300 10200 3315
rect 10300 3785 10350 3800
rect 10300 3765 10315 3785
rect 10335 3765 10350 3785
rect 10300 3735 10350 3765
rect 10300 3715 10315 3735
rect 10335 3715 10350 3735
rect 10300 3685 10350 3715
rect 10300 3665 10315 3685
rect 10335 3665 10350 3685
rect 10300 3635 10350 3665
rect 10300 3615 10315 3635
rect 10335 3615 10350 3635
rect 10300 3585 10350 3615
rect 10300 3565 10315 3585
rect 10335 3565 10350 3585
rect 10300 3535 10350 3565
rect 10300 3515 10315 3535
rect 10335 3515 10350 3535
rect 10300 3485 10350 3515
rect 10300 3465 10315 3485
rect 10335 3465 10350 3485
rect 10300 3435 10350 3465
rect 10300 3415 10315 3435
rect 10335 3415 10350 3435
rect 10300 3385 10350 3415
rect 10300 3365 10315 3385
rect 10335 3365 10350 3385
rect 10300 3335 10350 3365
rect 10300 3315 10315 3335
rect 10335 3315 10350 3335
rect 10300 3300 10350 3315
rect 10450 3785 10500 3800
rect 10450 3765 10465 3785
rect 10485 3765 10500 3785
rect 10450 3735 10500 3765
rect 10450 3715 10465 3735
rect 10485 3715 10500 3735
rect 10450 3685 10500 3715
rect 10450 3665 10465 3685
rect 10485 3665 10500 3685
rect 10450 3635 10500 3665
rect 10450 3615 10465 3635
rect 10485 3615 10500 3635
rect 10450 3585 10500 3615
rect 10450 3565 10465 3585
rect 10485 3565 10500 3585
rect 10450 3535 10500 3565
rect 10450 3515 10465 3535
rect 10485 3515 10500 3535
rect 10450 3485 10500 3515
rect 10450 3465 10465 3485
rect 10485 3465 10500 3485
rect 10450 3435 10500 3465
rect 10450 3415 10465 3435
rect 10485 3415 10500 3435
rect 10450 3385 10500 3415
rect 10450 3365 10465 3385
rect 10485 3365 10500 3385
rect 10450 3335 10500 3365
rect 10450 3315 10465 3335
rect 10485 3315 10500 3335
rect 10450 3300 10500 3315
rect 10600 3785 10650 3800
rect 10600 3765 10615 3785
rect 10635 3765 10650 3785
rect 10600 3735 10650 3765
rect 10600 3715 10615 3735
rect 10635 3715 10650 3735
rect 10600 3685 10650 3715
rect 10600 3665 10615 3685
rect 10635 3665 10650 3685
rect 10600 3635 10650 3665
rect 10600 3615 10615 3635
rect 10635 3615 10650 3635
rect 10600 3585 10650 3615
rect 10600 3565 10615 3585
rect 10635 3565 10650 3585
rect 10600 3535 10650 3565
rect 10600 3515 10615 3535
rect 10635 3515 10650 3535
rect 10600 3485 10650 3515
rect 10600 3465 10615 3485
rect 10635 3465 10650 3485
rect 10600 3435 10650 3465
rect 10600 3415 10615 3435
rect 10635 3415 10650 3435
rect 10600 3385 10650 3415
rect 10600 3365 10615 3385
rect 10635 3365 10650 3385
rect 10600 3335 10650 3365
rect 10600 3315 10615 3335
rect 10635 3315 10650 3335
rect 10600 3300 10650 3315
rect 10750 3785 10800 3800
rect 10750 3765 10765 3785
rect 10785 3765 10800 3785
rect 10750 3735 10800 3765
rect 10750 3715 10765 3735
rect 10785 3715 10800 3735
rect 10750 3685 10800 3715
rect 10750 3665 10765 3685
rect 10785 3665 10800 3685
rect 10750 3635 10800 3665
rect 10750 3615 10765 3635
rect 10785 3615 10800 3635
rect 10750 3585 10800 3615
rect 10750 3565 10765 3585
rect 10785 3565 10800 3585
rect 10750 3535 10800 3565
rect 10750 3515 10765 3535
rect 10785 3515 10800 3535
rect 10750 3485 10800 3515
rect 10750 3465 10765 3485
rect 10785 3465 10800 3485
rect 10750 3435 10800 3465
rect 10750 3415 10765 3435
rect 10785 3415 10800 3435
rect 10750 3385 10800 3415
rect 10750 3365 10765 3385
rect 10785 3365 10800 3385
rect 10750 3335 10800 3365
rect 10750 3315 10765 3335
rect 10785 3315 10800 3335
rect 10750 3300 10800 3315
rect 10900 3300 10950 3800
rect 11050 3300 11100 3800
rect 11200 3300 11250 3800
rect 11350 3785 11400 3800
rect 11350 3765 11365 3785
rect 11385 3765 11400 3785
rect 11350 3735 11400 3765
rect 11350 3715 11365 3735
rect 11385 3715 11400 3735
rect 11350 3685 11400 3715
rect 11350 3665 11365 3685
rect 11385 3665 11400 3685
rect 11350 3635 11400 3665
rect 11350 3615 11365 3635
rect 11385 3615 11400 3635
rect 11350 3585 11400 3615
rect 11350 3565 11365 3585
rect 11385 3565 11400 3585
rect 11350 3535 11400 3565
rect 11350 3515 11365 3535
rect 11385 3515 11400 3535
rect 11350 3485 11400 3515
rect 11350 3465 11365 3485
rect 11385 3465 11400 3485
rect 11350 3435 11400 3465
rect 11350 3415 11365 3435
rect 11385 3415 11400 3435
rect 11350 3385 11400 3415
rect 11350 3365 11365 3385
rect 11385 3365 11400 3385
rect 11350 3335 11400 3365
rect 11350 3315 11365 3335
rect 11385 3315 11400 3335
rect 11350 3300 11400 3315
rect 11500 3300 11550 3800
rect 11650 3300 11700 3800
rect 11800 3300 11850 3800
rect 11950 3785 12000 3800
rect 11950 3765 11965 3785
rect 11985 3765 12000 3785
rect 11950 3735 12000 3765
rect 11950 3715 11965 3735
rect 11985 3715 12000 3735
rect 11950 3685 12000 3715
rect 11950 3665 11965 3685
rect 11985 3665 12000 3685
rect 11950 3635 12000 3665
rect 11950 3615 11965 3635
rect 11985 3615 12000 3635
rect 11950 3585 12000 3615
rect 11950 3565 11965 3585
rect 11985 3565 12000 3585
rect 11950 3535 12000 3565
rect 11950 3515 11965 3535
rect 11985 3515 12000 3535
rect 11950 3485 12000 3515
rect 11950 3465 11965 3485
rect 11985 3465 12000 3485
rect 11950 3435 12000 3465
rect 11950 3415 11965 3435
rect 11985 3415 12000 3435
rect 11950 3385 12000 3415
rect 11950 3365 11965 3385
rect 11985 3365 12000 3385
rect 11950 3335 12000 3365
rect 11950 3315 11965 3335
rect 11985 3315 12000 3335
rect 11950 3300 12000 3315
rect 12100 3300 12150 3800
rect 12250 3300 12300 3800
rect 12400 3300 12450 3800
rect 12550 3785 12600 3800
rect 12550 3765 12565 3785
rect 12585 3765 12600 3785
rect 12550 3735 12600 3765
rect 12550 3715 12565 3735
rect 12585 3715 12600 3735
rect 12550 3685 12600 3715
rect 12550 3665 12565 3685
rect 12585 3665 12600 3685
rect 12550 3635 12600 3665
rect 12550 3615 12565 3635
rect 12585 3615 12600 3635
rect 12550 3585 12600 3615
rect 12550 3565 12565 3585
rect 12585 3565 12600 3585
rect 12550 3535 12600 3565
rect 12550 3515 12565 3535
rect 12585 3515 12600 3535
rect 12550 3485 12600 3515
rect 12550 3465 12565 3485
rect 12585 3465 12600 3485
rect 12550 3435 12600 3465
rect 12550 3415 12565 3435
rect 12585 3415 12600 3435
rect 12550 3385 12600 3415
rect 12550 3365 12565 3385
rect 12585 3365 12600 3385
rect 12550 3335 12600 3365
rect 12550 3315 12565 3335
rect 12585 3315 12600 3335
rect 12550 3300 12600 3315
rect 12700 3300 12750 3800
rect 12850 3300 12900 3800
rect 13000 3300 13050 3800
rect 13150 3785 13200 3800
rect 13150 3765 13165 3785
rect 13185 3765 13200 3785
rect 13150 3735 13200 3765
rect 13150 3715 13165 3735
rect 13185 3715 13200 3735
rect 13150 3685 13200 3715
rect 13150 3665 13165 3685
rect 13185 3665 13200 3685
rect 13150 3635 13200 3665
rect 13150 3615 13165 3635
rect 13185 3615 13200 3635
rect 13150 3585 13200 3615
rect 13150 3565 13165 3585
rect 13185 3565 13200 3585
rect 13150 3535 13200 3565
rect 13150 3515 13165 3535
rect 13185 3515 13200 3535
rect 13150 3485 13200 3515
rect 13150 3465 13165 3485
rect 13185 3465 13200 3485
rect 13150 3435 13200 3465
rect 13150 3415 13165 3435
rect 13185 3415 13200 3435
rect 13150 3385 13200 3415
rect 13150 3365 13165 3385
rect 13185 3365 13200 3385
rect 13150 3335 13200 3365
rect 13150 3315 13165 3335
rect 13185 3315 13200 3335
rect 13150 3300 13200 3315
rect 13300 3300 13350 3800
rect 13450 3300 13500 3800
rect 13600 3300 13650 3800
rect 13750 3785 13800 3800
rect 13750 3765 13765 3785
rect 13785 3765 13800 3785
rect 13750 3735 13800 3765
rect 13750 3715 13765 3735
rect 13785 3715 13800 3735
rect 13750 3685 13800 3715
rect 13750 3665 13765 3685
rect 13785 3665 13800 3685
rect 13750 3635 13800 3665
rect 13750 3615 13765 3635
rect 13785 3615 13800 3635
rect 13750 3585 13800 3615
rect 13750 3565 13765 3585
rect 13785 3565 13800 3585
rect 13750 3535 13800 3565
rect 13750 3515 13765 3535
rect 13785 3515 13800 3535
rect 13750 3485 13800 3515
rect 13750 3465 13765 3485
rect 13785 3465 13800 3485
rect 13750 3435 13800 3465
rect 13750 3415 13765 3435
rect 13785 3415 13800 3435
rect 13750 3385 13800 3415
rect 13750 3365 13765 3385
rect 13785 3365 13800 3385
rect 13750 3335 13800 3365
rect 13750 3315 13765 3335
rect 13785 3315 13800 3335
rect 13750 3300 13800 3315
rect 13900 3300 13950 3800
rect 14050 3300 14100 3800
rect 14200 3300 14250 3800
rect 14350 3785 14400 3800
rect 14350 3765 14365 3785
rect 14385 3765 14400 3785
rect 14350 3735 14400 3765
rect 14350 3715 14365 3735
rect 14385 3715 14400 3735
rect 14350 3685 14400 3715
rect 14350 3665 14365 3685
rect 14385 3665 14400 3685
rect 14350 3635 14400 3665
rect 14350 3615 14365 3635
rect 14385 3615 14400 3635
rect 14350 3585 14400 3615
rect 14350 3565 14365 3585
rect 14385 3565 14400 3585
rect 14350 3535 14400 3565
rect 14350 3515 14365 3535
rect 14385 3515 14400 3535
rect 14350 3485 14400 3515
rect 14350 3465 14365 3485
rect 14385 3465 14400 3485
rect 14350 3435 14400 3465
rect 14350 3415 14365 3435
rect 14385 3415 14400 3435
rect 14350 3385 14400 3415
rect 14350 3365 14365 3385
rect 14385 3365 14400 3385
rect 14350 3335 14400 3365
rect 14350 3315 14365 3335
rect 14385 3315 14400 3335
rect 14350 3300 14400 3315
rect 14500 3300 14550 3800
rect 14650 3300 14700 3800
rect 14800 3300 14850 3800
rect 14950 3785 15000 3800
rect 14950 3765 14965 3785
rect 14985 3765 15000 3785
rect 14950 3735 15000 3765
rect 14950 3715 14965 3735
rect 14985 3715 15000 3735
rect 14950 3685 15000 3715
rect 14950 3665 14965 3685
rect 14985 3665 15000 3685
rect 14950 3635 15000 3665
rect 14950 3615 14965 3635
rect 14985 3615 15000 3635
rect 14950 3585 15000 3615
rect 14950 3565 14965 3585
rect 14985 3565 15000 3585
rect 14950 3535 15000 3565
rect 14950 3515 14965 3535
rect 14985 3515 15000 3535
rect 14950 3485 15000 3515
rect 14950 3465 14965 3485
rect 14985 3465 15000 3485
rect 14950 3435 15000 3465
rect 14950 3415 14965 3435
rect 14985 3415 15000 3435
rect 14950 3385 15000 3415
rect 14950 3365 14965 3385
rect 14985 3365 15000 3385
rect 14950 3335 15000 3365
rect 14950 3315 14965 3335
rect 14985 3315 15000 3335
rect 14950 3300 15000 3315
rect 15100 3300 15150 3800
rect 15250 3300 15300 3800
rect 15400 3300 15450 3800
rect 15550 3785 15600 3800
rect 15550 3765 15565 3785
rect 15585 3765 15600 3785
rect 15550 3735 15600 3765
rect 15550 3715 15565 3735
rect 15585 3715 15600 3735
rect 15550 3685 15600 3715
rect 15550 3665 15565 3685
rect 15585 3665 15600 3685
rect 15550 3635 15600 3665
rect 15550 3615 15565 3635
rect 15585 3615 15600 3635
rect 15550 3585 15600 3615
rect 15550 3565 15565 3585
rect 15585 3565 15600 3585
rect 15550 3535 15600 3565
rect 15550 3515 15565 3535
rect 15585 3515 15600 3535
rect 15550 3485 15600 3515
rect 15550 3465 15565 3485
rect 15585 3465 15600 3485
rect 15550 3435 15600 3465
rect 15550 3415 15565 3435
rect 15585 3415 15600 3435
rect 15550 3385 15600 3415
rect 15550 3365 15565 3385
rect 15585 3365 15600 3385
rect 15550 3335 15600 3365
rect 15550 3315 15565 3335
rect 15585 3315 15600 3335
rect 15550 3300 15600 3315
rect 15700 3300 15750 3800
rect 15850 3300 15900 3800
rect 16000 3300 16050 3800
rect 16150 3785 16200 3800
rect 16150 3765 16165 3785
rect 16185 3765 16200 3785
rect 16150 3735 16200 3765
rect 16150 3715 16165 3735
rect 16185 3715 16200 3735
rect 16150 3685 16200 3715
rect 16150 3665 16165 3685
rect 16185 3665 16200 3685
rect 16150 3635 16200 3665
rect 16150 3615 16165 3635
rect 16185 3615 16200 3635
rect 16150 3585 16200 3615
rect 16150 3565 16165 3585
rect 16185 3565 16200 3585
rect 16150 3535 16200 3565
rect 16150 3515 16165 3535
rect 16185 3515 16200 3535
rect 16150 3485 16200 3515
rect 16150 3465 16165 3485
rect 16185 3465 16200 3485
rect 16150 3435 16200 3465
rect 16150 3415 16165 3435
rect 16185 3415 16200 3435
rect 16150 3385 16200 3415
rect 16150 3365 16165 3385
rect 16185 3365 16200 3385
rect 16150 3335 16200 3365
rect 16150 3315 16165 3335
rect 16185 3315 16200 3335
rect 16150 3300 16200 3315
rect 16300 3785 16350 3800
rect 16300 3765 16315 3785
rect 16335 3765 16350 3785
rect 16300 3735 16350 3765
rect 16300 3715 16315 3735
rect 16335 3715 16350 3735
rect 16300 3685 16350 3715
rect 16300 3665 16315 3685
rect 16335 3665 16350 3685
rect 16300 3635 16350 3665
rect 16300 3615 16315 3635
rect 16335 3615 16350 3635
rect 16300 3585 16350 3615
rect 16300 3565 16315 3585
rect 16335 3565 16350 3585
rect 16300 3535 16350 3565
rect 16300 3515 16315 3535
rect 16335 3515 16350 3535
rect 16300 3485 16350 3515
rect 16300 3465 16315 3485
rect 16335 3465 16350 3485
rect 16300 3435 16350 3465
rect 16300 3415 16315 3435
rect 16335 3415 16350 3435
rect 16300 3385 16350 3415
rect 16300 3365 16315 3385
rect 16335 3365 16350 3385
rect 16300 3335 16350 3365
rect 16300 3315 16315 3335
rect 16335 3315 16350 3335
rect 16300 3300 16350 3315
rect 16450 3785 16500 3800
rect 16450 3765 16465 3785
rect 16485 3765 16500 3785
rect 16450 3735 16500 3765
rect 16450 3715 16465 3735
rect 16485 3715 16500 3735
rect 16450 3685 16500 3715
rect 16450 3665 16465 3685
rect 16485 3665 16500 3685
rect 16450 3635 16500 3665
rect 16450 3615 16465 3635
rect 16485 3615 16500 3635
rect 16450 3585 16500 3615
rect 16450 3565 16465 3585
rect 16485 3565 16500 3585
rect 16450 3535 16500 3565
rect 16450 3515 16465 3535
rect 16485 3515 16500 3535
rect 16450 3485 16500 3515
rect 16450 3465 16465 3485
rect 16485 3465 16500 3485
rect 16450 3435 16500 3465
rect 16450 3415 16465 3435
rect 16485 3415 16500 3435
rect 16450 3385 16500 3415
rect 16450 3365 16465 3385
rect 16485 3365 16500 3385
rect 16450 3335 16500 3365
rect 16450 3315 16465 3335
rect 16485 3315 16500 3335
rect 16450 3300 16500 3315
rect 16600 3785 16650 3800
rect 16600 3765 16615 3785
rect 16635 3765 16650 3785
rect 16600 3735 16650 3765
rect 16600 3715 16615 3735
rect 16635 3715 16650 3735
rect 16600 3685 16650 3715
rect 16600 3665 16615 3685
rect 16635 3665 16650 3685
rect 16600 3635 16650 3665
rect 16600 3615 16615 3635
rect 16635 3615 16650 3635
rect 16600 3585 16650 3615
rect 16600 3565 16615 3585
rect 16635 3565 16650 3585
rect 16600 3535 16650 3565
rect 16600 3515 16615 3535
rect 16635 3515 16650 3535
rect 16600 3485 16650 3515
rect 16600 3465 16615 3485
rect 16635 3465 16650 3485
rect 16600 3435 16650 3465
rect 16600 3415 16615 3435
rect 16635 3415 16650 3435
rect 16600 3385 16650 3415
rect 16600 3365 16615 3385
rect 16635 3365 16650 3385
rect 16600 3335 16650 3365
rect 16600 3315 16615 3335
rect 16635 3315 16650 3335
rect 16600 3300 16650 3315
rect 16750 3785 16800 3800
rect 16750 3765 16765 3785
rect 16785 3765 16800 3785
rect 16750 3735 16800 3765
rect 16750 3715 16765 3735
rect 16785 3715 16800 3735
rect 16750 3685 16800 3715
rect 16750 3665 16765 3685
rect 16785 3665 16800 3685
rect 16750 3635 16800 3665
rect 16750 3615 16765 3635
rect 16785 3615 16800 3635
rect 16750 3585 16800 3615
rect 16750 3565 16765 3585
rect 16785 3565 16800 3585
rect 16750 3535 16800 3565
rect 16750 3515 16765 3535
rect 16785 3515 16800 3535
rect 16750 3485 16800 3515
rect 16750 3465 16765 3485
rect 16785 3465 16800 3485
rect 16750 3435 16800 3465
rect 16750 3415 16765 3435
rect 16785 3415 16800 3435
rect 16750 3385 16800 3415
rect 16750 3365 16765 3385
rect 16785 3365 16800 3385
rect 16750 3335 16800 3365
rect 16750 3315 16765 3335
rect 16785 3315 16800 3335
rect 16750 3300 16800 3315
rect 16900 3785 16950 3800
rect 16900 3765 16915 3785
rect 16935 3765 16950 3785
rect 16900 3735 16950 3765
rect 16900 3715 16915 3735
rect 16935 3715 16950 3735
rect 16900 3685 16950 3715
rect 16900 3665 16915 3685
rect 16935 3665 16950 3685
rect 16900 3635 16950 3665
rect 16900 3615 16915 3635
rect 16935 3615 16950 3635
rect 16900 3585 16950 3615
rect 16900 3565 16915 3585
rect 16935 3565 16950 3585
rect 16900 3535 16950 3565
rect 16900 3515 16915 3535
rect 16935 3515 16950 3535
rect 16900 3485 16950 3515
rect 16900 3465 16915 3485
rect 16935 3465 16950 3485
rect 16900 3435 16950 3465
rect 16900 3415 16915 3435
rect 16935 3415 16950 3435
rect 16900 3385 16950 3415
rect 16900 3365 16915 3385
rect 16935 3365 16950 3385
rect 16900 3335 16950 3365
rect 16900 3315 16915 3335
rect 16935 3315 16950 3335
rect 16900 3300 16950 3315
rect 17050 3785 17100 3800
rect 17050 3765 17065 3785
rect 17085 3765 17100 3785
rect 17050 3735 17100 3765
rect 17050 3715 17065 3735
rect 17085 3715 17100 3735
rect 17050 3685 17100 3715
rect 17050 3665 17065 3685
rect 17085 3665 17100 3685
rect 17050 3635 17100 3665
rect 17050 3615 17065 3635
rect 17085 3615 17100 3635
rect 17050 3585 17100 3615
rect 17050 3565 17065 3585
rect 17085 3565 17100 3585
rect 17050 3535 17100 3565
rect 17050 3515 17065 3535
rect 17085 3515 17100 3535
rect 17050 3485 17100 3515
rect 17050 3465 17065 3485
rect 17085 3465 17100 3485
rect 17050 3435 17100 3465
rect 17050 3415 17065 3435
rect 17085 3415 17100 3435
rect 17050 3385 17100 3415
rect 17050 3365 17065 3385
rect 17085 3365 17100 3385
rect 17050 3335 17100 3365
rect 17050 3315 17065 3335
rect 17085 3315 17100 3335
rect 17050 3300 17100 3315
rect 17200 3785 17250 3800
rect 17200 3765 17215 3785
rect 17235 3765 17250 3785
rect 17200 3735 17250 3765
rect 17200 3715 17215 3735
rect 17235 3715 17250 3735
rect 17200 3685 17250 3715
rect 17200 3665 17215 3685
rect 17235 3665 17250 3685
rect 17200 3635 17250 3665
rect 17200 3615 17215 3635
rect 17235 3615 17250 3635
rect 17200 3585 17250 3615
rect 17200 3565 17215 3585
rect 17235 3565 17250 3585
rect 17200 3535 17250 3565
rect 17200 3515 17215 3535
rect 17235 3515 17250 3535
rect 17200 3485 17250 3515
rect 17200 3465 17215 3485
rect 17235 3465 17250 3485
rect 17200 3435 17250 3465
rect 17200 3415 17215 3435
rect 17235 3415 17250 3435
rect 17200 3385 17250 3415
rect 17200 3365 17215 3385
rect 17235 3365 17250 3385
rect 17200 3335 17250 3365
rect 17200 3315 17215 3335
rect 17235 3315 17250 3335
rect 17200 3300 17250 3315
rect 17350 3785 17400 3800
rect 17350 3765 17365 3785
rect 17385 3765 17400 3785
rect 17350 3735 17400 3765
rect 17350 3715 17365 3735
rect 17385 3715 17400 3735
rect 17350 3685 17400 3715
rect 17350 3665 17365 3685
rect 17385 3665 17400 3685
rect 17350 3635 17400 3665
rect 17350 3615 17365 3635
rect 17385 3615 17400 3635
rect 17350 3585 17400 3615
rect 17350 3565 17365 3585
rect 17385 3565 17400 3585
rect 17350 3535 17400 3565
rect 17350 3515 17365 3535
rect 17385 3515 17400 3535
rect 17350 3485 17400 3515
rect 17350 3465 17365 3485
rect 17385 3465 17400 3485
rect 17350 3435 17400 3465
rect 17350 3415 17365 3435
rect 17385 3415 17400 3435
rect 17350 3385 17400 3415
rect 17350 3365 17365 3385
rect 17385 3365 17400 3385
rect 17350 3335 17400 3365
rect 17350 3315 17365 3335
rect 17385 3315 17400 3335
rect 17350 3300 17400 3315
rect 17500 3300 17550 3800
rect 17650 3300 17700 3800
rect 17800 3300 17850 3800
rect 17950 3785 18000 3800
rect 17950 3765 17965 3785
rect 17985 3765 18000 3785
rect 17950 3735 18000 3765
rect 17950 3715 17965 3735
rect 17985 3715 18000 3735
rect 17950 3685 18000 3715
rect 17950 3665 17965 3685
rect 17985 3665 18000 3685
rect 17950 3635 18000 3665
rect 17950 3615 17965 3635
rect 17985 3615 18000 3635
rect 17950 3585 18000 3615
rect 17950 3565 17965 3585
rect 17985 3565 18000 3585
rect 17950 3535 18000 3565
rect 17950 3515 17965 3535
rect 17985 3515 18000 3535
rect 17950 3485 18000 3515
rect 17950 3465 17965 3485
rect 17985 3465 18000 3485
rect 17950 3435 18000 3465
rect 17950 3415 17965 3435
rect 17985 3415 18000 3435
rect 17950 3385 18000 3415
rect 17950 3365 17965 3385
rect 17985 3365 18000 3385
rect 17950 3335 18000 3365
rect 17950 3315 17965 3335
rect 17985 3315 18000 3335
rect 17950 3300 18000 3315
rect 18100 3300 18150 3800
rect 18250 3300 18300 3800
rect 18400 3300 18450 3800
rect 18550 3785 18600 3800
rect 18550 3765 18565 3785
rect 18585 3765 18600 3785
rect 18550 3735 18600 3765
rect 18550 3715 18565 3735
rect 18585 3715 18600 3735
rect 18550 3685 18600 3715
rect 18550 3665 18565 3685
rect 18585 3665 18600 3685
rect 18550 3635 18600 3665
rect 18550 3615 18565 3635
rect 18585 3615 18600 3635
rect 18550 3585 18600 3615
rect 18550 3565 18565 3585
rect 18585 3565 18600 3585
rect 18550 3535 18600 3565
rect 18550 3515 18565 3535
rect 18585 3515 18600 3535
rect 18550 3485 18600 3515
rect 18550 3465 18565 3485
rect 18585 3465 18600 3485
rect 18550 3435 18600 3465
rect 18550 3415 18565 3435
rect 18585 3415 18600 3435
rect 18550 3385 18600 3415
rect 18550 3365 18565 3385
rect 18585 3365 18600 3385
rect 18550 3335 18600 3365
rect 18550 3315 18565 3335
rect 18585 3315 18600 3335
rect 18550 3300 18600 3315
rect 18700 3785 18750 3800
rect 18700 3765 18715 3785
rect 18735 3765 18750 3785
rect 18700 3735 18750 3765
rect 18700 3715 18715 3735
rect 18735 3715 18750 3735
rect 18700 3685 18750 3715
rect 18700 3665 18715 3685
rect 18735 3665 18750 3685
rect 18700 3635 18750 3665
rect 18700 3615 18715 3635
rect 18735 3615 18750 3635
rect 18700 3585 18750 3615
rect 18700 3565 18715 3585
rect 18735 3565 18750 3585
rect 18700 3535 18750 3565
rect 18700 3515 18715 3535
rect 18735 3515 18750 3535
rect 18700 3485 18750 3515
rect 18700 3465 18715 3485
rect 18735 3465 18750 3485
rect 18700 3435 18750 3465
rect 18700 3415 18715 3435
rect 18735 3415 18750 3435
rect 18700 3385 18750 3415
rect 18700 3365 18715 3385
rect 18735 3365 18750 3385
rect 18700 3335 18750 3365
rect 18700 3315 18715 3335
rect 18735 3315 18750 3335
rect 18700 3300 18750 3315
rect 18850 3785 18900 3800
rect 18850 3765 18865 3785
rect 18885 3765 18900 3785
rect 18850 3735 18900 3765
rect 18850 3715 18865 3735
rect 18885 3715 18900 3735
rect 18850 3685 18900 3715
rect 18850 3665 18865 3685
rect 18885 3665 18900 3685
rect 18850 3635 18900 3665
rect 18850 3615 18865 3635
rect 18885 3615 18900 3635
rect 18850 3585 18900 3615
rect 18850 3565 18865 3585
rect 18885 3565 18900 3585
rect 18850 3535 18900 3565
rect 18850 3515 18865 3535
rect 18885 3515 18900 3535
rect 18850 3485 18900 3515
rect 18850 3465 18865 3485
rect 18885 3465 18900 3485
rect 18850 3435 18900 3465
rect 18850 3415 18865 3435
rect 18885 3415 18900 3435
rect 18850 3385 18900 3415
rect 18850 3365 18865 3385
rect 18885 3365 18900 3385
rect 18850 3335 18900 3365
rect 18850 3315 18865 3335
rect 18885 3315 18900 3335
rect 18850 3300 18900 3315
rect 19000 3785 19050 3800
rect 19000 3765 19015 3785
rect 19035 3765 19050 3785
rect 19000 3735 19050 3765
rect 19000 3715 19015 3735
rect 19035 3715 19050 3735
rect 19000 3685 19050 3715
rect 19000 3665 19015 3685
rect 19035 3665 19050 3685
rect 19000 3635 19050 3665
rect 19000 3615 19015 3635
rect 19035 3615 19050 3635
rect 19000 3585 19050 3615
rect 19000 3565 19015 3585
rect 19035 3565 19050 3585
rect 19000 3535 19050 3565
rect 19000 3515 19015 3535
rect 19035 3515 19050 3535
rect 19000 3485 19050 3515
rect 19000 3465 19015 3485
rect 19035 3465 19050 3485
rect 19000 3435 19050 3465
rect 19000 3415 19015 3435
rect 19035 3415 19050 3435
rect 19000 3385 19050 3415
rect 19000 3365 19015 3385
rect 19035 3365 19050 3385
rect 19000 3335 19050 3365
rect 19000 3315 19015 3335
rect 19035 3315 19050 3335
rect 19000 3300 19050 3315
rect 19150 3785 19200 3800
rect 19150 3765 19165 3785
rect 19185 3765 19200 3785
rect 19150 3735 19200 3765
rect 19150 3715 19165 3735
rect 19185 3715 19200 3735
rect 19150 3685 19200 3715
rect 19150 3665 19165 3685
rect 19185 3665 19200 3685
rect 19150 3635 19200 3665
rect 19150 3615 19165 3635
rect 19185 3615 19200 3635
rect 19150 3585 19200 3615
rect 19150 3565 19165 3585
rect 19185 3565 19200 3585
rect 19150 3535 19200 3565
rect 19150 3515 19165 3535
rect 19185 3515 19200 3535
rect 19150 3485 19200 3515
rect 19150 3465 19165 3485
rect 19185 3465 19200 3485
rect 19150 3435 19200 3465
rect 19150 3415 19165 3435
rect 19185 3415 19200 3435
rect 19150 3385 19200 3415
rect 19150 3365 19165 3385
rect 19185 3365 19200 3385
rect 19150 3335 19200 3365
rect 19150 3315 19165 3335
rect 19185 3315 19200 3335
rect 19150 3300 19200 3315
rect 19300 3785 19350 3800
rect 19300 3765 19315 3785
rect 19335 3765 19350 3785
rect 19300 3735 19350 3765
rect 19300 3715 19315 3735
rect 19335 3715 19350 3735
rect 19300 3685 19350 3715
rect 19300 3665 19315 3685
rect 19335 3665 19350 3685
rect 19300 3635 19350 3665
rect 19300 3615 19315 3635
rect 19335 3615 19350 3635
rect 19300 3585 19350 3615
rect 19300 3565 19315 3585
rect 19335 3565 19350 3585
rect 19300 3535 19350 3565
rect 19300 3515 19315 3535
rect 19335 3515 19350 3535
rect 19300 3485 19350 3515
rect 19300 3465 19315 3485
rect 19335 3465 19350 3485
rect 19300 3435 19350 3465
rect 19300 3415 19315 3435
rect 19335 3415 19350 3435
rect 19300 3385 19350 3415
rect 19300 3365 19315 3385
rect 19335 3365 19350 3385
rect 19300 3335 19350 3365
rect 19300 3315 19315 3335
rect 19335 3315 19350 3335
rect 19300 3300 19350 3315
rect 19450 3785 19500 3800
rect 19450 3765 19465 3785
rect 19485 3765 19500 3785
rect 19450 3735 19500 3765
rect 19450 3715 19465 3735
rect 19485 3715 19500 3735
rect 19450 3685 19500 3715
rect 19450 3665 19465 3685
rect 19485 3665 19500 3685
rect 19450 3635 19500 3665
rect 19450 3615 19465 3635
rect 19485 3615 19500 3635
rect 19450 3585 19500 3615
rect 19450 3565 19465 3585
rect 19485 3565 19500 3585
rect 19450 3535 19500 3565
rect 19450 3515 19465 3535
rect 19485 3515 19500 3535
rect 19450 3485 19500 3515
rect 19450 3465 19465 3485
rect 19485 3465 19500 3485
rect 19450 3435 19500 3465
rect 19450 3415 19465 3435
rect 19485 3415 19500 3435
rect 19450 3385 19500 3415
rect 19450 3365 19465 3385
rect 19485 3365 19500 3385
rect 19450 3335 19500 3365
rect 19450 3315 19465 3335
rect 19485 3315 19500 3335
rect 19450 3300 19500 3315
rect 19600 3785 19650 3800
rect 19600 3765 19615 3785
rect 19635 3765 19650 3785
rect 19600 3735 19650 3765
rect 19600 3715 19615 3735
rect 19635 3715 19650 3735
rect 19600 3685 19650 3715
rect 19600 3665 19615 3685
rect 19635 3665 19650 3685
rect 19600 3635 19650 3665
rect 19600 3615 19615 3635
rect 19635 3615 19650 3635
rect 19600 3585 19650 3615
rect 19600 3565 19615 3585
rect 19635 3565 19650 3585
rect 19600 3535 19650 3565
rect 19600 3515 19615 3535
rect 19635 3515 19650 3535
rect 19600 3485 19650 3515
rect 19600 3465 19615 3485
rect 19635 3465 19650 3485
rect 19600 3435 19650 3465
rect 19600 3415 19615 3435
rect 19635 3415 19650 3435
rect 19600 3385 19650 3415
rect 19600 3365 19615 3385
rect 19635 3365 19650 3385
rect 19600 3335 19650 3365
rect 19600 3315 19615 3335
rect 19635 3315 19650 3335
rect 19600 3300 19650 3315
rect 19750 3785 19800 3800
rect 19750 3765 19765 3785
rect 19785 3765 19800 3785
rect 19750 3735 19800 3765
rect 19750 3715 19765 3735
rect 19785 3715 19800 3735
rect 19750 3685 19800 3715
rect 19750 3665 19765 3685
rect 19785 3665 19800 3685
rect 19750 3635 19800 3665
rect 19750 3615 19765 3635
rect 19785 3615 19800 3635
rect 19750 3585 19800 3615
rect 19750 3565 19765 3585
rect 19785 3565 19800 3585
rect 19750 3535 19800 3565
rect 19750 3515 19765 3535
rect 19785 3515 19800 3535
rect 19750 3485 19800 3515
rect 19750 3465 19765 3485
rect 19785 3465 19800 3485
rect 19750 3435 19800 3465
rect 19750 3415 19765 3435
rect 19785 3415 19800 3435
rect 19750 3385 19800 3415
rect 19750 3365 19765 3385
rect 19785 3365 19800 3385
rect 19750 3335 19800 3365
rect 19750 3315 19765 3335
rect 19785 3315 19800 3335
rect 19750 3300 19800 3315
rect 19900 3300 19950 3800
rect 20050 3300 20100 3800
rect 20200 3300 20250 3800
rect 20350 3785 20400 3800
rect 20350 3765 20365 3785
rect 20385 3765 20400 3785
rect 20350 3735 20400 3765
rect 20350 3715 20365 3735
rect 20385 3715 20400 3735
rect 20350 3685 20400 3715
rect 20350 3665 20365 3685
rect 20385 3665 20400 3685
rect 20350 3635 20400 3665
rect 20350 3615 20365 3635
rect 20385 3615 20400 3635
rect 20350 3585 20400 3615
rect 20350 3565 20365 3585
rect 20385 3565 20400 3585
rect 20350 3535 20400 3565
rect 20350 3515 20365 3535
rect 20385 3515 20400 3535
rect 20350 3485 20400 3515
rect 20350 3465 20365 3485
rect 20385 3465 20400 3485
rect 20350 3435 20400 3465
rect 20350 3415 20365 3435
rect 20385 3415 20400 3435
rect 20350 3385 20400 3415
rect 20350 3365 20365 3385
rect 20385 3365 20400 3385
rect 20350 3335 20400 3365
rect 20350 3315 20365 3335
rect 20385 3315 20400 3335
rect 20350 3300 20400 3315
rect -650 3135 -600 3150
rect -650 3115 -635 3135
rect -615 3115 -600 3135
rect -650 3085 -600 3115
rect -650 3065 -635 3085
rect -615 3065 -600 3085
rect -650 3035 -600 3065
rect -650 3015 -635 3035
rect -615 3015 -600 3035
rect -650 2985 -600 3015
rect -650 2965 -635 2985
rect -615 2965 -600 2985
rect -650 2935 -600 2965
rect -650 2915 -635 2935
rect -615 2915 -600 2935
rect -650 2885 -600 2915
rect -650 2865 -635 2885
rect -615 2865 -600 2885
rect -650 2835 -600 2865
rect -650 2815 -635 2835
rect -615 2815 -600 2835
rect -650 2785 -600 2815
rect -650 2765 -635 2785
rect -615 2765 -600 2785
rect -650 2735 -600 2765
rect -650 2715 -635 2735
rect -615 2715 -600 2735
rect -650 2685 -600 2715
rect -650 2665 -635 2685
rect -615 2665 -600 2685
rect -650 2650 -600 2665
rect -500 3135 -450 3150
rect -500 3115 -485 3135
rect -465 3115 -450 3135
rect -500 3085 -450 3115
rect -500 3065 -485 3085
rect -465 3065 -450 3085
rect -500 3035 -450 3065
rect -500 3015 -485 3035
rect -465 3015 -450 3035
rect -500 2985 -450 3015
rect -500 2965 -485 2985
rect -465 2965 -450 2985
rect -500 2935 -450 2965
rect -500 2915 -485 2935
rect -465 2915 -450 2935
rect -500 2885 -450 2915
rect -500 2865 -485 2885
rect -465 2865 -450 2885
rect -500 2835 -450 2865
rect -500 2815 -485 2835
rect -465 2815 -450 2835
rect -500 2785 -450 2815
rect -500 2765 -485 2785
rect -465 2765 -450 2785
rect -500 2735 -450 2765
rect -500 2715 -485 2735
rect -465 2715 -450 2735
rect -500 2685 -450 2715
rect -500 2665 -485 2685
rect -465 2665 -450 2685
rect -500 2650 -450 2665
rect -350 3135 -300 3150
rect -350 3115 -335 3135
rect -315 3115 -300 3135
rect -350 3085 -300 3115
rect -350 3065 -335 3085
rect -315 3065 -300 3085
rect -350 3035 -300 3065
rect -350 3015 -335 3035
rect -315 3015 -300 3035
rect -350 2985 -300 3015
rect -350 2965 -335 2985
rect -315 2965 -300 2985
rect -350 2935 -300 2965
rect -350 2915 -335 2935
rect -315 2915 -300 2935
rect -350 2885 -300 2915
rect -350 2865 -335 2885
rect -315 2865 -300 2885
rect -350 2835 -300 2865
rect -350 2815 -335 2835
rect -315 2815 -300 2835
rect -350 2785 -300 2815
rect -350 2765 -335 2785
rect -315 2765 -300 2785
rect -350 2735 -300 2765
rect -350 2715 -335 2735
rect -315 2715 -300 2735
rect -350 2685 -300 2715
rect -350 2665 -335 2685
rect -315 2665 -300 2685
rect -350 2650 -300 2665
rect -200 3135 -150 3150
rect -200 3115 -185 3135
rect -165 3115 -150 3135
rect -200 3085 -150 3115
rect -200 3065 -185 3085
rect -165 3065 -150 3085
rect -200 3035 -150 3065
rect -200 3015 -185 3035
rect -165 3015 -150 3035
rect -200 2985 -150 3015
rect -200 2965 -185 2985
rect -165 2965 -150 2985
rect -200 2935 -150 2965
rect -200 2915 -185 2935
rect -165 2915 -150 2935
rect -200 2885 -150 2915
rect -200 2865 -185 2885
rect -165 2865 -150 2885
rect -200 2835 -150 2865
rect -200 2815 -185 2835
rect -165 2815 -150 2835
rect -200 2785 -150 2815
rect -200 2765 -185 2785
rect -165 2765 -150 2785
rect -200 2735 -150 2765
rect -200 2715 -185 2735
rect -165 2715 -150 2735
rect -200 2685 -150 2715
rect -200 2665 -185 2685
rect -165 2665 -150 2685
rect -200 2650 -150 2665
rect -50 3135 0 3150
rect -50 3115 -35 3135
rect -15 3115 0 3135
rect -50 3085 0 3115
rect -50 3065 -35 3085
rect -15 3065 0 3085
rect -50 3035 0 3065
rect -50 3015 -35 3035
rect -15 3015 0 3035
rect -50 2985 0 3015
rect -50 2965 -35 2985
rect -15 2965 0 2985
rect -50 2935 0 2965
rect -50 2915 -35 2935
rect -15 2915 0 2935
rect -50 2885 0 2915
rect -50 2865 -35 2885
rect -15 2865 0 2885
rect -50 2835 0 2865
rect -50 2815 -35 2835
rect -15 2815 0 2835
rect -50 2785 0 2815
rect -50 2765 -35 2785
rect -15 2765 0 2785
rect -50 2735 0 2765
rect -50 2715 -35 2735
rect -15 2715 0 2735
rect -50 2685 0 2715
rect -50 2665 -35 2685
rect -15 2665 0 2685
rect -50 2650 0 2665
rect 100 2650 150 3150
rect 250 2650 300 3150
rect 400 2650 450 3150
rect 550 3135 600 3150
rect 550 3115 565 3135
rect 585 3115 600 3135
rect 550 3085 600 3115
rect 550 3065 565 3085
rect 585 3065 600 3085
rect 550 3035 600 3065
rect 550 3015 565 3035
rect 585 3015 600 3035
rect 550 2985 600 3015
rect 550 2965 565 2985
rect 585 2965 600 2985
rect 550 2935 600 2965
rect 550 2915 565 2935
rect 585 2915 600 2935
rect 550 2885 600 2915
rect 550 2865 565 2885
rect 585 2865 600 2885
rect 550 2835 600 2865
rect 550 2815 565 2835
rect 585 2815 600 2835
rect 550 2785 600 2815
rect 550 2765 565 2785
rect 585 2765 600 2785
rect 550 2735 600 2765
rect 550 2715 565 2735
rect 585 2715 600 2735
rect 550 2685 600 2715
rect 550 2665 565 2685
rect 585 2665 600 2685
rect 550 2650 600 2665
rect 700 3135 750 3150
rect 700 3115 715 3135
rect 735 3115 750 3135
rect 700 3085 750 3115
rect 700 3065 715 3085
rect 735 3065 750 3085
rect 700 3035 750 3065
rect 700 3015 715 3035
rect 735 3015 750 3035
rect 700 2985 750 3015
rect 700 2965 715 2985
rect 735 2965 750 2985
rect 700 2935 750 2965
rect 700 2915 715 2935
rect 735 2915 750 2935
rect 700 2885 750 2915
rect 700 2865 715 2885
rect 735 2865 750 2885
rect 700 2835 750 2865
rect 700 2815 715 2835
rect 735 2815 750 2835
rect 700 2785 750 2815
rect 700 2765 715 2785
rect 735 2765 750 2785
rect 700 2735 750 2765
rect 700 2715 715 2735
rect 735 2715 750 2735
rect 700 2685 750 2715
rect 700 2665 715 2685
rect 735 2665 750 2685
rect 700 2650 750 2665
rect 850 3135 900 3150
rect 850 3115 865 3135
rect 885 3115 900 3135
rect 850 3085 900 3115
rect 850 3065 865 3085
rect 885 3065 900 3085
rect 850 3035 900 3065
rect 850 3015 865 3035
rect 885 3015 900 3035
rect 850 2985 900 3015
rect 850 2965 865 2985
rect 885 2965 900 2985
rect 850 2935 900 2965
rect 850 2915 865 2935
rect 885 2915 900 2935
rect 850 2885 900 2915
rect 850 2865 865 2885
rect 885 2865 900 2885
rect 850 2835 900 2865
rect 850 2815 865 2835
rect 885 2815 900 2835
rect 850 2785 900 2815
rect 850 2765 865 2785
rect 885 2765 900 2785
rect 850 2735 900 2765
rect 850 2715 865 2735
rect 885 2715 900 2735
rect 850 2685 900 2715
rect 850 2665 865 2685
rect 885 2665 900 2685
rect 850 2650 900 2665
rect 1000 3135 1050 3150
rect 1000 3115 1015 3135
rect 1035 3115 1050 3135
rect 1000 3085 1050 3115
rect 1000 3065 1015 3085
rect 1035 3065 1050 3085
rect 1000 3035 1050 3065
rect 1000 3015 1015 3035
rect 1035 3015 1050 3035
rect 1000 2985 1050 3015
rect 1000 2965 1015 2985
rect 1035 2965 1050 2985
rect 1000 2935 1050 2965
rect 1000 2915 1015 2935
rect 1035 2915 1050 2935
rect 1000 2885 1050 2915
rect 1000 2865 1015 2885
rect 1035 2865 1050 2885
rect 1000 2835 1050 2865
rect 1000 2815 1015 2835
rect 1035 2815 1050 2835
rect 1000 2785 1050 2815
rect 1000 2765 1015 2785
rect 1035 2765 1050 2785
rect 1000 2735 1050 2765
rect 1000 2715 1015 2735
rect 1035 2715 1050 2735
rect 1000 2685 1050 2715
rect 1000 2665 1015 2685
rect 1035 2665 1050 2685
rect 1000 2650 1050 2665
rect 1150 3135 1200 3150
rect 1150 3115 1165 3135
rect 1185 3115 1200 3135
rect 1150 3085 1200 3115
rect 1150 3065 1165 3085
rect 1185 3065 1200 3085
rect 1150 3035 1200 3065
rect 1150 3015 1165 3035
rect 1185 3015 1200 3035
rect 1150 2985 1200 3015
rect 1150 2965 1165 2985
rect 1185 2965 1200 2985
rect 1150 2935 1200 2965
rect 1150 2915 1165 2935
rect 1185 2915 1200 2935
rect 1150 2885 1200 2915
rect 1150 2865 1165 2885
rect 1185 2865 1200 2885
rect 1150 2835 1200 2865
rect 1150 2815 1165 2835
rect 1185 2815 1200 2835
rect 1150 2785 1200 2815
rect 1150 2765 1165 2785
rect 1185 2765 1200 2785
rect 1150 2735 1200 2765
rect 1150 2715 1165 2735
rect 1185 2715 1200 2735
rect 1150 2685 1200 2715
rect 1150 2665 1165 2685
rect 1185 2665 1200 2685
rect 1150 2650 1200 2665
rect 1300 3135 1350 3150
rect 1300 3115 1315 3135
rect 1335 3115 1350 3135
rect 1300 3085 1350 3115
rect 1300 3065 1315 3085
rect 1335 3065 1350 3085
rect 1300 3035 1350 3065
rect 1300 3015 1315 3035
rect 1335 3015 1350 3035
rect 1300 2985 1350 3015
rect 1300 2965 1315 2985
rect 1335 2965 1350 2985
rect 1300 2935 1350 2965
rect 1300 2915 1315 2935
rect 1335 2915 1350 2935
rect 1300 2885 1350 2915
rect 1300 2865 1315 2885
rect 1335 2865 1350 2885
rect 1300 2835 1350 2865
rect 1300 2815 1315 2835
rect 1335 2815 1350 2835
rect 1300 2785 1350 2815
rect 1300 2765 1315 2785
rect 1335 2765 1350 2785
rect 1300 2735 1350 2765
rect 1300 2715 1315 2735
rect 1335 2715 1350 2735
rect 1300 2685 1350 2715
rect 1300 2665 1315 2685
rect 1335 2665 1350 2685
rect 1300 2650 1350 2665
rect 1450 3135 1500 3150
rect 1450 3115 1465 3135
rect 1485 3115 1500 3135
rect 1450 3085 1500 3115
rect 1450 3065 1465 3085
rect 1485 3065 1500 3085
rect 1450 3035 1500 3065
rect 1450 3015 1465 3035
rect 1485 3015 1500 3035
rect 1450 2985 1500 3015
rect 1450 2965 1465 2985
rect 1485 2965 1500 2985
rect 1450 2935 1500 2965
rect 1450 2915 1465 2935
rect 1485 2915 1500 2935
rect 1450 2885 1500 2915
rect 1450 2865 1465 2885
rect 1485 2865 1500 2885
rect 1450 2835 1500 2865
rect 1450 2815 1465 2835
rect 1485 2815 1500 2835
rect 1450 2785 1500 2815
rect 1450 2765 1465 2785
rect 1485 2765 1500 2785
rect 1450 2735 1500 2765
rect 1450 2715 1465 2735
rect 1485 2715 1500 2735
rect 1450 2685 1500 2715
rect 1450 2665 1465 2685
rect 1485 2665 1500 2685
rect 1450 2650 1500 2665
rect 1600 3135 1650 3150
rect 1600 3115 1615 3135
rect 1635 3115 1650 3135
rect 1600 3085 1650 3115
rect 1600 3065 1615 3085
rect 1635 3065 1650 3085
rect 1600 3035 1650 3065
rect 1600 3015 1615 3035
rect 1635 3015 1650 3035
rect 1600 2985 1650 3015
rect 1600 2965 1615 2985
rect 1635 2965 1650 2985
rect 1600 2935 1650 2965
rect 1600 2915 1615 2935
rect 1635 2915 1650 2935
rect 1600 2885 1650 2915
rect 1600 2865 1615 2885
rect 1635 2865 1650 2885
rect 1600 2835 1650 2865
rect 1600 2815 1615 2835
rect 1635 2815 1650 2835
rect 1600 2785 1650 2815
rect 1600 2765 1615 2785
rect 1635 2765 1650 2785
rect 1600 2735 1650 2765
rect 1600 2715 1615 2735
rect 1635 2715 1650 2735
rect 1600 2685 1650 2715
rect 1600 2665 1615 2685
rect 1635 2665 1650 2685
rect 1600 2650 1650 2665
rect 1750 3135 1800 3150
rect 1750 3115 1765 3135
rect 1785 3115 1800 3135
rect 1750 3085 1800 3115
rect 1750 3065 1765 3085
rect 1785 3065 1800 3085
rect 1750 3035 1800 3065
rect 1750 3015 1765 3035
rect 1785 3015 1800 3035
rect 1750 2985 1800 3015
rect 1750 2965 1765 2985
rect 1785 2965 1800 2985
rect 1750 2935 1800 2965
rect 1750 2915 1765 2935
rect 1785 2915 1800 2935
rect 1750 2885 1800 2915
rect 1750 2865 1765 2885
rect 1785 2865 1800 2885
rect 1750 2835 1800 2865
rect 1750 2815 1765 2835
rect 1785 2815 1800 2835
rect 1750 2785 1800 2815
rect 1750 2765 1765 2785
rect 1785 2765 1800 2785
rect 1750 2735 1800 2765
rect 1750 2715 1765 2735
rect 1785 2715 1800 2735
rect 1750 2685 1800 2715
rect 1750 2665 1765 2685
rect 1785 2665 1800 2685
rect 1750 2650 1800 2665
rect 1900 3135 1950 3150
rect 1900 3115 1915 3135
rect 1935 3115 1950 3135
rect 1900 3085 1950 3115
rect 1900 3065 1915 3085
rect 1935 3065 1950 3085
rect 1900 3035 1950 3065
rect 1900 3015 1915 3035
rect 1935 3015 1950 3035
rect 1900 2985 1950 3015
rect 1900 2965 1915 2985
rect 1935 2965 1950 2985
rect 1900 2935 1950 2965
rect 1900 2915 1915 2935
rect 1935 2915 1950 2935
rect 1900 2885 1950 2915
rect 1900 2865 1915 2885
rect 1935 2865 1950 2885
rect 1900 2835 1950 2865
rect 1900 2815 1915 2835
rect 1935 2815 1950 2835
rect 1900 2785 1950 2815
rect 1900 2765 1915 2785
rect 1935 2765 1950 2785
rect 1900 2735 1950 2765
rect 1900 2715 1915 2735
rect 1935 2715 1950 2735
rect 1900 2685 1950 2715
rect 1900 2665 1915 2685
rect 1935 2665 1950 2685
rect 1900 2650 1950 2665
rect 2050 3135 2100 3150
rect 2050 3115 2065 3135
rect 2085 3115 2100 3135
rect 2050 3085 2100 3115
rect 2050 3065 2065 3085
rect 2085 3065 2100 3085
rect 2050 3035 2100 3065
rect 2050 3015 2065 3035
rect 2085 3015 2100 3035
rect 2050 2985 2100 3015
rect 2050 2965 2065 2985
rect 2085 2965 2100 2985
rect 2050 2935 2100 2965
rect 2050 2915 2065 2935
rect 2085 2915 2100 2935
rect 2050 2885 2100 2915
rect 2050 2865 2065 2885
rect 2085 2865 2100 2885
rect 2050 2835 2100 2865
rect 2050 2815 2065 2835
rect 2085 2815 2100 2835
rect 2050 2785 2100 2815
rect 2050 2765 2065 2785
rect 2085 2765 2100 2785
rect 2050 2735 2100 2765
rect 2050 2715 2065 2735
rect 2085 2715 2100 2735
rect 2050 2685 2100 2715
rect 2050 2665 2065 2685
rect 2085 2665 2100 2685
rect 2050 2650 2100 2665
rect 2200 3135 2250 3150
rect 2200 3115 2215 3135
rect 2235 3115 2250 3135
rect 2200 3085 2250 3115
rect 2200 3065 2215 3085
rect 2235 3065 2250 3085
rect 2200 3035 2250 3065
rect 2200 3015 2215 3035
rect 2235 3015 2250 3035
rect 2200 2985 2250 3015
rect 2200 2965 2215 2985
rect 2235 2965 2250 2985
rect 2200 2935 2250 2965
rect 2200 2915 2215 2935
rect 2235 2915 2250 2935
rect 2200 2885 2250 2915
rect 2200 2865 2215 2885
rect 2235 2865 2250 2885
rect 2200 2835 2250 2865
rect 2200 2815 2215 2835
rect 2235 2815 2250 2835
rect 2200 2785 2250 2815
rect 2200 2765 2215 2785
rect 2235 2765 2250 2785
rect 2200 2735 2250 2765
rect 2200 2715 2215 2735
rect 2235 2715 2250 2735
rect 2200 2685 2250 2715
rect 2200 2665 2215 2685
rect 2235 2665 2250 2685
rect 2200 2650 2250 2665
rect 2350 3135 2400 3150
rect 2350 3115 2365 3135
rect 2385 3115 2400 3135
rect 2350 3085 2400 3115
rect 2350 3065 2365 3085
rect 2385 3065 2400 3085
rect 2350 3035 2400 3065
rect 2350 3015 2365 3035
rect 2385 3015 2400 3035
rect 2350 2985 2400 3015
rect 2350 2965 2365 2985
rect 2385 2965 2400 2985
rect 2350 2935 2400 2965
rect 2350 2915 2365 2935
rect 2385 2915 2400 2935
rect 2350 2885 2400 2915
rect 2350 2865 2365 2885
rect 2385 2865 2400 2885
rect 2350 2835 2400 2865
rect 2350 2815 2365 2835
rect 2385 2815 2400 2835
rect 2350 2785 2400 2815
rect 2350 2765 2365 2785
rect 2385 2765 2400 2785
rect 2350 2735 2400 2765
rect 2350 2715 2365 2735
rect 2385 2715 2400 2735
rect 2350 2685 2400 2715
rect 2350 2665 2365 2685
rect 2385 2665 2400 2685
rect 2350 2650 2400 2665
rect 2500 3135 2550 3150
rect 2500 3115 2515 3135
rect 2535 3115 2550 3135
rect 2500 3085 2550 3115
rect 2500 3065 2515 3085
rect 2535 3065 2550 3085
rect 2500 3035 2550 3065
rect 2500 3015 2515 3035
rect 2535 3015 2550 3035
rect 2500 2985 2550 3015
rect 2500 2965 2515 2985
rect 2535 2965 2550 2985
rect 2500 2935 2550 2965
rect 2500 2915 2515 2935
rect 2535 2915 2550 2935
rect 2500 2885 2550 2915
rect 2500 2865 2515 2885
rect 2535 2865 2550 2885
rect 2500 2835 2550 2865
rect 2500 2815 2515 2835
rect 2535 2815 2550 2835
rect 2500 2785 2550 2815
rect 2500 2765 2515 2785
rect 2535 2765 2550 2785
rect 2500 2735 2550 2765
rect 2500 2715 2515 2735
rect 2535 2715 2550 2735
rect 2500 2685 2550 2715
rect 2500 2665 2515 2685
rect 2535 2665 2550 2685
rect 2500 2650 2550 2665
rect 2650 3135 2700 3150
rect 2650 3115 2665 3135
rect 2685 3115 2700 3135
rect 2650 3085 2700 3115
rect 2650 3065 2665 3085
rect 2685 3065 2700 3085
rect 2650 3035 2700 3065
rect 2650 3015 2665 3035
rect 2685 3015 2700 3035
rect 2650 2985 2700 3015
rect 2650 2965 2665 2985
rect 2685 2965 2700 2985
rect 2650 2935 2700 2965
rect 2650 2915 2665 2935
rect 2685 2915 2700 2935
rect 2650 2885 2700 2915
rect 2650 2865 2665 2885
rect 2685 2865 2700 2885
rect 2650 2835 2700 2865
rect 2650 2815 2665 2835
rect 2685 2815 2700 2835
rect 2650 2785 2700 2815
rect 2650 2765 2665 2785
rect 2685 2765 2700 2785
rect 2650 2735 2700 2765
rect 2650 2715 2665 2735
rect 2685 2715 2700 2735
rect 2650 2685 2700 2715
rect 2650 2665 2665 2685
rect 2685 2665 2700 2685
rect 2650 2650 2700 2665
rect 2800 3135 2850 3150
rect 2800 3115 2815 3135
rect 2835 3115 2850 3135
rect 2800 3085 2850 3115
rect 2800 3065 2815 3085
rect 2835 3065 2850 3085
rect 2800 3035 2850 3065
rect 2800 3015 2815 3035
rect 2835 3015 2850 3035
rect 2800 2985 2850 3015
rect 2800 2965 2815 2985
rect 2835 2965 2850 2985
rect 2800 2935 2850 2965
rect 2800 2915 2815 2935
rect 2835 2915 2850 2935
rect 2800 2885 2850 2915
rect 2800 2865 2815 2885
rect 2835 2865 2850 2885
rect 2800 2835 2850 2865
rect 2800 2815 2815 2835
rect 2835 2815 2850 2835
rect 2800 2785 2850 2815
rect 2800 2765 2815 2785
rect 2835 2765 2850 2785
rect 2800 2735 2850 2765
rect 2800 2715 2815 2735
rect 2835 2715 2850 2735
rect 2800 2685 2850 2715
rect 2800 2665 2815 2685
rect 2835 2665 2850 2685
rect 2800 2650 2850 2665
rect 2950 3135 3000 3150
rect 2950 3115 2965 3135
rect 2985 3115 3000 3135
rect 2950 3085 3000 3115
rect 2950 3065 2965 3085
rect 2985 3065 3000 3085
rect 2950 3035 3000 3065
rect 2950 3015 2965 3035
rect 2985 3015 3000 3035
rect 2950 2985 3000 3015
rect 2950 2965 2965 2985
rect 2985 2965 3000 2985
rect 2950 2935 3000 2965
rect 2950 2915 2965 2935
rect 2985 2915 3000 2935
rect 2950 2885 3000 2915
rect 2950 2865 2965 2885
rect 2985 2865 3000 2885
rect 2950 2835 3000 2865
rect 2950 2815 2965 2835
rect 2985 2815 3000 2835
rect 2950 2785 3000 2815
rect 2950 2765 2965 2785
rect 2985 2765 3000 2785
rect 2950 2735 3000 2765
rect 2950 2715 2965 2735
rect 2985 2715 3000 2735
rect 2950 2685 3000 2715
rect 2950 2665 2965 2685
rect 2985 2665 3000 2685
rect 2950 2650 3000 2665
rect 3100 3135 3150 3150
rect 3100 3115 3115 3135
rect 3135 3115 3150 3135
rect 3100 3085 3150 3115
rect 3100 3065 3115 3085
rect 3135 3065 3150 3085
rect 3100 3035 3150 3065
rect 3100 3015 3115 3035
rect 3135 3015 3150 3035
rect 3100 2985 3150 3015
rect 3100 2965 3115 2985
rect 3135 2965 3150 2985
rect 3100 2935 3150 2965
rect 3100 2915 3115 2935
rect 3135 2915 3150 2935
rect 3100 2885 3150 2915
rect 3100 2865 3115 2885
rect 3135 2865 3150 2885
rect 3100 2835 3150 2865
rect 3100 2815 3115 2835
rect 3135 2815 3150 2835
rect 3100 2785 3150 2815
rect 3100 2765 3115 2785
rect 3135 2765 3150 2785
rect 3100 2735 3150 2765
rect 3100 2715 3115 2735
rect 3135 2715 3150 2735
rect 3100 2685 3150 2715
rect 3100 2665 3115 2685
rect 3135 2665 3150 2685
rect 3100 2650 3150 2665
rect 3250 3135 3300 3150
rect 3250 3115 3265 3135
rect 3285 3115 3300 3135
rect 3250 3085 3300 3115
rect 3250 3065 3265 3085
rect 3285 3065 3300 3085
rect 3250 3035 3300 3065
rect 3250 3015 3265 3035
rect 3285 3015 3300 3035
rect 3250 2985 3300 3015
rect 3250 2965 3265 2985
rect 3285 2965 3300 2985
rect 3250 2935 3300 2965
rect 3250 2915 3265 2935
rect 3285 2915 3300 2935
rect 3250 2885 3300 2915
rect 3250 2865 3265 2885
rect 3285 2865 3300 2885
rect 3250 2835 3300 2865
rect 3250 2815 3265 2835
rect 3285 2815 3300 2835
rect 3250 2785 3300 2815
rect 3250 2765 3265 2785
rect 3285 2765 3300 2785
rect 3250 2735 3300 2765
rect 3250 2715 3265 2735
rect 3285 2715 3300 2735
rect 3250 2685 3300 2715
rect 3250 2665 3265 2685
rect 3285 2665 3300 2685
rect 3250 2650 3300 2665
rect 3400 3135 3450 3150
rect 3400 3115 3415 3135
rect 3435 3115 3450 3135
rect 3400 3085 3450 3115
rect 3400 3065 3415 3085
rect 3435 3065 3450 3085
rect 3400 3035 3450 3065
rect 3400 3015 3415 3035
rect 3435 3015 3450 3035
rect 3400 2985 3450 3015
rect 3400 2965 3415 2985
rect 3435 2965 3450 2985
rect 3400 2935 3450 2965
rect 3400 2915 3415 2935
rect 3435 2915 3450 2935
rect 3400 2885 3450 2915
rect 3400 2865 3415 2885
rect 3435 2865 3450 2885
rect 3400 2835 3450 2865
rect 3400 2815 3415 2835
rect 3435 2815 3450 2835
rect 3400 2785 3450 2815
rect 3400 2765 3415 2785
rect 3435 2765 3450 2785
rect 3400 2735 3450 2765
rect 3400 2715 3415 2735
rect 3435 2715 3450 2735
rect 3400 2685 3450 2715
rect 3400 2665 3415 2685
rect 3435 2665 3450 2685
rect 3400 2650 3450 2665
rect 3550 3135 3600 3150
rect 3550 3115 3565 3135
rect 3585 3115 3600 3135
rect 3550 3085 3600 3115
rect 3550 3065 3565 3085
rect 3585 3065 3600 3085
rect 3550 3035 3600 3065
rect 3550 3015 3565 3035
rect 3585 3015 3600 3035
rect 3550 2985 3600 3015
rect 3550 2965 3565 2985
rect 3585 2965 3600 2985
rect 3550 2935 3600 2965
rect 3550 2915 3565 2935
rect 3585 2915 3600 2935
rect 3550 2885 3600 2915
rect 3550 2865 3565 2885
rect 3585 2865 3600 2885
rect 3550 2835 3600 2865
rect 3550 2815 3565 2835
rect 3585 2815 3600 2835
rect 3550 2785 3600 2815
rect 3550 2765 3565 2785
rect 3585 2765 3600 2785
rect 3550 2735 3600 2765
rect 3550 2715 3565 2735
rect 3585 2715 3600 2735
rect 3550 2685 3600 2715
rect 3550 2665 3565 2685
rect 3585 2665 3600 2685
rect 3550 2650 3600 2665
rect 3700 2650 3750 3150
rect 3850 2650 3900 3150
rect 4000 2650 4050 3150
rect 4150 3135 4200 3150
rect 4150 3115 4165 3135
rect 4185 3115 4200 3135
rect 4150 3085 4200 3115
rect 4150 3065 4165 3085
rect 4185 3065 4200 3085
rect 4150 3035 4200 3065
rect 4150 3015 4165 3035
rect 4185 3015 4200 3035
rect 4150 2985 4200 3015
rect 4150 2965 4165 2985
rect 4185 2965 4200 2985
rect 4150 2935 4200 2965
rect 4150 2915 4165 2935
rect 4185 2915 4200 2935
rect 4150 2885 4200 2915
rect 4150 2865 4165 2885
rect 4185 2865 4200 2885
rect 4150 2835 4200 2865
rect 4150 2815 4165 2835
rect 4185 2815 4200 2835
rect 4150 2785 4200 2815
rect 4150 2765 4165 2785
rect 4185 2765 4200 2785
rect 4150 2735 4200 2765
rect 4150 2715 4165 2735
rect 4185 2715 4200 2735
rect 4150 2685 4200 2715
rect 4150 2665 4165 2685
rect 4185 2665 4200 2685
rect 4150 2650 4200 2665
rect 4300 2650 4350 3150
rect 4450 2650 4500 3150
rect 4600 2650 4650 3150
rect 4750 3135 4800 3150
rect 4750 3115 4765 3135
rect 4785 3115 4800 3135
rect 4750 3085 4800 3115
rect 4750 3065 4765 3085
rect 4785 3065 4800 3085
rect 4750 3035 4800 3065
rect 4750 3015 4765 3035
rect 4785 3015 4800 3035
rect 4750 2985 4800 3015
rect 4750 2965 4765 2985
rect 4785 2965 4800 2985
rect 4750 2935 4800 2965
rect 4750 2915 4765 2935
rect 4785 2915 4800 2935
rect 4750 2885 4800 2915
rect 4750 2865 4765 2885
rect 4785 2865 4800 2885
rect 4750 2835 4800 2865
rect 4750 2815 4765 2835
rect 4785 2815 4800 2835
rect 4750 2785 4800 2815
rect 4750 2765 4765 2785
rect 4785 2765 4800 2785
rect 4750 2735 4800 2765
rect 4750 2715 4765 2735
rect 4785 2715 4800 2735
rect 4750 2685 4800 2715
rect 4750 2665 4765 2685
rect 4785 2665 4800 2685
rect 4750 2650 4800 2665
rect 4900 3135 4950 3150
rect 4900 3115 4915 3135
rect 4935 3115 4950 3135
rect 4900 3085 4950 3115
rect 4900 3065 4915 3085
rect 4935 3065 4950 3085
rect 4900 3035 4950 3065
rect 4900 3015 4915 3035
rect 4935 3015 4950 3035
rect 4900 2985 4950 3015
rect 4900 2965 4915 2985
rect 4935 2965 4950 2985
rect 4900 2935 4950 2965
rect 4900 2915 4915 2935
rect 4935 2915 4950 2935
rect 4900 2885 4950 2915
rect 4900 2865 4915 2885
rect 4935 2865 4950 2885
rect 4900 2835 4950 2865
rect 4900 2815 4915 2835
rect 4935 2815 4950 2835
rect 4900 2785 4950 2815
rect 4900 2765 4915 2785
rect 4935 2765 4950 2785
rect 4900 2735 4950 2765
rect 4900 2715 4915 2735
rect 4935 2715 4950 2735
rect 4900 2685 4950 2715
rect 4900 2665 4915 2685
rect 4935 2665 4950 2685
rect 4900 2650 4950 2665
rect 5050 3135 5100 3150
rect 5050 3115 5065 3135
rect 5085 3115 5100 3135
rect 5050 3085 5100 3115
rect 5050 3065 5065 3085
rect 5085 3065 5100 3085
rect 5050 3035 5100 3065
rect 5050 3015 5065 3035
rect 5085 3015 5100 3035
rect 5050 2985 5100 3015
rect 5050 2965 5065 2985
rect 5085 2965 5100 2985
rect 5050 2935 5100 2965
rect 5050 2915 5065 2935
rect 5085 2915 5100 2935
rect 5050 2885 5100 2915
rect 5050 2865 5065 2885
rect 5085 2865 5100 2885
rect 5050 2835 5100 2865
rect 5050 2815 5065 2835
rect 5085 2815 5100 2835
rect 5050 2785 5100 2815
rect 5050 2765 5065 2785
rect 5085 2765 5100 2785
rect 5050 2735 5100 2765
rect 5050 2715 5065 2735
rect 5085 2715 5100 2735
rect 5050 2685 5100 2715
rect 5050 2665 5065 2685
rect 5085 2665 5100 2685
rect 5050 2650 5100 2665
rect 5200 3135 5250 3150
rect 5200 3115 5215 3135
rect 5235 3115 5250 3135
rect 5200 3085 5250 3115
rect 5200 3065 5215 3085
rect 5235 3065 5250 3085
rect 5200 3035 5250 3065
rect 5200 3015 5215 3035
rect 5235 3015 5250 3035
rect 5200 2985 5250 3015
rect 5200 2965 5215 2985
rect 5235 2965 5250 2985
rect 5200 2935 5250 2965
rect 5200 2915 5215 2935
rect 5235 2915 5250 2935
rect 5200 2885 5250 2915
rect 5200 2865 5215 2885
rect 5235 2865 5250 2885
rect 5200 2835 5250 2865
rect 5200 2815 5215 2835
rect 5235 2815 5250 2835
rect 5200 2785 5250 2815
rect 5200 2765 5215 2785
rect 5235 2765 5250 2785
rect 5200 2735 5250 2765
rect 5200 2715 5215 2735
rect 5235 2715 5250 2735
rect 5200 2685 5250 2715
rect 5200 2665 5215 2685
rect 5235 2665 5250 2685
rect 5200 2650 5250 2665
rect 5350 3135 5400 3150
rect 5350 3115 5365 3135
rect 5385 3115 5400 3135
rect 5350 3085 5400 3115
rect 5350 3065 5365 3085
rect 5385 3065 5400 3085
rect 5350 3035 5400 3065
rect 5350 3015 5365 3035
rect 5385 3015 5400 3035
rect 5350 2985 5400 3015
rect 5350 2965 5365 2985
rect 5385 2965 5400 2985
rect 5350 2935 5400 2965
rect 5350 2915 5365 2935
rect 5385 2915 5400 2935
rect 5350 2885 5400 2915
rect 5350 2865 5365 2885
rect 5385 2865 5400 2885
rect 5350 2835 5400 2865
rect 5350 2815 5365 2835
rect 5385 2815 5400 2835
rect 5350 2785 5400 2815
rect 5350 2765 5365 2785
rect 5385 2765 5400 2785
rect 5350 2735 5400 2765
rect 5350 2715 5365 2735
rect 5385 2715 5400 2735
rect 5350 2685 5400 2715
rect 5350 2665 5365 2685
rect 5385 2665 5400 2685
rect 5350 2650 5400 2665
rect 5500 3135 5550 3150
rect 5500 3115 5515 3135
rect 5535 3115 5550 3135
rect 5500 3085 5550 3115
rect 5500 3065 5515 3085
rect 5535 3065 5550 3085
rect 5500 3035 5550 3065
rect 5500 3015 5515 3035
rect 5535 3015 5550 3035
rect 5500 2985 5550 3015
rect 5500 2965 5515 2985
rect 5535 2965 5550 2985
rect 5500 2935 5550 2965
rect 5500 2915 5515 2935
rect 5535 2915 5550 2935
rect 5500 2885 5550 2915
rect 5500 2865 5515 2885
rect 5535 2865 5550 2885
rect 5500 2835 5550 2865
rect 5500 2815 5515 2835
rect 5535 2815 5550 2835
rect 5500 2785 5550 2815
rect 5500 2765 5515 2785
rect 5535 2765 5550 2785
rect 5500 2735 5550 2765
rect 5500 2715 5515 2735
rect 5535 2715 5550 2735
rect 5500 2685 5550 2715
rect 5500 2665 5515 2685
rect 5535 2665 5550 2685
rect 5500 2650 5550 2665
rect 5650 3135 5700 3150
rect 5650 3115 5665 3135
rect 5685 3115 5700 3135
rect 5650 3085 5700 3115
rect 5650 3065 5665 3085
rect 5685 3065 5700 3085
rect 5650 3035 5700 3065
rect 5650 3015 5665 3035
rect 5685 3015 5700 3035
rect 5650 2985 5700 3015
rect 5650 2965 5665 2985
rect 5685 2965 5700 2985
rect 5650 2935 5700 2965
rect 5650 2915 5665 2935
rect 5685 2915 5700 2935
rect 5650 2885 5700 2915
rect 5650 2865 5665 2885
rect 5685 2865 5700 2885
rect 5650 2835 5700 2865
rect 5650 2815 5665 2835
rect 5685 2815 5700 2835
rect 5650 2785 5700 2815
rect 5650 2765 5665 2785
rect 5685 2765 5700 2785
rect 5650 2735 5700 2765
rect 5650 2715 5665 2735
rect 5685 2715 5700 2735
rect 5650 2685 5700 2715
rect 5650 2665 5665 2685
rect 5685 2665 5700 2685
rect 5650 2650 5700 2665
rect 5800 3135 5850 3150
rect 5800 3115 5815 3135
rect 5835 3115 5850 3135
rect 5800 3085 5850 3115
rect 5800 3065 5815 3085
rect 5835 3065 5850 3085
rect 5800 3035 5850 3065
rect 5800 3015 5815 3035
rect 5835 3015 5850 3035
rect 5800 2985 5850 3015
rect 5800 2965 5815 2985
rect 5835 2965 5850 2985
rect 5800 2935 5850 2965
rect 5800 2915 5815 2935
rect 5835 2915 5850 2935
rect 5800 2885 5850 2915
rect 5800 2865 5815 2885
rect 5835 2865 5850 2885
rect 5800 2835 5850 2865
rect 5800 2815 5815 2835
rect 5835 2815 5850 2835
rect 5800 2785 5850 2815
rect 5800 2765 5815 2785
rect 5835 2765 5850 2785
rect 5800 2735 5850 2765
rect 5800 2715 5815 2735
rect 5835 2715 5850 2735
rect 5800 2685 5850 2715
rect 5800 2665 5815 2685
rect 5835 2665 5850 2685
rect 5800 2650 5850 2665
rect 5950 3135 6000 3150
rect 5950 3115 5965 3135
rect 5985 3115 6000 3135
rect 5950 3085 6000 3115
rect 5950 3065 5965 3085
rect 5985 3065 6000 3085
rect 5950 3035 6000 3065
rect 5950 3015 5965 3035
rect 5985 3015 6000 3035
rect 5950 2985 6000 3015
rect 5950 2965 5965 2985
rect 5985 2965 6000 2985
rect 5950 2935 6000 2965
rect 5950 2915 5965 2935
rect 5985 2915 6000 2935
rect 5950 2885 6000 2915
rect 5950 2865 5965 2885
rect 5985 2865 6000 2885
rect 5950 2835 6000 2865
rect 5950 2815 5965 2835
rect 5985 2815 6000 2835
rect 5950 2785 6000 2815
rect 5950 2765 5965 2785
rect 5985 2765 6000 2785
rect 5950 2735 6000 2765
rect 5950 2715 5965 2735
rect 5985 2715 6000 2735
rect 5950 2685 6000 2715
rect 5950 2665 5965 2685
rect 5985 2665 6000 2685
rect 5950 2650 6000 2665
rect 6100 3135 6150 3150
rect 6100 3115 6115 3135
rect 6135 3115 6150 3135
rect 6100 3085 6150 3115
rect 6100 3065 6115 3085
rect 6135 3065 6150 3085
rect 6100 3035 6150 3065
rect 6100 3015 6115 3035
rect 6135 3015 6150 3035
rect 6100 2985 6150 3015
rect 6100 2965 6115 2985
rect 6135 2965 6150 2985
rect 6100 2935 6150 2965
rect 6100 2915 6115 2935
rect 6135 2915 6150 2935
rect 6100 2885 6150 2915
rect 6100 2865 6115 2885
rect 6135 2865 6150 2885
rect 6100 2835 6150 2865
rect 6100 2815 6115 2835
rect 6135 2815 6150 2835
rect 6100 2785 6150 2815
rect 6100 2765 6115 2785
rect 6135 2765 6150 2785
rect 6100 2735 6150 2765
rect 6100 2715 6115 2735
rect 6135 2715 6150 2735
rect 6100 2685 6150 2715
rect 6100 2665 6115 2685
rect 6135 2665 6150 2685
rect 6100 2650 6150 2665
rect 6250 3135 6300 3150
rect 6250 3115 6265 3135
rect 6285 3115 6300 3135
rect 6250 3085 6300 3115
rect 6250 3065 6265 3085
rect 6285 3065 6300 3085
rect 6250 3035 6300 3065
rect 6250 3015 6265 3035
rect 6285 3015 6300 3035
rect 6250 2985 6300 3015
rect 6250 2965 6265 2985
rect 6285 2965 6300 2985
rect 6250 2935 6300 2965
rect 6250 2915 6265 2935
rect 6285 2915 6300 2935
rect 6250 2885 6300 2915
rect 6250 2865 6265 2885
rect 6285 2865 6300 2885
rect 6250 2835 6300 2865
rect 6250 2815 6265 2835
rect 6285 2815 6300 2835
rect 6250 2785 6300 2815
rect 6250 2765 6265 2785
rect 6285 2765 6300 2785
rect 6250 2735 6300 2765
rect 6250 2715 6265 2735
rect 6285 2715 6300 2735
rect 6250 2685 6300 2715
rect 6250 2665 6265 2685
rect 6285 2665 6300 2685
rect 6250 2650 6300 2665
rect 6400 3135 6450 3150
rect 6400 3115 6415 3135
rect 6435 3115 6450 3135
rect 6400 3085 6450 3115
rect 6400 3065 6415 3085
rect 6435 3065 6450 3085
rect 6400 3035 6450 3065
rect 6400 3015 6415 3035
rect 6435 3015 6450 3035
rect 6400 2985 6450 3015
rect 6400 2965 6415 2985
rect 6435 2965 6450 2985
rect 6400 2935 6450 2965
rect 6400 2915 6415 2935
rect 6435 2915 6450 2935
rect 6400 2885 6450 2915
rect 6400 2865 6415 2885
rect 6435 2865 6450 2885
rect 6400 2835 6450 2865
rect 6400 2815 6415 2835
rect 6435 2815 6450 2835
rect 6400 2785 6450 2815
rect 6400 2765 6415 2785
rect 6435 2765 6450 2785
rect 6400 2735 6450 2765
rect 6400 2715 6415 2735
rect 6435 2715 6450 2735
rect 6400 2685 6450 2715
rect 6400 2665 6415 2685
rect 6435 2665 6450 2685
rect 6400 2650 6450 2665
rect 6550 3135 6600 3150
rect 6550 3115 6565 3135
rect 6585 3115 6600 3135
rect 6550 3085 6600 3115
rect 6550 3065 6565 3085
rect 6585 3065 6600 3085
rect 6550 3035 6600 3065
rect 6550 3015 6565 3035
rect 6585 3015 6600 3035
rect 6550 2985 6600 3015
rect 6550 2965 6565 2985
rect 6585 2965 6600 2985
rect 6550 2935 6600 2965
rect 6550 2915 6565 2935
rect 6585 2915 6600 2935
rect 6550 2885 6600 2915
rect 6550 2865 6565 2885
rect 6585 2865 6600 2885
rect 6550 2835 6600 2865
rect 6550 2815 6565 2835
rect 6585 2815 6600 2835
rect 6550 2785 6600 2815
rect 6550 2765 6565 2785
rect 6585 2765 6600 2785
rect 6550 2735 6600 2765
rect 6550 2715 6565 2735
rect 6585 2715 6600 2735
rect 6550 2685 6600 2715
rect 6550 2665 6565 2685
rect 6585 2665 6600 2685
rect 6550 2650 6600 2665
rect 6700 3135 6750 3150
rect 6700 3115 6715 3135
rect 6735 3115 6750 3135
rect 6700 3085 6750 3115
rect 6700 3065 6715 3085
rect 6735 3065 6750 3085
rect 6700 3035 6750 3065
rect 6700 3015 6715 3035
rect 6735 3015 6750 3035
rect 6700 2985 6750 3015
rect 6700 2965 6715 2985
rect 6735 2965 6750 2985
rect 6700 2935 6750 2965
rect 6700 2915 6715 2935
rect 6735 2915 6750 2935
rect 6700 2885 6750 2915
rect 6700 2865 6715 2885
rect 6735 2865 6750 2885
rect 6700 2835 6750 2865
rect 6700 2815 6715 2835
rect 6735 2815 6750 2835
rect 6700 2785 6750 2815
rect 6700 2765 6715 2785
rect 6735 2765 6750 2785
rect 6700 2735 6750 2765
rect 6700 2715 6715 2735
rect 6735 2715 6750 2735
rect 6700 2685 6750 2715
rect 6700 2665 6715 2685
rect 6735 2665 6750 2685
rect 6700 2650 6750 2665
rect 6850 3135 6900 3150
rect 6850 3115 6865 3135
rect 6885 3115 6900 3135
rect 6850 3085 6900 3115
rect 6850 3065 6865 3085
rect 6885 3065 6900 3085
rect 6850 3035 6900 3065
rect 6850 3015 6865 3035
rect 6885 3015 6900 3035
rect 6850 2985 6900 3015
rect 6850 2965 6865 2985
rect 6885 2965 6900 2985
rect 6850 2935 6900 2965
rect 6850 2915 6865 2935
rect 6885 2915 6900 2935
rect 6850 2885 6900 2915
rect 6850 2865 6865 2885
rect 6885 2865 6900 2885
rect 6850 2835 6900 2865
rect 6850 2815 6865 2835
rect 6885 2815 6900 2835
rect 6850 2785 6900 2815
rect 6850 2765 6865 2785
rect 6885 2765 6900 2785
rect 6850 2735 6900 2765
rect 6850 2715 6865 2735
rect 6885 2715 6900 2735
rect 6850 2685 6900 2715
rect 6850 2665 6865 2685
rect 6885 2665 6900 2685
rect 6850 2650 6900 2665
rect 7000 3135 7050 3150
rect 7000 3115 7015 3135
rect 7035 3115 7050 3135
rect 7000 3085 7050 3115
rect 7000 3065 7015 3085
rect 7035 3065 7050 3085
rect 7000 3035 7050 3065
rect 7000 3015 7015 3035
rect 7035 3015 7050 3035
rect 7000 2985 7050 3015
rect 7000 2965 7015 2985
rect 7035 2965 7050 2985
rect 7000 2935 7050 2965
rect 7000 2915 7015 2935
rect 7035 2915 7050 2935
rect 7000 2885 7050 2915
rect 7000 2865 7015 2885
rect 7035 2865 7050 2885
rect 7000 2835 7050 2865
rect 7000 2815 7015 2835
rect 7035 2815 7050 2835
rect 7000 2785 7050 2815
rect 7000 2765 7015 2785
rect 7035 2765 7050 2785
rect 7000 2735 7050 2765
rect 7000 2715 7015 2735
rect 7035 2715 7050 2735
rect 7000 2685 7050 2715
rect 7000 2665 7015 2685
rect 7035 2665 7050 2685
rect 7000 2650 7050 2665
rect 7150 3135 7200 3150
rect 7150 3115 7165 3135
rect 7185 3115 7200 3135
rect 7150 3085 7200 3115
rect 7150 3065 7165 3085
rect 7185 3065 7200 3085
rect 7150 3035 7200 3065
rect 7150 3015 7165 3035
rect 7185 3015 7200 3035
rect 7150 2985 7200 3015
rect 7150 2965 7165 2985
rect 7185 2965 7200 2985
rect 7150 2935 7200 2965
rect 7150 2915 7165 2935
rect 7185 2915 7200 2935
rect 7150 2885 7200 2915
rect 7150 2865 7165 2885
rect 7185 2865 7200 2885
rect 7150 2835 7200 2865
rect 7150 2815 7165 2835
rect 7185 2815 7200 2835
rect 7150 2785 7200 2815
rect 7150 2765 7165 2785
rect 7185 2765 7200 2785
rect 7150 2735 7200 2765
rect 7150 2715 7165 2735
rect 7185 2715 7200 2735
rect 7150 2685 7200 2715
rect 7150 2665 7165 2685
rect 7185 2665 7200 2685
rect 7150 2650 7200 2665
rect 7300 3135 7350 3150
rect 7300 3115 7315 3135
rect 7335 3115 7350 3135
rect 7300 3085 7350 3115
rect 7300 3065 7315 3085
rect 7335 3065 7350 3085
rect 7300 3035 7350 3065
rect 7300 3015 7315 3035
rect 7335 3015 7350 3035
rect 7300 2985 7350 3015
rect 7300 2965 7315 2985
rect 7335 2965 7350 2985
rect 7300 2935 7350 2965
rect 7300 2915 7315 2935
rect 7335 2915 7350 2935
rect 7300 2885 7350 2915
rect 7300 2865 7315 2885
rect 7335 2865 7350 2885
rect 7300 2835 7350 2865
rect 7300 2815 7315 2835
rect 7335 2815 7350 2835
rect 7300 2785 7350 2815
rect 7300 2765 7315 2785
rect 7335 2765 7350 2785
rect 7300 2735 7350 2765
rect 7300 2715 7315 2735
rect 7335 2715 7350 2735
rect 7300 2685 7350 2715
rect 7300 2665 7315 2685
rect 7335 2665 7350 2685
rect 7300 2650 7350 2665
rect 7450 3135 7500 3150
rect 7450 3115 7465 3135
rect 7485 3115 7500 3135
rect 7450 3085 7500 3115
rect 7450 3065 7465 3085
rect 7485 3065 7500 3085
rect 7450 3035 7500 3065
rect 7450 3015 7465 3035
rect 7485 3015 7500 3035
rect 7450 2985 7500 3015
rect 7450 2965 7465 2985
rect 7485 2965 7500 2985
rect 7450 2935 7500 2965
rect 7450 2915 7465 2935
rect 7485 2915 7500 2935
rect 7450 2885 7500 2915
rect 7450 2865 7465 2885
rect 7485 2865 7500 2885
rect 7450 2835 7500 2865
rect 7450 2815 7465 2835
rect 7485 2815 7500 2835
rect 7450 2785 7500 2815
rect 7450 2765 7465 2785
rect 7485 2765 7500 2785
rect 7450 2735 7500 2765
rect 7450 2715 7465 2735
rect 7485 2715 7500 2735
rect 7450 2685 7500 2715
rect 7450 2665 7465 2685
rect 7485 2665 7500 2685
rect 7450 2650 7500 2665
rect 7600 3135 7650 3150
rect 7600 3115 7615 3135
rect 7635 3115 7650 3135
rect 7600 3085 7650 3115
rect 7600 3065 7615 3085
rect 7635 3065 7650 3085
rect 7600 3035 7650 3065
rect 7600 3015 7615 3035
rect 7635 3015 7650 3035
rect 7600 2985 7650 3015
rect 7600 2965 7615 2985
rect 7635 2965 7650 2985
rect 7600 2935 7650 2965
rect 7600 2915 7615 2935
rect 7635 2915 7650 2935
rect 7600 2885 7650 2915
rect 7600 2865 7615 2885
rect 7635 2865 7650 2885
rect 7600 2835 7650 2865
rect 7600 2815 7615 2835
rect 7635 2815 7650 2835
rect 7600 2785 7650 2815
rect 7600 2765 7615 2785
rect 7635 2765 7650 2785
rect 7600 2735 7650 2765
rect 7600 2715 7615 2735
rect 7635 2715 7650 2735
rect 7600 2685 7650 2715
rect 7600 2665 7615 2685
rect 7635 2665 7650 2685
rect 7600 2650 7650 2665
rect 7750 3135 7800 3150
rect 7750 3115 7765 3135
rect 7785 3115 7800 3135
rect 7750 3085 7800 3115
rect 7750 3065 7765 3085
rect 7785 3065 7800 3085
rect 7750 3035 7800 3065
rect 7750 3015 7765 3035
rect 7785 3015 7800 3035
rect 7750 2985 7800 3015
rect 7750 2965 7765 2985
rect 7785 2965 7800 2985
rect 7750 2935 7800 2965
rect 7750 2915 7765 2935
rect 7785 2915 7800 2935
rect 7750 2885 7800 2915
rect 7750 2865 7765 2885
rect 7785 2865 7800 2885
rect 7750 2835 7800 2865
rect 7750 2815 7765 2835
rect 7785 2815 7800 2835
rect 7750 2785 7800 2815
rect 7750 2765 7765 2785
rect 7785 2765 7800 2785
rect 7750 2735 7800 2765
rect 7750 2715 7765 2735
rect 7785 2715 7800 2735
rect 7750 2685 7800 2715
rect 7750 2665 7765 2685
rect 7785 2665 7800 2685
rect 7750 2650 7800 2665
rect 7900 2650 7950 3150
rect 8050 2650 8100 3150
rect 8200 2650 8250 3150
rect 8350 3135 8400 3150
rect 8350 3115 8365 3135
rect 8385 3115 8400 3135
rect 8350 3085 8400 3115
rect 8350 3065 8365 3085
rect 8385 3065 8400 3085
rect 8350 3035 8400 3065
rect 8350 3015 8365 3035
rect 8385 3015 8400 3035
rect 8350 2985 8400 3015
rect 8350 2965 8365 2985
rect 8385 2965 8400 2985
rect 8350 2935 8400 2965
rect 8350 2915 8365 2935
rect 8385 2915 8400 2935
rect 8350 2885 8400 2915
rect 8350 2865 8365 2885
rect 8385 2865 8400 2885
rect 8350 2835 8400 2865
rect 8350 2815 8365 2835
rect 8385 2815 8400 2835
rect 8350 2785 8400 2815
rect 8350 2765 8365 2785
rect 8385 2765 8400 2785
rect 8350 2735 8400 2765
rect 8350 2715 8365 2735
rect 8385 2715 8400 2735
rect 8350 2685 8400 2715
rect 8350 2665 8365 2685
rect 8385 2665 8400 2685
rect 8350 2650 8400 2665
rect 8500 3135 8550 3150
rect 8500 3115 8515 3135
rect 8535 3115 8550 3135
rect 8500 3085 8550 3115
rect 8500 3065 8515 3085
rect 8535 3065 8550 3085
rect 8500 3035 8550 3065
rect 8500 3015 8515 3035
rect 8535 3015 8550 3035
rect 8500 2985 8550 3015
rect 8500 2965 8515 2985
rect 8535 2965 8550 2985
rect 8500 2935 8550 2965
rect 8500 2915 8515 2935
rect 8535 2915 8550 2935
rect 8500 2885 8550 2915
rect 8500 2865 8515 2885
rect 8535 2865 8550 2885
rect 8500 2835 8550 2865
rect 8500 2815 8515 2835
rect 8535 2815 8550 2835
rect 8500 2785 8550 2815
rect 8500 2765 8515 2785
rect 8535 2765 8550 2785
rect 8500 2735 8550 2765
rect 8500 2715 8515 2735
rect 8535 2715 8550 2735
rect 8500 2685 8550 2715
rect 8500 2665 8515 2685
rect 8535 2665 8550 2685
rect 8500 2650 8550 2665
rect 8650 3135 8700 3150
rect 8650 3115 8665 3135
rect 8685 3115 8700 3135
rect 8650 3085 8700 3115
rect 8650 3065 8665 3085
rect 8685 3065 8700 3085
rect 8650 3035 8700 3065
rect 8650 3015 8665 3035
rect 8685 3015 8700 3035
rect 8650 2985 8700 3015
rect 8650 2965 8665 2985
rect 8685 2965 8700 2985
rect 8650 2935 8700 2965
rect 8650 2915 8665 2935
rect 8685 2915 8700 2935
rect 8650 2885 8700 2915
rect 8650 2865 8665 2885
rect 8685 2865 8700 2885
rect 8650 2835 8700 2865
rect 8650 2815 8665 2835
rect 8685 2815 8700 2835
rect 8650 2785 8700 2815
rect 8650 2765 8665 2785
rect 8685 2765 8700 2785
rect 8650 2735 8700 2765
rect 8650 2715 8665 2735
rect 8685 2715 8700 2735
rect 8650 2685 8700 2715
rect 8650 2665 8665 2685
rect 8685 2665 8700 2685
rect 8650 2650 8700 2665
rect 8800 3135 8850 3150
rect 8800 3115 8815 3135
rect 8835 3115 8850 3135
rect 8800 3085 8850 3115
rect 8800 3065 8815 3085
rect 8835 3065 8850 3085
rect 8800 3035 8850 3065
rect 8800 3015 8815 3035
rect 8835 3015 8850 3035
rect 8800 2985 8850 3015
rect 8800 2965 8815 2985
rect 8835 2965 8850 2985
rect 8800 2935 8850 2965
rect 8800 2915 8815 2935
rect 8835 2915 8850 2935
rect 8800 2885 8850 2915
rect 8800 2865 8815 2885
rect 8835 2865 8850 2885
rect 8800 2835 8850 2865
rect 8800 2815 8815 2835
rect 8835 2815 8850 2835
rect 8800 2785 8850 2815
rect 8800 2765 8815 2785
rect 8835 2765 8850 2785
rect 8800 2735 8850 2765
rect 8800 2715 8815 2735
rect 8835 2715 8850 2735
rect 8800 2685 8850 2715
rect 8800 2665 8815 2685
rect 8835 2665 8850 2685
rect 8800 2650 8850 2665
rect 8950 3135 9000 3150
rect 8950 3115 8965 3135
rect 8985 3115 9000 3135
rect 8950 3085 9000 3115
rect 8950 3065 8965 3085
rect 8985 3065 9000 3085
rect 8950 3035 9000 3065
rect 8950 3015 8965 3035
rect 8985 3015 9000 3035
rect 8950 2985 9000 3015
rect 8950 2965 8965 2985
rect 8985 2965 9000 2985
rect 8950 2935 9000 2965
rect 8950 2915 8965 2935
rect 8985 2915 9000 2935
rect 8950 2885 9000 2915
rect 8950 2865 8965 2885
rect 8985 2865 9000 2885
rect 8950 2835 9000 2865
rect 8950 2815 8965 2835
rect 8985 2815 9000 2835
rect 8950 2785 9000 2815
rect 8950 2765 8965 2785
rect 8985 2765 9000 2785
rect 8950 2735 9000 2765
rect 8950 2715 8965 2735
rect 8985 2715 9000 2735
rect 8950 2685 9000 2715
rect 8950 2665 8965 2685
rect 8985 2665 9000 2685
rect 8950 2650 9000 2665
rect 9100 3135 9150 3150
rect 9100 3115 9115 3135
rect 9135 3115 9150 3135
rect 9100 3085 9150 3115
rect 9100 3065 9115 3085
rect 9135 3065 9150 3085
rect 9100 3035 9150 3065
rect 9100 3015 9115 3035
rect 9135 3015 9150 3035
rect 9100 2985 9150 3015
rect 9100 2965 9115 2985
rect 9135 2965 9150 2985
rect 9100 2935 9150 2965
rect 9100 2915 9115 2935
rect 9135 2915 9150 2935
rect 9100 2885 9150 2915
rect 9100 2865 9115 2885
rect 9135 2865 9150 2885
rect 9100 2835 9150 2865
rect 9100 2815 9115 2835
rect 9135 2815 9150 2835
rect 9100 2785 9150 2815
rect 9100 2765 9115 2785
rect 9135 2765 9150 2785
rect 9100 2735 9150 2765
rect 9100 2715 9115 2735
rect 9135 2715 9150 2735
rect 9100 2685 9150 2715
rect 9100 2665 9115 2685
rect 9135 2665 9150 2685
rect 9100 2650 9150 2665
rect 9250 3135 9300 3150
rect 9250 3115 9265 3135
rect 9285 3115 9300 3135
rect 9250 3085 9300 3115
rect 9250 3065 9265 3085
rect 9285 3065 9300 3085
rect 9250 3035 9300 3065
rect 9250 3015 9265 3035
rect 9285 3015 9300 3035
rect 9250 2985 9300 3015
rect 9250 2965 9265 2985
rect 9285 2965 9300 2985
rect 9250 2935 9300 2965
rect 9250 2915 9265 2935
rect 9285 2915 9300 2935
rect 9250 2885 9300 2915
rect 9250 2865 9265 2885
rect 9285 2865 9300 2885
rect 9250 2835 9300 2865
rect 9250 2815 9265 2835
rect 9285 2815 9300 2835
rect 9250 2785 9300 2815
rect 9250 2765 9265 2785
rect 9285 2765 9300 2785
rect 9250 2735 9300 2765
rect 9250 2715 9265 2735
rect 9285 2715 9300 2735
rect 9250 2685 9300 2715
rect 9250 2665 9265 2685
rect 9285 2665 9300 2685
rect 9250 2650 9300 2665
rect 9400 3135 9450 3150
rect 9400 3115 9415 3135
rect 9435 3115 9450 3135
rect 9400 3085 9450 3115
rect 9400 3065 9415 3085
rect 9435 3065 9450 3085
rect 9400 3035 9450 3065
rect 9400 3015 9415 3035
rect 9435 3015 9450 3035
rect 9400 2985 9450 3015
rect 9400 2965 9415 2985
rect 9435 2965 9450 2985
rect 9400 2935 9450 2965
rect 9400 2915 9415 2935
rect 9435 2915 9450 2935
rect 9400 2885 9450 2915
rect 9400 2865 9415 2885
rect 9435 2865 9450 2885
rect 9400 2835 9450 2865
rect 9400 2815 9415 2835
rect 9435 2815 9450 2835
rect 9400 2785 9450 2815
rect 9400 2765 9415 2785
rect 9435 2765 9450 2785
rect 9400 2735 9450 2765
rect 9400 2715 9415 2735
rect 9435 2715 9450 2735
rect 9400 2685 9450 2715
rect 9400 2665 9415 2685
rect 9435 2665 9450 2685
rect 9400 2650 9450 2665
rect 9550 3135 9600 3150
rect 9550 3115 9565 3135
rect 9585 3115 9600 3135
rect 9550 3085 9600 3115
rect 9550 3065 9565 3085
rect 9585 3065 9600 3085
rect 9550 3035 9600 3065
rect 9550 3015 9565 3035
rect 9585 3015 9600 3035
rect 9550 2985 9600 3015
rect 9550 2965 9565 2985
rect 9585 2965 9600 2985
rect 9550 2935 9600 2965
rect 9550 2915 9565 2935
rect 9585 2915 9600 2935
rect 9550 2885 9600 2915
rect 9550 2865 9565 2885
rect 9585 2865 9600 2885
rect 9550 2835 9600 2865
rect 9550 2815 9565 2835
rect 9585 2815 9600 2835
rect 9550 2785 9600 2815
rect 9550 2765 9565 2785
rect 9585 2765 9600 2785
rect 9550 2735 9600 2765
rect 9550 2715 9565 2735
rect 9585 2715 9600 2735
rect 9550 2685 9600 2715
rect 9550 2665 9565 2685
rect 9585 2665 9600 2685
rect 9550 2650 9600 2665
rect 9700 3135 9750 3150
rect 9700 3115 9715 3135
rect 9735 3115 9750 3135
rect 9700 3085 9750 3115
rect 9700 3065 9715 3085
rect 9735 3065 9750 3085
rect 9700 3035 9750 3065
rect 9700 3015 9715 3035
rect 9735 3015 9750 3035
rect 9700 2985 9750 3015
rect 9700 2965 9715 2985
rect 9735 2965 9750 2985
rect 9700 2935 9750 2965
rect 9700 2915 9715 2935
rect 9735 2915 9750 2935
rect 9700 2885 9750 2915
rect 9700 2865 9715 2885
rect 9735 2865 9750 2885
rect 9700 2835 9750 2865
rect 9700 2815 9715 2835
rect 9735 2815 9750 2835
rect 9700 2785 9750 2815
rect 9700 2765 9715 2785
rect 9735 2765 9750 2785
rect 9700 2735 9750 2765
rect 9700 2715 9715 2735
rect 9735 2715 9750 2735
rect 9700 2685 9750 2715
rect 9700 2665 9715 2685
rect 9735 2665 9750 2685
rect 9700 2650 9750 2665
rect 9850 3135 9900 3150
rect 9850 3115 9865 3135
rect 9885 3115 9900 3135
rect 9850 3085 9900 3115
rect 9850 3065 9865 3085
rect 9885 3065 9900 3085
rect 9850 3035 9900 3065
rect 9850 3015 9865 3035
rect 9885 3015 9900 3035
rect 9850 2985 9900 3015
rect 9850 2965 9865 2985
rect 9885 2965 9900 2985
rect 9850 2935 9900 2965
rect 9850 2915 9865 2935
rect 9885 2915 9900 2935
rect 9850 2885 9900 2915
rect 9850 2865 9865 2885
rect 9885 2865 9900 2885
rect 9850 2835 9900 2865
rect 9850 2815 9865 2835
rect 9885 2815 9900 2835
rect 9850 2785 9900 2815
rect 9850 2765 9865 2785
rect 9885 2765 9900 2785
rect 9850 2735 9900 2765
rect 9850 2715 9865 2735
rect 9885 2715 9900 2735
rect 9850 2685 9900 2715
rect 9850 2665 9865 2685
rect 9885 2665 9900 2685
rect 9850 2650 9900 2665
rect 10000 3135 10050 3150
rect 10000 3115 10015 3135
rect 10035 3115 10050 3135
rect 10000 3085 10050 3115
rect 10000 3065 10015 3085
rect 10035 3065 10050 3085
rect 10000 3035 10050 3065
rect 10000 3015 10015 3035
rect 10035 3015 10050 3035
rect 10000 2985 10050 3015
rect 10000 2965 10015 2985
rect 10035 2965 10050 2985
rect 10000 2935 10050 2965
rect 10000 2915 10015 2935
rect 10035 2915 10050 2935
rect 10000 2885 10050 2915
rect 10000 2865 10015 2885
rect 10035 2865 10050 2885
rect 10000 2835 10050 2865
rect 10000 2815 10015 2835
rect 10035 2815 10050 2835
rect 10000 2785 10050 2815
rect 10000 2765 10015 2785
rect 10035 2765 10050 2785
rect 10000 2735 10050 2765
rect 10000 2715 10015 2735
rect 10035 2715 10050 2735
rect 10000 2685 10050 2715
rect 10000 2665 10015 2685
rect 10035 2665 10050 2685
rect 10000 2650 10050 2665
rect 10150 3135 10200 3150
rect 10150 3115 10165 3135
rect 10185 3115 10200 3135
rect 10150 3085 10200 3115
rect 10150 3065 10165 3085
rect 10185 3065 10200 3085
rect 10150 3035 10200 3065
rect 10150 3015 10165 3035
rect 10185 3015 10200 3035
rect 10150 2985 10200 3015
rect 10150 2965 10165 2985
rect 10185 2965 10200 2985
rect 10150 2935 10200 2965
rect 10150 2915 10165 2935
rect 10185 2915 10200 2935
rect 10150 2885 10200 2915
rect 10150 2865 10165 2885
rect 10185 2865 10200 2885
rect 10150 2835 10200 2865
rect 10150 2815 10165 2835
rect 10185 2815 10200 2835
rect 10150 2785 10200 2815
rect 10150 2765 10165 2785
rect 10185 2765 10200 2785
rect 10150 2735 10200 2765
rect 10150 2715 10165 2735
rect 10185 2715 10200 2735
rect 10150 2685 10200 2715
rect 10150 2665 10165 2685
rect 10185 2665 10200 2685
rect 10150 2650 10200 2665
rect 10300 3135 10350 3150
rect 10300 3115 10315 3135
rect 10335 3115 10350 3135
rect 10300 3085 10350 3115
rect 10300 3065 10315 3085
rect 10335 3065 10350 3085
rect 10300 3035 10350 3065
rect 10300 3015 10315 3035
rect 10335 3015 10350 3035
rect 10300 2985 10350 3015
rect 10300 2965 10315 2985
rect 10335 2965 10350 2985
rect 10300 2935 10350 2965
rect 10300 2915 10315 2935
rect 10335 2915 10350 2935
rect 10300 2885 10350 2915
rect 10300 2865 10315 2885
rect 10335 2865 10350 2885
rect 10300 2835 10350 2865
rect 10300 2815 10315 2835
rect 10335 2815 10350 2835
rect 10300 2785 10350 2815
rect 10300 2765 10315 2785
rect 10335 2765 10350 2785
rect 10300 2735 10350 2765
rect 10300 2715 10315 2735
rect 10335 2715 10350 2735
rect 10300 2685 10350 2715
rect 10300 2665 10315 2685
rect 10335 2665 10350 2685
rect 10300 2650 10350 2665
rect 10450 3135 10500 3150
rect 10450 3115 10465 3135
rect 10485 3115 10500 3135
rect 10450 3085 10500 3115
rect 10450 3065 10465 3085
rect 10485 3065 10500 3085
rect 10450 3035 10500 3065
rect 10450 3015 10465 3035
rect 10485 3015 10500 3035
rect 10450 2985 10500 3015
rect 10450 2965 10465 2985
rect 10485 2965 10500 2985
rect 10450 2935 10500 2965
rect 10450 2915 10465 2935
rect 10485 2915 10500 2935
rect 10450 2885 10500 2915
rect 10450 2865 10465 2885
rect 10485 2865 10500 2885
rect 10450 2835 10500 2865
rect 10450 2815 10465 2835
rect 10485 2815 10500 2835
rect 10450 2785 10500 2815
rect 10450 2765 10465 2785
rect 10485 2765 10500 2785
rect 10450 2735 10500 2765
rect 10450 2715 10465 2735
rect 10485 2715 10500 2735
rect 10450 2685 10500 2715
rect 10450 2665 10465 2685
rect 10485 2665 10500 2685
rect 10450 2650 10500 2665
rect 10600 3135 10650 3150
rect 10600 3115 10615 3135
rect 10635 3115 10650 3135
rect 10600 3085 10650 3115
rect 10600 3065 10615 3085
rect 10635 3065 10650 3085
rect 10600 3035 10650 3065
rect 10600 3015 10615 3035
rect 10635 3015 10650 3035
rect 10600 2985 10650 3015
rect 10600 2965 10615 2985
rect 10635 2965 10650 2985
rect 10600 2935 10650 2965
rect 10600 2915 10615 2935
rect 10635 2915 10650 2935
rect 10600 2885 10650 2915
rect 10600 2865 10615 2885
rect 10635 2865 10650 2885
rect 10600 2835 10650 2865
rect 10600 2815 10615 2835
rect 10635 2815 10650 2835
rect 10600 2785 10650 2815
rect 10600 2765 10615 2785
rect 10635 2765 10650 2785
rect 10600 2735 10650 2765
rect 10600 2715 10615 2735
rect 10635 2715 10650 2735
rect 10600 2685 10650 2715
rect 10600 2665 10615 2685
rect 10635 2665 10650 2685
rect 10600 2650 10650 2665
rect 10750 3135 10800 3150
rect 10750 3115 10765 3135
rect 10785 3115 10800 3135
rect 10750 3085 10800 3115
rect 10750 3065 10765 3085
rect 10785 3065 10800 3085
rect 10750 3035 10800 3065
rect 10750 3015 10765 3035
rect 10785 3015 10800 3035
rect 10750 2985 10800 3015
rect 10750 2965 10765 2985
rect 10785 2965 10800 2985
rect 10750 2935 10800 2965
rect 10750 2915 10765 2935
rect 10785 2915 10800 2935
rect 10750 2885 10800 2915
rect 10750 2865 10765 2885
rect 10785 2865 10800 2885
rect 10750 2835 10800 2865
rect 10750 2815 10765 2835
rect 10785 2815 10800 2835
rect 10750 2785 10800 2815
rect 10750 2765 10765 2785
rect 10785 2765 10800 2785
rect 10750 2735 10800 2765
rect 10750 2715 10765 2735
rect 10785 2715 10800 2735
rect 10750 2685 10800 2715
rect 10750 2665 10765 2685
rect 10785 2665 10800 2685
rect 10750 2650 10800 2665
rect 10900 2650 10950 3150
rect 11050 2650 11100 3150
rect 11200 2650 11250 3150
rect 11350 3135 11400 3150
rect 11350 3115 11365 3135
rect 11385 3115 11400 3135
rect 11350 3085 11400 3115
rect 11350 3065 11365 3085
rect 11385 3065 11400 3085
rect 11350 3035 11400 3065
rect 11350 3015 11365 3035
rect 11385 3015 11400 3035
rect 11350 2985 11400 3015
rect 11350 2965 11365 2985
rect 11385 2965 11400 2985
rect 11350 2935 11400 2965
rect 11350 2915 11365 2935
rect 11385 2915 11400 2935
rect 11350 2885 11400 2915
rect 11350 2865 11365 2885
rect 11385 2865 11400 2885
rect 11350 2835 11400 2865
rect 11350 2815 11365 2835
rect 11385 2815 11400 2835
rect 11350 2785 11400 2815
rect 11350 2765 11365 2785
rect 11385 2765 11400 2785
rect 11350 2735 11400 2765
rect 11350 2715 11365 2735
rect 11385 2715 11400 2735
rect 11350 2685 11400 2715
rect 11350 2665 11365 2685
rect 11385 2665 11400 2685
rect 11350 2650 11400 2665
rect 11500 2650 11550 3150
rect 11650 2650 11700 3150
rect 11800 2650 11850 3150
rect 11950 3135 12000 3150
rect 11950 3115 11965 3135
rect 11985 3115 12000 3135
rect 11950 3085 12000 3115
rect 11950 3065 11965 3085
rect 11985 3065 12000 3085
rect 11950 3035 12000 3065
rect 11950 3015 11965 3035
rect 11985 3015 12000 3035
rect 11950 2985 12000 3015
rect 11950 2965 11965 2985
rect 11985 2965 12000 2985
rect 11950 2935 12000 2965
rect 11950 2915 11965 2935
rect 11985 2915 12000 2935
rect 11950 2885 12000 2915
rect 11950 2865 11965 2885
rect 11985 2865 12000 2885
rect 11950 2835 12000 2865
rect 11950 2815 11965 2835
rect 11985 2815 12000 2835
rect 11950 2785 12000 2815
rect 11950 2765 11965 2785
rect 11985 2765 12000 2785
rect 11950 2735 12000 2765
rect 11950 2715 11965 2735
rect 11985 2715 12000 2735
rect 11950 2685 12000 2715
rect 11950 2665 11965 2685
rect 11985 2665 12000 2685
rect 11950 2650 12000 2665
rect 12100 2650 12150 3150
rect 12250 2650 12300 3150
rect 12400 2650 12450 3150
rect 12550 3135 12600 3150
rect 12550 3115 12565 3135
rect 12585 3115 12600 3135
rect 12550 3085 12600 3115
rect 12550 3065 12565 3085
rect 12585 3065 12600 3085
rect 12550 3035 12600 3065
rect 12550 3015 12565 3035
rect 12585 3015 12600 3035
rect 12550 2985 12600 3015
rect 12550 2965 12565 2985
rect 12585 2965 12600 2985
rect 12550 2935 12600 2965
rect 12550 2915 12565 2935
rect 12585 2915 12600 2935
rect 12550 2885 12600 2915
rect 12550 2865 12565 2885
rect 12585 2865 12600 2885
rect 12550 2835 12600 2865
rect 12550 2815 12565 2835
rect 12585 2815 12600 2835
rect 12550 2785 12600 2815
rect 12550 2765 12565 2785
rect 12585 2765 12600 2785
rect 12550 2735 12600 2765
rect 12550 2715 12565 2735
rect 12585 2715 12600 2735
rect 12550 2685 12600 2715
rect 12550 2665 12565 2685
rect 12585 2665 12600 2685
rect 12550 2650 12600 2665
rect 12700 2650 12750 3150
rect 12850 2650 12900 3150
rect 13000 2650 13050 3150
rect 13150 3135 13200 3150
rect 13150 3115 13165 3135
rect 13185 3115 13200 3135
rect 13150 3085 13200 3115
rect 13150 3065 13165 3085
rect 13185 3065 13200 3085
rect 13150 3035 13200 3065
rect 13150 3015 13165 3035
rect 13185 3015 13200 3035
rect 13150 2985 13200 3015
rect 13150 2965 13165 2985
rect 13185 2965 13200 2985
rect 13150 2935 13200 2965
rect 13150 2915 13165 2935
rect 13185 2915 13200 2935
rect 13150 2885 13200 2915
rect 13150 2865 13165 2885
rect 13185 2865 13200 2885
rect 13150 2835 13200 2865
rect 13150 2815 13165 2835
rect 13185 2815 13200 2835
rect 13150 2785 13200 2815
rect 13150 2765 13165 2785
rect 13185 2765 13200 2785
rect 13150 2735 13200 2765
rect 13150 2715 13165 2735
rect 13185 2715 13200 2735
rect 13150 2685 13200 2715
rect 13150 2665 13165 2685
rect 13185 2665 13200 2685
rect 13150 2650 13200 2665
rect 13300 2650 13350 3150
rect 13450 2650 13500 3150
rect 13600 2650 13650 3150
rect 13750 3135 13800 3150
rect 13750 3115 13765 3135
rect 13785 3115 13800 3135
rect 13750 3085 13800 3115
rect 13750 3065 13765 3085
rect 13785 3065 13800 3085
rect 13750 3035 13800 3065
rect 13750 3015 13765 3035
rect 13785 3015 13800 3035
rect 13750 2985 13800 3015
rect 13750 2965 13765 2985
rect 13785 2965 13800 2985
rect 13750 2935 13800 2965
rect 13750 2915 13765 2935
rect 13785 2915 13800 2935
rect 13750 2885 13800 2915
rect 13750 2865 13765 2885
rect 13785 2865 13800 2885
rect 13750 2835 13800 2865
rect 13750 2815 13765 2835
rect 13785 2815 13800 2835
rect 13750 2785 13800 2815
rect 13750 2765 13765 2785
rect 13785 2765 13800 2785
rect 13750 2735 13800 2765
rect 13750 2715 13765 2735
rect 13785 2715 13800 2735
rect 13750 2685 13800 2715
rect 13750 2665 13765 2685
rect 13785 2665 13800 2685
rect 13750 2650 13800 2665
rect 13900 2650 13950 3150
rect 14050 2650 14100 3150
rect 14200 2650 14250 3150
rect 14350 3135 14400 3150
rect 14350 3115 14365 3135
rect 14385 3115 14400 3135
rect 14350 3085 14400 3115
rect 14350 3065 14365 3085
rect 14385 3065 14400 3085
rect 14350 3035 14400 3065
rect 14350 3015 14365 3035
rect 14385 3015 14400 3035
rect 14350 2985 14400 3015
rect 14350 2965 14365 2985
rect 14385 2965 14400 2985
rect 14350 2935 14400 2965
rect 14350 2915 14365 2935
rect 14385 2915 14400 2935
rect 14350 2885 14400 2915
rect 14350 2865 14365 2885
rect 14385 2865 14400 2885
rect 14350 2835 14400 2865
rect 14350 2815 14365 2835
rect 14385 2815 14400 2835
rect 14350 2785 14400 2815
rect 14350 2765 14365 2785
rect 14385 2765 14400 2785
rect 14350 2735 14400 2765
rect 14350 2715 14365 2735
rect 14385 2715 14400 2735
rect 14350 2685 14400 2715
rect 14350 2665 14365 2685
rect 14385 2665 14400 2685
rect 14350 2650 14400 2665
rect 14500 2650 14550 3150
rect 14650 2650 14700 3150
rect 14800 2650 14850 3150
rect 14950 3135 15000 3150
rect 14950 3115 14965 3135
rect 14985 3115 15000 3135
rect 14950 3085 15000 3115
rect 14950 3065 14965 3085
rect 14985 3065 15000 3085
rect 14950 3035 15000 3065
rect 14950 3015 14965 3035
rect 14985 3015 15000 3035
rect 14950 2985 15000 3015
rect 14950 2965 14965 2985
rect 14985 2965 15000 2985
rect 14950 2935 15000 2965
rect 14950 2915 14965 2935
rect 14985 2915 15000 2935
rect 14950 2885 15000 2915
rect 14950 2865 14965 2885
rect 14985 2865 15000 2885
rect 14950 2835 15000 2865
rect 14950 2815 14965 2835
rect 14985 2815 15000 2835
rect 14950 2785 15000 2815
rect 14950 2765 14965 2785
rect 14985 2765 15000 2785
rect 14950 2735 15000 2765
rect 14950 2715 14965 2735
rect 14985 2715 15000 2735
rect 14950 2685 15000 2715
rect 14950 2665 14965 2685
rect 14985 2665 15000 2685
rect 14950 2650 15000 2665
rect 15100 2650 15150 3150
rect 15250 2650 15300 3150
rect 15400 2650 15450 3150
rect 15550 3135 15600 3150
rect 15550 3115 15565 3135
rect 15585 3115 15600 3135
rect 15550 3085 15600 3115
rect 15550 3065 15565 3085
rect 15585 3065 15600 3085
rect 15550 3035 15600 3065
rect 15550 3015 15565 3035
rect 15585 3015 15600 3035
rect 15550 2985 15600 3015
rect 15550 2965 15565 2985
rect 15585 2965 15600 2985
rect 15550 2935 15600 2965
rect 15550 2915 15565 2935
rect 15585 2915 15600 2935
rect 15550 2885 15600 2915
rect 15550 2865 15565 2885
rect 15585 2865 15600 2885
rect 15550 2835 15600 2865
rect 15550 2815 15565 2835
rect 15585 2815 15600 2835
rect 15550 2785 15600 2815
rect 15550 2765 15565 2785
rect 15585 2765 15600 2785
rect 15550 2735 15600 2765
rect 15550 2715 15565 2735
rect 15585 2715 15600 2735
rect 15550 2685 15600 2715
rect 15550 2665 15565 2685
rect 15585 2665 15600 2685
rect 15550 2650 15600 2665
rect 15700 2650 15750 3150
rect 15850 2650 15900 3150
rect 16000 2650 16050 3150
rect 16150 3135 16200 3150
rect 16150 3115 16165 3135
rect 16185 3115 16200 3135
rect 16150 3085 16200 3115
rect 16150 3065 16165 3085
rect 16185 3065 16200 3085
rect 16150 3035 16200 3065
rect 16150 3015 16165 3035
rect 16185 3015 16200 3035
rect 16150 2985 16200 3015
rect 16150 2965 16165 2985
rect 16185 2965 16200 2985
rect 16150 2935 16200 2965
rect 16150 2915 16165 2935
rect 16185 2915 16200 2935
rect 16150 2885 16200 2915
rect 16150 2865 16165 2885
rect 16185 2865 16200 2885
rect 16150 2835 16200 2865
rect 16150 2815 16165 2835
rect 16185 2815 16200 2835
rect 16150 2785 16200 2815
rect 16150 2765 16165 2785
rect 16185 2765 16200 2785
rect 16150 2735 16200 2765
rect 16150 2715 16165 2735
rect 16185 2715 16200 2735
rect 16150 2685 16200 2715
rect 16150 2665 16165 2685
rect 16185 2665 16200 2685
rect 16150 2650 16200 2665
rect 16300 3135 16350 3150
rect 16300 3115 16315 3135
rect 16335 3115 16350 3135
rect 16300 3085 16350 3115
rect 16300 3065 16315 3085
rect 16335 3065 16350 3085
rect 16300 3035 16350 3065
rect 16300 3015 16315 3035
rect 16335 3015 16350 3035
rect 16300 2985 16350 3015
rect 16300 2965 16315 2985
rect 16335 2965 16350 2985
rect 16300 2935 16350 2965
rect 16300 2915 16315 2935
rect 16335 2915 16350 2935
rect 16300 2885 16350 2915
rect 16300 2865 16315 2885
rect 16335 2865 16350 2885
rect 16300 2835 16350 2865
rect 16300 2815 16315 2835
rect 16335 2815 16350 2835
rect 16300 2785 16350 2815
rect 16300 2765 16315 2785
rect 16335 2765 16350 2785
rect 16300 2735 16350 2765
rect 16300 2715 16315 2735
rect 16335 2715 16350 2735
rect 16300 2685 16350 2715
rect 16300 2665 16315 2685
rect 16335 2665 16350 2685
rect 16300 2650 16350 2665
rect 16450 3135 16500 3150
rect 16450 3115 16465 3135
rect 16485 3115 16500 3135
rect 16450 3085 16500 3115
rect 16450 3065 16465 3085
rect 16485 3065 16500 3085
rect 16450 3035 16500 3065
rect 16450 3015 16465 3035
rect 16485 3015 16500 3035
rect 16450 2985 16500 3015
rect 16450 2965 16465 2985
rect 16485 2965 16500 2985
rect 16450 2935 16500 2965
rect 16450 2915 16465 2935
rect 16485 2915 16500 2935
rect 16450 2885 16500 2915
rect 16450 2865 16465 2885
rect 16485 2865 16500 2885
rect 16450 2835 16500 2865
rect 16450 2815 16465 2835
rect 16485 2815 16500 2835
rect 16450 2785 16500 2815
rect 16450 2765 16465 2785
rect 16485 2765 16500 2785
rect 16450 2735 16500 2765
rect 16450 2715 16465 2735
rect 16485 2715 16500 2735
rect 16450 2685 16500 2715
rect 16450 2665 16465 2685
rect 16485 2665 16500 2685
rect 16450 2650 16500 2665
rect 16600 3135 16650 3150
rect 16600 3115 16615 3135
rect 16635 3115 16650 3135
rect 16600 3085 16650 3115
rect 16600 3065 16615 3085
rect 16635 3065 16650 3085
rect 16600 3035 16650 3065
rect 16600 3015 16615 3035
rect 16635 3015 16650 3035
rect 16600 2985 16650 3015
rect 16600 2965 16615 2985
rect 16635 2965 16650 2985
rect 16600 2935 16650 2965
rect 16600 2915 16615 2935
rect 16635 2915 16650 2935
rect 16600 2885 16650 2915
rect 16600 2865 16615 2885
rect 16635 2865 16650 2885
rect 16600 2835 16650 2865
rect 16600 2815 16615 2835
rect 16635 2815 16650 2835
rect 16600 2785 16650 2815
rect 16600 2765 16615 2785
rect 16635 2765 16650 2785
rect 16600 2735 16650 2765
rect 16600 2715 16615 2735
rect 16635 2715 16650 2735
rect 16600 2685 16650 2715
rect 16600 2665 16615 2685
rect 16635 2665 16650 2685
rect 16600 2650 16650 2665
rect 16750 3135 16800 3150
rect 16750 3115 16765 3135
rect 16785 3115 16800 3135
rect 16750 3085 16800 3115
rect 16750 3065 16765 3085
rect 16785 3065 16800 3085
rect 16750 3035 16800 3065
rect 16750 3015 16765 3035
rect 16785 3015 16800 3035
rect 16750 2985 16800 3015
rect 16750 2965 16765 2985
rect 16785 2965 16800 2985
rect 16750 2935 16800 2965
rect 16750 2915 16765 2935
rect 16785 2915 16800 2935
rect 16750 2885 16800 2915
rect 16750 2865 16765 2885
rect 16785 2865 16800 2885
rect 16750 2835 16800 2865
rect 16750 2815 16765 2835
rect 16785 2815 16800 2835
rect 16750 2785 16800 2815
rect 16750 2765 16765 2785
rect 16785 2765 16800 2785
rect 16750 2735 16800 2765
rect 16750 2715 16765 2735
rect 16785 2715 16800 2735
rect 16750 2685 16800 2715
rect 16750 2665 16765 2685
rect 16785 2665 16800 2685
rect 16750 2650 16800 2665
rect 16900 3135 16950 3150
rect 16900 3115 16915 3135
rect 16935 3115 16950 3135
rect 16900 3085 16950 3115
rect 16900 3065 16915 3085
rect 16935 3065 16950 3085
rect 16900 3035 16950 3065
rect 16900 3015 16915 3035
rect 16935 3015 16950 3035
rect 16900 2985 16950 3015
rect 16900 2965 16915 2985
rect 16935 2965 16950 2985
rect 16900 2935 16950 2965
rect 16900 2915 16915 2935
rect 16935 2915 16950 2935
rect 16900 2885 16950 2915
rect 16900 2865 16915 2885
rect 16935 2865 16950 2885
rect 16900 2835 16950 2865
rect 16900 2815 16915 2835
rect 16935 2815 16950 2835
rect 16900 2785 16950 2815
rect 16900 2765 16915 2785
rect 16935 2765 16950 2785
rect 16900 2735 16950 2765
rect 16900 2715 16915 2735
rect 16935 2715 16950 2735
rect 16900 2685 16950 2715
rect 16900 2665 16915 2685
rect 16935 2665 16950 2685
rect 16900 2650 16950 2665
rect 17050 3135 17100 3150
rect 17050 3115 17065 3135
rect 17085 3115 17100 3135
rect 17050 3085 17100 3115
rect 17050 3065 17065 3085
rect 17085 3065 17100 3085
rect 17050 3035 17100 3065
rect 17050 3015 17065 3035
rect 17085 3015 17100 3035
rect 17050 2985 17100 3015
rect 17050 2965 17065 2985
rect 17085 2965 17100 2985
rect 17050 2935 17100 2965
rect 17050 2915 17065 2935
rect 17085 2915 17100 2935
rect 17050 2885 17100 2915
rect 17050 2865 17065 2885
rect 17085 2865 17100 2885
rect 17050 2835 17100 2865
rect 17050 2815 17065 2835
rect 17085 2815 17100 2835
rect 17050 2785 17100 2815
rect 17050 2765 17065 2785
rect 17085 2765 17100 2785
rect 17050 2735 17100 2765
rect 17050 2715 17065 2735
rect 17085 2715 17100 2735
rect 17050 2685 17100 2715
rect 17050 2665 17065 2685
rect 17085 2665 17100 2685
rect 17050 2650 17100 2665
rect 17200 3135 17250 3150
rect 17200 3115 17215 3135
rect 17235 3115 17250 3135
rect 17200 3085 17250 3115
rect 17200 3065 17215 3085
rect 17235 3065 17250 3085
rect 17200 3035 17250 3065
rect 17200 3015 17215 3035
rect 17235 3015 17250 3035
rect 17200 2985 17250 3015
rect 17200 2965 17215 2985
rect 17235 2965 17250 2985
rect 17200 2935 17250 2965
rect 17200 2915 17215 2935
rect 17235 2915 17250 2935
rect 17200 2885 17250 2915
rect 17200 2865 17215 2885
rect 17235 2865 17250 2885
rect 17200 2835 17250 2865
rect 17200 2815 17215 2835
rect 17235 2815 17250 2835
rect 17200 2785 17250 2815
rect 17200 2765 17215 2785
rect 17235 2765 17250 2785
rect 17200 2735 17250 2765
rect 17200 2715 17215 2735
rect 17235 2715 17250 2735
rect 17200 2685 17250 2715
rect 17200 2665 17215 2685
rect 17235 2665 17250 2685
rect 17200 2650 17250 2665
rect 17350 3135 17400 3150
rect 17350 3115 17365 3135
rect 17385 3115 17400 3135
rect 17350 3085 17400 3115
rect 17350 3065 17365 3085
rect 17385 3065 17400 3085
rect 17350 3035 17400 3065
rect 17350 3015 17365 3035
rect 17385 3015 17400 3035
rect 17350 2985 17400 3015
rect 17350 2965 17365 2985
rect 17385 2965 17400 2985
rect 17350 2935 17400 2965
rect 17350 2915 17365 2935
rect 17385 2915 17400 2935
rect 17350 2885 17400 2915
rect 17350 2865 17365 2885
rect 17385 2865 17400 2885
rect 17350 2835 17400 2865
rect 17350 2815 17365 2835
rect 17385 2815 17400 2835
rect 17350 2785 17400 2815
rect 17350 2765 17365 2785
rect 17385 2765 17400 2785
rect 17350 2735 17400 2765
rect 17350 2715 17365 2735
rect 17385 2715 17400 2735
rect 17350 2685 17400 2715
rect 17350 2665 17365 2685
rect 17385 2665 17400 2685
rect 17350 2650 17400 2665
rect 17500 2650 17550 3150
rect 17650 2650 17700 3150
rect 17800 2650 17850 3150
rect 17950 3135 18000 3150
rect 17950 3115 17965 3135
rect 17985 3115 18000 3135
rect 17950 3085 18000 3115
rect 17950 3065 17965 3085
rect 17985 3065 18000 3085
rect 17950 3035 18000 3065
rect 17950 3015 17965 3035
rect 17985 3015 18000 3035
rect 17950 2985 18000 3015
rect 17950 2965 17965 2985
rect 17985 2965 18000 2985
rect 17950 2935 18000 2965
rect 17950 2915 17965 2935
rect 17985 2915 18000 2935
rect 17950 2885 18000 2915
rect 17950 2865 17965 2885
rect 17985 2865 18000 2885
rect 17950 2835 18000 2865
rect 17950 2815 17965 2835
rect 17985 2815 18000 2835
rect 17950 2785 18000 2815
rect 17950 2765 17965 2785
rect 17985 2765 18000 2785
rect 17950 2735 18000 2765
rect 17950 2715 17965 2735
rect 17985 2715 18000 2735
rect 17950 2685 18000 2715
rect 17950 2665 17965 2685
rect 17985 2665 18000 2685
rect 17950 2650 18000 2665
rect 18100 2650 18150 3150
rect 18250 2650 18300 3150
rect 18400 2650 18450 3150
rect 18550 3135 18600 3150
rect 18550 3115 18565 3135
rect 18585 3115 18600 3135
rect 18550 3085 18600 3115
rect 18550 3065 18565 3085
rect 18585 3065 18600 3085
rect 18550 3035 18600 3065
rect 18550 3015 18565 3035
rect 18585 3015 18600 3035
rect 18550 2985 18600 3015
rect 18550 2965 18565 2985
rect 18585 2965 18600 2985
rect 18550 2935 18600 2965
rect 18550 2915 18565 2935
rect 18585 2915 18600 2935
rect 18550 2885 18600 2915
rect 18550 2865 18565 2885
rect 18585 2865 18600 2885
rect 18550 2835 18600 2865
rect 18550 2815 18565 2835
rect 18585 2815 18600 2835
rect 18550 2785 18600 2815
rect 18550 2765 18565 2785
rect 18585 2765 18600 2785
rect 18550 2735 18600 2765
rect 18550 2715 18565 2735
rect 18585 2715 18600 2735
rect 18550 2685 18600 2715
rect 18550 2665 18565 2685
rect 18585 2665 18600 2685
rect 18550 2650 18600 2665
rect 18700 3135 18750 3150
rect 18700 3115 18715 3135
rect 18735 3115 18750 3135
rect 18700 3085 18750 3115
rect 18700 3065 18715 3085
rect 18735 3065 18750 3085
rect 18700 3035 18750 3065
rect 18700 3015 18715 3035
rect 18735 3015 18750 3035
rect 18700 2985 18750 3015
rect 18700 2965 18715 2985
rect 18735 2965 18750 2985
rect 18700 2935 18750 2965
rect 18700 2915 18715 2935
rect 18735 2915 18750 2935
rect 18700 2885 18750 2915
rect 18700 2865 18715 2885
rect 18735 2865 18750 2885
rect 18700 2835 18750 2865
rect 18700 2815 18715 2835
rect 18735 2815 18750 2835
rect 18700 2785 18750 2815
rect 18700 2765 18715 2785
rect 18735 2765 18750 2785
rect 18700 2735 18750 2765
rect 18700 2715 18715 2735
rect 18735 2715 18750 2735
rect 18700 2685 18750 2715
rect 18700 2665 18715 2685
rect 18735 2665 18750 2685
rect 18700 2650 18750 2665
rect 18850 3135 18900 3150
rect 18850 3115 18865 3135
rect 18885 3115 18900 3135
rect 18850 3085 18900 3115
rect 18850 3065 18865 3085
rect 18885 3065 18900 3085
rect 18850 3035 18900 3065
rect 18850 3015 18865 3035
rect 18885 3015 18900 3035
rect 18850 2985 18900 3015
rect 18850 2965 18865 2985
rect 18885 2965 18900 2985
rect 18850 2935 18900 2965
rect 18850 2915 18865 2935
rect 18885 2915 18900 2935
rect 18850 2885 18900 2915
rect 18850 2865 18865 2885
rect 18885 2865 18900 2885
rect 18850 2835 18900 2865
rect 18850 2815 18865 2835
rect 18885 2815 18900 2835
rect 18850 2785 18900 2815
rect 18850 2765 18865 2785
rect 18885 2765 18900 2785
rect 18850 2735 18900 2765
rect 18850 2715 18865 2735
rect 18885 2715 18900 2735
rect 18850 2685 18900 2715
rect 18850 2665 18865 2685
rect 18885 2665 18900 2685
rect 18850 2650 18900 2665
rect 19000 3135 19050 3150
rect 19000 3115 19015 3135
rect 19035 3115 19050 3135
rect 19000 3085 19050 3115
rect 19000 3065 19015 3085
rect 19035 3065 19050 3085
rect 19000 3035 19050 3065
rect 19000 3015 19015 3035
rect 19035 3015 19050 3035
rect 19000 2985 19050 3015
rect 19000 2965 19015 2985
rect 19035 2965 19050 2985
rect 19000 2935 19050 2965
rect 19000 2915 19015 2935
rect 19035 2915 19050 2935
rect 19000 2885 19050 2915
rect 19000 2865 19015 2885
rect 19035 2865 19050 2885
rect 19000 2835 19050 2865
rect 19000 2815 19015 2835
rect 19035 2815 19050 2835
rect 19000 2785 19050 2815
rect 19000 2765 19015 2785
rect 19035 2765 19050 2785
rect 19000 2735 19050 2765
rect 19000 2715 19015 2735
rect 19035 2715 19050 2735
rect 19000 2685 19050 2715
rect 19000 2665 19015 2685
rect 19035 2665 19050 2685
rect 19000 2650 19050 2665
rect 19150 3135 19200 3150
rect 19150 3115 19165 3135
rect 19185 3115 19200 3135
rect 19150 3085 19200 3115
rect 19150 3065 19165 3085
rect 19185 3065 19200 3085
rect 19150 3035 19200 3065
rect 19150 3015 19165 3035
rect 19185 3015 19200 3035
rect 19150 2985 19200 3015
rect 19150 2965 19165 2985
rect 19185 2965 19200 2985
rect 19150 2935 19200 2965
rect 19150 2915 19165 2935
rect 19185 2915 19200 2935
rect 19150 2885 19200 2915
rect 19150 2865 19165 2885
rect 19185 2865 19200 2885
rect 19150 2835 19200 2865
rect 19150 2815 19165 2835
rect 19185 2815 19200 2835
rect 19150 2785 19200 2815
rect 19150 2765 19165 2785
rect 19185 2765 19200 2785
rect 19150 2735 19200 2765
rect 19150 2715 19165 2735
rect 19185 2715 19200 2735
rect 19150 2685 19200 2715
rect 19150 2665 19165 2685
rect 19185 2665 19200 2685
rect 19150 2650 19200 2665
rect 19300 3135 19350 3150
rect 19300 3115 19315 3135
rect 19335 3115 19350 3135
rect 19300 3085 19350 3115
rect 19300 3065 19315 3085
rect 19335 3065 19350 3085
rect 19300 3035 19350 3065
rect 19300 3015 19315 3035
rect 19335 3015 19350 3035
rect 19300 2985 19350 3015
rect 19300 2965 19315 2985
rect 19335 2965 19350 2985
rect 19300 2935 19350 2965
rect 19300 2915 19315 2935
rect 19335 2915 19350 2935
rect 19300 2885 19350 2915
rect 19300 2865 19315 2885
rect 19335 2865 19350 2885
rect 19300 2835 19350 2865
rect 19300 2815 19315 2835
rect 19335 2815 19350 2835
rect 19300 2785 19350 2815
rect 19300 2765 19315 2785
rect 19335 2765 19350 2785
rect 19300 2735 19350 2765
rect 19300 2715 19315 2735
rect 19335 2715 19350 2735
rect 19300 2685 19350 2715
rect 19300 2665 19315 2685
rect 19335 2665 19350 2685
rect 19300 2650 19350 2665
rect 19450 3135 19500 3150
rect 19450 3115 19465 3135
rect 19485 3115 19500 3135
rect 19450 3085 19500 3115
rect 19450 3065 19465 3085
rect 19485 3065 19500 3085
rect 19450 3035 19500 3065
rect 19450 3015 19465 3035
rect 19485 3015 19500 3035
rect 19450 2985 19500 3015
rect 19450 2965 19465 2985
rect 19485 2965 19500 2985
rect 19450 2935 19500 2965
rect 19450 2915 19465 2935
rect 19485 2915 19500 2935
rect 19450 2885 19500 2915
rect 19450 2865 19465 2885
rect 19485 2865 19500 2885
rect 19450 2835 19500 2865
rect 19450 2815 19465 2835
rect 19485 2815 19500 2835
rect 19450 2785 19500 2815
rect 19450 2765 19465 2785
rect 19485 2765 19500 2785
rect 19450 2735 19500 2765
rect 19450 2715 19465 2735
rect 19485 2715 19500 2735
rect 19450 2685 19500 2715
rect 19450 2665 19465 2685
rect 19485 2665 19500 2685
rect 19450 2650 19500 2665
rect 19600 3135 19650 3150
rect 19600 3115 19615 3135
rect 19635 3115 19650 3135
rect 19600 3085 19650 3115
rect 19600 3065 19615 3085
rect 19635 3065 19650 3085
rect 19600 3035 19650 3065
rect 19600 3015 19615 3035
rect 19635 3015 19650 3035
rect 19600 2985 19650 3015
rect 19600 2965 19615 2985
rect 19635 2965 19650 2985
rect 19600 2935 19650 2965
rect 19600 2915 19615 2935
rect 19635 2915 19650 2935
rect 19600 2885 19650 2915
rect 19600 2865 19615 2885
rect 19635 2865 19650 2885
rect 19600 2835 19650 2865
rect 19600 2815 19615 2835
rect 19635 2815 19650 2835
rect 19600 2785 19650 2815
rect 19600 2765 19615 2785
rect 19635 2765 19650 2785
rect 19600 2735 19650 2765
rect 19600 2715 19615 2735
rect 19635 2715 19650 2735
rect 19600 2685 19650 2715
rect 19600 2665 19615 2685
rect 19635 2665 19650 2685
rect 19600 2650 19650 2665
rect 19750 3135 19800 3150
rect 19750 3115 19765 3135
rect 19785 3115 19800 3135
rect 19750 3085 19800 3115
rect 19750 3065 19765 3085
rect 19785 3065 19800 3085
rect 19750 3035 19800 3065
rect 19750 3015 19765 3035
rect 19785 3015 19800 3035
rect 19750 2985 19800 3015
rect 19750 2965 19765 2985
rect 19785 2965 19800 2985
rect 19750 2935 19800 2965
rect 19750 2915 19765 2935
rect 19785 2915 19800 2935
rect 19750 2885 19800 2915
rect 19750 2865 19765 2885
rect 19785 2865 19800 2885
rect 19750 2835 19800 2865
rect 19750 2815 19765 2835
rect 19785 2815 19800 2835
rect 19750 2785 19800 2815
rect 19750 2765 19765 2785
rect 19785 2765 19800 2785
rect 19750 2735 19800 2765
rect 19750 2715 19765 2735
rect 19785 2715 19800 2735
rect 19750 2685 19800 2715
rect 19750 2665 19765 2685
rect 19785 2665 19800 2685
rect 19750 2650 19800 2665
rect 19900 2650 19950 3150
rect 20050 2650 20100 3150
rect 20200 2650 20250 3150
rect 20350 3135 20400 3150
rect 20350 3115 20365 3135
rect 20385 3115 20400 3135
rect 20350 3085 20400 3115
rect 20350 3065 20365 3085
rect 20385 3065 20400 3085
rect 20350 3035 20400 3065
rect 20350 3015 20365 3035
rect 20385 3015 20400 3035
rect 20350 2985 20400 3015
rect 20350 2965 20365 2985
rect 20385 2965 20400 2985
rect 20350 2935 20400 2965
rect 20350 2915 20365 2935
rect 20385 2915 20400 2935
rect 20350 2885 20400 2915
rect 20350 2865 20365 2885
rect 20385 2865 20400 2885
rect 20350 2835 20400 2865
rect 20350 2815 20365 2835
rect 20385 2815 20400 2835
rect 20350 2785 20400 2815
rect 20350 2765 20365 2785
rect 20385 2765 20400 2785
rect 20350 2735 20400 2765
rect 20350 2715 20365 2735
rect 20385 2715 20400 2735
rect 20350 2685 20400 2715
rect 20350 2665 20365 2685
rect 20385 2665 20400 2685
rect 20350 2650 20400 2665
<< mvndiffc >>
rect -635 1565 -615 1585
rect -635 1515 -615 1535
rect -635 1465 -615 1485
rect -635 1415 -615 1435
rect -635 1365 -615 1385
rect -635 1315 -615 1335
rect -635 1265 -615 1285
rect -635 1215 -615 1235
rect -635 1165 -615 1185
rect -635 1115 -615 1135
rect -635 1065 -615 1085
rect -635 1015 -615 1035
rect -635 965 -615 985
rect -635 915 -615 935
rect -485 1565 -465 1585
rect -485 1515 -465 1535
rect -485 1465 -465 1485
rect -485 1415 -465 1435
rect -485 1365 -465 1385
rect -485 1315 -465 1335
rect -485 1265 -465 1285
rect -485 1215 -465 1235
rect -485 1165 -465 1185
rect -485 1115 -465 1135
rect -485 1065 -465 1085
rect -485 1015 -465 1035
rect -485 965 -465 985
rect -485 915 -465 935
rect -335 1565 -315 1585
rect -335 1515 -315 1535
rect -335 1465 -315 1485
rect -335 1415 -315 1435
rect -335 1365 -315 1385
rect -335 1315 -315 1335
rect -335 1265 -315 1285
rect -335 1215 -315 1235
rect -335 1165 -315 1185
rect -335 1115 -315 1135
rect -335 1065 -315 1085
rect -335 1015 -315 1035
rect -335 965 -315 985
rect -335 915 -315 935
rect -185 1565 -165 1585
rect -185 1515 -165 1535
rect -185 1465 -165 1485
rect -185 1415 -165 1435
rect -185 1365 -165 1385
rect -185 1315 -165 1335
rect -185 1265 -165 1285
rect -185 1215 -165 1235
rect -185 1165 -165 1185
rect -185 1115 -165 1135
rect -185 1065 -165 1085
rect -185 1015 -165 1035
rect -185 965 -165 985
rect -185 915 -165 935
rect -35 1565 -15 1585
rect -35 1515 -15 1535
rect -35 1465 -15 1485
rect -35 1415 -15 1435
rect -35 1365 -15 1385
rect -35 1315 -15 1335
rect -35 1265 -15 1285
rect -35 1215 -15 1235
rect -35 1165 -15 1185
rect -35 1115 -15 1135
rect -35 1065 -15 1085
rect -35 1015 -15 1035
rect -35 965 -15 985
rect -35 915 -15 935
rect 1165 1565 1185 1585
rect 1165 1515 1185 1535
rect 1165 1465 1185 1485
rect 1165 1415 1185 1435
rect 1165 1365 1185 1385
rect 1165 1315 1185 1335
rect 1165 1265 1185 1285
rect 1165 1215 1185 1235
rect 1165 1165 1185 1185
rect 1165 1115 1185 1135
rect 1165 1065 1185 1085
rect 1165 1015 1185 1035
rect 1165 965 1185 985
rect 1165 915 1185 935
rect 1465 1565 1485 1585
rect 1465 1515 1485 1535
rect 1465 1465 1485 1485
rect 1465 1415 1485 1435
rect 1465 1365 1485 1385
rect 1465 1315 1485 1335
rect 1465 1265 1485 1285
rect 1465 1215 1485 1235
rect 1465 1165 1485 1185
rect 1465 1115 1485 1135
rect 1465 1065 1485 1085
rect 1465 1015 1485 1035
rect 1465 965 1485 985
rect 1465 915 1485 935
rect 1765 1565 1785 1585
rect 1765 1515 1785 1535
rect 1765 1465 1785 1485
rect 1765 1415 1785 1435
rect 1765 1365 1785 1385
rect 1765 1315 1785 1335
rect 1765 1265 1785 1285
rect 1765 1215 1785 1235
rect 1765 1165 1785 1185
rect 1765 1115 1785 1135
rect 1765 1065 1785 1085
rect 1765 1015 1785 1035
rect 1765 965 1785 985
rect 1765 915 1785 935
rect 2065 1565 2085 1585
rect 2065 1515 2085 1535
rect 2065 1465 2085 1485
rect 2065 1415 2085 1435
rect 2065 1365 2085 1385
rect 2065 1315 2085 1335
rect 2065 1265 2085 1285
rect 2065 1215 2085 1235
rect 2065 1165 2085 1185
rect 2065 1115 2085 1135
rect 2065 1065 2085 1085
rect 2065 1015 2085 1035
rect 2065 965 2085 985
rect 2065 915 2085 935
rect 2365 1565 2385 1585
rect 2365 1515 2385 1535
rect 2365 1465 2385 1485
rect 2365 1415 2385 1435
rect 2365 1365 2385 1385
rect 2365 1315 2385 1335
rect 2365 1265 2385 1285
rect 2365 1215 2385 1235
rect 2365 1165 2385 1185
rect 2365 1115 2385 1135
rect 2365 1065 2385 1085
rect 2365 1015 2385 1035
rect 2365 965 2385 985
rect 2365 915 2385 935
rect 2665 1565 2685 1585
rect 2665 1515 2685 1535
rect 2665 1465 2685 1485
rect 2665 1415 2685 1435
rect 2665 1365 2685 1385
rect 2665 1315 2685 1335
rect 2665 1265 2685 1285
rect 2665 1215 2685 1235
rect 2665 1165 2685 1185
rect 2665 1115 2685 1135
rect 2665 1065 2685 1085
rect 2665 1015 2685 1035
rect 2665 965 2685 985
rect 2665 915 2685 935
rect 2965 1565 2985 1585
rect 2965 1515 2985 1535
rect 2965 1465 2985 1485
rect 2965 1415 2985 1435
rect 2965 1365 2985 1385
rect 2965 1315 2985 1335
rect 2965 1265 2985 1285
rect 2965 1215 2985 1235
rect 2965 1165 2985 1185
rect 2965 1115 2985 1135
rect 2965 1065 2985 1085
rect 2965 1015 2985 1035
rect 2965 965 2985 985
rect 2965 915 2985 935
rect 3265 1565 3285 1585
rect 3265 1515 3285 1535
rect 3265 1465 3285 1485
rect 3265 1415 3285 1435
rect 3265 1365 3285 1385
rect 3265 1315 3285 1335
rect 3265 1265 3285 1285
rect 3265 1215 3285 1235
rect 3265 1165 3285 1185
rect 3265 1115 3285 1135
rect 3265 1065 3285 1085
rect 3265 1015 3285 1035
rect 3265 965 3285 985
rect 3265 915 3285 935
rect 3565 1565 3585 1585
rect 3565 1515 3585 1535
rect 3565 1465 3585 1485
rect 3565 1415 3585 1435
rect 3565 1365 3585 1385
rect 3565 1315 3585 1335
rect 3565 1265 3585 1285
rect 3565 1215 3585 1235
rect 3565 1165 3585 1185
rect 3565 1115 3585 1135
rect 3565 1065 3585 1085
rect 3565 1015 3585 1035
rect 3565 965 3585 985
rect 3565 915 3585 935
rect 3715 1565 3735 1585
rect 3715 1515 3735 1535
rect 3715 1465 3735 1485
rect 3715 1415 3735 1435
rect 3715 1365 3735 1385
rect 3715 1315 3735 1335
rect 3715 1265 3735 1285
rect 3715 1215 3735 1235
rect 3715 1165 3735 1185
rect 3715 1115 3735 1135
rect 3715 1065 3735 1085
rect 3715 1015 3735 1035
rect 3715 965 3735 985
rect 3715 915 3735 935
rect 3865 1565 3885 1585
rect 3865 1515 3885 1535
rect 3865 1465 3885 1485
rect 3865 1415 3885 1435
rect 3865 1365 3885 1385
rect 3865 1315 3885 1335
rect 3865 1265 3885 1285
rect 3865 1215 3885 1235
rect 3865 1165 3885 1185
rect 3865 1115 3885 1135
rect 3865 1065 3885 1085
rect 3865 1015 3885 1035
rect 3865 965 3885 985
rect 3865 915 3885 935
rect 4015 1565 4035 1585
rect 4015 1515 4035 1535
rect 4015 1465 4035 1485
rect 4015 1415 4035 1435
rect 4015 1365 4035 1385
rect 4015 1315 4035 1335
rect 4015 1265 4035 1285
rect 4015 1215 4035 1235
rect 4015 1165 4035 1185
rect 4015 1115 4035 1135
rect 4015 1065 4035 1085
rect 4015 1015 4035 1035
rect 4015 965 4035 985
rect 4015 915 4035 935
rect 4165 1565 4185 1585
rect 4165 1515 4185 1535
rect 4165 1465 4185 1485
rect 4165 1415 4185 1435
rect 4165 1365 4185 1385
rect 4165 1315 4185 1335
rect 4165 1265 4185 1285
rect 4165 1215 4185 1235
rect 4165 1165 4185 1185
rect 4165 1115 4185 1135
rect 4165 1065 4185 1085
rect 4165 1015 4185 1035
rect 4165 965 4185 985
rect 4165 915 4185 935
rect 4315 1565 4335 1585
rect 4315 1515 4335 1535
rect 4315 1465 4335 1485
rect 4315 1415 4335 1435
rect 4315 1365 4335 1385
rect 4315 1315 4335 1335
rect 4315 1265 4335 1285
rect 4315 1215 4335 1235
rect 4315 1165 4335 1185
rect 4315 1115 4335 1135
rect 4315 1065 4335 1085
rect 4315 1015 4335 1035
rect 4315 965 4335 985
rect 4315 915 4335 935
rect 4465 1565 4485 1585
rect 4465 1515 4485 1535
rect 4465 1465 4485 1485
rect 4465 1415 4485 1435
rect 4465 1365 4485 1385
rect 4465 1315 4485 1335
rect 4465 1265 4485 1285
rect 4465 1215 4485 1235
rect 4465 1165 4485 1185
rect 4465 1115 4485 1135
rect 4465 1065 4485 1085
rect 4465 1015 4485 1035
rect 4465 965 4485 985
rect 4465 915 4485 935
rect 4615 1565 4635 1585
rect 4615 1515 4635 1535
rect 4615 1465 4635 1485
rect 4615 1415 4635 1435
rect 4615 1365 4635 1385
rect 4615 1315 4635 1335
rect 4615 1265 4635 1285
rect 4615 1215 4635 1235
rect 4615 1165 4635 1185
rect 4615 1115 4635 1135
rect 4615 1065 4635 1085
rect 4615 1015 4635 1035
rect 4615 965 4635 985
rect 4615 915 4635 935
rect 4765 1565 4785 1585
rect 4765 1515 4785 1535
rect 4765 1465 4785 1485
rect 4765 1415 4785 1435
rect 4765 1365 4785 1385
rect 4765 1315 4785 1335
rect 4765 1265 4785 1285
rect 4765 1215 4785 1235
rect 4765 1165 4785 1185
rect 4765 1115 4785 1135
rect 4765 1065 4785 1085
rect 4765 1015 4785 1035
rect 4765 965 4785 985
rect 4765 915 4785 935
rect 5065 1565 5085 1585
rect 5065 1515 5085 1535
rect 5065 1465 5085 1485
rect 5065 1415 5085 1435
rect 5065 1365 5085 1385
rect 5065 1315 5085 1335
rect 5065 1265 5085 1285
rect 5065 1215 5085 1235
rect 5065 1165 5085 1185
rect 5065 1115 5085 1135
rect 5065 1065 5085 1085
rect 5065 1015 5085 1035
rect 5065 965 5085 985
rect 5065 915 5085 935
rect 5365 1565 5385 1585
rect 5365 1515 5385 1535
rect 5365 1465 5385 1485
rect 5365 1415 5385 1435
rect 5365 1365 5385 1385
rect 5365 1315 5385 1335
rect 5365 1265 5385 1285
rect 5365 1215 5385 1235
rect 5365 1165 5385 1185
rect 5365 1115 5385 1135
rect 5365 1065 5385 1085
rect 5365 1015 5385 1035
rect 5365 965 5385 985
rect 5365 915 5385 935
rect 5665 1565 5685 1585
rect 5665 1515 5685 1535
rect 5665 1465 5685 1485
rect 5665 1415 5685 1435
rect 5665 1365 5685 1385
rect 5665 1315 5685 1335
rect 5665 1265 5685 1285
rect 5665 1215 5685 1235
rect 5665 1165 5685 1185
rect 5665 1115 5685 1135
rect 5665 1065 5685 1085
rect 5665 1015 5685 1035
rect 5665 965 5685 985
rect 5665 915 5685 935
rect 5965 1565 5985 1585
rect 5965 1515 5985 1535
rect 5965 1465 5985 1485
rect 5965 1415 5985 1435
rect 5965 1365 5985 1385
rect 5965 1315 5985 1335
rect 5965 1265 5985 1285
rect 5965 1215 5985 1235
rect 5965 1165 5985 1185
rect 5965 1115 5985 1135
rect 5965 1065 5985 1085
rect 5965 1015 5985 1035
rect 5965 965 5985 985
rect 5965 915 5985 935
rect 6265 1565 6285 1585
rect 6265 1515 6285 1535
rect 6265 1465 6285 1485
rect 6265 1415 6285 1435
rect 6265 1365 6285 1385
rect 6265 1315 6285 1335
rect 6265 1265 6285 1285
rect 6265 1215 6285 1235
rect 6265 1165 6285 1185
rect 6265 1115 6285 1135
rect 6265 1065 6285 1085
rect 6265 1015 6285 1035
rect 6265 965 6285 985
rect 6265 915 6285 935
rect 6565 1565 6585 1585
rect 6565 1515 6585 1535
rect 6565 1465 6585 1485
rect 6565 1415 6585 1435
rect 6565 1365 6585 1385
rect 6565 1315 6585 1335
rect 6565 1265 6585 1285
rect 6565 1215 6585 1235
rect 6565 1165 6585 1185
rect 6565 1115 6585 1135
rect 6565 1065 6585 1085
rect 6565 1015 6585 1035
rect 6565 965 6585 985
rect 6565 915 6585 935
rect 6865 1565 6885 1585
rect 6865 1515 6885 1535
rect 6865 1465 6885 1485
rect 6865 1415 6885 1435
rect 6865 1365 6885 1385
rect 6865 1315 6885 1335
rect 6865 1265 6885 1285
rect 6865 1215 6885 1235
rect 6865 1165 6885 1185
rect 6865 1115 6885 1135
rect 6865 1065 6885 1085
rect 6865 1015 6885 1035
rect 6865 965 6885 985
rect 6865 915 6885 935
rect 7165 1565 7185 1585
rect 7165 1515 7185 1535
rect 7165 1465 7185 1485
rect 7165 1415 7185 1435
rect 7165 1365 7185 1385
rect 7165 1315 7185 1335
rect 7165 1265 7185 1285
rect 7165 1215 7185 1235
rect 7165 1165 7185 1185
rect 7165 1115 7185 1135
rect 7165 1065 7185 1085
rect 7165 1015 7185 1035
rect 7165 965 7185 985
rect 7165 915 7185 935
rect 8365 1565 8385 1585
rect 8365 1515 8385 1535
rect 8365 1465 8385 1485
rect 8365 1415 8385 1435
rect 8365 1365 8385 1385
rect 8365 1315 8385 1335
rect 8365 1265 8385 1285
rect 8365 1215 8385 1235
rect 8365 1165 8385 1185
rect 8365 1115 8385 1135
rect 8365 1065 8385 1085
rect 8365 1015 8385 1035
rect 8365 965 8385 985
rect 8365 915 8385 935
rect 9565 1565 9585 1585
rect 9565 1515 9585 1535
rect 9565 1465 9585 1485
rect 9565 1415 9585 1435
rect 9565 1365 9585 1385
rect 9565 1315 9585 1335
rect 9565 1265 9585 1285
rect 9565 1215 9585 1235
rect 9565 1165 9585 1185
rect 9565 1115 9585 1135
rect 9565 1065 9585 1085
rect 9565 1015 9585 1035
rect 9565 965 9585 985
rect 9565 915 9585 935
rect 10765 1565 10785 1585
rect 10765 1515 10785 1535
rect 10765 1465 10785 1485
rect 10765 1415 10785 1435
rect 10765 1365 10785 1385
rect 10765 1315 10785 1335
rect 10765 1265 10785 1285
rect 10765 1215 10785 1235
rect 10765 1165 10785 1185
rect 10765 1115 10785 1135
rect 10765 1065 10785 1085
rect 10765 1015 10785 1035
rect 10765 965 10785 985
rect 10765 915 10785 935
rect 11965 1565 11985 1585
rect 11965 1515 11985 1535
rect 11965 1465 11985 1485
rect 11965 1415 11985 1435
rect 11965 1365 11985 1385
rect 11965 1315 11985 1335
rect 11965 1265 11985 1285
rect 11965 1215 11985 1235
rect 11965 1165 11985 1185
rect 11965 1115 11985 1135
rect 11965 1065 11985 1085
rect 11965 1015 11985 1035
rect 11965 965 11985 985
rect 11965 915 11985 935
rect 12265 1565 12285 1585
rect 12265 1515 12285 1535
rect 12265 1465 12285 1485
rect 12265 1415 12285 1435
rect 12265 1365 12285 1385
rect 12265 1315 12285 1335
rect 12265 1265 12285 1285
rect 12265 1215 12285 1235
rect 12265 1165 12285 1185
rect 12265 1115 12285 1135
rect 12265 1065 12285 1085
rect 12265 1015 12285 1035
rect 12265 965 12285 985
rect 12265 915 12285 935
rect 12565 1565 12585 1585
rect 12565 1515 12585 1535
rect 12565 1465 12585 1485
rect 12565 1415 12585 1435
rect 12565 1365 12585 1385
rect 12565 1315 12585 1335
rect 12565 1265 12585 1285
rect 12565 1215 12585 1235
rect 12565 1165 12585 1185
rect 12565 1115 12585 1135
rect 12565 1065 12585 1085
rect 12565 1015 12585 1035
rect 12565 965 12585 985
rect 12565 915 12585 935
rect 12865 1565 12885 1585
rect 12865 1515 12885 1535
rect 12865 1465 12885 1485
rect 12865 1415 12885 1435
rect 12865 1365 12885 1385
rect 12865 1315 12885 1335
rect 12865 1265 12885 1285
rect 12865 1215 12885 1235
rect 12865 1165 12885 1185
rect 12865 1115 12885 1135
rect 12865 1065 12885 1085
rect 12865 1015 12885 1035
rect 12865 965 12885 985
rect 12865 915 12885 935
rect 13165 1565 13185 1585
rect 13165 1515 13185 1535
rect 13165 1465 13185 1485
rect 13165 1415 13185 1435
rect 13165 1365 13185 1385
rect 13165 1315 13185 1335
rect 13165 1265 13185 1285
rect 13165 1215 13185 1235
rect 13165 1165 13185 1185
rect 13165 1115 13185 1135
rect 13165 1065 13185 1085
rect 13165 1015 13185 1035
rect 13165 965 13185 985
rect 13165 915 13185 935
rect 13465 1565 13485 1585
rect 13465 1515 13485 1535
rect 13465 1465 13485 1485
rect 13465 1415 13485 1435
rect 13465 1365 13485 1385
rect 13465 1315 13485 1335
rect 13465 1265 13485 1285
rect 13465 1215 13485 1235
rect 13465 1165 13485 1185
rect 13465 1115 13485 1135
rect 13465 1065 13485 1085
rect 13465 1015 13485 1035
rect 13465 965 13485 985
rect 13465 915 13485 935
rect 13765 1565 13785 1585
rect 13765 1515 13785 1535
rect 13765 1465 13785 1485
rect 13765 1415 13785 1435
rect 13765 1365 13785 1385
rect 13765 1315 13785 1335
rect 13765 1265 13785 1285
rect 13765 1215 13785 1235
rect 13765 1165 13785 1185
rect 13765 1115 13785 1135
rect 13765 1065 13785 1085
rect 13765 1015 13785 1035
rect 13765 965 13785 985
rect 13765 915 13785 935
rect 14065 1565 14085 1585
rect 14065 1515 14085 1535
rect 14065 1465 14085 1485
rect 14065 1415 14085 1435
rect 14065 1365 14085 1385
rect 14065 1315 14085 1335
rect 14065 1265 14085 1285
rect 14065 1215 14085 1235
rect 14065 1165 14085 1185
rect 14065 1115 14085 1135
rect 14065 1065 14085 1085
rect 14065 1015 14085 1035
rect 14065 965 14085 985
rect 14065 915 14085 935
rect 14365 1565 14385 1585
rect 14365 1515 14385 1535
rect 14365 1465 14385 1485
rect 14365 1415 14385 1435
rect 14365 1365 14385 1385
rect 14365 1315 14385 1335
rect 14365 1265 14385 1285
rect 14365 1215 14385 1235
rect 14365 1165 14385 1185
rect 14365 1115 14385 1135
rect 14365 1065 14385 1085
rect 14365 1015 14385 1035
rect 14365 965 14385 985
rect 14365 915 14385 935
rect 15565 1565 15585 1585
rect 15565 1515 15585 1535
rect 15565 1465 15585 1485
rect 15565 1415 15585 1435
rect 15565 1365 15585 1385
rect 15565 1315 15585 1335
rect 15565 1265 15585 1285
rect 15565 1215 15585 1235
rect 15565 1165 15585 1185
rect 15565 1115 15585 1135
rect 15565 1065 15585 1085
rect 15565 1015 15585 1035
rect 15565 965 15585 985
rect 15565 915 15585 935
rect 16765 1565 16785 1585
rect 16765 1515 16785 1535
rect 16765 1465 16785 1485
rect 16765 1415 16785 1435
rect 16765 1365 16785 1385
rect 16765 1315 16785 1335
rect 16765 1265 16785 1285
rect 16765 1215 16785 1235
rect 16765 1165 16785 1185
rect 16765 1115 16785 1135
rect 16765 1065 16785 1085
rect 16765 1015 16785 1035
rect 16765 965 16785 985
rect 16765 915 16785 935
rect 17965 1565 17985 1585
rect 17965 1515 17985 1535
rect 17965 1465 17985 1485
rect 17965 1415 17985 1435
rect 17965 1365 17985 1385
rect 17965 1315 17985 1335
rect 17965 1265 17985 1285
rect 17965 1215 17985 1235
rect 17965 1165 17985 1185
rect 17965 1115 17985 1135
rect 17965 1065 17985 1085
rect 17965 1015 17985 1035
rect 17965 965 17985 985
rect 17965 915 17985 935
rect 19165 1565 19185 1585
rect 19165 1515 19185 1535
rect 19165 1465 19185 1485
rect 19165 1415 19185 1435
rect 19165 1365 19185 1385
rect 19165 1315 19185 1335
rect 19165 1265 19185 1285
rect 19165 1215 19185 1235
rect 19165 1165 19185 1185
rect 19165 1115 19185 1135
rect 19165 1065 19185 1085
rect 19165 1015 19185 1035
rect 19165 965 19185 985
rect 19165 915 19185 935
rect 20365 1565 20385 1585
rect 20365 1515 20385 1535
rect 20365 1465 20385 1485
rect 20365 1415 20385 1435
rect 20365 1365 20385 1385
rect 20365 1315 20385 1335
rect 20365 1265 20385 1285
rect 20365 1215 20385 1235
rect 20365 1165 20385 1185
rect 20365 1115 20385 1135
rect 20365 1065 20385 1085
rect 20365 1015 20385 1035
rect 20365 965 20385 985
rect 20365 915 20385 935
rect -635 715 -615 735
rect -635 665 -615 685
rect -635 615 -615 635
rect -635 565 -615 585
rect -635 515 -615 535
rect -635 465 -615 485
rect -635 415 -615 435
rect -635 365 -615 385
rect -635 315 -615 335
rect -635 265 -615 285
rect -635 215 -615 235
rect -635 165 -615 185
rect -635 115 -615 135
rect -635 65 -615 85
rect -485 715 -465 735
rect -485 665 -465 685
rect -485 615 -465 635
rect -485 565 -465 585
rect -485 515 -465 535
rect -485 465 -465 485
rect -485 415 -465 435
rect -485 365 -465 385
rect -485 315 -465 335
rect -485 265 -465 285
rect -485 215 -465 235
rect -485 165 -465 185
rect -485 115 -465 135
rect -485 65 -465 85
rect -335 715 -315 735
rect -335 665 -315 685
rect -335 615 -315 635
rect -335 565 -315 585
rect -335 515 -315 535
rect -335 465 -315 485
rect -335 415 -315 435
rect -335 365 -315 385
rect -335 315 -315 335
rect -335 265 -315 285
rect -335 215 -315 235
rect -335 165 -315 185
rect -335 115 -315 135
rect -335 65 -315 85
rect -185 715 -165 735
rect -185 665 -165 685
rect -185 615 -165 635
rect -185 565 -165 585
rect -185 515 -165 535
rect -185 465 -165 485
rect -185 415 -165 435
rect -185 365 -165 385
rect -185 315 -165 335
rect -185 265 -165 285
rect -185 215 -165 235
rect -185 165 -165 185
rect -185 115 -165 135
rect -185 65 -165 85
rect -35 715 -15 735
rect -35 665 -15 685
rect -35 615 -15 635
rect -35 565 -15 585
rect -35 515 -15 535
rect -35 465 -15 485
rect -35 415 -15 435
rect -35 365 -15 385
rect -35 315 -15 335
rect -35 265 -15 285
rect -35 215 -15 235
rect -35 165 -15 185
rect -35 115 -15 135
rect -35 65 -15 85
rect 1165 715 1185 735
rect 1165 665 1185 685
rect 1165 615 1185 635
rect 1165 565 1185 585
rect 1165 515 1185 535
rect 1165 465 1185 485
rect 1165 415 1185 435
rect 1165 365 1185 385
rect 1165 315 1185 335
rect 1165 265 1185 285
rect 1165 215 1185 235
rect 1165 165 1185 185
rect 1165 115 1185 135
rect 1165 65 1185 85
rect 1465 715 1485 735
rect 1465 665 1485 685
rect 1465 615 1485 635
rect 1465 565 1485 585
rect 1465 515 1485 535
rect 1465 465 1485 485
rect 1465 415 1485 435
rect 1465 365 1485 385
rect 1465 315 1485 335
rect 1465 265 1485 285
rect 1465 215 1485 235
rect 1465 165 1485 185
rect 1465 115 1485 135
rect 1465 65 1485 85
rect 1765 715 1785 735
rect 1765 665 1785 685
rect 1765 615 1785 635
rect 1765 565 1785 585
rect 1765 515 1785 535
rect 1765 465 1785 485
rect 1765 415 1785 435
rect 1765 365 1785 385
rect 1765 315 1785 335
rect 1765 265 1785 285
rect 1765 215 1785 235
rect 1765 165 1785 185
rect 1765 115 1785 135
rect 1765 65 1785 85
rect 2065 715 2085 735
rect 2065 665 2085 685
rect 2065 615 2085 635
rect 2065 565 2085 585
rect 2065 515 2085 535
rect 2065 465 2085 485
rect 2065 415 2085 435
rect 2065 365 2085 385
rect 2065 315 2085 335
rect 2065 265 2085 285
rect 2065 215 2085 235
rect 2065 165 2085 185
rect 2065 115 2085 135
rect 2065 65 2085 85
rect 2365 715 2385 735
rect 2365 665 2385 685
rect 2365 615 2385 635
rect 2365 565 2385 585
rect 2365 515 2385 535
rect 2365 465 2385 485
rect 2365 415 2385 435
rect 2365 365 2385 385
rect 2365 315 2385 335
rect 2365 265 2385 285
rect 2365 215 2385 235
rect 2365 165 2385 185
rect 2365 115 2385 135
rect 2365 65 2385 85
rect 2665 715 2685 735
rect 2665 665 2685 685
rect 2665 615 2685 635
rect 2665 565 2685 585
rect 2665 515 2685 535
rect 2665 465 2685 485
rect 2665 415 2685 435
rect 2665 365 2685 385
rect 2665 315 2685 335
rect 2665 265 2685 285
rect 2665 215 2685 235
rect 2665 165 2685 185
rect 2665 115 2685 135
rect 2665 65 2685 85
rect 2965 715 2985 735
rect 2965 665 2985 685
rect 2965 615 2985 635
rect 2965 565 2985 585
rect 2965 515 2985 535
rect 2965 465 2985 485
rect 2965 415 2985 435
rect 2965 365 2985 385
rect 2965 315 2985 335
rect 2965 265 2985 285
rect 2965 215 2985 235
rect 2965 165 2985 185
rect 2965 115 2985 135
rect 2965 65 2985 85
rect 3265 715 3285 735
rect 3265 665 3285 685
rect 3265 615 3285 635
rect 3265 565 3285 585
rect 3265 515 3285 535
rect 3265 465 3285 485
rect 3265 415 3285 435
rect 3265 365 3285 385
rect 3265 315 3285 335
rect 3265 265 3285 285
rect 3265 215 3285 235
rect 3265 165 3285 185
rect 3265 115 3285 135
rect 3265 65 3285 85
rect 3565 715 3585 735
rect 3565 665 3585 685
rect 3565 615 3585 635
rect 3565 565 3585 585
rect 3565 515 3585 535
rect 3565 465 3585 485
rect 3565 415 3585 435
rect 3565 365 3585 385
rect 3565 315 3585 335
rect 3565 265 3585 285
rect 3565 215 3585 235
rect 3565 165 3585 185
rect 3565 115 3585 135
rect 3565 65 3585 85
rect 3715 715 3735 735
rect 3715 665 3735 685
rect 3715 615 3735 635
rect 3715 565 3735 585
rect 3715 515 3735 535
rect 3715 465 3735 485
rect 3715 415 3735 435
rect 3715 365 3735 385
rect 3715 315 3735 335
rect 3715 265 3735 285
rect 3715 215 3735 235
rect 3715 165 3735 185
rect 3715 115 3735 135
rect 3715 65 3735 85
rect 3865 715 3885 735
rect 3865 665 3885 685
rect 3865 615 3885 635
rect 3865 565 3885 585
rect 3865 515 3885 535
rect 3865 465 3885 485
rect 3865 415 3885 435
rect 3865 365 3885 385
rect 3865 315 3885 335
rect 3865 265 3885 285
rect 3865 215 3885 235
rect 3865 165 3885 185
rect 3865 115 3885 135
rect 3865 65 3885 85
rect 4015 715 4035 735
rect 4015 665 4035 685
rect 4015 615 4035 635
rect 4015 565 4035 585
rect 4015 515 4035 535
rect 4015 465 4035 485
rect 4015 415 4035 435
rect 4015 365 4035 385
rect 4015 315 4035 335
rect 4015 265 4035 285
rect 4015 215 4035 235
rect 4015 165 4035 185
rect 4015 115 4035 135
rect 4015 65 4035 85
rect 4165 715 4185 735
rect 4165 665 4185 685
rect 4165 615 4185 635
rect 4165 565 4185 585
rect 4165 515 4185 535
rect 4165 465 4185 485
rect 4165 415 4185 435
rect 4165 365 4185 385
rect 4165 315 4185 335
rect 4165 265 4185 285
rect 4165 215 4185 235
rect 4165 165 4185 185
rect 4165 115 4185 135
rect 4165 65 4185 85
rect 4315 715 4335 735
rect 4315 665 4335 685
rect 4315 615 4335 635
rect 4315 565 4335 585
rect 4315 515 4335 535
rect 4315 465 4335 485
rect 4315 415 4335 435
rect 4315 365 4335 385
rect 4315 315 4335 335
rect 4315 265 4335 285
rect 4315 215 4335 235
rect 4315 165 4335 185
rect 4315 115 4335 135
rect 4315 65 4335 85
rect 4465 715 4485 735
rect 4465 665 4485 685
rect 4465 615 4485 635
rect 4465 565 4485 585
rect 4465 515 4485 535
rect 4465 465 4485 485
rect 4465 415 4485 435
rect 4465 365 4485 385
rect 4465 315 4485 335
rect 4465 265 4485 285
rect 4465 215 4485 235
rect 4465 165 4485 185
rect 4465 115 4485 135
rect 4465 65 4485 85
rect 4615 715 4635 735
rect 4615 665 4635 685
rect 4615 615 4635 635
rect 4615 565 4635 585
rect 4615 515 4635 535
rect 4615 465 4635 485
rect 4615 415 4635 435
rect 4615 365 4635 385
rect 4615 315 4635 335
rect 4615 265 4635 285
rect 4615 215 4635 235
rect 4615 165 4635 185
rect 4615 115 4635 135
rect 4615 65 4635 85
rect 4765 715 4785 735
rect 4765 665 4785 685
rect 4765 615 4785 635
rect 4765 565 4785 585
rect 4765 515 4785 535
rect 4765 465 4785 485
rect 4765 415 4785 435
rect 4765 365 4785 385
rect 4765 315 4785 335
rect 4765 265 4785 285
rect 4765 215 4785 235
rect 4765 165 4785 185
rect 4765 115 4785 135
rect 4765 65 4785 85
rect 5065 715 5085 735
rect 5065 665 5085 685
rect 5065 615 5085 635
rect 5065 565 5085 585
rect 5065 515 5085 535
rect 5065 465 5085 485
rect 5065 415 5085 435
rect 5065 365 5085 385
rect 5065 315 5085 335
rect 5065 265 5085 285
rect 5065 215 5085 235
rect 5065 165 5085 185
rect 5065 115 5085 135
rect 5065 65 5085 85
rect 5365 715 5385 735
rect 5365 665 5385 685
rect 5365 615 5385 635
rect 5365 565 5385 585
rect 5365 515 5385 535
rect 5365 465 5385 485
rect 5365 415 5385 435
rect 5365 365 5385 385
rect 5365 315 5385 335
rect 5365 265 5385 285
rect 5365 215 5385 235
rect 5365 165 5385 185
rect 5365 115 5385 135
rect 5365 65 5385 85
rect 5665 715 5685 735
rect 5665 665 5685 685
rect 5665 615 5685 635
rect 5665 565 5685 585
rect 5665 515 5685 535
rect 5665 465 5685 485
rect 5665 415 5685 435
rect 5665 365 5685 385
rect 5665 315 5685 335
rect 5665 265 5685 285
rect 5665 215 5685 235
rect 5665 165 5685 185
rect 5665 115 5685 135
rect 5665 65 5685 85
rect 5965 715 5985 735
rect 5965 665 5985 685
rect 5965 615 5985 635
rect 5965 565 5985 585
rect 5965 515 5985 535
rect 5965 465 5985 485
rect 5965 415 5985 435
rect 5965 365 5985 385
rect 5965 315 5985 335
rect 5965 265 5985 285
rect 5965 215 5985 235
rect 5965 165 5985 185
rect 5965 115 5985 135
rect 5965 65 5985 85
rect 6265 715 6285 735
rect 6265 665 6285 685
rect 6265 615 6285 635
rect 6265 565 6285 585
rect 6265 515 6285 535
rect 6265 465 6285 485
rect 6265 415 6285 435
rect 6265 365 6285 385
rect 6265 315 6285 335
rect 6265 265 6285 285
rect 6265 215 6285 235
rect 6265 165 6285 185
rect 6265 115 6285 135
rect 6265 65 6285 85
rect 6565 715 6585 735
rect 6565 665 6585 685
rect 6565 615 6585 635
rect 6565 565 6585 585
rect 6565 515 6585 535
rect 6565 465 6585 485
rect 6565 415 6585 435
rect 6565 365 6585 385
rect 6565 315 6585 335
rect 6565 265 6585 285
rect 6565 215 6585 235
rect 6565 165 6585 185
rect 6565 115 6585 135
rect 6565 65 6585 85
rect 6865 715 6885 735
rect 6865 665 6885 685
rect 6865 615 6885 635
rect 6865 565 6885 585
rect 6865 515 6885 535
rect 6865 465 6885 485
rect 6865 415 6885 435
rect 6865 365 6885 385
rect 6865 315 6885 335
rect 6865 265 6885 285
rect 6865 215 6885 235
rect 6865 165 6885 185
rect 6865 115 6885 135
rect 6865 65 6885 85
rect 7165 715 7185 735
rect 7165 665 7185 685
rect 7165 615 7185 635
rect 7165 565 7185 585
rect 7165 515 7185 535
rect 7165 465 7185 485
rect 7165 415 7185 435
rect 7165 365 7185 385
rect 7165 315 7185 335
rect 7165 265 7185 285
rect 7165 215 7185 235
rect 7165 165 7185 185
rect 7165 115 7185 135
rect 7165 65 7185 85
rect 8365 715 8385 735
rect 8365 665 8385 685
rect 8365 615 8385 635
rect 8365 565 8385 585
rect 8365 515 8385 535
rect 8365 465 8385 485
rect 8365 415 8385 435
rect 8365 365 8385 385
rect 8365 315 8385 335
rect 8365 265 8385 285
rect 8365 215 8385 235
rect 8365 165 8385 185
rect 8365 115 8385 135
rect 8365 65 8385 85
rect 9565 715 9585 735
rect 9565 665 9585 685
rect 9565 615 9585 635
rect 9565 565 9585 585
rect 9565 515 9585 535
rect 9565 465 9585 485
rect 9565 415 9585 435
rect 9565 365 9585 385
rect 9565 315 9585 335
rect 9565 265 9585 285
rect 9565 215 9585 235
rect 9565 165 9585 185
rect 9565 115 9585 135
rect 9565 65 9585 85
rect 10765 715 10785 735
rect 10765 665 10785 685
rect 10765 615 10785 635
rect 10765 565 10785 585
rect 10765 515 10785 535
rect 10765 465 10785 485
rect 10765 415 10785 435
rect 10765 365 10785 385
rect 10765 315 10785 335
rect 10765 265 10785 285
rect 10765 215 10785 235
rect 10765 165 10785 185
rect 10765 115 10785 135
rect 10765 65 10785 85
rect 11965 715 11985 735
rect 11965 665 11985 685
rect 11965 615 11985 635
rect 11965 565 11985 585
rect 11965 515 11985 535
rect 11965 465 11985 485
rect 11965 415 11985 435
rect 11965 365 11985 385
rect 11965 315 11985 335
rect 11965 265 11985 285
rect 11965 215 11985 235
rect 11965 165 11985 185
rect 11965 115 11985 135
rect 11965 65 11985 85
rect 12265 715 12285 735
rect 12265 665 12285 685
rect 12265 615 12285 635
rect 12265 565 12285 585
rect 12265 515 12285 535
rect 12265 465 12285 485
rect 12265 415 12285 435
rect 12265 365 12285 385
rect 12265 315 12285 335
rect 12265 265 12285 285
rect 12265 215 12285 235
rect 12265 165 12285 185
rect 12265 115 12285 135
rect 12265 65 12285 85
rect 12565 715 12585 735
rect 12565 665 12585 685
rect 12565 615 12585 635
rect 12565 565 12585 585
rect 12565 515 12585 535
rect 12565 465 12585 485
rect 12565 415 12585 435
rect 12565 365 12585 385
rect 12565 315 12585 335
rect 12565 265 12585 285
rect 12565 215 12585 235
rect 12565 165 12585 185
rect 12565 115 12585 135
rect 12565 65 12585 85
rect 12865 715 12885 735
rect 12865 665 12885 685
rect 12865 615 12885 635
rect 12865 565 12885 585
rect 12865 515 12885 535
rect 12865 465 12885 485
rect 12865 415 12885 435
rect 12865 365 12885 385
rect 12865 315 12885 335
rect 12865 265 12885 285
rect 12865 215 12885 235
rect 12865 165 12885 185
rect 12865 115 12885 135
rect 12865 65 12885 85
rect 13165 715 13185 735
rect 13165 665 13185 685
rect 13165 615 13185 635
rect 13165 565 13185 585
rect 13165 515 13185 535
rect 13165 465 13185 485
rect 13165 415 13185 435
rect 13165 365 13185 385
rect 13165 315 13185 335
rect 13165 265 13185 285
rect 13165 215 13185 235
rect 13165 165 13185 185
rect 13165 115 13185 135
rect 13165 65 13185 85
rect 13465 715 13485 735
rect 13465 665 13485 685
rect 13465 615 13485 635
rect 13465 565 13485 585
rect 13465 515 13485 535
rect 13465 465 13485 485
rect 13465 415 13485 435
rect 13465 365 13485 385
rect 13465 315 13485 335
rect 13465 265 13485 285
rect 13465 215 13485 235
rect 13465 165 13485 185
rect 13465 115 13485 135
rect 13465 65 13485 85
rect 13765 715 13785 735
rect 13765 665 13785 685
rect 13765 615 13785 635
rect 13765 565 13785 585
rect 13765 515 13785 535
rect 13765 465 13785 485
rect 13765 415 13785 435
rect 13765 365 13785 385
rect 13765 315 13785 335
rect 13765 265 13785 285
rect 13765 215 13785 235
rect 13765 165 13785 185
rect 13765 115 13785 135
rect 13765 65 13785 85
rect 14065 715 14085 735
rect 14065 665 14085 685
rect 14065 615 14085 635
rect 14065 565 14085 585
rect 14065 515 14085 535
rect 14065 465 14085 485
rect 14065 415 14085 435
rect 14065 365 14085 385
rect 14065 315 14085 335
rect 14065 265 14085 285
rect 14065 215 14085 235
rect 14065 165 14085 185
rect 14065 115 14085 135
rect 14065 65 14085 85
rect 14365 715 14385 735
rect 14365 665 14385 685
rect 14365 615 14385 635
rect 14365 565 14385 585
rect 14365 515 14385 535
rect 14365 465 14385 485
rect 14365 415 14385 435
rect 14365 365 14385 385
rect 14365 315 14385 335
rect 14365 265 14385 285
rect 14365 215 14385 235
rect 14365 165 14385 185
rect 14365 115 14385 135
rect 14365 65 14385 85
rect 15565 715 15585 735
rect 15565 665 15585 685
rect 15565 615 15585 635
rect 15565 565 15585 585
rect 15565 515 15585 535
rect 15565 465 15585 485
rect 15565 415 15585 435
rect 15565 365 15585 385
rect 15565 315 15585 335
rect 15565 265 15585 285
rect 15565 215 15585 235
rect 15565 165 15585 185
rect 15565 115 15585 135
rect 15565 65 15585 85
rect 16765 715 16785 735
rect 16765 665 16785 685
rect 16765 615 16785 635
rect 16765 565 16785 585
rect 16765 515 16785 535
rect 16765 465 16785 485
rect 16765 415 16785 435
rect 16765 365 16785 385
rect 16765 315 16785 335
rect 16765 265 16785 285
rect 16765 215 16785 235
rect 16765 165 16785 185
rect 16765 115 16785 135
rect 16765 65 16785 85
rect 17965 715 17985 735
rect 17965 665 17985 685
rect 17965 615 17985 635
rect 17965 565 17985 585
rect 17965 515 17985 535
rect 17965 465 17985 485
rect 17965 415 17985 435
rect 17965 365 17985 385
rect 17965 315 17985 335
rect 17965 265 17985 285
rect 17965 215 17985 235
rect 17965 165 17985 185
rect 17965 115 17985 135
rect 17965 65 17985 85
rect 19165 715 19185 735
rect 19165 665 19185 685
rect 19165 615 19185 635
rect 19165 565 19185 585
rect 19165 515 19185 535
rect 19165 465 19185 485
rect 19165 415 19185 435
rect 19165 365 19185 385
rect 19165 315 19185 335
rect 19165 265 19185 285
rect 19165 215 19185 235
rect 19165 165 19185 185
rect 19165 115 19185 135
rect 19165 65 19185 85
rect 20365 715 20385 735
rect 20365 665 20385 685
rect 20365 615 20385 635
rect 20365 565 20385 585
rect 20365 515 20385 535
rect 20365 465 20385 485
rect 20365 415 20385 435
rect 20365 365 20385 385
rect 20365 315 20385 335
rect 20365 265 20385 285
rect 20365 215 20385 235
rect 20365 165 20385 185
rect 20365 115 20385 135
rect 20365 65 20385 85
rect -635 -135 -615 -115
rect -635 -185 -615 -165
rect -635 -235 -615 -215
rect -635 -285 -615 -265
rect -635 -335 -615 -315
rect -635 -385 -615 -365
rect -635 -435 -615 -415
rect -635 -485 -615 -465
rect -635 -535 -615 -515
rect -635 -585 -615 -565
rect -635 -635 -615 -615
rect -635 -685 -615 -665
rect -635 -735 -615 -715
rect -635 -785 -615 -765
rect -485 -135 -465 -115
rect -485 -185 -465 -165
rect -485 -235 -465 -215
rect -485 -285 -465 -265
rect -485 -335 -465 -315
rect -485 -385 -465 -365
rect -485 -435 -465 -415
rect -485 -485 -465 -465
rect -485 -535 -465 -515
rect -485 -585 -465 -565
rect -485 -635 -465 -615
rect -485 -685 -465 -665
rect -485 -735 -465 -715
rect -485 -785 -465 -765
rect -335 -135 -315 -115
rect -335 -185 -315 -165
rect -335 -235 -315 -215
rect -335 -285 -315 -265
rect -335 -335 -315 -315
rect -335 -385 -315 -365
rect -335 -435 -315 -415
rect -335 -485 -315 -465
rect -335 -535 -315 -515
rect -335 -585 -315 -565
rect -335 -635 -315 -615
rect -335 -685 -315 -665
rect -335 -735 -315 -715
rect -335 -785 -315 -765
rect -185 -135 -165 -115
rect -185 -185 -165 -165
rect -185 -235 -165 -215
rect -185 -285 -165 -265
rect -185 -335 -165 -315
rect -185 -385 -165 -365
rect -185 -435 -165 -415
rect -185 -485 -165 -465
rect -185 -535 -165 -515
rect -185 -585 -165 -565
rect -185 -635 -165 -615
rect -185 -685 -165 -665
rect -185 -735 -165 -715
rect -185 -785 -165 -765
rect -35 -135 -15 -115
rect -35 -185 -15 -165
rect -35 -235 -15 -215
rect -35 -285 -15 -265
rect -35 -335 -15 -315
rect -35 -385 -15 -365
rect -35 -435 -15 -415
rect -35 -485 -15 -465
rect -35 -535 -15 -515
rect -35 -585 -15 -565
rect -35 -635 -15 -615
rect -35 -685 -15 -665
rect -35 -735 -15 -715
rect -35 -785 -15 -765
rect 1165 -135 1185 -115
rect 1165 -185 1185 -165
rect 1165 -235 1185 -215
rect 1165 -285 1185 -265
rect 1165 -335 1185 -315
rect 1165 -385 1185 -365
rect 1165 -435 1185 -415
rect 1165 -485 1185 -465
rect 1165 -535 1185 -515
rect 1165 -585 1185 -565
rect 1165 -635 1185 -615
rect 1165 -685 1185 -665
rect 1165 -735 1185 -715
rect 1165 -785 1185 -765
rect 1465 -135 1485 -115
rect 1465 -185 1485 -165
rect 1465 -235 1485 -215
rect 1465 -285 1485 -265
rect 1465 -335 1485 -315
rect 1465 -385 1485 -365
rect 1465 -435 1485 -415
rect 1465 -485 1485 -465
rect 1465 -535 1485 -515
rect 1465 -585 1485 -565
rect 1465 -635 1485 -615
rect 1465 -685 1485 -665
rect 1465 -735 1485 -715
rect 1465 -785 1485 -765
rect 1765 -135 1785 -115
rect 1765 -185 1785 -165
rect 1765 -235 1785 -215
rect 1765 -285 1785 -265
rect 1765 -335 1785 -315
rect 1765 -385 1785 -365
rect 1765 -435 1785 -415
rect 1765 -485 1785 -465
rect 1765 -535 1785 -515
rect 1765 -585 1785 -565
rect 1765 -635 1785 -615
rect 1765 -685 1785 -665
rect 1765 -735 1785 -715
rect 1765 -785 1785 -765
rect 2065 -135 2085 -115
rect 2065 -185 2085 -165
rect 2065 -235 2085 -215
rect 2065 -285 2085 -265
rect 2065 -335 2085 -315
rect 2065 -385 2085 -365
rect 2065 -435 2085 -415
rect 2065 -485 2085 -465
rect 2065 -535 2085 -515
rect 2065 -585 2085 -565
rect 2065 -635 2085 -615
rect 2065 -685 2085 -665
rect 2065 -735 2085 -715
rect 2065 -785 2085 -765
rect 2365 -135 2385 -115
rect 2365 -185 2385 -165
rect 2365 -235 2385 -215
rect 2365 -285 2385 -265
rect 2365 -335 2385 -315
rect 2365 -385 2385 -365
rect 2365 -435 2385 -415
rect 2365 -485 2385 -465
rect 2365 -535 2385 -515
rect 2365 -585 2385 -565
rect 2365 -635 2385 -615
rect 2365 -685 2385 -665
rect 2365 -735 2385 -715
rect 2365 -785 2385 -765
rect 2665 -135 2685 -115
rect 2665 -185 2685 -165
rect 2665 -235 2685 -215
rect 2665 -285 2685 -265
rect 2665 -335 2685 -315
rect 2665 -385 2685 -365
rect 2665 -435 2685 -415
rect 2665 -485 2685 -465
rect 2665 -535 2685 -515
rect 2665 -585 2685 -565
rect 2665 -635 2685 -615
rect 2665 -685 2685 -665
rect 2665 -735 2685 -715
rect 2665 -785 2685 -765
rect 2965 -135 2985 -115
rect 2965 -185 2985 -165
rect 2965 -235 2985 -215
rect 2965 -285 2985 -265
rect 2965 -335 2985 -315
rect 2965 -385 2985 -365
rect 2965 -435 2985 -415
rect 2965 -485 2985 -465
rect 2965 -535 2985 -515
rect 2965 -585 2985 -565
rect 2965 -635 2985 -615
rect 2965 -685 2985 -665
rect 2965 -735 2985 -715
rect 2965 -785 2985 -765
rect 3265 -135 3285 -115
rect 3265 -185 3285 -165
rect 3265 -235 3285 -215
rect 3265 -285 3285 -265
rect 3265 -335 3285 -315
rect 3265 -385 3285 -365
rect 3265 -435 3285 -415
rect 3265 -485 3285 -465
rect 3265 -535 3285 -515
rect 3265 -585 3285 -565
rect 3265 -635 3285 -615
rect 3265 -685 3285 -665
rect 3265 -735 3285 -715
rect 3265 -785 3285 -765
rect 3565 -135 3585 -115
rect 3565 -185 3585 -165
rect 3565 -235 3585 -215
rect 3565 -285 3585 -265
rect 3565 -335 3585 -315
rect 3565 -385 3585 -365
rect 3565 -435 3585 -415
rect 3565 -485 3585 -465
rect 3565 -535 3585 -515
rect 3565 -585 3585 -565
rect 3565 -635 3585 -615
rect 3565 -685 3585 -665
rect 3565 -735 3585 -715
rect 3565 -785 3585 -765
rect 3715 -135 3735 -115
rect 3715 -185 3735 -165
rect 3715 -235 3735 -215
rect 3715 -285 3735 -265
rect 3715 -335 3735 -315
rect 3715 -385 3735 -365
rect 3715 -435 3735 -415
rect 3715 -485 3735 -465
rect 3715 -535 3735 -515
rect 3715 -585 3735 -565
rect 3715 -635 3735 -615
rect 3715 -685 3735 -665
rect 3715 -735 3735 -715
rect 3715 -785 3735 -765
rect 3865 -135 3885 -115
rect 3865 -185 3885 -165
rect 3865 -235 3885 -215
rect 3865 -285 3885 -265
rect 3865 -335 3885 -315
rect 3865 -385 3885 -365
rect 3865 -435 3885 -415
rect 3865 -485 3885 -465
rect 3865 -535 3885 -515
rect 3865 -585 3885 -565
rect 3865 -635 3885 -615
rect 3865 -685 3885 -665
rect 3865 -735 3885 -715
rect 3865 -785 3885 -765
rect 4015 -135 4035 -115
rect 4015 -185 4035 -165
rect 4015 -235 4035 -215
rect 4015 -285 4035 -265
rect 4015 -335 4035 -315
rect 4015 -385 4035 -365
rect 4015 -435 4035 -415
rect 4015 -485 4035 -465
rect 4015 -535 4035 -515
rect 4015 -585 4035 -565
rect 4015 -635 4035 -615
rect 4015 -685 4035 -665
rect 4015 -735 4035 -715
rect 4015 -785 4035 -765
rect 4165 -135 4185 -115
rect 4165 -185 4185 -165
rect 4165 -235 4185 -215
rect 4165 -285 4185 -265
rect 4165 -335 4185 -315
rect 4165 -385 4185 -365
rect 4165 -435 4185 -415
rect 4165 -485 4185 -465
rect 4165 -535 4185 -515
rect 4165 -585 4185 -565
rect 4165 -635 4185 -615
rect 4165 -685 4185 -665
rect 4165 -735 4185 -715
rect 4165 -785 4185 -765
rect 4315 -135 4335 -115
rect 4315 -185 4335 -165
rect 4315 -235 4335 -215
rect 4315 -285 4335 -265
rect 4315 -335 4335 -315
rect 4315 -385 4335 -365
rect 4315 -435 4335 -415
rect 4315 -485 4335 -465
rect 4315 -535 4335 -515
rect 4315 -585 4335 -565
rect 4315 -635 4335 -615
rect 4315 -685 4335 -665
rect 4315 -735 4335 -715
rect 4315 -785 4335 -765
rect 4465 -135 4485 -115
rect 4465 -185 4485 -165
rect 4465 -235 4485 -215
rect 4465 -285 4485 -265
rect 4465 -335 4485 -315
rect 4465 -385 4485 -365
rect 4465 -435 4485 -415
rect 4465 -485 4485 -465
rect 4465 -535 4485 -515
rect 4465 -585 4485 -565
rect 4465 -635 4485 -615
rect 4465 -685 4485 -665
rect 4465 -735 4485 -715
rect 4465 -785 4485 -765
rect 4615 -135 4635 -115
rect 4615 -185 4635 -165
rect 4615 -235 4635 -215
rect 4615 -285 4635 -265
rect 4615 -335 4635 -315
rect 4615 -385 4635 -365
rect 4615 -435 4635 -415
rect 4615 -485 4635 -465
rect 4615 -535 4635 -515
rect 4615 -585 4635 -565
rect 4615 -635 4635 -615
rect 4615 -685 4635 -665
rect 4615 -735 4635 -715
rect 4615 -785 4635 -765
rect 4765 -135 4785 -115
rect 4765 -185 4785 -165
rect 4765 -235 4785 -215
rect 4765 -285 4785 -265
rect 4765 -335 4785 -315
rect 4765 -385 4785 -365
rect 4765 -435 4785 -415
rect 4765 -485 4785 -465
rect 4765 -535 4785 -515
rect 4765 -585 4785 -565
rect 4765 -635 4785 -615
rect 4765 -685 4785 -665
rect 4765 -735 4785 -715
rect 4765 -785 4785 -765
rect 5065 -135 5085 -115
rect 5065 -185 5085 -165
rect 5065 -235 5085 -215
rect 5065 -285 5085 -265
rect 5065 -335 5085 -315
rect 5065 -385 5085 -365
rect 5065 -435 5085 -415
rect 5065 -485 5085 -465
rect 5065 -535 5085 -515
rect 5065 -585 5085 -565
rect 5065 -635 5085 -615
rect 5065 -685 5085 -665
rect 5065 -735 5085 -715
rect 5065 -785 5085 -765
rect 5365 -135 5385 -115
rect 5365 -185 5385 -165
rect 5365 -235 5385 -215
rect 5365 -285 5385 -265
rect 5365 -335 5385 -315
rect 5365 -385 5385 -365
rect 5365 -435 5385 -415
rect 5365 -485 5385 -465
rect 5365 -535 5385 -515
rect 5365 -585 5385 -565
rect 5365 -635 5385 -615
rect 5365 -685 5385 -665
rect 5365 -735 5385 -715
rect 5365 -785 5385 -765
rect 5665 -135 5685 -115
rect 5665 -185 5685 -165
rect 5665 -235 5685 -215
rect 5665 -285 5685 -265
rect 5665 -335 5685 -315
rect 5665 -385 5685 -365
rect 5665 -435 5685 -415
rect 5665 -485 5685 -465
rect 5665 -535 5685 -515
rect 5665 -585 5685 -565
rect 5665 -635 5685 -615
rect 5665 -685 5685 -665
rect 5665 -735 5685 -715
rect 5665 -785 5685 -765
rect 5965 -135 5985 -115
rect 5965 -185 5985 -165
rect 5965 -235 5985 -215
rect 5965 -285 5985 -265
rect 5965 -335 5985 -315
rect 5965 -385 5985 -365
rect 5965 -435 5985 -415
rect 5965 -485 5985 -465
rect 5965 -535 5985 -515
rect 5965 -585 5985 -565
rect 5965 -635 5985 -615
rect 5965 -685 5985 -665
rect 5965 -735 5985 -715
rect 5965 -785 5985 -765
rect 6265 -135 6285 -115
rect 6265 -185 6285 -165
rect 6265 -235 6285 -215
rect 6265 -285 6285 -265
rect 6265 -335 6285 -315
rect 6265 -385 6285 -365
rect 6265 -435 6285 -415
rect 6265 -485 6285 -465
rect 6265 -535 6285 -515
rect 6265 -585 6285 -565
rect 6265 -635 6285 -615
rect 6265 -685 6285 -665
rect 6265 -735 6285 -715
rect 6265 -785 6285 -765
rect 6565 -135 6585 -115
rect 6565 -185 6585 -165
rect 6565 -235 6585 -215
rect 6565 -285 6585 -265
rect 6565 -335 6585 -315
rect 6565 -385 6585 -365
rect 6565 -435 6585 -415
rect 6565 -485 6585 -465
rect 6565 -535 6585 -515
rect 6565 -585 6585 -565
rect 6565 -635 6585 -615
rect 6565 -685 6585 -665
rect 6565 -735 6585 -715
rect 6565 -785 6585 -765
rect 6865 -135 6885 -115
rect 6865 -185 6885 -165
rect 6865 -235 6885 -215
rect 6865 -285 6885 -265
rect 6865 -335 6885 -315
rect 6865 -385 6885 -365
rect 6865 -435 6885 -415
rect 6865 -485 6885 -465
rect 6865 -535 6885 -515
rect 6865 -585 6885 -565
rect 6865 -635 6885 -615
rect 6865 -685 6885 -665
rect 6865 -735 6885 -715
rect 6865 -785 6885 -765
rect 7165 -135 7185 -115
rect 7165 -185 7185 -165
rect 7165 -235 7185 -215
rect 7165 -285 7185 -265
rect 7165 -335 7185 -315
rect 7165 -385 7185 -365
rect 7165 -435 7185 -415
rect 7165 -485 7185 -465
rect 7165 -535 7185 -515
rect 7165 -585 7185 -565
rect 7165 -635 7185 -615
rect 7165 -685 7185 -665
rect 7165 -735 7185 -715
rect 7165 -785 7185 -765
rect 8365 -135 8385 -115
rect 8365 -185 8385 -165
rect 8365 -235 8385 -215
rect 8365 -285 8385 -265
rect 8365 -335 8385 -315
rect 8365 -385 8385 -365
rect 8365 -435 8385 -415
rect 8365 -485 8385 -465
rect 8365 -535 8385 -515
rect 8365 -585 8385 -565
rect 8365 -635 8385 -615
rect 8365 -685 8385 -665
rect 8365 -735 8385 -715
rect 8365 -785 8385 -765
rect 9565 -135 9585 -115
rect 9565 -185 9585 -165
rect 9565 -235 9585 -215
rect 9565 -285 9585 -265
rect 9565 -335 9585 -315
rect 9565 -385 9585 -365
rect 9565 -435 9585 -415
rect 9565 -485 9585 -465
rect 9565 -535 9585 -515
rect 9565 -585 9585 -565
rect 9565 -635 9585 -615
rect 9565 -685 9585 -665
rect 9565 -735 9585 -715
rect 9565 -785 9585 -765
rect 10765 -135 10785 -115
rect 10765 -185 10785 -165
rect 10765 -235 10785 -215
rect 10765 -285 10785 -265
rect 10765 -335 10785 -315
rect 10765 -385 10785 -365
rect 10765 -435 10785 -415
rect 10765 -485 10785 -465
rect 10765 -535 10785 -515
rect 10765 -585 10785 -565
rect 10765 -635 10785 -615
rect 10765 -685 10785 -665
rect 10765 -735 10785 -715
rect 10765 -785 10785 -765
rect 11965 -135 11985 -115
rect 11965 -185 11985 -165
rect 11965 -235 11985 -215
rect 11965 -285 11985 -265
rect 11965 -335 11985 -315
rect 11965 -385 11985 -365
rect 11965 -435 11985 -415
rect 11965 -485 11985 -465
rect 11965 -535 11985 -515
rect 11965 -585 11985 -565
rect 11965 -635 11985 -615
rect 11965 -685 11985 -665
rect 11965 -735 11985 -715
rect 11965 -785 11985 -765
rect 12265 -135 12285 -115
rect 12265 -185 12285 -165
rect 12265 -235 12285 -215
rect 12265 -285 12285 -265
rect 12265 -335 12285 -315
rect 12265 -385 12285 -365
rect 12265 -435 12285 -415
rect 12265 -485 12285 -465
rect 12265 -535 12285 -515
rect 12265 -585 12285 -565
rect 12265 -635 12285 -615
rect 12265 -685 12285 -665
rect 12265 -735 12285 -715
rect 12265 -785 12285 -765
rect 12565 -135 12585 -115
rect 12565 -185 12585 -165
rect 12565 -235 12585 -215
rect 12565 -285 12585 -265
rect 12565 -335 12585 -315
rect 12565 -385 12585 -365
rect 12565 -435 12585 -415
rect 12565 -485 12585 -465
rect 12565 -535 12585 -515
rect 12565 -585 12585 -565
rect 12565 -635 12585 -615
rect 12565 -685 12585 -665
rect 12565 -735 12585 -715
rect 12565 -785 12585 -765
rect 12865 -135 12885 -115
rect 12865 -185 12885 -165
rect 12865 -235 12885 -215
rect 12865 -285 12885 -265
rect 12865 -335 12885 -315
rect 12865 -385 12885 -365
rect 12865 -435 12885 -415
rect 12865 -485 12885 -465
rect 12865 -535 12885 -515
rect 12865 -585 12885 -565
rect 12865 -635 12885 -615
rect 12865 -685 12885 -665
rect 12865 -735 12885 -715
rect 12865 -785 12885 -765
rect 13165 -135 13185 -115
rect 13165 -185 13185 -165
rect 13165 -235 13185 -215
rect 13165 -285 13185 -265
rect 13165 -335 13185 -315
rect 13165 -385 13185 -365
rect 13165 -435 13185 -415
rect 13165 -485 13185 -465
rect 13165 -535 13185 -515
rect 13165 -585 13185 -565
rect 13165 -635 13185 -615
rect 13165 -685 13185 -665
rect 13165 -735 13185 -715
rect 13165 -785 13185 -765
rect 13465 -135 13485 -115
rect 13465 -185 13485 -165
rect 13465 -235 13485 -215
rect 13465 -285 13485 -265
rect 13465 -335 13485 -315
rect 13465 -385 13485 -365
rect 13465 -435 13485 -415
rect 13465 -485 13485 -465
rect 13465 -535 13485 -515
rect 13465 -585 13485 -565
rect 13465 -635 13485 -615
rect 13465 -685 13485 -665
rect 13465 -735 13485 -715
rect 13465 -785 13485 -765
rect 13765 -135 13785 -115
rect 13765 -185 13785 -165
rect 13765 -235 13785 -215
rect 13765 -285 13785 -265
rect 13765 -335 13785 -315
rect 13765 -385 13785 -365
rect 13765 -435 13785 -415
rect 13765 -485 13785 -465
rect 13765 -535 13785 -515
rect 13765 -585 13785 -565
rect 13765 -635 13785 -615
rect 13765 -685 13785 -665
rect 13765 -735 13785 -715
rect 13765 -785 13785 -765
rect 14065 -135 14085 -115
rect 14065 -185 14085 -165
rect 14065 -235 14085 -215
rect 14065 -285 14085 -265
rect 14065 -335 14085 -315
rect 14065 -385 14085 -365
rect 14065 -435 14085 -415
rect 14065 -485 14085 -465
rect 14065 -535 14085 -515
rect 14065 -585 14085 -565
rect 14065 -635 14085 -615
rect 14065 -685 14085 -665
rect 14065 -735 14085 -715
rect 14065 -785 14085 -765
rect 14365 -135 14385 -115
rect 14365 -185 14385 -165
rect 14365 -235 14385 -215
rect 14365 -285 14385 -265
rect 14365 -335 14385 -315
rect 14365 -385 14385 -365
rect 14365 -435 14385 -415
rect 14365 -485 14385 -465
rect 14365 -535 14385 -515
rect 14365 -585 14385 -565
rect 14365 -635 14385 -615
rect 14365 -685 14385 -665
rect 14365 -735 14385 -715
rect 14365 -785 14385 -765
rect 15565 -135 15585 -115
rect 15565 -185 15585 -165
rect 15565 -235 15585 -215
rect 15565 -285 15585 -265
rect 15565 -335 15585 -315
rect 15565 -385 15585 -365
rect 15565 -435 15585 -415
rect 15565 -485 15585 -465
rect 15565 -535 15585 -515
rect 15565 -585 15585 -565
rect 15565 -635 15585 -615
rect 15565 -685 15585 -665
rect 15565 -735 15585 -715
rect 15565 -785 15585 -765
rect 16765 -135 16785 -115
rect 16765 -185 16785 -165
rect 16765 -235 16785 -215
rect 16765 -285 16785 -265
rect 16765 -335 16785 -315
rect 16765 -385 16785 -365
rect 16765 -435 16785 -415
rect 16765 -485 16785 -465
rect 16765 -535 16785 -515
rect 16765 -585 16785 -565
rect 16765 -635 16785 -615
rect 16765 -685 16785 -665
rect 16765 -735 16785 -715
rect 16765 -785 16785 -765
rect 17965 -135 17985 -115
rect 17965 -185 17985 -165
rect 17965 -235 17985 -215
rect 17965 -285 17985 -265
rect 17965 -335 17985 -315
rect 17965 -385 17985 -365
rect 17965 -435 17985 -415
rect 17965 -485 17985 -465
rect 17965 -535 17985 -515
rect 17965 -585 17985 -565
rect 17965 -635 17985 -615
rect 17965 -685 17985 -665
rect 17965 -735 17985 -715
rect 17965 -785 17985 -765
rect 19165 -135 19185 -115
rect 19165 -185 19185 -165
rect 19165 -235 19185 -215
rect 19165 -285 19185 -265
rect 19165 -335 19185 -315
rect 19165 -385 19185 -365
rect 19165 -435 19185 -415
rect 19165 -485 19185 -465
rect 19165 -535 19185 -515
rect 19165 -585 19185 -565
rect 19165 -635 19185 -615
rect 19165 -685 19185 -665
rect 19165 -735 19185 -715
rect 19165 -785 19185 -765
rect 20365 -135 20385 -115
rect 20365 -185 20385 -165
rect 20365 -235 20385 -215
rect 20365 -285 20385 -265
rect 20365 -335 20385 -315
rect 20365 -385 20385 -365
rect 20365 -435 20385 -415
rect 20365 -485 20385 -465
rect 20365 -535 20385 -515
rect 20365 -585 20385 -565
rect 20365 -635 20385 -615
rect 20365 -685 20385 -665
rect 20365 -735 20385 -715
rect 20365 -785 20385 -765
rect -635 -985 -615 -965
rect -635 -1035 -615 -1015
rect -635 -1085 -615 -1065
rect -635 -1135 -615 -1115
rect -635 -1185 -615 -1165
rect -635 -1235 -615 -1215
rect -635 -1285 -615 -1265
rect -635 -1335 -615 -1315
rect -635 -1385 -615 -1365
rect -635 -1435 -615 -1415
rect -635 -1485 -615 -1465
rect -635 -1535 -615 -1515
rect -635 -1585 -615 -1565
rect -635 -1635 -615 -1615
rect -485 -985 -465 -965
rect -485 -1035 -465 -1015
rect -485 -1085 -465 -1065
rect -485 -1135 -465 -1115
rect -485 -1185 -465 -1165
rect -485 -1235 -465 -1215
rect -485 -1285 -465 -1265
rect -485 -1335 -465 -1315
rect -485 -1385 -465 -1365
rect -485 -1435 -465 -1415
rect -485 -1485 -465 -1465
rect -485 -1535 -465 -1515
rect -485 -1585 -465 -1565
rect -485 -1635 -465 -1615
rect -335 -985 -315 -965
rect -335 -1035 -315 -1015
rect -335 -1085 -315 -1065
rect -335 -1135 -315 -1115
rect -335 -1185 -315 -1165
rect -335 -1235 -315 -1215
rect -335 -1285 -315 -1265
rect -335 -1335 -315 -1315
rect -335 -1385 -315 -1365
rect -335 -1435 -315 -1415
rect -335 -1485 -315 -1465
rect -335 -1535 -315 -1515
rect -335 -1585 -315 -1565
rect -335 -1635 -315 -1615
rect -185 -985 -165 -965
rect -185 -1035 -165 -1015
rect -185 -1085 -165 -1065
rect -185 -1135 -165 -1115
rect -185 -1185 -165 -1165
rect -185 -1235 -165 -1215
rect -185 -1285 -165 -1265
rect -185 -1335 -165 -1315
rect -185 -1385 -165 -1365
rect -185 -1435 -165 -1415
rect -185 -1485 -165 -1465
rect -185 -1535 -165 -1515
rect -185 -1585 -165 -1565
rect -185 -1635 -165 -1615
rect -35 -985 -15 -965
rect -35 -1035 -15 -1015
rect -35 -1085 -15 -1065
rect -35 -1135 -15 -1115
rect -35 -1185 -15 -1165
rect -35 -1235 -15 -1215
rect -35 -1285 -15 -1265
rect -35 -1335 -15 -1315
rect -35 -1385 -15 -1365
rect -35 -1435 -15 -1415
rect -35 -1485 -15 -1465
rect -35 -1535 -15 -1515
rect -35 -1585 -15 -1565
rect -35 -1635 -15 -1615
rect 1165 -985 1185 -965
rect 1165 -1035 1185 -1015
rect 1165 -1085 1185 -1065
rect 1165 -1135 1185 -1115
rect 1165 -1185 1185 -1165
rect 1165 -1235 1185 -1215
rect 1165 -1285 1185 -1265
rect 1165 -1335 1185 -1315
rect 1165 -1385 1185 -1365
rect 1165 -1435 1185 -1415
rect 1165 -1485 1185 -1465
rect 1165 -1535 1185 -1515
rect 1165 -1585 1185 -1565
rect 1165 -1635 1185 -1615
rect 1465 -985 1485 -965
rect 1465 -1035 1485 -1015
rect 1465 -1085 1485 -1065
rect 1465 -1135 1485 -1115
rect 1465 -1185 1485 -1165
rect 1465 -1235 1485 -1215
rect 1465 -1285 1485 -1265
rect 1465 -1335 1485 -1315
rect 1465 -1385 1485 -1365
rect 1465 -1435 1485 -1415
rect 1465 -1485 1485 -1465
rect 1465 -1535 1485 -1515
rect 1465 -1585 1485 -1565
rect 1465 -1635 1485 -1615
rect 1765 -985 1785 -965
rect 1765 -1035 1785 -1015
rect 1765 -1085 1785 -1065
rect 1765 -1135 1785 -1115
rect 1765 -1185 1785 -1165
rect 1765 -1235 1785 -1215
rect 1765 -1285 1785 -1265
rect 1765 -1335 1785 -1315
rect 1765 -1385 1785 -1365
rect 1765 -1435 1785 -1415
rect 1765 -1485 1785 -1465
rect 1765 -1535 1785 -1515
rect 1765 -1585 1785 -1565
rect 1765 -1635 1785 -1615
rect 2065 -985 2085 -965
rect 2065 -1035 2085 -1015
rect 2065 -1085 2085 -1065
rect 2065 -1135 2085 -1115
rect 2065 -1185 2085 -1165
rect 2065 -1235 2085 -1215
rect 2065 -1285 2085 -1265
rect 2065 -1335 2085 -1315
rect 2065 -1385 2085 -1365
rect 2065 -1435 2085 -1415
rect 2065 -1485 2085 -1465
rect 2065 -1535 2085 -1515
rect 2065 -1585 2085 -1565
rect 2065 -1635 2085 -1615
rect 2365 -985 2385 -965
rect 2365 -1035 2385 -1015
rect 2365 -1085 2385 -1065
rect 2365 -1135 2385 -1115
rect 2365 -1185 2385 -1165
rect 2365 -1235 2385 -1215
rect 2365 -1285 2385 -1265
rect 2365 -1335 2385 -1315
rect 2365 -1385 2385 -1365
rect 2365 -1435 2385 -1415
rect 2365 -1485 2385 -1465
rect 2365 -1535 2385 -1515
rect 2365 -1585 2385 -1565
rect 2365 -1635 2385 -1615
rect 2665 -985 2685 -965
rect 2665 -1035 2685 -1015
rect 2665 -1085 2685 -1065
rect 2665 -1135 2685 -1115
rect 2665 -1185 2685 -1165
rect 2665 -1235 2685 -1215
rect 2665 -1285 2685 -1265
rect 2665 -1335 2685 -1315
rect 2665 -1385 2685 -1365
rect 2665 -1435 2685 -1415
rect 2665 -1485 2685 -1465
rect 2665 -1535 2685 -1515
rect 2665 -1585 2685 -1565
rect 2665 -1635 2685 -1615
rect 2965 -985 2985 -965
rect 2965 -1035 2985 -1015
rect 2965 -1085 2985 -1065
rect 2965 -1135 2985 -1115
rect 2965 -1185 2985 -1165
rect 2965 -1235 2985 -1215
rect 2965 -1285 2985 -1265
rect 2965 -1335 2985 -1315
rect 2965 -1385 2985 -1365
rect 2965 -1435 2985 -1415
rect 2965 -1485 2985 -1465
rect 2965 -1535 2985 -1515
rect 2965 -1585 2985 -1565
rect 2965 -1635 2985 -1615
rect 3265 -985 3285 -965
rect 3265 -1035 3285 -1015
rect 3265 -1085 3285 -1065
rect 3265 -1135 3285 -1115
rect 3265 -1185 3285 -1165
rect 3265 -1235 3285 -1215
rect 3265 -1285 3285 -1265
rect 3265 -1335 3285 -1315
rect 3265 -1385 3285 -1365
rect 3265 -1435 3285 -1415
rect 3265 -1485 3285 -1465
rect 3265 -1535 3285 -1515
rect 3265 -1585 3285 -1565
rect 3265 -1635 3285 -1615
rect 3565 -985 3585 -965
rect 3565 -1035 3585 -1015
rect 3565 -1085 3585 -1065
rect 3565 -1135 3585 -1115
rect 3565 -1185 3585 -1165
rect 3565 -1235 3585 -1215
rect 3565 -1285 3585 -1265
rect 3565 -1335 3585 -1315
rect 3565 -1385 3585 -1365
rect 3565 -1435 3585 -1415
rect 3565 -1485 3585 -1465
rect 3565 -1535 3585 -1515
rect 3565 -1585 3585 -1565
rect 3565 -1635 3585 -1615
rect 3715 -985 3735 -965
rect 3715 -1035 3735 -1015
rect 3715 -1085 3735 -1065
rect 3715 -1135 3735 -1115
rect 3715 -1185 3735 -1165
rect 3715 -1235 3735 -1215
rect 3715 -1285 3735 -1265
rect 3715 -1335 3735 -1315
rect 3715 -1385 3735 -1365
rect 3715 -1435 3735 -1415
rect 3715 -1485 3735 -1465
rect 3715 -1535 3735 -1515
rect 3715 -1585 3735 -1565
rect 3715 -1635 3735 -1615
rect 3865 -985 3885 -965
rect 3865 -1035 3885 -1015
rect 3865 -1085 3885 -1065
rect 3865 -1135 3885 -1115
rect 3865 -1185 3885 -1165
rect 3865 -1235 3885 -1215
rect 3865 -1285 3885 -1265
rect 3865 -1335 3885 -1315
rect 3865 -1385 3885 -1365
rect 3865 -1435 3885 -1415
rect 3865 -1485 3885 -1465
rect 3865 -1535 3885 -1515
rect 3865 -1585 3885 -1565
rect 3865 -1635 3885 -1615
rect 4015 -985 4035 -965
rect 4015 -1035 4035 -1015
rect 4015 -1085 4035 -1065
rect 4015 -1135 4035 -1115
rect 4015 -1185 4035 -1165
rect 4015 -1235 4035 -1215
rect 4015 -1285 4035 -1265
rect 4015 -1335 4035 -1315
rect 4015 -1385 4035 -1365
rect 4015 -1435 4035 -1415
rect 4015 -1485 4035 -1465
rect 4015 -1535 4035 -1515
rect 4015 -1585 4035 -1565
rect 4015 -1635 4035 -1615
rect 4165 -985 4185 -965
rect 4165 -1035 4185 -1015
rect 4165 -1085 4185 -1065
rect 4165 -1135 4185 -1115
rect 4165 -1185 4185 -1165
rect 4165 -1235 4185 -1215
rect 4165 -1285 4185 -1265
rect 4165 -1335 4185 -1315
rect 4165 -1385 4185 -1365
rect 4165 -1435 4185 -1415
rect 4165 -1485 4185 -1465
rect 4165 -1535 4185 -1515
rect 4165 -1585 4185 -1565
rect 4165 -1635 4185 -1615
rect 4315 -985 4335 -965
rect 4315 -1035 4335 -1015
rect 4315 -1085 4335 -1065
rect 4315 -1135 4335 -1115
rect 4315 -1185 4335 -1165
rect 4315 -1235 4335 -1215
rect 4315 -1285 4335 -1265
rect 4315 -1335 4335 -1315
rect 4315 -1385 4335 -1365
rect 4315 -1435 4335 -1415
rect 4315 -1485 4335 -1465
rect 4315 -1535 4335 -1515
rect 4315 -1585 4335 -1565
rect 4315 -1635 4335 -1615
rect 4465 -985 4485 -965
rect 4465 -1035 4485 -1015
rect 4465 -1085 4485 -1065
rect 4465 -1135 4485 -1115
rect 4465 -1185 4485 -1165
rect 4465 -1235 4485 -1215
rect 4465 -1285 4485 -1265
rect 4465 -1335 4485 -1315
rect 4465 -1385 4485 -1365
rect 4465 -1435 4485 -1415
rect 4465 -1485 4485 -1465
rect 4465 -1535 4485 -1515
rect 4465 -1585 4485 -1565
rect 4465 -1635 4485 -1615
rect 4615 -985 4635 -965
rect 4615 -1035 4635 -1015
rect 4615 -1085 4635 -1065
rect 4615 -1135 4635 -1115
rect 4615 -1185 4635 -1165
rect 4615 -1235 4635 -1215
rect 4615 -1285 4635 -1265
rect 4615 -1335 4635 -1315
rect 4615 -1385 4635 -1365
rect 4615 -1435 4635 -1415
rect 4615 -1485 4635 -1465
rect 4615 -1535 4635 -1515
rect 4615 -1585 4635 -1565
rect 4615 -1635 4635 -1615
rect 4765 -985 4785 -965
rect 4765 -1035 4785 -1015
rect 4765 -1085 4785 -1065
rect 4765 -1135 4785 -1115
rect 4765 -1185 4785 -1165
rect 4765 -1235 4785 -1215
rect 4765 -1285 4785 -1265
rect 4765 -1335 4785 -1315
rect 4765 -1385 4785 -1365
rect 4765 -1435 4785 -1415
rect 4765 -1485 4785 -1465
rect 4765 -1535 4785 -1515
rect 4765 -1585 4785 -1565
rect 4765 -1635 4785 -1615
rect 5065 -985 5085 -965
rect 5065 -1035 5085 -1015
rect 5065 -1085 5085 -1065
rect 5065 -1135 5085 -1115
rect 5065 -1185 5085 -1165
rect 5065 -1235 5085 -1215
rect 5065 -1285 5085 -1265
rect 5065 -1335 5085 -1315
rect 5065 -1385 5085 -1365
rect 5065 -1435 5085 -1415
rect 5065 -1485 5085 -1465
rect 5065 -1535 5085 -1515
rect 5065 -1585 5085 -1565
rect 5065 -1635 5085 -1615
rect 5365 -985 5385 -965
rect 5365 -1035 5385 -1015
rect 5365 -1085 5385 -1065
rect 5365 -1135 5385 -1115
rect 5365 -1185 5385 -1165
rect 5365 -1235 5385 -1215
rect 5365 -1285 5385 -1265
rect 5365 -1335 5385 -1315
rect 5365 -1385 5385 -1365
rect 5365 -1435 5385 -1415
rect 5365 -1485 5385 -1465
rect 5365 -1535 5385 -1515
rect 5365 -1585 5385 -1565
rect 5365 -1635 5385 -1615
rect 5665 -985 5685 -965
rect 5665 -1035 5685 -1015
rect 5665 -1085 5685 -1065
rect 5665 -1135 5685 -1115
rect 5665 -1185 5685 -1165
rect 5665 -1235 5685 -1215
rect 5665 -1285 5685 -1265
rect 5665 -1335 5685 -1315
rect 5665 -1385 5685 -1365
rect 5665 -1435 5685 -1415
rect 5665 -1485 5685 -1465
rect 5665 -1535 5685 -1515
rect 5665 -1585 5685 -1565
rect 5665 -1635 5685 -1615
rect 5965 -985 5985 -965
rect 5965 -1035 5985 -1015
rect 5965 -1085 5985 -1065
rect 5965 -1135 5985 -1115
rect 5965 -1185 5985 -1165
rect 5965 -1235 5985 -1215
rect 5965 -1285 5985 -1265
rect 5965 -1335 5985 -1315
rect 5965 -1385 5985 -1365
rect 5965 -1435 5985 -1415
rect 5965 -1485 5985 -1465
rect 5965 -1535 5985 -1515
rect 5965 -1585 5985 -1565
rect 5965 -1635 5985 -1615
rect 6265 -985 6285 -965
rect 6265 -1035 6285 -1015
rect 6265 -1085 6285 -1065
rect 6265 -1135 6285 -1115
rect 6265 -1185 6285 -1165
rect 6265 -1235 6285 -1215
rect 6265 -1285 6285 -1265
rect 6265 -1335 6285 -1315
rect 6265 -1385 6285 -1365
rect 6265 -1435 6285 -1415
rect 6265 -1485 6285 -1465
rect 6265 -1535 6285 -1515
rect 6265 -1585 6285 -1565
rect 6265 -1635 6285 -1615
rect 6565 -985 6585 -965
rect 6565 -1035 6585 -1015
rect 6565 -1085 6585 -1065
rect 6565 -1135 6585 -1115
rect 6565 -1185 6585 -1165
rect 6565 -1235 6585 -1215
rect 6565 -1285 6585 -1265
rect 6565 -1335 6585 -1315
rect 6565 -1385 6585 -1365
rect 6565 -1435 6585 -1415
rect 6565 -1485 6585 -1465
rect 6565 -1535 6585 -1515
rect 6565 -1585 6585 -1565
rect 6565 -1635 6585 -1615
rect 6865 -985 6885 -965
rect 6865 -1035 6885 -1015
rect 6865 -1085 6885 -1065
rect 6865 -1135 6885 -1115
rect 6865 -1185 6885 -1165
rect 6865 -1235 6885 -1215
rect 6865 -1285 6885 -1265
rect 6865 -1335 6885 -1315
rect 6865 -1385 6885 -1365
rect 6865 -1435 6885 -1415
rect 6865 -1485 6885 -1465
rect 6865 -1535 6885 -1515
rect 6865 -1585 6885 -1565
rect 6865 -1635 6885 -1615
rect 7165 -985 7185 -965
rect 7165 -1035 7185 -1015
rect 7165 -1085 7185 -1065
rect 7165 -1135 7185 -1115
rect 7165 -1185 7185 -1165
rect 7165 -1235 7185 -1215
rect 7165 -1285 7185 -1265
rect 7165 -1335 7185 -1315
rect 7165 -1385 7185 -1365
rect 7165 -1435 7185 -1415
rect 7165 -1485 7185 -1465
rect 7165 -1535 7185 -1515
rect 7165 -1585 7185 -1565
rect 7165 -1635 7185 -1615
rect 8365 -985 8385 -965
rect 8365 -1035 8385 -1015
rect 8365 -1085 8385 -1065
rect 8365 -1135 8385 -1115
rect 8365 -1185 8385 -1165
rect 8365 -1235 8385 -1215
rect 8365 -1285 8385 -1265
rect 8365 -1335 8385 -1315
rect 8365 -1385 8385 -1365
rect 8365 -1435 8385 -1415
rect 8365 -1485 8385 -1465
rect 8365 -1535 8385 -1515
rect 8365 -1585 8385 -1565
rect 8365 -1635 8385 -1615
rect 9565 -985 9585 -965
rect 9565 -1035 9585 -1015
rect 9565 -1085 9585 -1065
rect 9565 -1135 9585 -1115
rect 9565 -1185 9585 -1165
rect 9565 -1235 9585 -1215
rect 9565 -1285 9585 -1265
rect 9565 -1335 9585 -1315
rect 9565 -1385 9585 -1365
rect 9565 -1435 9585 -1415
rect 9565 -1485 9585 -1465
rect 9565 -1535 9585 -1515
rect 9565 -1585 9585 -1565
rect 9565 -1635 9585 -1615
rect 10765 -985 10785 -965
rect 10765 -1035 10785 -1015
rect 10765 -1085 10785 -1065
rect 10765 -1135 10785 -1115
rect 10765 -1185 10785 -1165
rect 10765 -1235 10785 -1215
rect 10765 -1285 10785 -1265
rect 10765 -1335 10785 -1315
rect 10765 -1385 10785 -1365
rect 10765 -1435 10785 -1415
rect 10765 -1485 10785 -1465
rect 10765 -1535 10785 -1515
rect 10765 -1585 10785 -1565
rect 10765 -1635 10785 -1615
rect 11965 -985 11985 -965
rect 11965 -1035 11985 -1015
rect 11965 -1085 11985 -1065
rect 11965 -1135 11985 -1115
rect 11965 -1185 11985 -1165
rect 11965 -1235 11985 -1215
rect 11965 -1285 11985 -1265
rect 11965 -1335 11985 -1315
rect 11965 -1385 11985 -1365
rect 11965 -1435 11985 -1415
rect 11965 -1485 11985 -1465
rect 11965 -1535 11985 -1515
rect 11965 -1585 11985 -1565
rect 11965 -1635 11985 -1615
rect 12265 -985 12285 -965
rect 12265 -1035 12285 -1015
rect 12265 -1085 12285 -1065
rect 12265 -1135 12285 -1115
rect 12265 -1185 12285 -1165
rect 12265 -1235 12285 -1215
rect 12265 -1285 12285 -1265
rect 12265 -1335 12285 -1315
rect 12265 -1385 12285 -1365
rect 12265 -1435 12285 -1415
rect 12265 -1485 12285 -1465
rect 12265 -1535 12285 -1515
rect 12265 -1585 12285 -1565
rect 12265 -1635 12285 -1615
rect 12565 -985 12585 -965
rect 12565 -1035 12585 -1015
rect 12565 -1085 12585 -1065
rect 12565 -1135 12585 -1115
rect 12565 -1185 12585 -1165
rect 12565 -1235 12585 -1215
rect 12565 -1285 12585 -1265
rect 12565 -1335 12585 -1315
rect 12565 -1385 12585 -1365
rect 12565 -1435 12585 -1415
rect 12565 -1485 12585 -1465
rect 12565 -1535 12585 -1515
rect 12565 -1585 12585 -1565
rect 12565 -1635 12585 -1615
rect 12865 -985 12885 -965
rect 12865 -1035 12885 -1015
rect 12865 -1085 12885 -1065
rect 12865 -1135 12885 -1115
rect 12865 -1185 12885 -1165
rect 12865 -1235 12885 -1215
rect 12865 -1285 12885 -1265
rect 12865 -1335 12885 -1315
rect 12865 -1385 12885 -1365
rect 12865 -1435 12885 -1415
rect 12865 -1485 12885 -1465
rect 12865 -1535 12885 -1515
rect 12865 -1585 12885 -1565
rect 12865 -1635 12885 -1615
rect 13165 -985 13185 -965
rect 13165 -1035 13185 -1015
rect 13165 -1085 13185 -1065
rect 13165 -1135 13185 -1115
rect 13165 -1185 13185 -1165
rect 13165 -1235 13185 -1215
rect 13165 -1285 13185 -1265
rect 13165 -1335 13185 -1315
rect 13165 -1385 13185 -1365
rect 13165 -1435 13185 -1415
rect 13165 -1485 13185 -1465
rect 13165 -1535 13185 -1515
rect 13165 -1585 13185 -1565
rect 13165 -1635 13185 -1615
rect 13465 -985 13485 -965
rect 13465 -1035 13485 -1015
rect 13465 -1085 13485 -1065
rect 13465 -1135 13485 -1115
rect 13465 -1185 13485 -1165
rect 13465 -1235 13485 -1215
rect 13465 -1285 13485 -1265
rect 13465 -1335 13485 -1315
rect 13465 -1385 13485 -1365
rect 13465 -1435 13485 -1415
rect 13465 -1485 13485 -1465
rect 13465 -1535 13485 -1515
rect 13465 -1585 13485 -1565
rect 13465 -1635 13485 -1615
rect 13765 -985 13785 -965
rect 13765 -1035 13785 -1015
rect 13765 -1085 13785 -1065
rect 13765 -1135 13785 -1115
rect 13765 -1185 13785 -1165
rect 13765 -1235 13785 -1215
rect 13765 -1285 13785 -1265
rect 13765 -1335 13785 -1315
rect 13765 -1385 13785 -1365
rect 13765 -1435 13785 -1415
rect 13765 -1485 13785 -1465
rect 13765 -1535 13785 -1515
rect 13765 -1585 13785 -1565
rect 13765 -1635 13785 -1615
rect 14065 -985 14085 -965
rect 14065 -1035 14085 -1015
rect 14065 -1085 14085 -1065
rect 14065 -1135 14085 -1115
rect 14065 -1185 14085 -1165
rect 14065 -1235 14085 -1215
rect 14065 -1285 14085 -1265
rect 14065 -1335 14085 -1315
rect 14065 -1385 14085 -1365
rect 14065 -1435 14085 -1415
rect 14065 -1485 14085 -1465
rect 14065 -1535 14085 -1515
rect 14065 -1585 14085 -1565
rect 14065 -1635 14085 -1615
rect 14365 -985 14385 -965
rect 14365 -1035 14385 -1015
rect 14365 -1085 14385 -1065
rect 14365 -1135 14385 -1115
rect 14365 -1185 14385 -1165
rect 14365 -1235 14385 -1215
rect 14365 -1285 14385 -1265
rect 14365 -1335 14385 -1315
rect 14365 -1385 14385 -1365
rect 14365 -1435 14385 -1415
rect 14365 -1485 14385 -1465
rect 14365 -1535 14385 -1515
rect 14365 -1585 14385 -1565
rect 14365 -1635 14385 -1615
rect 15565 -985 15585 -965
rect 15565 -1035 15585 -1015
rect 15565 -1085 15585 -1065
rect 15565 -1135 15585 -1115
rect 15565 -1185 15585 -1165
rect 15565 -1235 15585 -1215
rect 15565 -1285 15585 -1265
rect 15565 -1335 15585 -1315
rect 15565 -1385 15585 -1365
rect 15565 -1435 15585 -1415
rect 15565 -1485 15585 -1465
rect 15565 -1535 15585 -1515
rect 15565 -1585 15585 -1565
rect 15565 -1635 15585 -1615
rect 16765 -985 16785 -965
rect 16765 -1035 16785 -1015
rect 16765 -1085 16785 -1065
rect 16765 -1135 16785 -1115
rect 16765 -1185 16785 -1165
rect 16765 -1235 16785 -1215
rect 16765 -1285 16785 -1265
rect 16765 -1335 16785 -1315
rect 16765 -1385 16785 -1365
rect 16765 -1435 16785 -1415
rect 16765 -1485 16785 -1465
rect 16765 -1535 16785 -1515
rect 16765 -1585 16785 -1565
rect 16765 -1635 16785 -1615
rect 17965 -985 17985 -965
rect 17965 -1035 17985 -1015
rect 17965 -1085 17985 -1065
rect 17965 -1135 17985 -1115
rect 17965 -1185 17985 -1165
rect 17965 -1235 17985 -1215
rect 17965 -1285 17985 -1265
rect 17965 -1335 17985 -1315
rect 17965 -1385 17985 -1365
rect 17965 -1435 17985 -1415
rect 17965 -1485 17985 -1465
rect 17965 -1535 17985 -1515
rect 17965 -1585 17985 -1565
rect 17965 -1635 17985 -1615
rect 19165 -985 19185 -965
rect 19165 -1035 19185 -1015
rect 19165 -1085 19185 -1065
rect 19165 -1135 19185 -1115
rect 19165 -1185 19185 -1165
rect 19165 -1235 19185 -1215
rect 19165 -1285 19185 -1265
rect 19165 -1335 19185 -1315
rect 19165 -1385 19185 -1365
rect 19165 -1435 19185 -1415
rect 19165 -1485 19185 -1465
rect 19165 -1535 19185 -1515
rect 19165 -1585 19185 -1565
rect 19165 -1635 19185 -1615
rect 20365 -985 20385 -965
rect 20365 -1035 20385 -1015
rect 20365 -1085 20385 -1065
rect 20365 -1135 20385 -1115
rect 20365 -1185 20385 -1165
rect 20365 -1235 20385 -1215
rect 20365 -1285 20385 -1265
rect 20365 -1335 20385 -1315
rect 20365 -1385 20385 -1365
rect 20365 -1435 20385 -1415
rect 20365 -1485 20385 -1465
rect 20365 -1535 20385 -1515
rect 20365 -1585 20385 -1565
rect 20365 -1635 20385 -1615
<< mvpdiffc >>
rect -635 5065 -615 5085
rect -635 5015 -615 5035
rect -635 4965 -615 4985
rect -635 4915 -615 4935
rect -635 4865 -615 4885
rect -635 4815 -615 4835
rect -635 4765 -615 4785
rect -635 4715 -615 4735
rect -635 4665 -615 4685
rect -635 4615 -615 4635
rect -485 5065 -465 5085
rect -485 5015 -465 5035
rect -485 4965 -465 4985
rect -485 4915 -465 4935
rect -485 4865 -465 4885
rect -485 4815 -465 4835
rect -485 4765 -465 4785
rect -485 4715 -465 4735
rect -485 4665 -465 4685
rect -485 4615 -465 4635
rect -335 5065 -315 5085
rect -335 5015 -315 5035
rect -335 4965 -315 4985
rect -335 4915 -315 4935
rect -335 4865 -315 4885
rect -335 4815 -315 4835
rect -335 4765 -315 4785
rect -335 4715 -315 4735
rect -335 4665 -315 4685
rect -335 4615 -315 4635
rect -185 5065 -165 5085
rect -185 5015 -165 5035
rect -185 4965 -165 4985
rect -185 4915 -165 4935
rect -185 4865 -165 4885
rect -185 4815 -165 4835
rect -185 4765 -165 4785
rect -185 4715 -165 4735
rect -185 4665 -165 4685
rect -185 4615 -165 4635
rect -35 5065 -15 5085
rect -35 5015 -15 5035
rect -35 4965 -15 4985
rect -35 4915 -15 4935
rect -35 4865 -15 4885
rect -35 4815 -15 4835
rect -35 4765 -15 4785
rect -35 4715 -15 4735
rect -35 4665 -15 4685
rect -35 4615 -15 4635
rect 565 5065 585 5085
rect 565 5015 585 5035
rect 565 4965 585 4985
rect 565 4915 585 4935
rect 565 4865 585 4885
rect 565 4815 585 4835
rect 565 4765 585 4785
rect 565 4715 585 4735
rect 565 4665 585 4685
rect 565 4615 585 4635
rect 715 5065 735 5085
rect 715 5015 735 5035
rect 715 4965 735 4985
rect 715 4915 735 4935
rect 715 4865 735 4885
rect 715 4815 735 4835
rect 715 4765 735 4785
rect 715 4715 735 4735
rect 715 4665 735 4685
rect 715 4615 735 4635
rect 865 5065 885 5085
rect 865 5015 885 5035
rect 865 4965 885 4985
rect 865 4915 885 4935
rect 865 4865 885 4885
rect 865 4815 885 4835
rect 865 4765 885 4785
rect 865 4715 885 4735
rect 865 4665 885 4685
rect 865 4615 885 4635
rect 1015 5065 1035 5085
rect 1015 5015 1035 5035
rect 1015 4965 1035 4985
rect 1015 4915 1035 4935
rect 1015 4865 1035 4885
rect 1015 4815 1035 4835
rect 1015 4765 1035 4785
rect 1015 4715 1035 4735
rect 1015 4665 1035 4685
rect 1015 4615 1035 4635
rect 1165 5065 1185 5085
rect 1165 5015 1185 5035
rect 1165 4965 1185 4985
rect 1165 4915 1185 4935
rect 1165 4865 1185 4885
rect 1165 4815 1185 4835
rect 1165 4765 1185 4785
rect 1165 4715 1185 4735
rect 1165 4665 1185 4685
rect 1165 4615 1185 4635
rect 1315 5065 1335 5085
rect 1315 5015 1335 5035
rect 1315 4965 1335 4985
rect 1315 4915 1335 4935
rect 1315 4865 1335 4885
rect 1315 4815 1335 4835
rect 1315 4765 1335 4785
rect 1315 4715 1335 4735
rect 1315 4665 1335 4685
rect 1315 4615 1335 4635
rect 1465 5065 1485 5085
rect 1465 5015 1485 5035
rect 1465 4965 1485 4985
rect 1465 4915 1485 4935
rect 1465 4865 1485 4885
rect 1465 4815 1485 4835
rect 1465 4765 1485 4785
rect 1465 4715 1485 4735
rect 1465 4665 1485 4685
rect 1465 4615 1485 4635
rect 1615 5065 1635 5085
rect 1615 5015 1635 5035
rect 1615 4965 1635 4985
rect 1615 4915 1635 4935
rect 1615 4865 1635 4885
rect 1615 4815 1635 4835
rect 1615 4765 1635 4785
rect 1615 4715 1635 4735
rect 1615 4665 1635 4685
rect 1615 4615 1635 4635
rect 1765 5065 1785 5085
rect 1765 5015 1785 5035
rect 1765 4965 1785 4985
rect 1765 4915 1785 4935
rect 1765 4865 1785 4885
rect 1765 4815 1785 4835
rect 1765 4765 1785 4785
rect 1765 4715 1785 4735
rect 1765 4665 1785 4685
rect 1765 4615 1785 4635
rect 1915 5065 1935 5085
rect 1915 5015 1935 5035
rect 1915 4965 1935 4985
rect 1915 4915 1935 4935
rect 1915 4865 1935 4885
rect 1915 4815 1935 4835
rect 1915 4765 1935 4785
rect 1915 4715 1935 4735
rect 1915 4665 1935 4685
rect 1915 4615 1935 4635
rect 2065 5065 2085 5085
rect 2065 5015 2085 5035
rect 2065 4965 2085 4985
rect 2065 4915 2085 4935
rect 2065 4865 2085 4885
rect 2065 4815 2085 4835
rect 2065 4765 2085 4785
rect 2065 4715 2085 4735
rect 2065 4665 2085 4685
rect 2065 4615 2085 4635
rect 2215 5065 2235 5085
rect 2215 5015 2235 5035
rect 2215 4965 2235 4985
rect 2215 4915 2235 4935
rect 2215 4865 2235 4885
rect 2215 4815 2235 4835
rect 2215 4765 2235 4785
rect 2215 4715 2235 4735
rect 2215 4665 2235 4685
rect 2215 4615 2235 4635
rect 2365 5065 2385 5085
rect 2365 5015 2385 5035
rect 2365 4965 2385 4985
rect 2365 4915 2385 4935
rect 2365 4865 2385 4885
rect 2365 4815 2385 4835
rect 2365 4765 2385 4785
rect 2365 4715 2385 4735
rect 2365 4665 2385 4685
rect 2365 4615 2385 4635
rect 2515 5065 2535 5085
rect 2515 5015 2535 5035
rect 2515 4965 2535 4985
rect 2515 4915 2535 4935
rect 2515 4865 2535 4885
rect 2515 4815 2535 4835
rect 2515 4765 2535 4785
rect 2515 4715 2535 4735
rect 2515 4665 2535 4685
rect 2515 4615 2535 4635
rect 2665 5065 2685 5085
rect 2665 5015 2685 5035
rect 2665 4965 2685 4985
rect 2665 4915 2685 4935
rect 2665 4865 2685 4885
rect 2665 4815 2685 4835
rect 2665 4765 2685 4785
rect 2665 4715 2685 4735
rect 2665 4665 2685 4685
rect 2665 4615 2685 4635
rect 2815 5065 2835 5085
rect 2815 5015 2835 5035
rect 2815 4965 2835 4985
rect 2815 4915 2835 4935
rect 2815 4865 2835 4885
rect 2815 4815 2835 4835
rect 2815 4765 2835 4785
rect 2815 4715 2835 4735
rect 2815 4665 2835 4685
rect 2815 4615 2835 4635
rect 2965 5065 2985 5085
rect 2965 5015 2985 5035
rect 2965 4965 2985 4985
rect 2965 4915 2985 4935
rect 2965 4865 2985 4885
rect 2965 4815 2985 4835
rect 2965 4765 2985 4785
rect 2965 4715 2985 4735
rect 2965 4665 2985 4685
rect 2965 4615 2985 4635
rect 3115 5065 3135 5085
rect 3115 5015 3135 5035
rect 3115 4965 3135 4985
rect 3115 4915 3135 4935
rect 3115 4865 3135 4885
rect 3115 4815 3135 4835
rect 3115 4765 3135 4785
rect 3115 4715 3135 4735
rect 3115 4665 3135 4685
rect 3115 4615 3135 4635
rect 3265 5065 3285 5085
rect 3265 5015 3285 5035
rect 3265 4965 3285 4985
rect 3265 4915 3285 4935
rect 3265 4865 3285 4885
rect 3265 4815 3285 4835
rect 3265 4765 3285 4785
rect 3265 4715 3285 4735
rect 3265 4665 3285 4685
rect 3265 4615 3285 4635
rect 3415 5065 3435 5085
rect 3415 5015 3435 5035
rect 3415 4965 3435 4985
rect 3415 4915 3435 4935
rect 3415 4865 3435 4885
rect 3415 4815 3435 4835
rect 3415 4765 3435 4785
rect 3415 4715 3435 4735
rect 3415 4665 3435 4685
rect 3415 4615 3435 4635
rect 3565 5065 3585 5085
rect 3565 5015 3585 5035
rect 3565 4965 3585 4985
rect 3565 4915 3585 4935
rect 3565 4865 3585 4885
rect 3565 4815 3585 4835
rect 3565 4765 3585 4785
rect 3565 4715 3585 4735
rect 3565 4665 3585 4685
rect 3565 4615 3585 4635
rect 4165 5065 4185 5085
rect 4165 5015 4185 5035
rect 4165 4965 4185 4985
rect 4165 4915 4185 4935
rect 4165 4865 4185 4885
rect 4165 4815 4185 4835
rect 4165 4765 4185 4785
rect 4165 4715 4185 4735
rect 4165 4665 4185 4685
rect 4165 4615 4185 4635
rect 4765 5065 4785 5085
rect 4765 5015 4785 5035
rect 4765 4965 4785 4985
rect 4765 4915 4785 4935
rect 4765 4865 4785 4885
rect 4765 4815 4785 4835
rect 4765 4765 4785 4785
rect 4765 4715 4785 4735
rect 4765 4665 4785 4685
rect 4765 4615 4785 4635
rect 4915 5065 4935 5085
rect 4915 5015 4935 5035
rect 4915 4965 4935 4985
rect 4915 4915 4935 4935
rect 4915 4865 4935 4885
rect 4915 4815 4935 4835
rect 4915 4765 4935 4785
rect 4915 4715 4935 4735
rect 4915 4665 4935 4685
rect 4915 4615 4935 4635
rect 5065 5065 5085 5085
rect 5065 5015 5085 5035
rect 5065 4965 5085 4985
rect 5065 4915 5085 4935
rect 5065 4865 5085 4885
rect 5065 4815 5085 4835
rect 5065 4765 5085 4785
rect 5065 4715 5085 4735
rect 5065 4665 5085 4685
rect 5065 4615 5085 4635
rect 5215 5065 5235 5085
rect 5215 5015 5235 5035
rect 5215 4965 5235 4985
rect 5215 4915 5235 4935
rect 5215 4865 5235 4885
rect 5215 4815 5235 4835
rect 5215 4765 5235 4785
rect 5215 4715 5235 4735
rect 5215 4665 5235 4685
rect 5215 4615 5235 4635
rect 5365 5065 5385 5085
rect 5365 5015 5385 5035
rect 5365 4965 5385 4985
rect 5365 4915 5385 4935
rect 5365 4865 5385 4885
rect 5365 4815 5385 4835
rect 5365 4765 5385 4785
rect 5365 4715 5385 4735
rect 5365 4665 5385 4685
rect 5365 4615 5385 4635
rect 5515 5065 5535 5085
rect 5515 5015 5535 5035
rect 5515 4965 5535 4985
rect 5515 4915 5535 4935
rect 5515 4865 5535 4885
rect 5515 4815 5535 4835
rect 5515 4765 5535 4785
rect 5515 4715 5535 4735
rect 5515 4665 5535 4685
rect 5515 4615 5535 4635
rect 5665 5065 5685 5085
rect 5665 5015 5685 5035
rect 5665 4965 5685 4985
rect 5665 4915 5685 4935
rect 5665 4865 5685 4885
rect 5665 4815 5685 4835
rect 5665 4765 5685 4785
rect 5665 4715 5685 4735
rect 5665 4665 5685 4685
rect 5665 4615 5685 4635
rect 5815 5065 5835 5085
rect 5815 5015 5835 5035
rect 5815 4965 5835 4985
rect 5815 4915 5835 4935
rect 5815 4865 5835 4885
rect 5815 4815 5835 4835
rect 5815 4765 5835 4785
rect 5815 4715 5835 4735
rect 5815 4665 5835 4685
rect 5815 4615 5835 4635
rect 5965 5065 5985 5085
rect 5965 5015 5985 5035
rect 5965 4965 5985 4985
rect 5965 4915 5985 4935
rect 5965 4865 5985 4885
rect 5965 4815 5985 4835
rect 5965 4765 5985 4785
rect 5965 4715 5985 4735
rect 5965 4665 5985 4685
rect 5965 4615 5985 4635
rect 6115 5065 6135 5085
rect 6115 5015 6135 5035
rect 6115 4965 6135 4985
rect 6115 4915 6135 4935
rect 6115 4865 6135 4885
rect 6115 4815 6135 4835
rect 6115 4765 6135 4785
rect 6115 4715 6135 4735
rect 6115 4665 6135 4685
rect 6115 4615 6135 4635
rect 6265 5065 6285 5085
rect 6265 5015 6285 5035
rect 6265 4965 6285 4985
rect 6265 4915 6285 4935
rect 6265 4865 6285 4885
rect 6265 4815 6285 4835
rect 6265 4765 6285 4785
rect 6265 4715 6285 4735
rect 6265 4665 6285 4685
rect 6265 4615 6285 4635
rect 6415 5065 6435 5085
rect 6415 5015 6435 5035
rect 6415 4965 6435 4985
rect 6415 4915 6435 4935
rect 6415 4865 6435 4885
rect 6415 4815 6435 4835
rect 6415 4765 6435 4785
rect 6415 4715 6435 4735
rect 6415 4665 6435 4685
rect 6415 4615 6435 4635
rect 6565 5065 6585 5085
rect 6565 5015 6585 5035
rect 6565 4965 6585 4985
rect 6565 4915 6585 4935
rect 6565 4865 6585 4885
rect 6565 4815 6585 4835
rect 6565 4765 6585 4785
rect 6565 4715 6585 4735
rect 6565 4665 6585 4685
rect 6565 4615 6585 4635
rect 6715 5065 6735 5085
rect 6715 5015 6735 5035
rect 6715 4965 6735 4985
rect 6715 4915 6735 4935
rect 6715 4865 6735 4885
rect 6715 4815 6735 4835
rect 6715 4765 6735 4785
rect 6715 4715 6735 4735
rect 6715 4665 6735 4685
rect 6715 4615 6735 4635
rect 6865 5065 6885 5085
rect 6865 5015 6885 5035
rect 6865 4965 6885 4985
rect 6865 4915 6885 4935
rect 6865 4865 6885 4885
rect 6865 4815 6885 4835
rect 6865 4765 6885 4785
rect 6865 4715 6885 4735
rect 6865 4665 6885 4685
rect 6865 4615 6885 4635
rect 7015 5065 7035 5085
rect 7015 5015 7035 5035
rect 7015 4965 7035 4985
rect 7015 4915 7035 4935
rect 7015 4865 7035 4885
rect 7015 4815 7035 4835
rect 7015 4765 7035 4785
rect 7015 4715 7035 4735
rect 7015 4665 7035 4685
rect 7015 4615 7035 4635
rect 7165 5065 7185 5085
rect 7165 5015 7185 5035
rect 7165 4965 7185 4985
rect 7165 4915 7185 4935
rect 7165 4865 7185 4885
rect 7165 4815 7185 4835
rect 7165 4765 7185 4785
rect 7165 4715 7185 4735
rect 7165 4665 7185 4685
rect 7165 4615 7185 4635
rect 7315 5065 7335 5085
rect 7315 5015 7335 5035
rect 7315 4965 7335 4985
rect 7315 4915 7335 4935
rect 7315 4865 7335 4885
rect 7315 4815 7335 4835
rect 7315 4765 7335 4785
rect 7315 4715 7335 4735
rect 7315 4665 7335 4685
rect 7315 4615 7335 4635
rect 7465 5065 7485 5085
rect 7465 5015 7485 5035
rect 7465 4965 7485 4985
rect 7465 4915 7485 4935
rect 7465 4865 7485 4885
rect 7465 4815 7485 4835
rect 7465 4765 7485 4785
rect 7465 4715 7485 4735
rect 7465 4665 7485 4685
rect 7465 4615 7485 4635
rect 7615 5065 7635 5085
rect 7615 5015 7635 5035
rect 7615 4965 7635 4985
rect 7615 4915 7635 4935
rect 7615 4865 7635 4885
rect 7615 4815 7635 4835
rect 7615 4765 7635 4785
rect 7615 4715 7635 4735
rect 7615 4665 7635 4685
rect 7615 4615 7635 4635
rect 7765 5065 7785 5085
rect 7765 5015 7785 5035
rect 7765 4965 7785 4985
rect 7765 4915 7785 4935
rect 7765 4865 7785 4885
rect 7765 4815 7785 4835
rect 7765 4765 7785 4785
rect 7765 4715 7785 4735
rect 7765 4665 7785 4685
rect 7765 4615 7785 4635
rect 8365 5065 8385 5085
rect 8365 5015 8385 5035
rect 8365 4965 8385 4985
rect 8365 4915 8385 4935
rect 8365 4865 8385 4885
rect 8365 4815 8385 4835
rect 8365 4765 8385 4785
rect 8365 4715 8385 4735
rect 8365 4665 8385 4685
rect 8365 4615 8385 4635
rect 8515 5065 8535 5085
rect 8515 5015 8535 5035
rect 8515 4965 8535 4985
rect 8515 4915 8535 4935
rect 8515 4865 8535 4885
rect 8515 4815 8535 4835
rect 8515 4765 8535 4785
rect 8515 4715 8535 4735
rect 8515 4665 8535 4685
rect 8515 4615 8535 4635
rect 8665 5065 8685 5085
rect 8665 5015 8685 5035
rect 8665 4965 8685 4985
rect 8665 4915 8685 4935
rect 8665 4865 8685 4885
rect 8665 4815 8685 4835
rect 8665 4765 8685 4785
rect 8665 4715 8685 4735
rect 8665 4665 8685 4685
rect 8665 4615 8685 4635
rect 8815 5065 8835 5085
rect 8815 5015 8835 5035
rect 8815 4965 8835 4985
rect 8815 4915 8835 4935
rect 8815 4865 8835 4885
rect 8815 4815 8835 4835
rect 8815 4765 8835 4785
rect 8815 4715 8835 4735
rect 8815 4665 8835 4685
rect 8815 4615 8835 4635
rect 8965 5065 8985 5085
rect 8965 5015 8985 5035
rect 8965 4965 8985 4985
rect 8965 4915 8985 4935
rect 8965 4865 8985 4885
rect 8965 4815 8985 4835
rect 8965 4765 8985 4785
rect 8965 4715 8985 4735
rect 8965 4665 8985 4685
rect 8965 4615 8985 4635
rect 9115 5065 9135 5085
rect 9115 5015 9135 5035
rect 9115 4965 9135 4985
rect 9115 4915 9135 4935
rect 9115 4865 9135 4885
rect 9115 4815 9135 4835
rect 9115 4765 9135 4785
rect 9115 4715 9135 4735
rect 9115 4665 9135 4685
rect 9115 4615 9135 4635
rect 9265 5065 9285 5085
rect 9265 5015 9285 5035
rect 9265 4965 9285 4985
rect 9265 4915 9285 4935
rect 9265 4865 9285 4885
rect 9265 4815 9285 4835
rect 9265 4765 9285 4785
rect 9265 4715 9285 4735
rect 9265 4665 9285 4685
rect 9265 4615 9285 4635
rect 9415 5065 9435 5085
rect 9415 5015 9435 5035
rect 9415 4965 9435 4985
rect 9415 4915 9435 4935
rect 9415 4865 9435 4885
rect 9415 4815 9435 4835
rect 9415 4765 9435 4785
rect 9415 4715 9435 4735
rect 9415 4665 9435 4685
rect 9415 4615 9435 4635
rect 9565 5065 9585 5085
rect 9565 5015 9585 5035
rect 9565 4965 9585 4985
rect 9565 4915 9585 4935
rect 9565 4865 9585 4885
rect 9565 4815 9585 4835
rect 9565 4765 9585 4785
rect 9565 4715 9585 4735
rect 9565 4665 9585 4685
rect 9565 4615 9585 4635
rect 9715 5065 9735 5085
rect 9715 5015 9735 5035
rect 9715 4965 9735 4985
rect 9715 4915 9735 4935
rect 9715 4865 9735 4885
rect 9715 4815 9735 4835
rect 9715 4765 9735 4785
rect 9715 4715 9735 4735
rect 9715 4665 9735 4685
rect 9715 4615 9735 4635
rect 9865 5065 9885 5085
rect 9865 5015 9885 5035
rect 9865 4965 9885 4985
rect 9865 4915 9885 4935
rect 9865 4865 9885 4885
rect 9865 4815 9885 4835
rect 9865 4765 9885 4785
rect 9865 4715 9885 4735
rect 9865 4665 9885 4685
rect 9865 4615 9885 4635
rect 10015 5065 10035 5085
rect 10015 5015 10035 5035
rect 10015 4965 10035 4985
rect 10015 4915 10035 4935
rect 10015 4865 10035 4885
rect 10015 4815 10035 4835
rect 10015 4765 10035 4785
rect 10015 4715 10035 4735
rect 10015 4665 10035 4685
rect 10015 4615 10035 4635
rect 10165 5065 10185 5085
rect 10165 5015 10185 5035
rect 10165 4965 10185 4985
rect 10165 4915 10185 4935
rect 10165 4865 10185 4885
rect 10165 4815 10185 4835
rect 10165 4765 10185 4785
rect 10165 4715 10185 4735
rect 10165 4665 10185 4685
rect 10165 4615 10185 4635
rect 10315 5065 10335 5085
rect 10315 5015 10335 5035
rect 10315 4965 10335 4985
rect 10315 4915 10335 4935
rect 10315 4865 10335 4885
rect 10315 4815 10335 4835
rect 10315 4765 10335 4785
rect 10315 4715 10335 4735
rect 10315 4665 10335 4685
rect 10315 4615 10335 4635
rect 10465 5065 10485 5085
rect 10465 5015 10485 5035
rect 10465 4965 10485 4985
rect 10465 4915 10485 4935
rect 10465 4865 10485 4885
rect 10465 4815 10485 4835
rect 10465 4765 10485 4785
rect 10465 4715 10485 4735
rect 10465 4665 10485 4685
rect 10465 4615 10485 4635
rect 10615 5065 10635 5085
rect 10615 5015 10635 5035
rect 10615 4965 10635 4985
rect 10615 4915 10635 4935
rect 10615 4865 10635 4885
rect 10615 4815 10635 4835
rect 10615 4765 10635 4785
rect 10615 4715 10635 4735
rect 10615 4665 10635 4685
rect 10615 4615 10635 4635
rect 10765 5065 10785 5085
rect 10765 5015 10785 5035
rect 10765 4965 10785 4985
rect 10765 4915 10785 4935
rect 10765 4865 10785 4885
rect 10765 4815 10785 4835
rect 10765 4765 10785 4785
rect 10765 4715 10785 4735
rect 10765 4665 10785 4685
rect 10765 4615 10785 4635
rect 11365 5065 11385 5085
rect 11365 5015 11385 5035
rect 11365 4965 11385 4985
rect 11365 4915 11385 4935
rect 11365 4865 11385 4885
rect 11365 4815 11385 4835
rect 11365 4765 11385 4785
rect 11365 4715 11385 4735
rect 11365 4665 11385 4685
rect 11365 4615 11385 4635
rect 11965 5065 11985 5085
rect 11965 5015 11985 5035
rect 11965 4965 11985 4985
rect 11965 4915 11985 4935
rect 11965 4865 11985 4885
rect 11965 4815 11985 4835
rect 11965 4765 11985 4785
rect 11965 4715 11985 4735
rect 11965 4665 11985 4685
rect 11965 4615 11985 4635
rect 12565 5065 12585 5085
rect 12565 5015 12585 5035
rect 12565 4965 12585 4985
rect 12565 4915 12585 4935
rect 12565 4865 12585 4885
rect 12565 4815 12585 4835
rect 12565 4765 12585 4785
rect 12565 4715 12585 4735
rect 12565 4665 12585 4685
rect 12565 4615 12585 4635
rect 13165 5065 13185 5085
rect 13165 5015 13185 5035
rect 13165 4965 13185 4985
rect 13165 4915 13185 4935
rect 13165 4865 13185 4885
rect 13165 4815 13185 4835
rect 13165 4765 13185 4785
rect 13165 4715 13185 4735
rect 13165 4665 13185 4685
rect 13165 4615 13185 4635
rect 13765 5065 13785 5085
rect 13765 5015 13785 5035
rect 13765 4965 13785 4985
rect 13765 4915 13785 4935
rect 13765 4865 13785 4885
rect 13765 4815 13785 4835
rect 13765 4765 13785 4785
rect 13765 4715 13785 4735
rect 13765 4665 13785 4685
rect 13765 4615 13785 4635
rect 14365 5065 14385 5085
rect 14365 5015 14385 5035
rect 14365 4965 14385 4985
rect 14365 4915 14385 4935
rect 14365 4865 14385 4885
rect 14365 4815 14385 4835
rect 14365 4765 14385 4785
rect 14365 4715 14385 4735
rect 14365 4665 14385 4685
rect 14365 4615 14385 4635
rect 14965 5065 14985 5085
rect 14965 5015 14985 5035
rect 14965 4965 14985 4985
rect 14965 4915 14985 4935
rect 14965 4865 14985 4885
rect 14965 4815 14985 4835
rect 14965 4765 14985 4785
rect 14965 4715 14985 4735
rect 14965 4665 14985 4685
rect 14965 4615 14985 4635
rect 15565 5065 15585 5085
rect 15565 5015 15585 5035
rect 15565 4965 15585 4985
rect 15565 4915 15585 4935
rect 15565 4865 15585 4885
rect 15565 4815 15585 4835
rect 15565 4765 15585 4785
rect 15565 4715 15585 4735
rect 15565 4665 15585 4685
rect 15565 4615 15585 4635
rect 16165 5065 16185 5085
rect 16165 5015 16185 5035
rect 16165 4965 16185 4985
rect 16165 4915 16185 4935
rect 16165 4865 16185 4885
rect 16165 4815 16185 4835
rect 16165 4765 16185 4785
rect 16165 4715 16185 4735
rect 16165 4665 16185 4685
rect 16165 4615 16185 4635
rect 16315 5065 16335 5085
rect 16315 5015 16335 5035
rect 16315 4965 16335 4985
rect 16315 4915 16335 4935
rect 16315 4865 16335 4885
rect 16315 4815 16335 4835
rect 16315 4765 16335 4785
rect 16315 4715 16335 4735
rect 16315 4665 16335 4685
rect 16315 4615 16335 4635
rect 16465 5065 16485 5085
rect 16465 5015 16485 5035
rect 16465 4965 16485 4985
rect 16465 4915 16485 4935
rect 16465 4865 16485 4885
rect 16465 4815 16485 4835
rect 16465 4765 16485 4785
rect 16465 4715 16485 4735
rect 16465 4665 16485 4685
rect 16465 4615 16485 4635
rect 16615 5065 16635 5085
rect 16615 5015 16635 5035
rect 16615 4965 16635 4985
rect 16615 4915 16635 4935
rect 16615 4865 16635 4885
rect 16615 4815 16635 4835
rect 16615 4765 16635 4785
rect 16615 4715 16635 4735
rect 16615 4665 16635 4685
rect 16615 4615 16635 4635
rect 16765 5065 16785 5085
rect 16765 5015 16785 5035
rect 16765 4965 16785 4985
rect 16765 4915 16785 4935
rect 16765 4865 16785 4885
rect 16765 4815 16785 4835
rect 16765 4765 16785 4785
rect 16765 4715 16785 4735
rect 16765 4665 16785 4685
rect 16765 4615 16785 4635
rect 16915 5065 16935 5085
rect 16915 5015 16935 5035
rect 16915 4965 16935 4985
rect 16915 4915 16935 4935
rect 16915 4865 16935 4885
rect 16915 4815 16935 4835
rect 16915 4765 16935 4785
rect 16915 4715 16935 4735
rect 16915 4665 16935 4685
rect 16915 4615 16935 4635
rect 17065 5065 17085 5085
rect 17065 5015 17085 5035
rect 17065 4965 17085 4985
rect 17065 4915 17085 4935
rect 17065 4865 17085 4885
rect 17065 4815 17085 4835
rect 17065 4765 17085 4785
rect 17065 4715 17085 4735
rect 17065 4665 17085 4685
rect 17065 4615 17085 4635
rect 17215 5065 17235 5085
rect 17215 5015 17235 5035
rect 17215 4965 17235 4985
rect 17215 4915 17235 4935
rect 17215 4865 17235 4885
rect 17215 4815 17235 4835
rect 17215 4765 17235 4785
rect 17215 4715 17235 4735
rect 17215 4665 17235 4685
rect 17215 4615 17235 4635
rect 17365 5065 17385 5085
rect 17365 5015 17385 5035
rect 17365 4965 17385 4985
rect 17365 4915 17385 4935
rect 17365 4865 17385 4885
rect 17365 4815 17385 4835
rect 17365 4765 17385 4785
rect 17365 4715 17385 4735
rect 17365 4665 17385 4685
rect 17365 4615 17385 4635
rect 17965 5065 17985 5085
rect 17965 5015 17985 5035
rect 17965 4965 17985 4985
rect 17965 4915 17985 4935
rect 17965 4865 17985 4885
rect 17965 4815 17985 4835
rect 17965 4765 17985 4785
rect 17965 4715 17985 4735
rect 17965 4665 17985 4685
rect 17965 4615 17985 4635
rect 18565 5065 18585 5085
rect 18565 5015 18585 5035
rect 18565 4965 18585 4985
rect 18565 4915 18585 4935
rect 18565 4865 18585 4885
rect 18565 4815 18585 4835
rect 18565 4765 18585 4785
rect 18565 4715 18585 4735
rect 18565 4665 18585 4685
rect 18565 4615 18585 4635
rect 18715 5065 18735 5085
rect 18715 5015 18735 5035
rect 18715 4965 18735 4985
rect 18715 4915 18735 4935
rect 18715 4865 18735 4885
rect 18715 4815 18735 4835
rect 18715 4765 18735 4785
rect 18715 4715 18735 4735
rect 18715 4665 18735 4685
rect 18715 4615 18735 4635
rect 18865 5065 18885 5085
rect 18865 5015 18885 5035
rect 18865 4965 18885 4985
rect 18865 4915 18885 4935
rect 18865 4865 18885 4885
rect 18865 4815 18885 4835
rect 18865 4765 18885 4785
rect 18865 4715 18885 4735
rect 18865 4665 18885 4685
rect 18865 4615 18885 4635
rect 19015 5065 19035 5085
rect 19015 5015 19035 5035
rect 19015 4965 19035 4985
rect 19015 4915 19035 4935
rect 19015 4865 19035 4885
rect 19015 4815 19035 4835
rect 19015 4765 19035 4785
rect 19015 4715 19035 4735
rect 19015 4665 19035 4685
rect 19015 4615 19035 4635
rect 19165 5065 19185 5085
rect 19165 5015 19185 5035
rect 19165 4965 19185 4985
rect 19165 4915 19185 4935
rect 19165 4865 19185 4885
rect 19165 4815 19185 4835
rect 19165 4765 19185 4785
rect 19165 4715 19185 4735
rect 19165 4665 19185 4685
rect 19165 4615 19185 4635
rect 19315 5065 19335 5085
rect 19315 5015 19335 5035
rect 19315 4965 19335 4985
rect 19315 4915 19335 4935
rect 19315 4865 19335 4885
rect 19315 4815 19335 4835
rect 19315 4765 19335 4785
rect 19315 4715 19335 4735
rect 19315 4665 19335 4685
rect 19315 4615 19335 4635
rect 19465 5065 19485 5085
rect 19465 5015 19485 5035
rect 19465 4965 19485 4985
rect 19465 4915 19485 4935
rect 19465 4865 19485 4885
rect 19465 4815 19485 4835
rect 19465 4765 19485 4785
rect 19465 4715 19485 4735
rect 19465 4665 19485 4685
rect 19465 4615 19485 4635
rect 19615 5065 19635 5085
rect 19615 5015 19635 5035
rect 19615 4965 19635 4985
rect 19615 4915 19635 4935
rect 19615 4865 19635 4885
rect 19615 4815 19635 4835
rect 19615 4765 19635 4785
rect 19615 4715 19635 4735
rect 19615 4665 19635 4685
rect 19615 4615 19635 4635
rect 19765 5065 19785 5085
rect 19765 5015 19785 5035
rect 19765 4965 19785 4985
rect 19765 4915 19785 4935
rect 19765 4865 19785 4885
rect 19765 4815 19785 4835
rect 19765 4765 19785 4785
rect 19765 4715 19785 4735
rect 19765 4665 19785 4685
rect 19765 4615 19785 4635
rect 20365 5065 20385 5085
rect 20365 5015 20385 5035
rect 20365 4965 20385 4985
rect 20365 4915 20385 4935
rect 20365 4865 20385 4885
rect 20365 4815 20385 4835
rect 20365 4765 20385 4785
rect 20365 4715 20385 4735
rect 20365 4665 20385 4685
rect 20365 4615 20385 4635
rect -635 4415 -615 4435
rect -635 4365 -615 4385
rect -635 4315 -615 4335
rect -635 4265 -615 4285
rect -635 4215 -615 4235
rect -635 4165 -615 4185
rect -635 4115 -615 4135
rect -635 4065 -615 4085
rect -635 4015 -615 4035
rect -635 3965 -615 3985
rect -485 4415 -465 4435
rect -485 4365 -465 4385
rect -485 4315 -465 4335
rect -485 4265 -465 4285
rect -485 4215 -465 4235
rect -485 4165 -465 4185
rect -485 4115 -465 4135
rect -485 4065 -465 4085
rect -485 4015 -465 4035
rect -485 3965 -465 3985
rect -335 4415 -315 4435
rect -335 4365 -315 4385
rect -335 4315 -315 4335
rect -335 4265 -315 4285
rect -335 4215 -315 4235
rect -335 4165 -315 4185
rect -335 4115 -315 4135
rect -335 4065 -315 4085
rect -335 4015 -315 4035
rect -335 3965 -315 3985
rect -185 4415 -165 4435
rect -185 4365 -165 4385
rect -185 4315 -165 4335
rect -185 4265 -165 4285
rect -185 4215 -165 4235
rect -185 4165 -165 4185
rect -185 4115 -165 4135
rect -185 4065 -165 4085
rect -185 4015 -165 4035
rect -185 3965 -165 3985
rect -35 4415 -15 4435
rect -35 4365 -15 4385
rect -35 4315 -15 4335
rect -35 4265 -15 4285
rect -35 4215 -15 4235
rect -35 4165 -15 4185
rect -35 4115 -15 4135
rect -35 4065 -15 4085
rect -35 4015 -15 4035
rect -35 3965 -15 3985
rect 565 4415 585 4435
rect 565 4365 585 4385
rect 565 4315 585 4335
rect 565 4265 585 4285
rect 565 4215 585 4235
rect 565 4165 585 4185
rect 565 4115 585 4135
rect 565 4065 585 4085
rect 565 4015 585 4035
rect 565 3965 585 3985
rect 715 4415 735 4435
rect 715 4365 735 4385
rect 715 4315 735 4335
rect 715 4265 735 4285
rect 715 4215 735 4235
rect 715 4165 735 4185
rect 715 4115 735 4135
rect 715 4065 735 4085
rect 715 4015 735 4035
rect 715 3965 735 3985
rect 865 4415 885 4435
rect 865 4365 885 4385
rect 865 4315 885 4335
rect 865 4265 885 4285
rect 865 4215 885 4235
rect 865 4165 885 4185
rect 865 4115 885 4135
rect 865 4065 885 4085
rect 865 4015 885 4035
rect 865 3965 885 3985
rect 1015 4415 1035 4435
rect 1015 4365 1035 4385
rect 1015 4315 1035 4335
rect 1015 4265 1035 4285
rect 1015 4215 1035 4235
rect 1015 4165 1035 4185
rect 1015 4115 1035 4135
rect 1015 4065 1035 4085
rect 1015 4015 1035 4035
rect 1015 3965 1035 3985
rect 1165 4415 1185 4435
rect 1165 4365 1185 4385
rect 1165 4315 1185 4335
rect 1165 4265 1185 4285
rect 1165 4215 1185 4235
rect 1165 4165 1185 4185
rect 1165 4115 1185 4135
rect 1165 4065 1185 4085
rect 1165 4015 1185 4035
rect 1165 3965 1185 3985
rect 1315 4415 1335 4435
rect 1315 4365 1335 4385
rect 1315 4315 1335 4335
rect 1315 4265 1335 4285
rect 1315 4215 1335 4235
rect 1315 4165 1335 4185
rect 1315 4115 1335 4135
rect 1315 4065 1335 4085
rect 1315 4015 1335 4035
rect 1315 3965 1335 3985
rect 1465 4415 1485 4435
rect 1465 4365 1485 4385
rect 1465 4315 1485 4335
rect 1465 4265 1485 4285
rect 1465 4215 1485 4235
rect 1465 4165 1485 4185
rect 1465 4115 1485 4135
rect 1465 4065 1485 4085
rect 1465 4015 1485 4035
rect 1465 3965 1485 3985
rect 1615 4415 1635 4435
rect 1615 4365 1635 4385
rect 1615 4315 1635 4335
rect 1615 4265 1635 4285
rect 1615 4215 1635 4235
rect 1615 4165 1635 4185
rect 1615 4115 1635 4135
rect 1615 4065 1635 4085
rect 1615 4015 1635 4035
rect 1615 3965 1635 3985
rect 1765 4415 1785 4435
rect 1765 4365 1785 4385
rect 1765 4315 1785 4335
rect 1765 4265 1785 4285
rect 1765 4215 1785 4235
rect 1765 4165 1785 4185
rect 1765 4115 1785 4135
rect 1765 4065 1785 4085
rect 1765 4015 1785 4035
rect 1765 3965 1785 3985
rect 1915 4415 1935 4435
rect 1915 4365 1935 4385
rect 1915 4315 1935 4335
rect 1915 4265 1935 4285
rect 1915 4215 1935 4235
rect 1915 4165 1935 4185
rect 1915 4115 1935 4135
rect 1915 4065 1935 4085
rect 1915 4015 1935 4035
rect 1915 3965 1935 3985
rect 2065 4415 2085 4435
rect 2065 4365 2085 4385
rect 2065 4315 2085 4335
rect 2065 4265 2085 4285
rect 2065 4215 2085 4235
rect 2065 4165 2085 4185
rect 2065 4115 2085 4135
rect 2065 4065 2085 4085
rect 2065 4015 2085 4035
rect 2065 3965 2085 3985
rect 2215 4415 2235 4435
rect 2215 4365 2235 4385
rect 2215 4315 2235 4335
rect 2215 4265 2235 4285
rect 2215 4215 2235 4235
rect 2215 4165 2235 4185
rect 2215 4115 2235 4135
rect 2215 4065 2235 4085
rect 2215 4015 2235 4035
rect 2215 3965 2235 3985
rect 2365 4415 2385 4435
rect 2365 4365 2385 4385
rect 2365 4315 2385 4335
rect 2365 4265 2385 4285
rect 2365 4215 2385 4235
rect 2365 4165 2385 4185
rect 2365 4115 2385 4135
rect 2365 4065 2385 4085
rect 2365 4015 2385 4035
rect 2365 3965 2385 3985
rect 2515 4415 2535 4435
rect 2515 4365 2535 4385
rect 2515 4315 2535 4335
rect 2515 4265 2535 4285
rect 2515 4215 2535 4235
rect 2515 4165 2535 4185
rect 2515 4115 2535 4135
rect 2515 4065 2535 4085
rect 2515 4015 2535 4035
rect 2515 3965 2535 3985
rect 2665 4415 2685 4435
rect 2665 4365 2685 4385
rect 2665 4315 2685 4335
rect 2665 4265 2685 4285
rect 2665 4215 2685 4235
rect 2665 4165 2685 4185
rect 2665 4115 2685 4135
rect 2665 4065 2685 4085
rect 2665 4015 2685 4035
rect 2665 3965 2685 3985
rect 2815 4415 2835 4435
rect 2815 4365 2835 4385
rect 2815 4315 2835 4335
rect 2815 4265 2835 4285
rect 2815 4215 2835 4235
rect 2815 4165 2835 4185
rect 2815 4115 2835 4135
rect 2815 4065 2835 4085
rect 2815 4015 2835 4035
rect 2815 3965 2835 3985
rect 2965 4415 2985 4435
rect 2965 4365 2985 4385
rect 2965 4315 2985 4335
rect 2965 4265 2985 4285
rect 2965 4215 2985 4235
rect 2965 4165 2985 4185
rect 2965 4115 2985 4135
rect 2965 4065 2985 4085
rect 2965 4015 2985 4035
rect 2965 3965 2985 3985
rect 3115 4415 3135 4435
rect 3115 4365 3135 4385
rect 3115 4315 3135 4335
rect 3115 4265 3135 4285
rect 3115 4215 3135 4235
rect 3115 4165 3135 4185
rect 3115 4115 3135 4135
rect 3115 4065 3135 4085
rect 3115 4015 3135 4035
rect 3115 3965 3135 3985
rect 3265 4415 3285 4435
rect 3265 4365 3285 4385
rect 3265 4315 3285 4335
rect 3265 4265 3285 4285
rect 3265 4215 3285 4235
rect 3265 4165 3285 4185
rect 3265 4115 3285 4135
rect 3265 4065 3285 4085
rect 3265 4015 3285 4035
rect 3265 3965 3285 3985
rect 3415 4415 3435 4435
rect 3415 4365 3435 4385
rect 3415 4315 3435 4335
rect 3415 4265 3435 4285
rect 3415 4215 3435 4235
rect 3415 4165 3435 4185
rect 3415 4115 3435 4135
rect 3415 4065 3435 4085
rect 3415 4015 3435 4035
rect 3415 3965 3435 3985
rect 3565 4415 3585 4435
rect 3565 4365 3585 4385
rect 3565 4315 3585 4335
rect 3565 4265 3585 4285
rect 3565 4215 3585 4235
rect 3565 4165 3585 4185
rect 3565 4115 3585 4135
rect 3565 4065 3585 4085
rect 3565 4015 3585 4035
rect 3565 3965 3585 3985
rect 4165 4415 4185 4435
rect 4165 4365 4185 4385
rect 4165 4315 4185 4335
rect 4165 4265 4185 4285
rect 4165 4215 4185 4235
rect 4165 4165 4185 4185
rect 4165 4115 4185 4135
rect 4165 4065 4185 4085
rect 4165 4015 4185 4035
rect 4165 3965 4185 3985
rect 4765 4415 4785 4435
rect 4765 4365 4785 4385
rect 4765 4315 4785 4335
rect 4765 4265 4785 4285
rect 4765 4215 4785 4235
rect 4765 4165 4785 4185
rect 4765 4115 4785 4135
rect 4765 4065 4785 4085
rect 4765 4015 4785 4035
rect 4765 3965 4785 3985
rect 4915 4415 4935 4435
rect 4915 4365 4935 4385
rect 4915 4315 4935 4335
rect 4915 4265 4935 4285
rect 4915 4215 4935 4235
rect 4915 4165 4935 4185
rect 4915 4115 4935 4135
rect 4915 4065 4935 4085
rect 4915 4015 4935 4035
rect 4915 3965 4935 3985
rect 5065 4415 5085 4435
rect 5065 4365 5085 4385
rect 5065 4315 5085 4335
rect 5065 4265 5085 4285
rect 5065 4215 5085 4235
rect 5065 4165 5085 4185
rect 5065 4115 5085 4135
rect 5065 4065 5085 4085
rect 5065 4015 5085 4035
rect 5065 3965 5085 3985
rect 5215 4415 5235 4435
rect 5215 4365 5235 4385
rect 5215 4315 5235 4335
rect 5215 4265 5235 4285
rect 5215 4215 5235 4235
rect 5215 4165 5235 4185
rect 5215 4115 5235 4135
rect 5215 4065 5235 4085
rect 5215 4015 5235 4035
rect 5215 3965 5235 3985
rect 5365 4415 5385 4435
rect 5365 4365 5385 4385
rect 5365 4315 5385 4335
rect 5365 4265 5385 4285
rect 5365 4215 5385 4235
rect 5365 4165 5385 4185
rect 5365 4115 5385 4135
rect 5365 4065 5385 4085
rect 5365 4015 5385 4035
rect 5365 3965 5385 3985
rect 5515 4415 5535 4435
rect 5515 4365 5535 4385
rect 5515 4315 5535 4335
rect 5515 4265 5535 4285
rect 5515 4215 5535 4235
rect 5515 4165 5535 4185
rect 5515 4115 5535 4135
rect 5515 4065 5535 4085
rect 5515 4015 5535 4035
rect 5515 3965 5535 3985
rect 5665 4415 5685 4435
rect 5665 4365 5685 4385
rect 5665 4315 5685 4335
rect 5665 4265 5685 4285
rect 5665 4215 5685 4235
rect 5665 4165 5685 4185
rect 5665 4115 5685 4135
rect 5665 4065 5685 4085
rect 5665 4015 5685 4035
rect 5665 3965 5685 3985
rect 5815 4415 5835 4435
rect 5815 4365 5835 4385
rect 5815 4315 5835 4335
rect 5815 4265 5835 4285
rect 5815 4215 5835 4235
rect 5815 4165 5835 4185
rect 5815 4115 5835 4135
rect 5815 4065 5835 4085
rect 5815 4015 5835 4035
rect 5815 3965 5835 3985
rect 5965 4415 5985 4435
rect 5965 4365 5985 4385
rect 5965 4315 5985 4335
rect 5965 4265 5985 4285
rect 5965 4215 5985 4235
rect 5965 4165 5985 4185
rect 5965 4115 5985 4135
rect 5965 4065 5985 4085
rect 5965 4015 5985 4035
rect 5965 3965 5985 3985
rect 6115 4415 6135 4435
rect 6115 4365 6135 4385
rect 6115 4315 6135 4335
rect 6115 4265 6135 4285
rect 6115 4215 6135 4235
rect 6115 4165 6135 4185
rect 6115 4115 6135 4135
rect 6115 4065 6135 4085
rect 6115 4015 6135 4035
rect 6115 3965 6135 3985
rect 6265 4415 6285 4435
rect 6265 4365 6285 4385
rect 6265 4315 6285 4335
rect 6265 4265 6285 4285
rect 6265 4215 6285 4235
rect 6265 4165 6285 4185
rect 6265 4115 6285 4135
rect 6265 4065 6285 4085
rect 6265 4015 6285 4035
rect 6265 3965 6285 3985
rect 6415 4415 6435 4435
rect 6415 4365 6435 4385
rect 6415 4315 6435 4335
rect 6415 4265 6435 4285
rect 6415 4215 6435 4235
rect 6415 4165 6435 4185
rect 6415 4115 6435 4135
rect 6415 4065 6435 4085
rect 6415 4015 6435 4035
rect 6415 3965 6435 3985
rect 6565 4415 6585 4435
rect 6565 4365 6585 4385
rect 6565 4315 6585 4335
rect 6565 4265 6585 4285
rect 6565 4215 6585 4235
rect 6565 4165 6585 4185
rect 6565 4115 6585 4135
rect 6565 4065 6585 4085
rect 6565 4015 6585 4035
rect 6565 3965 6585 3985
rect 6715 4415 6735 4435
rect 6715 4365 6735 4385
rect 6715 4315 6735 4335
rect 6715 4265 6735 4285
rect 6715 4215 6735 4235
rect 6715 4165 6735 4185
rect 6715 4115 6735 4135
rect 6715 4065 6735 4085
rect 6715 4015 6735 4035
rect 6715 3965 6735 3985
rect 6865 4415 6885 4435
rect 6865 4365 6885 4385
rect 6865 4315 6885 4335
rect 6865 4265 6885 4285
rect 6865 4215 6885 4235
rect 6865 4165 6885 4185
rect 6865 4115 6885 4135
rect 6865 4065 6885 4085
rect 6865 4015 6885 4035
rect 6865 3965 6885 3985
rect 7015 4415 7035 4435
rect 7015 4365 7035 4385
rect 7015 4315 7035 4335
rect 7015 4265 7035 4285
rect 7015 4215 7035 4235
rect 7015 4165 7035 4185
rect 7015 4115 7035 4135
rect 7015 4065 7035 4085
rect 7015 4015 7035 4035
rect 7015 3965 7035 3985
rect 7165 4415 7185 4435
rect 7165 4365 7185 4385
rect 7165 4315 7185 4335
rect 7165 4265 7185 4285
rect 7165 4215 7185 4235
rect 7165 4165 7185 4185
rect 7165 4115 7185 4135
rect 7165 4065 7185 4085
rect 7165 4015 7185 4035
rect 7165 3965 7185 3985
rect 7315 4415 7335 4435
rect 7315 4365 7335 4385
rect 7315 4315 7335 4335
rect 7315 4265 7335 4285
rect 7315 4215 7335 4235
rect 7315 4165 7335 4185
rect 7315 4115 7335 4135
rect 7315 4065 7335 4085
rect 7315 4015 7335 4035
rect 7315 3965 7335 3985
rect 7465 4415 7485 4435
rect 7465 4365 7485 4385
rect 7465 4315 7485 4335
rect 7465 4265 7485 4285
rect 7465 4215 7485 4235
rect 7465 4165 7485 4185
rect 7465 4115 7485 4135
rect 7465 4065 7485 4085
rect 7465 4015 7485 4035
rect 7465 3965 7485 3985
rect 7615 4415 7635 4435
rect 7615 4365 7635 4385
rect 7615 4315 7635 4335
rect 7615 4265 7635 4285
rect 7615 4215 7635 4235
rect 7615 4165 7635 4185
rect 7615 4115 7635 4135
rect 7615 4065 7635 4085
rect 7615 4015 7635 4035
rect 7615 3965 7635 3985
rect 7765 4415 7785 4435
rect 7765 4365 7785 4385
rect 7765 4315 7785 4335
rect 7765 4265 7785 4285
rect 7765 4215 7785 4235
rect 7765 4165 7785 4185
rect 7765 4115 7785 4135
rect 7765 4065 7785 4085
rect 7765 4015 7785 4035
rect 7765 3965 7785 3985
rect 8365 4415 8385 4435
rect 8365 4365 8385 4385
rect 8365 4315 8385 4335
rect 8365 4265 8385 4285
rect 8365 4215 8385 4235
rect 8365 4165 8385 4185
rect 8365 4115 8385 4135
rect 8365 4065 8385 4085
rect 8365 4015 8385 4035
rect 8365 3965 8385 3985
rect 8515 4415 8535 4435
rect 8515 4365 8535 4385
rect 8515 4315 8535 4335
rect 8515 4265 8535 4285
rect 8515 4215 8535 4235
rect 8515 4165 8535 4185
rect 8515 4115 8535 4135
rect 8515 4065 8535 4085
rect 8515 4015 8535 4035
rect 8515 3965 8535 3985
rect 8665 4415 8685 4435
rect 8665 4365 8685 4385
rect 8665 4315 8685 4335
rect 8665 4265 8685 4285
rect 8665 4215 8685 4235
rect 8665 4165 8685 4185
rect 8665 4115 8685 4135
rect 8665 4065 8685 4085
rect 8665 4015 8685 4035
rect 8665 3965 8685 3985
rect 8815 4415 8835 4435
rect 8815 4365 8835 4385
rect 8815 4315 8835 4335
rect 8815 4265 8835 4285
rect 8815 4215 8835 4235
rect 8815 4165 8835 4185
rect 8815 4115 8835 4135
rect 8815 4065 8835 4085
rect 8815 4015 8835 4035
rect 8815 3965 8835 3985
rect 8965 4415 8985 4435
rect 8965 4365 8985 4385
rect 8965 4315 8985 4335
rect 8965 4265 8985 4285
rect 8965 4215 8985 4235
rect 8965 4165 8985 4185
rect 8965 4115 8985 4135
rect 8965 4065 8985 4085
rect 8965 4015 8985 4035
rect 8965 3965 8985 3985
rect 9115 4415 9135 4435
rect 9115 4365 9135 4385
rect 9115 4315 9135 4335
rect 9115 4265 9135 4285
rect 9115 4215 9135 4235
rect 9115 4165 9135 4185
rect 9115 4115 9135 4135
rect 9115 4065 9135 4085
rect 9115 4015 9135 4035
rect 9115 3965 9135 3985
rect 9265 4415 9285 4435
rect 9265 4365 9285 4385
rect 9265 4315 9285 4335
rect 9265 4265 9285 4285
rect 9265 4215 9285 4235
rect 9265 4165 9285 4185
rect 9265 4115 9285 4135
rect 9265 4065 9285 4085
rect 9265 4015 9285 4035
rect 9265 3965 9285 3985
rect 9415 4415 9435 4435
rect 9415 4365 9435 4385
rect 9415 4315 9435 4335
rect 9415 4265 9435 4285
rect 9415 4215 9435 4235
rect 9415 4165 9435 4185
rect 9415 4115 9435 4135
rect 9415 4065 9435 4085
rect 9415 4015 9435 4035
rect 9415 3965 9435 3985
rect 9565 4415 9585 4435
rect 9565 4365 9585 4385
rect 9565 4315 9585 4335
rect 9565 4265 9585 4285
rect 9565 4215 9585 4235
rect 9565 4165 9585 4185
rect 9565 4115 9585 4135
rect 9565 4065 9585 4085
rect 9565 4015 9585 4035
rect 9565 3965 9585 3985
rect 9715 4415 9735 4435
rect 9715 4365 9735 4385
rect 9715 4315 9735 4335
rect 9715 4265 9735 4285
rect 9715 4215 9735 4235
rect 9715 4165 9735 4185
rect 9715 4115 9735 4135
rect 9715 4065 9735 4085
rect 9715 4015 9735 4035
rect 9715 3965 9735 3985
rect 9865 4415 9885 4435
rect 9865 4365 9885 4385
rect 9865 4315 9885 4335
rect 9865 4265 9885 4285
rect 9865 4215 9885 4235
rect 9865 4165 9885 4185
rect 9865 4115 9885 4135
rect 9865 4065 9885 4085
rect 9865 4015 9885 4035
rect 9865 3965 9885 3985
rect 10015 4415 10035 4435
rect 10015 4365 10035 4385
rect 10015 4315 10035 4335
rect 10015 4265 10035 4285
rect 10015 4215 10035 4235
rect 10015 4165 10035 4185
rect 10015 4115 10035 4135
rect 10015 4065 10035 4085
rect 10015 4015 10035 4035
rect 10015 3965 10035 3985
rect 10165 4415 10185 4435
rect 10165 4365 10185 4385
rect 10165 4315 10185 4335
rect 10165 4265 10185 4285
rect 10165 4215 10185 4235
rect 10165 4165 10185 4185
rect 10165 4115 10185 4135
rect 10165 4065 10185 4085
rect 10165 4015 10185 4035
rect 10165 3965 10185 3985
rect 10315 4415 10335 4435
rect 10315 4365 10335 4385
rect 10315 4315 10335 4335
rect 10315 4265 10335 4285
rect 10315 4215 10335 4235
rect 10315 4165 10335 4185
rect 10315 4115 10335 4135
rect 10315 4065 10335 4085
rect 10315 4015 10335 4035
rect 10315 3965 10335 3985
rect 10465 4415 10485 4435
rect 10465 4365 10485 4385
rect 10465 4315 10485 4335
rect 10465 4265 10485 4285
rect 10465 4215 10485 4235
rect 10465 4165 10485 4185
rect 10465 4115 10485 4135
rect 10465 4065 10485 4085
rect 10465 4015 10485 4035
rect 10465 3965 10485 3985
rect 10615 4415 10635 4435
rect 10615 4365 10635 4385
rect 10615 4315 10635 4335
rect 10615 4265 10635 4285
rect 10615 4215 10635 4235
rect 10615 4165 10635 4185
rect 10615 4115 10635 4135
rect 10615 4065 10635 4085
rect 10615 4015 10635 4035
rect 10615 3965 10635 3985
rect 10765 4415 10785 4435
rect 10765 4365 10785 4385
rect 10765 4315 10785 4335
rect 10765 4265 10785 4285
rect 10765 4215 10785 4235
rect 10765 4165 10785 4185
rect 10765 4115 10785 4135
rect 10765 4065 10785 4085
rect 10765 4015 10785 4035
rect 10765 3965 10785 3985
rect 11365 4415 11385 4435
rect 11365 4365 11385 4385
rect 11365 4315 11385 4335
rect 11365 4265 11385 4285
rect 11365 4215 11385 4235
rect 11365 4165 11385 4185
rect 11365 4115 11385 4135
rect 11365 4065 11385 4085
rect 11365 4015 11385 4035
rect 11365 3965 11385 3985
rect 11965 4415 11985 4435
rect 11965 4365 11985 4385
rect 11965 4315 11985 4335
rect 11965 4265 11985 4285
rect 11965 4215 11985 4235
rect 11965 4165 11985 4185
rect 11965 4115 11985 4135
rect 11965 4065 11985 4085
rect 11965 4015 11985 4035
rect 11965 3965 11985 3985
rect 12565 4415 12585 4435
rect 12565 4365 12585 4385
rect 12565 4315 12585 4335
rect 12565 4265 12585 4285
rect 12565 4215 12585 4235
rect 12565 4165 12585 4185
rect 12565 4115 12585 4135
rect 12565 4065 12585 4085
rect 12565 4015 12585 4035
rect 12565 3965 12585 3985
rect 13165 4415 13185 4435
rect 13165 4365 13185 4385
rect 13165 4315 13185 4335
rect 13165 4265 13185 4285
rect 13165 4215 13185 4235
rect 13165 4165 13185 4185
rect 13165 4115 13185 4135
rect 13165 4065 13185 4085
rect 13165 4015 13185 4035
rect 13165 3965 13185 3985
rect 13765 4415 13785 4435
rect 13765 4365 13785 4385
rect 13765 4315 13785 4335
rect 13765 4265 13785 4285
rect 13765 4215 13785 4235
rect 13765 4165 13785 4185
rect 13765 4115 13785 4135
rect 13765 4065 13785 4085
rect 13765 4015 13785 4035
rect 13765 3965 13785 3985
rect 14365 4415 14385 4435
rect 14365 4365 14385 4385
rect 14365 4315 14385 4335
rect 14365 4265 14385 4285
rect 14365 4215 14385 4235
rect 14365 4165 14385 4185
rect 14365 4115 14385 4135
rect 14365 4065 14385 4085
rect 14365 4015 14385 4035
rect 14365 3965 14385 3985
rect 14965 4415 14985 4435
rect 14965 4365 14985 4385
rect 14965 4315 14985 4335
rect 14965 4265 14985 4285
rect 14965 4215 14985 4235
rect 14965 4165 14985 4185
rect 14965 4115 14985 4135
rect 14965 4065 14985 4085
rect 14965 4015 14985 4035
rect 14965 3965 14985 3985
rect 15565 4415 15585 4435
rect 15565 4365 15585 4385
rect 15565 4315 15585 4335
rect 15565 4265 15585 4285
rect 15565 4215 15585 4235
rect 15565 4165 15585 4185
rect 15565 4115 15585 4135
rect 15565 4065 15585 4085
rect 15565 4015 15585 4035
rect 15565 3965 15585 3985
rect 16165 4415 16185 4435
rect 16165 4365 16185 4385
rect 16165 4315 16185 4335
rect 16165 4265 16185 4285
rect 16165 4215 16185 4235
rect 16165 4165 16185 4185
rect 16165 4115 16185 4135
rect 16165 4065 16185 4085
rect 16165 4015 16185 4035
rect 16165 3965 16185 3985
rect 16315 4415 16335 4435
rect 16315 4365 16335 4385
rect 16315 4315 16335 4335
rect 16315 4265 16335 4285
rect 16315 4215 16335 4235
rect 16315 4165 16335 4185
rect 16315 4115 16335 4135
rect 16315 4065 16335 4085
rect 16315 4015 16335 4035
rect 16315 3965 16335 3985
rect 16465 4415 16485 4435
rect 16465 4365 16485 4385
rect 16465 4315 16485 4335
rect 16465 4265 16485 4285
rect 16465 4215 16485 4235
rect 16465 4165 16485 4185
rect 16465 4115 16485 4135
rect 16465 4065 16485 4085
rect 16465 4015 16485 4035
rect 16465 3965 16485 3985
rect 16615 4415 16635 4435
rect 16615 4365 16635 4385
rect 16615 4315 16635 4335
rect 16615 4265 16635 4285
rect 16615 4215 16635 4235
rect 16615 4165 16635 4185
rect 16615 4115 16635 4135
rect 16615 4065 16635 4085
rect 16615 4015 16635 4035
rect 16615 3965 16635 3985
rect 16765 4415 16785 4435
rect 16765 4365 16785 4385
rect 16765 4315 16785 4335
rect 16765 4265 16785 4285
rect 16765 4215 16785 4235
rect 16765 4165 16785 4185
rect 16765 4115 16785 4135
rect 16765 4065 16785 4085
rect 16765 4015 16785 4035
rect 16765 3965 16785 3985
rect 16915 4415 16935 4435
rect 16915 4365 16935 4385
rect 16915 4315 16935 4335
rect 16915 4265 16935 4285
rect 16915 4215 16935 4235
rect 16915 4165 16935 4185
rect 16915 4115 16935 4135
rect 16915 4065 16935 4085
rect 16915 4015 16935 4035
rect 16915 3965 16935 3985
rect 17065 4415 17085 4435
rect 17065 4365 17085 4385
rect 17065 4315 17085 4335
rect 17065 4265 17085 4285
rect 17065 4215 17085 4235
rect 17065 4165 17085 4185
rect 17065 4115 17085 4135
rect 17065 4065 17085 4085
rect 17065 4015 17085 4035
rect 17065 3965 17085 3985
rect 17215 4415 17235 4435
rect 17215 4365 17235 4385
rect 17215 4315 17235 4335
rect 17215 4265 17235 4285
rect 17215 4215 17235 4235
rect 17215 4165 17235 4185
rect 17215 4115 17235 4135
rect 17215 4065 17235 4085
rect 17215 4015 17235 4035
rect 17215 3965 17235 3985
rect 17365 4415 17385 4435
rect 17365 4365 17385 4385
rect 17365 4315 17385 4335
rect 17365 4265 17385 4285
rect 17365 4215 17385 4235
rect 17365 4165 17385 4185
rect 17365 4115 17385 4135
rect 17365 4065 17385 4085
rect 17365 4015 17385 4035
rect 17365 3965 17385 3985
rect 17965 4415 17985 4435
rect 17965 4365 17985 4385
rect 17965 4315 17985 4335
rect 17965 4265 17985 4285
rect 17965 4215 17985 4235
rect 17965 4165 17985 4185
rect 17965 4115 17985 4135
rect 17965 4065 17985 4085
rect 17965 4015 17985 4035
rect 17965 3965 17985 3985
rect 18565 4415 18585 4435
rect 18565 4365 18585 4385
rect 18565 4315 18585 4335
rect 18565 4265 18585 4285
rect 18565 4215 18585 4235
rect 18565 4165 18585 4185
rect 18565 4115 18585 4135
rect 18565 4065 18585 4085
rect 18565 4015 18585 4035
rect 18565 3965 18585 3985
rect 18715 4415 18735 4435
rect 18715 4365 18735 4385
rect 18715 4315 18735 4335
rect 18715 4265 18735 4285
rect 18715 4215 18735 4235
rect 18715 4165 18735 4185
rect 18715 4115 18735 4135
rect 18715 4065 18735 4085
rect 18715 4015 18735 4035
rect 18715 3965 18735 3985
rect 18865 4415 18885 4435
rect 18865 4365 18885 4385
rect 18865 4315 18885 4335
rect 18865 4265 18885 4285
rect 18865 4215 18885 4235
rect 18865 4165 18885 4185
rect 18865 4115 18885 4135
rect 18865 4065 18885 4085
rect 18865 4015 18885 4035
rect 18865 3965 18885 3985
rect 19015 4415 19035 4435
rect 19015 4365 19035 4385
rect 19015 4315 19035 4335
rect 19015 4265 19035 4285
rect 19015 4215 19035 4235
rect 19015 4165 19035 4185
rect 19015 4115 19035 4135
rect 19015 4065 19035 4085
rect 19015 4015 19035 4035
rect 19015 3965 19035 3985
rect 19165 4415 19185 4435
rect 19165 4365 19185 4385
rect 19165 4315 19185 4335
rect 19165 4265 19185 4285
rect 19165 4215 19185 4235
rect 19165 4165 19185 4185
rect 19165 4115 19185 4135
rect 19165 4065 19185 4085
rect 19165 4015 19185 4035
rect 19165 3965 19185 3985
rect 19315 4415 19335 4435
rect 19315 4365 19335 4385
rect 19315 4315 19335 4335
rect 19315 4265 19335 4285
rect 19315 4215 19335 4235
rect 19315 4165 19335 4185
rect 19315 4115 19335 4135
rect 19315 4065 19335 4085
rect 19315 4015 19335 4035
rect 19315 3965 19335 3985
rect 19465 4415 19485 4435
rect 19465 4365 19485 4385
rect 19465 4315 19485 4335
rect 19465 4265 19485 4285
rect 19465 4215 19485 4235
rect 19465 4165 19485 4185
rect 19465 4115 19485 4135
rect 19465 4065 19485 4085
rect 19465 4015 19485 4035
rect 19465 3965 19485 3985
rect 19615 4415 19635 4435
rect 19615 4365 19635 4385
rect 19615 4315 19635 4335
rect 19615 4265 19635 4285
rect 19615 4215 19635 4235
rect 19615 4165 19635 4185
rect 19615 4115 19635 4135
rect 19615 4065 19635 4085
rect 19615 4015 19635 4035
rect 19615 3965 19635 3985
rect 19765 4415 19785 4435
rect 19765 4365 19785 4385
rect 19765 4315 19785 4335
rect 19765 4265 19785 4285
rect 19765 4215 19785 4235
rect 19765 4165 19785 4185
rect 19765 4115 19785 4135
rect 19765 4065 19785 4085
rect 19765 4015 19785 4035
rect 19765 3965 19785 3985
rect 20365 4415 20385 4435
rect 20365 4365 20385 4385
rect 20365 4315 20385 4335
rect 20365 4265 20385 4285
rect 20365 4215 20385 4235
rect 20365 4165 20385 4185
rect 20365 4115 20385 4135
rect 20365 4065 20385 4085
rect 20365 4015 20385 4035
rect 20365 3965 20385 3985
rect -635 3765 -615 3785
rect -635 3715 -615 3735
rect -635 3665 -615 3685
rect -635 3615 -615 3635
rect -635 3565 -615 3585
rect -635 3515 -615 3535
rect -635 3465 -615 3485
rect -635 3415 -615 3435
rect -635 3365 -615 3385
rect -635 3315 -615 3335
rect -485 3765 -465 3785
rect -485 3715 -465 3735
rect -485 3665 -465 3685
rect -485 3615 -465 3635
rect -485 3565 -465 3585
rect -485 3515 -465 3535
rect -485 3465 -465 3485
rect -485 3415 -465 3435
rect -485 3365 -465 3385
rect -485 3315 -465 3335
rect -335 3765 -315 3785
rect -335 3715 -315 3735
rect -335 3665 -315 3685
rect -335 3615 -315 3635
rect -335 3565 -315 3585
rect -335 3515 -315 3535
rect -335 3465 -315 3485
rect -335 3415 -315 3435
rect -335 3365 -315 3385
rect -335 3315 -315 3335
rect -185 3765 -165 3785
rect -185 3715 -165 3735
rect -185 3665 -165 3685
rect -185 3615 -165 3635
rect -185 3565 -165 3585
rect -185 3515 -165 3535
rect -185 3465 -165 3485
rect -185 3415 -165 3435
rect -185 3365 -165 3385
rect -185 3315 -165 3335
rect -35 3765 -15 3785
rect -35 3715 -15 3735
rect -35 3665 -15 3685
rect -35 3615 -15 3635
rect -35 3565 -15 3585
rect -35 3515 -15 3535
rect -35 3465 -15 3485
rect -35 3415 -15 3435
rect -35 3365 -15 3385
rect -35 3315 -15 3335
rect 565 3765 585 3785
rect 565 3715 585 3735
rect 565 3665 585 3685
rect 565 3615 585 3635
rect 565 3565 585 3585
rect 565 3515 585 3535
rect 565 3465 585 3485
rect 565 3415 585 3435
rect 565 3365 585 3385
rect 565 3315 585 3335
rect 715 3765 735 3785
rect 715 3715 735 3735
rect 715 3665 735 3685
rect 715 3615 735 3635
rect 715 3565 735 3585
rect 715 3515 735 3535
rect 715 3465 735 3485
rect 715 3415 735 3435
rect 715 3365 735 3385
rect 715 3315 735 3335
rect 865 3765 885 3785
rect 865 3715 885 3735
rect 865 3665 885 3685
rect 865 3615 885 3635
rect 865 3565 885 3585
rect 865 3515 885 3535
rect 865 3465 885 3485
rect 865 3415 885 3435
rect 865 3365 885 3385
rect 865 3315 885 3335
rect 1015 3765 1035 3785
rect 1015 3715 1035 3735
rect 1015 3665 1035 3685
rect 1015 3615 1035 3635
rect 1015 3565 1035 3585
rect 1015 3515 1035 3535
rect 1015 3465 1035 3485
rect 1015 3415 1035 3435
rect 1015 3365 1035 3385
rect 1015 3315 1035 3335
rect 1165 3765 1185 3785
rect 1165 3715 1185 3735
rect 1165 3665 1185 3685
rect 1165 3615 1185 3635
rect 1165 3565 1185 3585
rect 1165 3515 1185 3535
rect 1165 3465 1185 3485
rect 1165 3415 1185 3435
rect 1165 3365 1185 3385
rect 1165 3315 1185 3335
rect 1315 3765 1335 3785
rect 1315 3715 1335 3735
rect 1315 3665 1335 3685
rect 1315 3615 1335 3635
rect 1315 3565 1335 3585
rect 1315 3515 1335 3535
rect 1315 3465 1335 3485
rect 1315 3415 1335 3435
rect 1315 3365 1335 3385
rect 1315 3315 1335 3335
rect 1465 3765 1485 3785
rect 1465 3715 1485 3735
rect 1465 3665 1485 3685
rect 1465 3615 1485 3635
rect 1465 3565 1485 3585
rect 1465 3515 1485 3535
rect 1465 3465 1485 3485
rect 1465 3415 1485 3435
rect 1465 3365 1485 3385
rect 1465 3315 1485 3335
rect 1615 3765 1635 3785
rect 1615 3715 1635 3735
rect 1615 3665 1635 3685
rect 1615 3615 1635 3635
rect 1615 3565 1635 3585
rect 1615 3515 1635 3535
rect 1615 3465 1635 3485
rect 1615 3415 1635 3435
rect 1615 3365 1635 3385
rect 1615 3315 1635 3335
rect 1765 3765 1785 3785
rect 1765 3715 1785 3735
rect 1765 3665 1785 3685
rect 1765 3615 1785 3635
rect 1765 3565 1785 3585
rect 1765 3515 1785 3535
rect 1765 3465 1785 3485
rect 1765 3415 1785 3435
rect 1765 3365 1785 3385
rect 1765 3315 1785 3335
rect 1915 3765 1935 3785
rect 1915 3715 1935 3735
rect 1915 3665 1935 3685
rect 1915 3615 1935 3635
rect 1915 3565 1935 3585
rect 1915 3515 1935 3535
rect 1915 3465 1935 3485
rect 1915 3415 1935 3435
rect 1915 3365 1935 3385
rect 1915 3315 1935 3335
rect 2065 3765 2085 3785
rect 2065 3715 2085 3735
rect 2065 3665 2085 3685
rect 2065 3615 2085 3635
rect 2065 3565 2085 3585
rect 2065 3515 2085 3535
rect 2065 3465 2085 3485
rect 2065 3415 2085 3435
rect 2065 3365 2085 3385
rect 2065 3315 2085 3335
rect 2215 3765 2235 3785
rect 2215 3715 2235 3735
rect 2215 3665 2235 3685
rect 2215 3615 2235 3635
rect 2215 3565 2235 3585
rect 2215 3515 2235 3535
rect 2215 3465 2235 3485
rect 2215 3415 2235 3435
rect 2215 3365 2235 3385
rect 2215 3315 2235 3335
rect 2365 3765 2385 3785
rect 2365 3715 2385 3735
rect 2365 3665 2385 3685
rect 2365 3615 2385 3635
rect 2365 3565 2385 3585
rect 2365 3515 2385 3535
rect 2365 3465 2385 3485
rect 2365 3415 2385 3435
rect 2365 3365 2385 3385
rect 2365 3315 2385 3335
rect 2515 3765 2535 3785
rect 2515 3715 2535 3735
rect 2515 3665 2535 3685
rect 2515 3615 2535 3635
rect 2515 3565 2535 3585
rect 2515 3515 2535 3535
rect 2515 3465 2535 3485
rect 2515 3415 2535 3435
rect 2515 3365 2535 3385
rect 2515 3315 2535 3335
rect 2665 3765 2685 3785
rect 2665 3715 2685 3735
rect 2665 3665 2685 3685
rect 2665 3615 2685 3635
rect 2665 3565 2685 3585
rect 2665 3515 2685 3535
rect 2665 3465 2685 3485
rect 2665 3415 2685 3435
rect 2665 3365 2685 3385
rect 2665 3315 2685 3335
rect 2815 3765 2835 3785
rect 2815 3715 2835 3735
rect 2815 3665 2835 3685
rect 2815 3615 2835 3635
rect 2815 3565 2835 3585
rect 2815 3515 2835 3535
rect 2815 3465 2835 3485
rect 2815 3415 2835 3435
rect 2815 3365 2835 3385
rect 2815 3315 2835 3335
rect 2965 3765 2985 3785
rect 2965 3715 2985 3735
rect 2965 3665 2985 3685
rect 2965 3615 2985 3635
rect 2965 3565 2985 3585
rect 2965 3515 2985 3535
rect 2965 3465 2985 3485
rect 2965 3415 2985 3435
rect 2965 3365 2985 3385
rect 2965 3315 2985 3335
rect 3115 3765 3135 3785
rect 3115 3715 3135 3735
rect 3115 3665 3135 3685
rect 3115 3615 3135 3635
rect 3115 3565 3135 3585
rect 3115 3515 3135 3535
rect 3115 3465 3135 3485
rect 3115 3415 3135 3435
rect 3115 3365 3135 3385
rect 3115 3315 3135 3335
rect 3265 3765 3285 3785
rect 3265 3715 3285 3735
rect 3265 3665 3285 3685
rect 3265 3615 3285 3635
rect 3265 3565 3285 3585
rect 3265 3515 3285 3535
rect 3265 3465 3285 3485
rect 3265 3415 3285 3435
rect 3265 3365 3285 3385
rect 3265 3315 3285 3335
rect 3415 3765 3435 3785
rect 3415 3715 3435 3735
rect 3415 3665 3435 3685
rect 3415 3615 3435 3635
rect 3415 3565 3435 3585
rect 3415 3515 3435 3535
rect 3415 3465 3435 3485
rect 3415 3415 3435 3435
rect 3415 3365 3435 3385
rect 3415 3315 3435 3335
rect 3565 3765 3585 3785
rect 3565 3715 3585 3735
rect 3565 3665 3585 3685
rect 3565 3615 3585 3635
rect 3565 3565 3585 3585
rect 3565 3515 3585 3535
rect 3565 3465 3585 3485
rect 3565 3415 3585 3435
rect 3565 3365 3585 3385
rect 3565 3315 3585 3335
rect 4165 3765 4185 3785
rect 4165 3715 4185 3735
rect 4165 3665 4185 3685
rect 4165 3615 4185 3635
rect 4165 3565 4185 3585
rect 4165 3515 4185 3535
rect 4165 3465 4185 3485
rect 4165 3415 4185 3435
rect 4165 3365 4185 3385
rect 4165 3315 4185 3335
rect 4765 3765 4785 3785
rect 4765 3715 4785 3735
rect 4765 3665 4785 3685
rect 4765 3615 4785 3635
rect 4765 3565 4785 3585
rect 4765 3515 4785 3535
rect 4765 3465 4785 3485
rect 4765 3415 4785 3435
rect 4765 3365 4785 3385
rect 4765 3315 4785 3335
rect 4915 3765 4935 3785
rect 4915 3715 4935 3735
rect 4915 3665 4935 3685
rect 4915 3615 4935 3635
rect 4915 3565 4935 3585
rect 4915 3515 4935 3535
rect 4915 3465 4935 3485
rect 4915 3415 4935 3435
rect 4915 3365 4935 3385
rect 4915 3315 4935 3335
rect 5065 3765 5085 3785
rect 5065 3715 5085 3735
rect 5065 3665 5085 3685
rect 5065 3615 5085 3635
rect 5065 3565 5085 3585
rect 5065 3515 5085 3535
rect 5065 3465 5085 3485
rect 5065 3415 5085 3435
rect 5065 3365 5085 3385
rect 5065 3315 5085 3335
rect 5215 3765 5235 3785
rect 5215 3715 5235 3735
rect 5215 3665 5235 3685
rect 5215 3615 5235 3635
rect 5215 3565 5235 3585
rect 5215 3515 5235 3535
rect 5215 3465 5235 3485
rect 5215 3415 5235 3435
rect 5215 3365 5235 3385
rect 5215 3315 5235 3335
rect 5365 3765 5385 3785
rect 5365 3715 5385 3735
rect 5365 3665 5385 3685
rect 5365 3615 5385 3635
rect 5365 3565 5385 3585
rect 5365 3515 5385 3535
rect 5365 3465 5385 3485
rect 5365 3415 5385 3435
rect 5365 3365 5385 3385
rect 5365 3315 5385 3335
rect 5515 3765 5535 3785
rect 5515 3715 5535 3735
rect 5515 3665 5535 3685
rect 5515 3615 5535 3635
rect 5515 3565 5535 3585
rect 5515 3515 5535 3535
rect 5515 3465 5535 3485
rect 5515 3415 5535 3435
rect 5515 3365 5535 3385
rect 5515 3315 5535 3335
rect 5665 3765 5685 3785
rect 5665 3715 5685 3735
rect 5665 3665 5685 3685
rect 5665 3615 5685 3635
rect 5665 3565 5685 3585
rect 5665 3515 5685 3535
rect 5665 3465 5685 3485
rect 5665 3415 5685 3435
rect 5665 3365 5685 3385
rect 5665 3315 5685 3335
rect 5815 3765 5835 3785
rect 5815 3715 5835 3735
rect 5815 3665 5835 3685
rect 5815 3615 5835 3635
rect 5815 3565 5835 3585
rect 5815 3515 5835 3535
rect 5815 3465 5835 3485
rect 5815 3415 5835 3435
rect 5815 3365 5835 3385
rect 5815 3315 5835 3335
rect 5965 3765 5985 3785
rect 5965 3715 5985 3735
rect 5965 3665 5985 3685
rect 5965 3615 5985 3635
rect 5965 3565 5985 3585
rect 5965 3515 5985 3535
rect 5965 3465 5985 3485
rect 5965 3415 5985 3435
rect 5965 3365 5985 3385
rect 5965 3315 5985 3335
rect 6115 3765 6135 3785
rect 6115 3715 6135 3735
rect 6115 3665 6135 3685
rect 6115 3615 6135 3635
rect 6115 3565 6135 3585
rect 6115 3515 6135 3535
rect 6115 3465 6135 3485
rect 6115 3415 6135 3435
rect 6115 3365 6135 3385
rect 6115 3315 6135 3335
rect 6265 3765 6285 3785
rect 6265 3715 6285 3735
rect 6265 3665 6285 3685
rect 6265 3615 6285 3635
rect 6265 3565 6285 3585
rect 6265 3515 6285 3535
rect 6265 3465 6285 3485
rect 6265 3415 6285 3435
rect 6265 3365 6285 3385
rect 6265 3315 6285 3335
rect 6415 3765 6435 3785
rect 6415 3715 6435 3735
rect 6415 3665 6435 3685
rect 6415 3615 6435 3635
rect 6415 3565 6435 3585
rect 6415 3515 6435 3535
rect 6415 3465 6435 3485
rect 6415 3415 6435 3435
rect 6415 3365 6435 3385
rect 6415 3315 6435 3335
rect 6565 3765 6585 3785
rect 6565 3715 6585 3735
rect 6565 3665 6585 3685
rect 6565 3615 6585 3635
rect 6565 3565 6585 3585
rect 6565 3515 6585 3535
rect 6565 3465 6585 3485
rect 6565 3415 6585 3435
rect 6565 3365 6585 3385
rect 6565 3315 6585 3335
rect 6715 3765 6735 3785
rect 6715 3715 6735 3735
rect 6715 3665 6735 3685
rect 6715 3615 6735 3635
rect 6715 3565 6735 3585
rect 6715 3515 6735 3535
rect 6715 3465 6735 3485
rect 6715 3415 6735 3435
rect 6715 3365 6735 3385
rect 6715 3315 6735 3335
rect 6865 3765 6885 3785
rect 6865 3715 6885 3735
rect 6865 3665 6885 3685
rect 6865 3615 6885 3635
rect 6865 3565 6885 3585
rect 6865 3515 6885 3535
rect 6865 3465 6885 3485
rect 6865 3415 6885 3435
rect 6865 3365 6885 3385
rect 6865 3315 6885 3335
rect 7015 3765 7035 3785
rect 7015 3715 7035 3735
rect 7015 3665 7035 3685
rect 7015 3615 7035 3635
rect 7015 3565 7035 3585
rect 7015 3515 7035 3535
rect 7015 3465 7035 3485
rect 7015 3415 7035 3435
rect 7015 3365 7035 3385
rect 7015 3315 7035 3335
rect 7165 3765 7185 3785
rect 7165 3715 7185 3735
rect 7165 3665 7185 3685
rect 7165 3615 7185 3635
rect 7165 3565 7185 3585
rect 7165 3515 7185 3535
rect 7165 3465 7185 3485
rect 7165 3415 7185 3435
rect 7165 3365 7185 3385
rect 7165 3315 7185 3335
rect 7315 3765 7335 3785
rect 7315 3715 7335 3735
rect 7315 3665 7335 3685
rect 7315 3615 7335 3635
rect 7315 3565 7335 3585
rect 7315 3515 7335 3535
rect 7315 3465 7335 3485
rect 7315 3415 7335 3435
rect 7315 3365 7335 3385
rect 7315 3315 7335 3335
rect 7465 3765 7485 3785
rect 7465 3715 7485 3735
rect 7465 3665 7485 3685
rect 7465 3615 7485 3635
rect 7465 3565 7485 3585
rect 7465 3515 7485 3535
rect 7465 3465 7485 3485
rect 7465 3415 7485 3435
rect 7465 3365 7485 3385
rect 7465 3315 7485 3335
rect 7615 3765 7635 3785
rect 7615 3715 7635 3735
rect 7615 3665 7635 3685
rect 7615 3615 7635 3635
rect 7615 3565 7635 3585
rect 7615 3515 7635 3535
rect 7615 3465 7635 3485
rect 7615 3415 7635 3435
rect 7615 3365 7635 3385
rect 7615 3315 7635 3335
rect 7765 3765 7785 3785
rect 7765 3715 7785 3735
rect 7765 3665 7785 3685
rect 7765 3615 7785 3635
rect 7765 3565 7785 3585
rect 7765 3515 7785 3535
rect 7765 3465 7785 3485
rect 7765 3415 7785 3435
rect 7765 3365 7785 3385
rect 7765 3315 7785 3335
rect 8365 3765 8385 3785
rect 8365 3715 8385 3735
rect 8365 3665 8385 3685
rect 8365 3615 8385 3635
rect 8365 3565 8385 3585
rect 8365 3515 8385 3535
rect 8365 3465 8385 3485
rect 8365 3415 8385 3435
rect 8365 3365 8385 3385
rect 8365 3315 8385 3335
rect 8515 3765 8535 3785
rect 8515 3715 8535 3735
rect 8515 3665 8535 3685
rect 8515 3615 8535 3635
rect 8515 3565 8535 3585
rect 8515 3515 8535 3535
rect 8515 3465 8535 3485
rect 8515 3415 8535 3435
rect 8515 3365 8535 3385
rect 8515 3315 8535 3335
rect 8665 3765 8685 3785
rect 8665 3715 8685 3735
rect 8665 3665 8685 3685
rect 8665 3615 8685 3635
rect 8665 3565 8685 3585
rect 8665 3515 8685 3535
rect 8665 3465 8685 3485
rect 8665 3415 8685 3435
rect 8665 3365 8685 3385
rect 8665 3315 8685 3335
rect 8815 3765 8835 3785
rect 8815 3715 8835 3735
rect 8815 3665 8835 3685
rect 8815 3615 8835 3635
rect 8815 3565 8835 3585
rect 8815 3515 8835 3535
rect 8815 3465 8835 3485
rect 8815 3415 8835 3435
rect 8815 3365 8835 3385
rect 8815 3315 8835 3335
rect 8965 3765 8985 3785
rect 8965 3715 8985 3735
rect 8965 3665 8985 3685
rect 8965 3615 8985 3635
rect 8965 3565 8985 3585
rect 8965 3515 8985 3535
rect 8965 3465 8985 3485
rect 8965 3415 8985 3435
rect 8965 3365 8985 3385
rect 8965 3315 8985 3335
rect 9115 3765 9135 3785
rect 9115 3715 9135 3735
rect 9115 3665 9135 3685
rect 9115 3615 9135 3635
rect 9115 3565 9135 3585
rect 9115 3515 9135 3535
rect 9115 3465 9135 3485
rect 9115 3415 9135 3435
rect 9115 3365 9135 3385
rect 9115 3315 9135 3335
rect 9265 3765 9285 3785
rect 9265 3715 9285 3735
rect 9265 3665 9285 3685
rect 9265 3615 9285 3635
rect 9265 3565 9285 3585
rect 9265 3515 9285 3535
rect 9265 3465 9285 3485
rect 9265 3415 9285 3435
rect 9265 3365 9285 3385
rect 9265 3315 9285 3335
rect 9415 3765 9435 3785
rect 9415 3715 9435 3735
rect 9415 3665 9435 3685
rect 9415 3615 9435 3635
rect 9415 3565 9435 3585
rect 9415 3515 9435 3535
rect 9415 3465 9435 3485
rect 9415 3415 9435 3435
rect 9415 3365 9435 3385
rect 9415 3315 9435 3335
rect 9565 3765 9585 3785
rect 9565 3715 9585 3735
rect 9565 3665 9585 3685
rect 9565 3615 9585 3635
rect 9565 3565 9585 3585
rect 9565 3515 9585 3535
rect 9565 3465 9585 3485
rect 9565 3415 9585 3435
rect 9565 3365 9585 3385
rect 9565 3315 9585 3335
rect 9715 3765 9735 3785
rect 9715 3715 9735 3735
rect 9715 3665 9735 3685
rect 9715 3615 9735 3635
rect 9715 3565 9735 3585
rect 9715 3515 9735 3535
rect 9715 3465 9735 3485
rect 9715 3415 9735 3435
rect 9715 3365 9735 3385
rect 9715 3315 9735 3335
rect 9865 3765 9885 3785
rect 9865 3715 9885 3735
rect 9865 3665 9885 3685
rect 9865 3615 9885 3635
rect 9865 3565 9885 3585
rect 9865 3515 9885 3535
rect 9865 3465 9885 3485
rect 9865 3415 9885 3435
rect 9865 3365 9885 3385
rect 9865 3315 9885 3335
rect 10015 3765 10035 3785
rect 10015 3715 10035 3735
rect 10015 3665 10035 3685
rect 10015 3615 10035 3635
rect 10015 3565 10035 3585
rect 10015 3515 10035 3535
rect 10015 3465 10035 3485
rect 10015 3415 10035 3435
rect 10015 3365 10035 3385
rect 10015 3315 10035 3335
rect 10165 3765 10185 3785
rect 10165 3715 10185 3735
rect 10165 3665 10185 3685
rect 10165 3615 10185 3635
rect 10165 3565 10185 3585
rect 10165 3515 10185 3535
rect 10165 3465 10185 3485
rect 10165 3415 10185 3435
rect 10165 3365 10185 3385
rect 10165 3315 10185 3335
rect 10315 3765 10335 3785
rect 10315 3715 10335 3735
rect 10315 3665 10335 3685
rect 10315 3615 10335 3635
rect 10315 3565 10335 3585
rect 10315 3515 10335 3535
rect 10315 3465 10335 3485
rect 10315 3415 10335 3435
rect 10315 3365 10335 3385
rect 10315 3315 10335 3335
rect 10465 3765 10485 3785
rect 10465 3715 10485 3735
rect 10465 3665 10485 3685
rect 10465 3615 10485 3635
rect 10465 3565 10485 3585
rect 10465 3515 10485 3535
rect 10465 3465 10485 3485
rect 10465 3415 10485 3435
rect 10465 3365 10485 3385
rect 10465 3315 10485 3335
rect 10615 3765 10635 3785
rect 10615 3715 10635 3735
rect 10615 3665 10635 3685
rect 10615 3615 10635 3635
rect 10615 3565 10635 3585
rect 10615 3515 10635 3535
rect 10615 3465 10635 3485
rect 10615 3415 10635 3435
rect 10615 3365 10635 3385
rect 10615 3315 10635 3335
rect 10765 3765 10785 3785
rect 10765 3715 10785 3735
rect 10765 3665 10785 3685
rect 10765 3615 10785 3635
rect 10765 3565 10785 3585
rect 10765 3515 10785 3535
rect 10765 3465 10785 3485
rect 10765 3415 10785 3435
rect 10765 3365 10785 3385
rect 10765 3315 10785 3335
rect 11365 3765 11385 3785
rect 11365 3715 11385 3735
rect 11365 3665 11385 3685
rect 11365 3615 11385 3635
rect 11365 3565 11385 3585
rect 11365 3515 11385 3535
rect 11365 3465 11385 3485
rect 11365 3415 11385 3435
rect 11365 3365 11385 3385
rect 11365 3315 11385 3335
rect 11965 3765 11985 3785
rect 11965 3715 11985 3735
rect 11965 3665 11985 3685
rect 11965 3615 11985 3635
rect 11965 3565 11985 3585
rect 11965 3515 11985 3535
rect 11965 3465 11985 3485
rect 11965 3415 11985 3435
rect 11965 3365 11985 3385
rect 11965 3315 11985 3335
rect 12565 3765 12585 3785
rect 12565 3715 12585 3735
rect 12565 3665 12585 3685
rect 12565 3615 12585 3635
rect 12565 3565 12585 3585
rect 12565 3515 12585 3535
rect 12565 3465 12585 3485
rect 12565 3415 12585 3435
rect 12565 3365 12585 3385
rect 12565 3315 12585 3335
rect 13165 3765 13185 3785
rect 13165 3715 13185 3735
rect 13165 3665 13185 3685
rect 13165 3615 13185 3635
rect 13165 3565 13185 3585
rect 13165 3515 13185 3535
rect 13165 3465 13185 3485
rect 13165 3415 13185 3435
rect 13165 3365 13185 3385
rect 13165 3315 13185 3335
rect 13765 3765 13785 3785
rect 13765 3715 13785 3735
rect 13765 3665 13785 3685
rect 13765 3615 13785 3635
rect 13765 3565 13785 3585
rect 13765 3515 13785 3535
rect 13765 3465 13785 3485
rect 13765 3415 13785 3435
rect 13765 3365 13785 3385
rect 13765 3315 13785 3335
rect 14365 3765 14385 3785
rect 14365 3715 14385 3735
rect 14365 3665 14385 3685
rect 14365 3615 14385 3635
rect 14365 3565 14385 3585
rect 14365 3515 14385 3535
rect 14365 3465 14385 3485
rect 14365 3415 14385 3435
rect 14365 3365 14385 3385
rect 14365 3315 14385 3335
rect 14965 3765 14985 3785
rect 14965 3715 14985 3735
rect 14965 3665 14985 3685
rect 14965 3615 14985 3635
rect 14965 3565 14985 3585
rect 14965 3515 14985 3535
rect 14965 3465 14985 3485
rect 14965 3415 14985 3435
rect 14965 3365 14985 3385
rect 14965 3315 14985 3335
rect 15565 3765 15585 3785
rect 15565 3715 15585 3735
rect 15565 3665 15585 3685
rect 15565 3615 15585 3635
rect 15565 3565 15585 3585
rect 15565 3515 15585 3535
rect 15565 3465 15585 3485
rect 15565 3415 15585 3435
rect 15565 3365 15585 3385
rect 15565 3315 15585 3335
rect 16165 3765 16185 3785
rect 16165 3715 16185 3735
rect 16165 3665 16185 3685
rect 16165 3615 16185 3635
rect 16165 3565 16185 3585
rect 16165 3515 16185 3535
rect 16165 3465 16185 3485
rect 16165 3415 16185 3435
rect 16165 3365 16185 3385
rect 16165 3315 16185 3335
rect 16315 3765 16335 3785
rect 16315 3715 16335 3735
rect 16315 3665 16335 3685
rect 16315 3615 16335 3635
rect 16315 3565 16335 3585
rect 16315 3515 16335 3535
rect 16315 3465 16335 3485
rect 16315 3415 16335 3435
rect 16315 3365 16335 3385
rect 16315 3315 16335 3335
rect 16465 3765 16485 3785
rect 16465 3715 16485 3735
rect 16465 3665 16485 3685
rect 16465 3615 16485 3635
rect 16465 3565 16485 3585
rect 16465 3515 16485 3535
rect 16465 3465 16485 3485
rect 16465 3415 16485 3435
rect 16465 3365 16485 3385
rect 16465 3315 16485 3335
rect 16615 3765 16635 3785
rect 16615 3715 16635 3735
rect 16615 3665 16635 3685
rect 16615 3615 16635 3635
rect 16615 3565 16635 3585
rect 16615 3515 16635 3535
rect 16615 3465 16635 3485
rect 16615 3415 16635 3435
rect 16615 3365 16635 3385
rect 16615 3315 16635 3335
rect 16765 3765 16785 3785
rect 16765 3715 16785 3735
rect 16765 3665 16785 3685
rect 16765 3615 16785 3635
rect 16765 3565 16785 3585
rect 16765 3515 16785 3535
rect 16765 3465 16785 3485
rect 16765 3415 16785 3435
rect 16765 3365 16785 3385
rect 16765 3315 16785 3335
rect 16915 3765 16935 3785
rect 16915 3715 16935 3735
rect 16915 3665 16935 3685
rect 16915 3615 16935 3635
rect 16915 3565 16935 3585
rect 16915 3515 16935 3535
rect 16915 3465 16935 3485
rect 16915 3415 16935 3435
rect 16915 3365 16935 3385
rect 16915 3315 16935 3335
rect 17065 3765 17085 3785
rect 17065 3715 17085 3735
rect 17065 3665 17085 3685
rect 17065 3615 17085 3635
rect 17065 3565 17085 3585
rect 17065 3515 17085 3535
rect 17065 3465 17085 3485
rect 17065 3415 17085 3435
rect 17065 3365 17085 3385
rect 17065 3315 17085 3335
rect 17215 3765 17235 3785
rect 17215 3715 17235 3735
rect 17215 3665 17235 3685
rect 17215 3615 17235 3635
rect 17215 3565 17235 3585
rect 17215 3515 17235 3535
rect 17215 3465 17235 3485
rect 17215 3415 17235 3435
rect 17215 3365 17235 3385
rect 17215 3315 17235 3335
rect 17365 3765 17385 3785
rect 17365 3715 17385 3735
rect 17365 3665 17385 3685
rect 17365 3615 17385 3635
rect 17365 3565 17385 3585
rect 17365 3515 17385 3535
rect 17365 3465 17385 3485
rect 17365 3415 17385 3435
rect 17365 3365 17385 3385
rect 17365 3315 17385 3335
rect 17965 3765 17985 3785
rect 17965 3715 17985 3735
rect 17965 3665 17985 3685
rect 17965 3615 17985 3635
rect 17965 3565 17985 3585
rect 17965 3515 17985 3535
rect 17965 3465 17985 3485
rect 17965 3415 17985 3435
rect 17965 3365 17985 3385
rect 17965 3315 17985 3335
rect 18565 3765 18585 3785
rect 18565 3715 18585 3735
rect 18565 3665 18585 3685
rect 18565 3615 18585 3635
rect 18565 3565 18585 3585
rect 18565 3515 18585 3535
rect 18565 3465 18585 3485
rect 18565 3415 18585 3435
rect 18565 3365 18585 3385
rect 18565 3315 18585 3335
rect 18715 3765 18735 3785
rect 18715 3715 18735 3735
rect 18715 3665 18735 3685
rect 18715 3615 18735 3635
rect 18715 3565 18735 3585
rect 18715 3515 18735 3535
rect 18715 3465 18735 3485
rect 18715 3415 18735 3435
rect 18715 3365 18735 3385
rect 18715 3315 18735 3335
rect 18865 3765 18885 3785
rect 18865 3715 18885 3735
rect 18865 3665 18885 3685
rect 18865 3615 18885 3635
rect 18865 3565 18885 3585
rect 18865 3515 18885 3535
rect 18865 3465 18885 3485
rect 18865 3415 18885 3435
rect 18865 3365 18885 3385
rect 18865 3315 18885 3335
rect 19015 3765 19035 3785
rect 19015 3715 19035 3735
rect 19015 3665 19035 3685
rect 19015 3615 19035 3635
rect 19015 3565 19035 3585
rect 19015 3515 19035 3535
rect 19015 3465 19035 3485
rect 19015 3415 19035 3435
rect 19015 3365 19035 3385
rect 19015 3315 19035 3335
rect 19165 3765 19185 3785
rect 19165 3715 19185 3735
rect 19165 3665 19185 3685
rect 19165 3615 19185 3635
rect 19165 3565 19185 3585
rect 19165 3515 19185 3535
rect 19165 3465 19185 3485
rect 19165 3415 19185 3435
rect 19165 3365 19185 3385
rect 19165 3315 19185 3335
rect 19315 3765 19335 3785
rect 19315 3715 19335 3735
rect 19315 3665 19335 3685
rect 19315 3615 19335 3635
rect 19315 3565 19335 3585
rect 19315 3515 19335 3535
rect 19315 3465 19335 3485
rect 19315 3415 19335 3435
rect 19315 3365 19335 3385
rect 19315 3315 19335 3335
rect 19465 3765 19485 3785
rect 19465 3715 19485 3735
rect 19465 3665 19485 3685
rect 19465 3615 19485 3635
rect 19465 3565 19485 3585
rect 19465 3515 19485 3535
rect 19465 3465 19485 3485
rect 19465 3415 19485 3435
rect 19465 3365 19485 3385
rect 19465 3315 19485 3335
rect 19615 3765 19635 3785
rect 19615 3715 19635 3735
rect 19615 3665 19635 3685
rect 19615 3615 19635 3635
rect 19615 3565 19635 3585
rect 19615 3515 19635 3535
rect 19615 3465 19635 3485
rect 19615 3415 19635 3435
rect 19615 3365 19635 3385
rect 19615 3315 19635 3335
rect 19765 3765 19785 3785
rect 19765 3715 19785 3735
rect 19765 3665 19785 3685
rect 19765 3615 19785 3635
rect 19765 3565 19785 3585
rect 19765 3515 19785 3535
rect 19765 3465 19785 3485
rect 19765 3415 19785 3435
rect 19765 3365 19785 3385
rect 19765 3315 19785 3335
rect 20365 3765 20385 3785
rect 20365 3715 20385 3735
rect 20365 3665 20385 3685
rect 20365 3615 20385 3635
rect 20365 3565 20385 3585
rect 20365 3515 20385 3535
rect 20365 3465 20385 3485
rect 20365 3415 20385 3435
rect 20365 3365 20385 3385
rect 20365 3315 20385 3335
rect -635 3115 -615 3135
rect -635 3065 -615 3085
rect -635 3015 -615 3035
rect -635 2965 -615 2985
rect -635 2915 -615 2935
rect -635 2865 -615 2885
rect -635 2815 -615 2835
rect -635 2765 -615 2785
rect -635 2715 -615 2735
rect -635 2665 -615 2685
rect -485 3115 -465 3135
rect -485 3065 -465 3085
rect -485 3015 -465 3035
rect -485 2965 -465 2985
rect -485 2915 -465 2935
rect -485 2865 -465 2885
rect -485 2815 -465 2835
rect -485 2765 -465 2785
rect -485 2715 -465 2735
rect -485 2665 -465 2685
rect -335 3115 -315 3135
rect -335 3065 -315 3085
rect -335 3015 -315 3035
rect -335 2965 -315 2985
rect -335 2915 -315 2935
rect -335 2865 -315 2885
rect -335 2815 -315 2835
rect -335 2765 -315 2785
rect -335 2715 -315 2735
rect -335 2665 -315 2685
rect -185 3115 -165 3135
rect -185 3065 -165 3085
rect -185 3015 -165 3035
rect -185 2965 -165 2985
rect -185 2915 -165 2935
rect -185 2865 -165 2885
rect -185 2815 -165 2835
rect -185 2765 -165 2785
rect -185 2715 -165 2735
rect -185 2665 -165 2685
rect -35 3115 -15 3135
rect -35 3065 -15 3085
rect -35 3015 -15 3035
rect -35 2965 -15 2985
rect -35 2915 -15 2935
rect -35 2865 -15 2885
rect -35 2815 -15 2835
rect -35 2765 -15 2785
rect -35 2715 -15 2735
rect -35 2665 -15 2685
rect 565 3115 585 3135
rect 565 3065 585 3085
rect 565 3015 585 3035
rect 565 2965 585 2985
rect 565 2915 585 2935
rect 565 2865 585 2885
rect 565 2815 585 2835
rect 565 2765 585 2785
rect 565 2715 585 2735
rect 565 2665 585 2685
rect 715 3115 735 3135
rect 715 3065 735 3085
rect 715 3015 735 3035
rect 715 2965 735 2985
rect 715 2915 735 2935
rect 715 2865 735 2885
rect 715 2815 735 2835
rect 715 2765 735 2785
rect 715 2715 735 2735
rect 715 2665 735 2685
rect 865 3115 885 3135
rect 865 3065 885 3085
rect 865 3015 885 3035
rect 865 2965 885 2985
rect 865 2915 885 2935
rect 865 2865 885 2885
rect 865 2815 885 2835
rect 865 2765 885 2785
rect 865 2715 885 2735
rect 865 2665 885 2685
rect 1015 3115 1035 3135
rect 1015 3065 1035 3085
rect 1015 3015 1035 3035
rect 1015 2965 1035 2985
rect 1015 2915 1035 2935
rect 1015 2865 1035 2885
rect 1015 2815 1035 2835
rect 1015 2765 1035 2785
rect 1015 2715 1035 2735
rect 1015 2665 1035 2685
rect 1165 3115 1185 3135
rect 1165 3065 1185 3085
rect 1165 3015 1185 3035
rect 1165 2965 1185 2985
rect 1165 2915 1185 2935
rect 1165 2865 1185 2885
rect 1165 2815 1185 2835
rect 1165 2765 1185 2785
rect 1165 2715 1185 2735
rect 1165 2665 1185 2685
rect 1315 3115 1335 3135
rect 1315 3065 1335 3085
rect 1315 3015 1335 3035
rect 1315 2965 1335 2985
rect 1315 2915 1335 2935
rect 1315 2865 1335 2885
rect 1315 2815 1335 2835
rect 1315 2765 1335 2785
rect 1315 2715 1335 2735
rect 1315 2665 1335 2685
rect 1465 3115 1485 3135
rect 1465 3065 1485 3085
rect 1465 3015 1485 3035
rect 1465 2965 1485 2985
rect 1465 2915 1485 2935
rect 1465 2865 1485 2885
rect 1465 2815 1485 2835
rect 1465 2765 1485 2785
rect 1465 2715 1485 2735
rect 1465 2665 1485 2685
rect 1615 3115 1635 3135
rect 1615 3065 1635 3085
rect 1615 3015 1635 3035
rect 1615 2965 1635 2985
rect 1615 2915 1635 2935
rect 1615 2865 1635 2885
rect 1615 2815 1635 2835
rect 1615 2765 1635 2785
rect 1615 2715 1635 2735
rect 1615 2665 1635 2685
rect 1765 3115 1785 3135
rect 1765 3065 1785 3085
rect 1765 3015 1785 3035
rect 1765 2965 1785 2985
rect 1765 2915 1785 2935
rect 1765 2865 1785 2885
rect 1765 2815 1785 2835
rect 1765 2765 1785 2785
rect 1765 2715 1785 2735
rect 1765 2665 1785 2685
rect 1915 3115 1935 3135
rect 1915 3065 1935 3085
rect 1915 3015 1935 3035
rect 1915 2965 1935 2985
rect 1915 2915 1935 2935
rect 1915 2865 1935 2885
rect 1915 2815 1935 2835
rect 1915 2765 1935 2785
rect 1915 2715 1935 2735
rect 1915 2665 1935 2685
rect 2065 3115 2085 3135
rect 2065 3065 2085 3085
rect 2065 3015 2085 3035
rect 2065 2965 2085 2985
rect 2065 2915 2085 2935
rect 2065 2865 2085 2885
rect 2065 2815 2085 2835
rect 2065 2765 2085 2785
rect 2065 2715 2085 2735
rect 2065 2665 2085 2685
rect 2215 3115 2235 3135
rect 2215 3065 2235 3085
rect 2215 3015 2235 3035
rect 2215 2965 2235 2985
rect 2215 2915 2235 2935
rect 2215 2865 2235 2885
rect 2215 2815 2235 2835
rect 2215 2765 2235 2785
rect 2215 2715 2235 2735
rect 2215 2665 2235 2685
rect 2365 3115 2385 3135
rect 2365 3065 2385 3085
rect 2365 3015 2385 3035
rect 2365 2965 2385 2985
rect 2365 2915 2385 2935
rect 2365 2865 2385 2885
rect 2365 2815 2385 2835
rect 2365 2765 2385 2785
rect 2365 2715 2385 2735
rect 2365 2665 2385 2685
rect 2515 3115 2535 3135
rect 2515 3065 2535 3085
rect 2515 3015 2535 3035
rect 2515 2965 2535 2985
rect 2515 2915 2535 2935
rect 2515 2865 2535 2885
rect 2515 2815 2535 2835
rect 2515 2765 2535 2785
rect 2515 2715 2535 2735
rect 2515 2665 2535 2685
rect 2665 3115 2685 3135
rect 2665 3065 2685 3085
rect 2665 3015 2685 3035
rect 2665 2965 2685 2985
rect 2665 2915 2685 2935
rect 2665 2865 2685 2885
rect 2665 2815 2685 2835
rect 2665 2765 2685 2785
rect 2665 2715 2685 2735
rect 2665 2665 2685 2685
rect 2815 3115 2835 3135
rect 2815 3065 2835 3085
rect 2815 3015 2835 3035
rect 2815 2965 2835 2985
rect 2815 2915 2835 2935
rect 2815 2865 2835 2885
rect 2815 2815 2835 2835
rect 2815 2765 2835 2785
rect 2815 2715 2835 2735
rect 2815 2665 2835 2685
rect 2965 3115 2985 3135
rect 2965 3065 2985 3085
rect 2965 3015 2985 3035
rect 2965 2965 2985 2985
rect 2965 2915 2985 2935
rect 2965 2865 2985 2885
rect 2965 2815 2985 2835
rect 2965 2765 2985 2785
rect 2965 2715 2985 2735
rect 2965 2665 2985 2685
rect 3115 3115 3135 3135
rect 3115 3065 3135 3085
rect 3115 3015 3135 3035
rect 3115 2965 3135 2985
rect 3115 2915 3135 2935
rect 3115 2865 3135 2885
rect 3115 2815 3135 2835
rect 3115 2765 3135 2785
rect 3115 2715 3135 2735
rect 3115 2665 3135 2685
rect 3265 3115 3285 3135
rect 3265 3065 3285 3085
rect 3265 3015 3285 3035
rect 3265 2965 3285 2985
rect 3265 2915 3285 2935
rect 3265 2865 3285 2885
rect 3265 2815 3285 2835
rect 3265 2765 3285 2785
rect 3265 2715 3285 2735
rect 3265 2665 3285 2685
rect 3415 3115 3435 3135
rect 3415 3065 3435 3085
rect 3415 3015 3435 3035
rect 3415 2965 3435 2985
rect 3415 2915 3435 2935
rect 3415 2865 3435 2885
rect 3415 2815 3435 2835
rect 3415 2765 3435 2785
rect 3415 2715 3435 2735
rect 3415 2665 3435 2685
rect 3565 3115 3585 3135
rect 3565 3065 3585 3085
rect 3565 3015 3585 3035
rect 3565 2965 3585 2985
rect 3565 2915 3585 2935
rect 3565 2865 3585 2885
rect 3565 2815 3585 2835
rect 3565 2765 3585 2785
rect 3565 2715 3585 2735
rect 3565 2665 3585 2685
rect 4165 3115 4185 3135
rect 4165 3065 4185 3085
rect 4165 3015 4185 3035
rect 4165 2965 4185 2985
rect 4165 2915 4185 2935
rect 4165 2865 4185 2885
rect 4165 2815 4185 2835
rect 4165 2765 4185 2785
rect 4165 2715 4185 2735
rect 4165 2665 4185 2685
rect 4765 3115 4785 3135
rect 4765 3065 4785 3085
rect 4765 3015 4785 3035
rect 4765 2965 4785 2985
rect 4765 2915 4785 2935
rect 4765 2865 4785 2885
rect 4765 2815 4785 2835
rect 4765 2765 4785 2785
rect 4765 2715 4785 2735
rect 4765 2665 4785 2685
rect 4915 3115 4935 3135
rect 4915 3065 4935 3085
rect 4915 3015 4935 3035
rect 4915 2965 4935 2985
rect 4915 2915 4935 2935
rect 4915 2865 4935 2885
rect 4915 2815 4935 2835
rect 4915 2765 4935 2785
rect 4915 2715 4935 2735
rect 4915 2665 4935 2685
rect 5065 3115 5085 3135
rect 5065 3065 5085 3085
rect 5065 3015 5085 3035
rect 5065 2965 5085 2985
rect 5065 2915 5085 2935
rect 5065 2865 5085 2885
rect 5065 2815 5085 2835
rect 5065 2765 5085 2785
rect 5065 2715 5085 2735
rect 5065 2665 5085 2685
rect 5215 3115 5235 3135
rect 5215 3065 5235 3085
rect 5215 3015 5235 3035
rect 5215 2965 5235 2985
rect 5215 2915 5235 2935
rect 5215 2865 5235 2885
rect 5215 2815 5235 2835
rect 5215 2765 5235 2785
rect 5215 2715 5235 2735
rect 5215 2665 5235 2685
rect 5365 3115 5385 3135
rect 5365 3065 5385 3085
rect 5365 3015 5385 3035
rect 5365 2965 5385 2985
rect 5365 2915 5385 2935
rect 5365 2865 5385 2885
rect 5365 2815 5385 2835
rect 5365 2765 5385 2785
rect 5365 2715 5385 2735
rect 5365 2665 5385 2685
rect 5515 3115 5535 3135
rect 5515 3065 5535 3085
rect 5515 3015 5535 3035
rect 5515 2965 5535 2985
rect 5515 2915 5535 2935
rect 5515 2865 5535 2885
rect 5515 2815 5535 2835
rect 5515 2765 5535 2785
rect 5515 2715 5535 2735
rect 5515 2665 5535 2685
rect 5665 3115 5685 3135
rect 5665 3065 5685 3085
rect 5665 3015 5685 3035
rect 5665 2965 5685 2985
rect 5665 2915 5685 2935
rect 5665 2865 5685 2885
rect 5665 2815 5685 2835
rect 5665 2765 5685 2785
rect 5665 2715 5685 2735
rect 5665 2665 5685 2685
rect 5815 3115 5835 3135
rect 5815 3065 5835 3085
rect 5815 3015 5835 3035
rect 5815 2965 5835 2985
rect 5815 2915 5835 2935
rect 5815 2865 5835 2885
rect 5815 2815 5835 2835
rect 5815 2765 5835 2785
rect 5815 2715 5835 2735
rect 5815 2665 5835 2685
rect 5965 3115 5985 3135
rect 5965 3065 5985 3085
rect 5965 3015 5985 3035
rect 5965 2965 5985 2985
rect 5965 2915 5985 2935
rect 5965 2865 5985 2885
rect 5965 2815 5985 2835
rect 5965 2765 5985 2785
rect 5965 2715 5985 2735
rect 5965 2665 5985 2685
rect 6115 3115 6135 3135
rect 6115 3065 6135 3085
rect 6115 3015 6135 3035
rect 6115 2965 6135 2985
rect 6115 2915 6135 2935
rect 6115 2865 6135 2885
rect 6115 2815 6135 2835
rect 6115 2765 6135 2785
rect 6115 2715 6135 2735
rect 6115 2665 6135 2685
rect 6265 3115 6285 3135
rect 6265 3065 6285 3085
rect 6265 3015 6285 3035
rect 6265 2965 6285 2985
rect 6265 2915 6285 2935
rect 6265 2865 6285 2885
rect 6265 2815 6285 2835
rect 6265 2765 6285 2785
rect 6265 2715 6285 2735
rect 6265 2665 6285 2685
rect 6415 3115 6435 3135
rect 6415 3065 6435 3085
rect 6415 3015 6435 3035
rect 6415 2965 6435 2985
rect 6415 2915 6435 2935
rect 6415 2865 6435 2885
rect 6415 2815 6435 2835
rect 6415 2765 6435 2785
rect 6415 2715 6435 2735
rect 6415 2665 6435 2685
rect 6565 3115 6585 3135
rect 6565 3065 6585 3085
rect 6565 3015 6585 3035
rect 6565 2965 6585 2985
rect 6565 2915 6585 2935
rect 6565 2865 6585 2885
rect 6565 2815 6585 2835
rect 6565 2765 6585 2785
rect 6565 2715 6585 2735
rect 6565 2665 6585 2685
rect 6715 3115 6735 3135
rect 6715 3065 6735 3085
rect 6715 3015 6735 3035
rect 6715 2965 6735 2985
rect 6715 2915 6735 2935
rect 6715 2865 6735 2885
rect 6715 2815 6735 2835
rect 6715 2765 6735 2785
rect 6715 2715 6735 2735
rect 6715 2665 6735 2685
rect 6865 3115 6885 3135
rect 6865 3065 6885 3085
rect 6865 3015 6885 3035
rect 6865 2965 6885 2985
rect 6865 2915 6885 2935
rect 6865 2865 6885 2885
rect 6865 2815 6885 2835
rect 6865 2765 6885 2785
rect 6865 2715 6885 2735
rect 6865 2665 6885 2685
rect 7015 3115 7035 3135
rect 7015 3065 7035 3085
rect 7015 3015 7035 3035
rect 7015 2965 7035 2985
rect 7015 2915 7035 2935
rect 7015 2865 7035 2885
rect 7015 2815 7035 2835
rect 7015 2765 7035 2785
rect 7015 2715 7035 2735
rect 7015 2665 7035 2685
rect 7165 3115 7185 3135
rect 7165 3065 7185 3085
rect 7165 3015 7185 3035
rect 7165 2965 7185 2985
rect 7165 2915 7185 2935
rect 7165 2865 7185 2885
rect 7165 2815 7185 2835
rect 7165 2765 7185 2785
rect 7165 2715 7185 2735
rect 7165 2665 7185 2685
rect 7315 3115 7335 3135
rect 7315 3065 7335 3085
rect 7315 3015 7335 3035
rect 7315 2965 7335 2985
rect 7315 2915 7335 2935
rect 7315 2865 7335 2885
rect 7315 2815 7335 2835
rect 7315 2765 7335 2785
rect 7315 2715 7335 2735
rect 7315 2665 7335 2685
rect 7465 3115 7485 3135
rect 7465 3065 7485 3085
rect 7465 3015 7485 3035
rect 7465 2965 7485 2985
rect 7465 2915 7485 2935
rect 7465 2865 7485 2885
rect 7465 2815 7485 2835
rect 7465 2765 7485 2785
rect 7465 2715 7485 2735
rect 7465 2665 7485 2685
rect 7615 3115 7635 3135
rect 7615 3065 7635 3085
rect 7615 3015 7635 3035
rect 7615 2965 7635 2985
rect 7615 2915 7635 2935
rect 7615 2865 7635 2885
rect 7615 2815 7635 2835
rect 7615 2765 7635 2785
rect 7615 2715 7635 2735
rect 7615 2665 7635 2685
rect 7765 3115 7785 3135
rect 7765 3065 7785 3085
rect 7765 3015 7785 3035
rect 7765 2965 7785 2985
rect 7765 2915 7785 2935
rect 7765 2865 7785 2885
rect 7765 2815 7785 2835
rect 7765 2765 7785 2785
rect 7765 2715 7785 2735
rect 7765 2665 7785 2685
rect 8365 3115 8385 3135
rect 8365 3065 8385 3085
rect 8365 3015 8385 3035
rect 8365 2965 8385 2985
rect 8365 2915 8385 2935
rect 8365 2865 8385 2885
rect 8365 2815 8385 2835
rect 8365 2765 8385 2785
rect 8365 2715 8385 2735
rect 8365 2665 8385 2685
rect 8515 3115 8535 3135
rect 8515 3065 8535 3085
rect 8515 3015 8535 3035
rect 8515 2965 8535 2985
rect 8515 2915 8535 2935
rect 8515 2865 8535 2885
rect 8515 2815 8535 2835
rect 8515 2765 8535 2785
rect 8515 2715 8535 2735
rect 8515 2665 8535 2685
rect 8665 3115 8685 3135
rect 8665 3065 8685 3085
rect 8665 3015 8685 3035
rect 8665 2965 8685 2985
rect 8665 2915 8685 2935
rect 8665 2865 8685 2885
rect 8665 2815 8685 2835
rect 8665 2765 8685 2785
rect 8665 2715 8685 2735
rect 8665 2665 8685 2685
rect 8815 3115 8835 3135
rect 8815 3065 8835 3085
rect 8815 3015 8835 3035
rect 8815 2965 8835 2985
rect 8815 2915 8835 2935
rect 8815 2865 8835 2885
rect 8815 2815 8835 2835
rect 8815 2765 8835 2785
rect 8815 2715 8835 2735
rect 8815 2665 8835 2685
rect 8965 3115 8985 3135
rect 8965 3065 8985 3085
rect 8965 3015 8985 3035
rect 8965 2965 8985 2985
rect 8965 2915 8985 2935
rect 8965 2865 8985 2885
rect 8965 2815 8985 2835
rect 8965 2765 8985 2785
rect 8965 2715 8985 2735
rect 8965 2665 8985 2685
rect 9115 3115 9135 3135
rect 9115 3065 9135 3085
rect 9115 3015 9135 3035
rect 9115 2965 9135 2985
rect 9115 2915 9135 2935
rect 9115 2865 9135 2885
rect 9115 2815 9135 2835
rect 9115 2765 9135 2785
rect 9115 2715 9135 2735
rect 9115 2665 9135 2685
rect 9265 3115 9285 3135
rect 9265 3065 9285 3085
rect 9265 3015 9285 3035
rect 9265 2965 9285 2985
rect 9265 2915 9285 2935
rect 9265 2865 9285 2885
rect 9265 2815 9285 2835
rect 9265 2765 9285 2785
rect 9265 2715 9285 2735
rect 9265 2665 9285 2685
rect 9415 3115 9435 3135
rect 9415 3065 9435 3085
rect 9415 3015 9435 3035
rect 9415 2965 9435 2985
rect 9415 2915 9435 2935
rect 9415 2865 9435 2885
rect 9415 2815 9435 2835
rect 9415 2765 9435 2785
rect 9415 2715 9435 2735
rect 9415 2665 9435 2685
rect 9565 3115 9585 3135
rect 9565 3065 9585 3085
rect 9565 3015 9585 3035
rect 9565 2965 9585 2985
rect 9565 2915 9585 2935
rect 9565 2865 9585 2885
rect 9565 2815 9585 2835
rect 9565 2765 9585 2785
rect 9565 2715 9585 2735
rect 9565 2665 9585 2685
rect 9715 3115 9735 3135
rect 9715 3065 9735 3085
rect 9715 3015 9735 3035
rect 9715 2965 9735 2985
rect 9715 2915 9735 2935
rect 9715 2865 9735 2885
rect 9715 2815 9735 2835
rect 9715 2765 9735 2785
rect 9715 2715 9735 2735
rect 9715 2665 9735 2685
rect 9865 3115 9885 3135
rect 9865 3065 9885 3085
rect 9865 3015 9885 3035
rect 9865 2965 9885 2985
rect 9865 2915 9885 2935
rect 9865 2865 9885 2885
rect 9865 2815 9885 2835
rect 9865 2765 9885 2785
rect 9865 2715 9885 2735
rect 9865 2665 9885 2685
rect 10015 3115 10035 3135
rect 10015 3065 10035 3085
rect 10015 3015 10035 3035
rect 10015 2965 10035 2985
rect 10015 2915 10035 2935
rect 10015 2865 10035 2885
rect 10015 2815 10035 2835
rect 10015 2765 10035 2785
rect 10015 2715 10035 2735
rect 10015 2665 10035 2685
rect 10165 3115 10185 3135
rect 10165 3065 10185 3085
rect 10165 3015 10185 3035
rect 10165 2965 10185 2985
rect 10165 2915 10185 2935
rect 10165 2865 10185 2885
rect 10165 2815 10185 2835
rect 10165 2765 10185 2785
rect 10165 2715 10185 2735
rect 10165 2665 10185 2685
rect 10315 3115 10335 3135
rect 10315 3065 10335 3085
rect 10315 3015 10335 3035
rect 10315 2965 10335 2985
rect 10315 2915 10335 2935
rect 10315 2865 10335 2885
rect 10315 2815 10335 2835
rect 10315 2765 10335 2785
rect 10315 2715 10335 2735
rect 10315 2665 10335 2685
rect 10465 3115 10485 3135
rect 10465 3065 10485 3085
rect 10465 3015 10485 3035
rect 10465 2965 10485 2985
rect 10465 2915 10485 2935
rect 10465 2865 10485 2885
rect 10465 2815 10485 2835
rect 10465 2765 10485 2785
rect 10465 2715 10485 2735
rect 10465 2665 10485 2685
rect 10615 3115 10635 3135
rect 10615 3065 10635 3085
rect 10615 3015 10635 3035
rect 10615 2965 10635 2985
rect 10615 2915 10635 2935
rect 10615 2865 10635 2885
rect 10615 2815 10635 2835
rect 10615 2765 10635 2785
rect 10615 2715 10635 2735
rect 10615 2665 10635 2685
rect 10765 3115 10785 3135
rect 10765 3065 10785 3085
rect 10765 3015 10785 3035
rect 10765 2965 10785 2985
rect 10765 2915 10785 2935
rect 10765 2865 10785 2885
rect 10765 2815 10785 2835
rect 10765 2765 10785 2785
rect 10765 2715 10785 2735
rect 10765 2665 10785 2685
rect 11365 3115 11385 3135
rect 11365 3065 11385 3085
rect 11365 3015 11385 3035
rect 11365 2965 11385 2985
rect 11365 2915 11385 2935
rect 11365 2865 11385 2885
rect 11365 2815 11385 2835
rect 11365 2765 11385 2785
rect 11365 2715 11385 2735
rect 11365 2665 11385 2685
rect 11965 3115 11985 3135
rect 11965 3065 11985 3085
rect 11965 3015 11985 3035
rect 11965 2965 11985 2985
rect 11965 2915 11985 2935
rect 11965 2865 11985 2885
rect 11965 2815 11985 2835
rect 11965 2765 11985 2785
rect 11965 2715 11985 2735
rect 11965 2665 11985 2685
rect 12565 3115 12585 3135
rect 12565 3065 12585 3085
rect 12565 3015 12585 3035
rect 12565 2965 12585 2985
rect 12565 2915 12585 2935
rect 12565 2865 12585 2885
rect 12565 2815 12585 2835
rect 12565 2765 12585 2785
rect 12565 2715 12585 2735
rect 12565 2665 12585 2685
rect 13165 3115 13185 3135
rect 13165 3065 13185 3085
rect 13165 3015 13185 3035
rect 13165 2965 13185 2985
rect 13165 2915 13185 2935
rect 13165 2865 13185 2885
rect 13165 2815 13185 2835
rect 13165 2765 13185 2785
rect 13165 2715 13185 2735
rect 13165 2665 13185 2685
rect 13765 3115 13785 3135
rect 13765 3065 13785 3085
rect 13765 3015 13785 3035
rect 13765 2965 13785 2985
rect 13765 2915 13785 2935
rect 13765 2865 13785 2885
rect 13765 2815 13785 2835
rect 13765 2765 13785 2785
rect 13765 2715 13785 2735
rect 13765 2665 13785 2685
rect 14365 3115 14385 3135
rect 14365 3065 14385 3085
rect 14365 3015 14385 3035
rect 14365 2965 14385 2985
rect 14365 2915 14385 2935
rect 14365 2865 14385 2885
rect 14365 2815 14385 2835
rect 14365 2765 14385 2785
rect 14365 2715 14385 2735
rect 14365 2665 14385 2685
rect 14965 3115 14985 3135
rect 14965 3065 14985 3085
rect 14965 3015 14985 3035
rect 14965 2965 14985 2985
rect 14965 2915 14985 2935
rect 14965 2865 14985 2885
rect 14965 2815 14985 2835
rect 14965 2765 14985 2785
rect 14965 2715 14985 2735
rect 14965 2665 14985 2685
rect 15565 3115 15585 3135
rect 15565 3065 15585 3085
rect 15565 3015 15585 3035
rect 15565 2965 15585 2985
rect 15565 2915 15585 2935
rect 15565 2865 15585 2885
rect 15565 2815 15585 2835
rect 15565 2765 15585 2785
rect 15565 2715 15585 2735
rect 15565 2665 15585 2685
rect 16165 3115 16185 3135
rect 16165 3065 16185 3085
rect 16165 3015 16185 3035
rect 16165 2965 16185 2985
rect 16165 2915 16185 2935
rect 16165 2865 16185 2885
rect 16165 2815 16185 2835
rect 16165 2765 16185 2785
rect 16165 2715 16185 2735
rect 16165 2665 16185 2685
rect 16315 3115 16335 3135
rect 16315 3065 16335 3085
rect 16315 3015 16335 3035
rect 16315 2965 16335 2985
rect 16315 2915 16335 2935
rect 16315 2865 16335 2885
rect 16315 2815 16335 2835
rect 16315 2765 16335 2785
rect 16315 2715 16335 2735
rect 16315 2665 16335 2685
rect 16465 3115 16485 3135
rect 16465 3065 16485 3085
rect 16465 3015 16485 3035
rect 16465 2965 16485 2985
rect 16465 2915 16485 2935
rect 16465 2865 16485 2885
rect 16465 2815 16485 2835
rect 16465 2765 16485 2785
rect 16465 2715 16485 2735
rect 16465 2665 16485 2685
rect 16615 3115 16635 3135
rect 16615 3065 16635 3085
rect 16615 3015 16635 3035
rect 16615 2965 16635 2985
rect 16615 2915 16635 2935
rect 16615 2865 16635 2885
rect 16615 2815 16635 2835
rect 16615 2765 16635 2785
rect 16615 2715 16635 2735
rect 16615 2665 16635 2685
rect 16765 3115 16785 3135
rect 16765 3065 16785 3085
rect 16765 3015 16785 3035
rect 16765 2965 16785 2985
rect 16765 2915 16785 2935
rect 16765 2865 16785 2885
rect 16765 2815 16785 2835
rect 16765 2765 16785 2785
rect 16765 2715 16785 2735
rect 16765 2665 16785 2685
rect 16915 3115 16935 3135
rect 16915 3065 16935 3085
rect 16915 3015 16935 3035
rect 16915 2965 16935 2985
rect 16915 2915 16935 2935
rect 16915 2865 16935 2885
rect 16915 2815 16935 2835
rect 16915 2765 16935 2785
rect 16915 2715 16935 2735
rect 16915 2665 16935 2685
rect 17065 3115 17085 3135
rect 17065 3065 17085 3085
rect 17065 3015 17085 3035
rect 17065 2965 17085 2985
rect 17065 2915 17085 2935
rect 17065 2865 17085 2885
rect 17065 2815 17085 2835
rect 17065 2765 17085 2785
rect 17065 2715 17085 2735
rect 17065 2665 17085 2685
rect 17215 3115 17235 3135
rect 17215 3065 17235 3085
rect 17215 3015 17235 3035
rect 17215 2965 17235 2985
rect 17215 2915 17235 2935
rect 17215 2865 17235 2885
rect 17215 2815 17235 2835
rect 17215 2765 17235 2785
rect 17215 2715 17235 2735
rect 17215 2665 17235 2685
rect 17365 3115 17385 3135
rect 17365 3065 17385 3085
rect 17365 3015 17385 3035
rect 17365 2965 17385 2985
rect 17365 2915 17385 2935
rect 17365 2865 17385 2885
rect 17365 2815 17385 2835
rect 17365 2765 17385 2785
rect 17365 2715 17385 2735
rect 17365 2665 17385 2685
rect 17965 3115 17985 3135
rect 17965 3065 17985 3085
rect 17965 3015 17985 3035
rect 17965 2965 17985 2985
rect 17965 2915 17985 2935
rect 17965 2865 17985 2885
rect 17965 2815 17985 2835
rect 17965 2765 17985 2785
rect 17965 2715 17985 2735
rect 17965 2665 17985 2685
rect 18565 3115 18585 3135
rect 18565 3065 18585 3085
rect 18565 3015 18585 3035
rect 18565 2965 18585 2985
rect 18565 2915 18585 2935
rect 18565 2865 18585 2885
rect 18565 2815 18585 2835
rect 18565 2765 18585 2785
rect 18565 2715 18585 2735
rect 18565 2665 18585 2685
rect 18715 3115 18735 3135
rect 18715 3065 18735 3085
rect 18715 3015 18735 3035
rect 18715 2965 18735 2985
rect 18715 2915 18735 2935
rect 18715 2865 18735 2885
rect 18715 2815 18735 2835
rect 18715 2765 18735 2785
rect 18715 2715 18735 2735
rect 18715 2665 18735 2685
rect 18865 3115 18885 3135
rect 18865 3065 18885 3085
rect 18865 3015 18885 3035
rect 18865 2965 18885 2985
rect 18865 2915 18885 2935
rect 18865 2865 18885 2885
rect 18865 2815 18885 2835
rect 18865 2765 18885 2785
rect 18865 2715 18885 2735
rect 18865 2665 18885 2685
rect 19015 3115 19035 3135
rect 19015 3065 19035 3085
rect 19015 3015 19035 3035
rect 19015 2965 19035 2985
rect 19015 2915 19035 2935
rect 19015 2865 19035 2885
rect 19015 2815 19035 2835
rect 19015 2765 19035 2785
rect 19015 2715 19035 2735
rect 19015 2665 19035 2685
rect 19165 3115 19185 3135
rect 19165 3065 19185 3085
rect 19165 3015 19185 3035
rect 19165 2965 19185 2985
rect 19165 2915 19185 2935
rect 19165 2865 19185 2885
rect 19165 2815 19185 2835
rect 19165 2765 19185 2785
rect 19165 2715 19185 2735
rect 19165 2665 19185 2685
rect 19315 3115 19335 3135
rect 19315 3065 19335 3085
rect 19315 3015 19335 3035
rect 19315 2965 19335 2985
rect 19315 2915 19335 2935
rect 19315 2865 19335 2885
rect 19315 2815 19335 2835
rect 19315 2765 19335 2785
rect 19315 2715 19335 2735
rect 19315 2665 19335 2685
rect 19465 3115 19485 3135
rect 19465 3065 19485 3085
rect 19465 3015 19485 3035
rect 19465 2965 19485 2985
rect 19465 2915 19485 2935
rect 19465 2865 19485 2885
rect 19465 2815 19485 2835
rect 19465 2765 19485 2785
rect 19465 2715 19485 2735
rect 19465 2665 19485 2685
rect 19615 3115 19635 3135
rect 19615 3065 19635 3085
rect 19615 3015 19635 3035
rect 19615 2965 19635 2985
rect 19615 2915 19635 2935
rect 19615 2865 19635 2885
rect 19615 2815 19635 2835
rect 19615 2765 19635 2785
rect 19615 2715 19635 2735
rect 19615 2665 19635 2685
rect 19765 3115 19785 3135
rect 19765 3065 19785 3085
rect 19765 3015 19785 3035
rect 19765 2965 19785 2985
rect 19765 2915 19785 2935
rect 19765 2865 19785 2885
rect 19765 2815 19785 2835
rect 19765 2765 19785 2785
rect 19765 2715 19785 2735
rect 19765 2665 19785 2685
rect 20365 3115 20385 3135
rect 20365 3065 20385 3085
rect 20365 3015 20385 3035
rect 20365 2965 20385 2985
rect 20365 2915 20385 2935
rect 20365 2865 20385 2885
rect 20365 2815 20385 2835
rect 20365 2765 20385 2785
rect 20365 2715 20385 2735
rect 20365 2665 20385 2685
<< mvpsubdiff >>
rect -900 2435 20400 2450
rect -900 2415 -885 2435
rect -865 2415 -835 2435
rect -815 2415 -785 2435
rect -765 2415 -735 2435
rect -715 2415 -685 2435
rect -665 2415 -635 2435
rect -615 2415 -585 2435
rect -565 2415 -535 2435
rect -515 2415 -485 2435
rect -465 2415 -435 2435
rect -415 2415 -385 2435
rect -365 2415 -335 2435
rect -315 2415 -285 2435
rect -265 2415 -235 2435
rect -215 2415 -185 2435
rect -165 2415 -135 2435
rect -115 2415 -85 2435
rect -65 2415 -35 2435
rect -15 2415 15 2435
rect 35 2415 65 2435
rect 85 2415 115 2435
rect 135 2415 165 2435
rect 185 2415 215 2435
rect 235 2415 265 2435
rect 285 2415 315 2435
rect 335 2415 365 2435
rect 385 2415 415 2435
rect 435 2415 465 2435
rect 485 2415 515 2435
rect 535 2415 565 2435
rect 585 2415 615 2435
rect 635 2415 665 2435
rect 685 2415 715 2435
rect 735 2415 765 2435
rect 785 2415 815 2435
rect 835 2415 865 2435
rect 885 2415 915 2435
rect 935 2415 965 2435
rect 985 2415 1015 2435
rect 1035 2415 1065 2435
rect 1085 2415 1115 2435
rect 1135 2415 1165 2435
rect 1185 2415 1215 2435
rect 1235 2415 1265 2435
rect 1285 2415 1315 2435
rect 1335 2415 1365 2435
rect 1385 2415 1415 2435
rect 1435 2415 1465 2435
rect 1485 2415 1515 2435
rect 1535 2415 1565 2435
rect 1585 2415 1615 2435
rect 1635 2415 1665 2435
rect 1685 2415 1715 2435
rect 1735 2415 1765 2435
rect 1785 2415 1815 2435
rect 1835 2415 1865 2435
rect 1885 2415 1915 2435
rect 1935 2415 1965 2435
rect 1985 2415 2015 2435
rect 2035 2415 2065 2435
rect 2085 2415 2115 2435
rect 2135 2415 2165 2435
rect 2185 2415 2215 2435
rect 2235 2415 2265 2435
rect 2285 2415 2315 2435
rect 2335 2415 2365 2435
rect 2385 2415 2415 2435
rect 2435 2415 2465 2435
rect 2485 2415 2515 2435
rect 2535 2415 2565 2435
rect 2585 2415 2615 2435
rect 2635 2415 2665 2435
rect 2685 2415 2715 2435
rect 2735 2415 2765 2435
rect 2785 2415 2815 2435
rect 2835 2415 2865 2435
rect 2885 2415 2915 2435
rect 2935 2415 2965 2435
rect 2985 2415 3015 2435
rect 3035 2415 3065 2435
rect 3085 2415 3115 2435
rect 3135 2415 3165 2435
rect 3185 2415 3215 2435
rect 3235 2415 3265 2435
rect 3285 2415 3315 2435
rect 3335 2415 3365 2435
rect 3385 2415 3415 2435
rect 3435 2415 3465 2435
rect 3485 2415 3515 2435
rect 3535 2415 3565 2435
rect 3585 2415 3615 2435
rect 3635 2415 3665 2435
rect 3685 2415 3715 2435
rect 3735 2415 3765 2435
rect 3785 2415 3815 2435
rect 3835 2415 3865 2435
rect 3885 2415 3915 2435
rect 3935 2415 3965 2435
rect 3985 2415 4015 2435
rect 4035 2415 4065 2435
rect 4085 2415 4115 2435
rect 4135 2415 4165 2435
rect 4185 2415 4215 2435
rect 4235 2415 4265 2435
rect 4285 2415 4315 2435
rect 4335 2415 4365 2435
rect 4385 2415 4415 2435
rect 4435 2415 4465 2435
rect 4485 2415 4515 2435
rect 4535 2415 4565 2435
rect 4585 2415 4615 2435
rect 4635 2415 4665 2435
rect 4685 2415 4715 2435
rect 4735 2415 4765 2435
rect 4785 2415 4815 2435
rect 4835 2415 4865 2435
rect 4885 2415 4915 2435
rect 4935 2415 4965 2435
rect 4985 2415 5015 2435
rect 5035 2415 5065 2435
rect 5085 2415 5115 2435
rect 5135 2415 5165 2435
rect 5185 2415 5215 2435
rect 5235 2415 5265 2435
rect 5285 2415 5315 2435
rect 5335 2415 5365 2435
rect 5385 2415 5415 2435
rect 5435 2415 5465 2435
rect 5485 2415 5515 2435
rect 5535 2415 5565 2435
rect 5585 2415 5615 2435
rect 5635 2415 5665 2435
rect 5685 2415 5715 2435
rect 5735 2415 5765 2435
rect 5785 2415 5815 2435
rect 5835 2415 5865 2435
rect 5885 2415 5915 2435
rect 5935 2415 5965 2435
rect 5985 2415 6015 2435
rect 6035 2415 6065 2435
rect 6085 2415 6115 2435
rect 6135 2415 6165 2435
rect 6185 2415 6215 2435
rect 6235 2415 6265 2435
rect 6285 2415 6315 2435
rect 6335 2415 6365 2435
rect 6385 2415 6415 2435
rect 6435 2415 6465 2435
rect 6485 2415 6515 2435
rect 6535 2415 6565 2435
rect 6585 2415 6615 2435
rect 6635 2415 6665 2435
rect 6685 2415 6715 2435
rect 6735 2415 6765 2435
rect 6785 2415 6815 2435
rect 6835 2415 6865 2435
rect 6885 2415 6915 2435
rect 6935 2415 6965 2435
rect 6985 2415 7015 2435
rect 7035 2415 7065 2435
rect 7085 2415 7115 2435
rect 7135 2415 7165 2435
rect 7185 2415 7215 2435
rect 7235 2415 7265 2435
rect 7285 2415 7315 2435
rect 7335 2415 7365 2435
rect 7385 2415 7415 2435
rect 7435 2415 7465 2435
rect 7485 2415 7515 2435
rect 7535 2415 7565 2435
rect 7585 2415 7615 2435
rect 7635 2415 7665 2435
rect 7685 2415 7715 2435
rect 7735 2415 7765 2435
rect 7785 2415 7815 2435
rect 7835 2415 7865 2435
rect 7885 2415 7915 2435
rect 7935 2415 7965 2435
rect 7985 2415 8015 2435
rect 8035 2415 8065 2435
rect 8085 2415 8115 2435
rect 8135 2415 8165 2435
rect 8185 2415 8215 2435
rect 8235 2415 8265 2435
rect 8285 2415 8315 2435
rect 8335 2415 8365 2435
rect 8385 2415 8415 2435
rect 8435 2415 8465 2435
rect 8485 2415 8515 2435
rect 8535 2415 8565 2435
rect 8585 2415 8615 2435
rect 8635 2415 8665 2435
rect 8685 2415 8715 2435
rect 8735 2415 8765 2435
rect 8785 2415 8815 2435
rect 8835 2415 8865 2435
rect 8885 2415 8915 2435
rect 8935 2415 8965 2435
rect 8985 2415 9015 2435
rect 9035 2415 9065 2435
rect 9085 2415 9115 2435
rect 9135 2415 9165 2435
rect 9185 2415 9215 2435
rect 9235 2415 9265 2435
rect 9285 2415 9315 2435
rect 9335 2415 9365 2435
rect 9385 2415 9415 2435
rect 9435 2415 9465 2435
rect 9485 2415 9515 2435
rect 9535 2415 9565 2435
rect 9585 2415 9615 2435
rect 9635 2415 9665 2435
rect 9685 2415 9715 2435
rect 9735 2415 9765 2435
rect 9785 2415 9815 2435
rect 9835 2415 9865 2435
rect 9885 2415 9915 2435
rect 9935 2415 9965 2435
rect 9985 2415 10015 2435
rect 10035 2415 10065 2435
rect 10085 2415 10115 2435
rect 10135 2415 10165 2435
rect 10185 2415 10215 2435
rect 10235 2415 10265 2435
rect 10285 2415 10315 2435
rect 10335 2415 10365 2435
rect 10385 2415 10415 2435
rect 10435 2415 10465 2435
rect 10485 2415 10515 2435
rect 10535 2415 10565 2435
rect 10585 2415 10615 2435
rect 10635 2415 10665 2435
rect 10685 2415 10715 2435
rect 10735 2415 10765 2435
rect 10785 2415 10815 2435
rect 10835 2415 10865 2435
rect 10885 2415 10915 2435
rect 10935 2415 10965 2435
rect 10985 2415 11015 2435
rect 11035 2415 11065 2435
rect 11085 2415 11115 2435
rect 11135 2415 11165 2435
rect 11185 2415 11215 2435
rect 11235 2415 11265 2435
rect 11285 2415 11315 2435
rect 11335 2415 11365 2435
rect 11385 2415 11415 2435
rect 11435 2415 11465 2435
rect 11485 2415 11515 2435
rect 11535 2415 11565 2435
rect 11585 2415 11615 2435
rect 11635 2415 11665 2435
rect 11685 2415 11715 2435
rect 11735 2415 11765 2435
rect 11785 2415 11815 2435
rect 11835 2415 11865 2435
rect 11885 2415 11915 2435
rect 11935 2415 11965 2435
rect 11985 2415 12015 2435
rect 12035 2415 12065 2435
rect 12085 2415 12115 2435
rect 12135 2415 12165 2435
rect 12185 2415 12215 2435
rect 12235 2415 12265 2435
rect 12285 2415 12315 2435
rect 12335 2415 12365 2435
rect 12385 2415 12415 2435
rect 12435 2415 12465 2435
rect 12485 2415 12515 2435
rect 12535 2415 12565 2435
rect 12585 2415 12615 2435
rect 12635 2415 12665 2435
rect 12685 2415 12715 2435
rect 12735 2415 12765 2435
rect 12785 2415 12815 2435
rect 12835 2415 12865 2435
rect 12885 2415 12915 2435
rect 12935 2415 12965 2435
rect 12985 2415 13015 2435
rect 13035 2415 13065 2435
rect 13085 2415 13115 2435
rect 13135 2415 13165 2435
rect 13185 2415 13215 2435
rect 13235 2415 13265 2435
rect 13285 2415 13315 2435
rect 13335 2415 13365 2435
rect 13385 2415 13415 2435
rect 13435 2415 13465 2435
rect 13485 2415 13515 2435
rect 13535 2415 13565 2435
rect 13585 2415 13615 2435
rect 13635 2415 13665 2435
rect 13685 2415 13715 2435
rect 13735 2415 13765 2435
rect 13785 2415 13815 2435
rect 13835 2415 13865 2435
rect 13885 2415 13915 2435
rect 13935 2415 13965 2435
rect 13985 2415 14015 2435
rect 14035 2415 14065 2435
rect 14085 2415 14115 2435
rect 14135 2415 14165 2435
rect 14185 2415 14215 2435
rect 14235 2415 14265 2435
rect 14285 2415 14315 2435
rect 14335 2415 14365 2435
rect 14385 2415 14415 2435
rect 14435 2415 14465 2435
rect 14485 2415 14515 2435
rect 14535 2415 14565 2435
rect 14585 2415 14615 2435
rect 14635 2415 14665 2435
rect 14685 2415 14715 2435
rect 14735 2415 14765 2435
rect 14785 2415 14815 2435
rect 14835 2415 14865 2435
rect 14885 2415 14915 2435
rect 14935 2415 14965 2435
rect 14985 2415 15015 2435
rect 15035 2415 15065 2435
rect 15085 2415 15115 2435
rect 15135 2415 15165 2435
rect 15185 2415 15215 2435
rect 15235 2415 15265 2435
rect 15285 2415 15315 2435
rect 15335 2415 15365 2435
rect 15385 2415 15415 2435
rect 15435 2415 15465 2435
rect 15485 2415 15515 2435
rect 15535 2415 15565 2435
rect 15585 2415 15615 2435
rect 15635 2415 15665 2435
rect 15685 2415 15715 2435
rect 15735 2415 15765 2435
rect 15785 2415 15815 2435
rect 15835 2415 15865 2435
rect 15885 2415 15915 2435
rect 15935 2415 15965 2435
rect 15985 2415 16015 2435
rect 16035 2415 16065 2435
rect 16085 2415 16115 2435
rect 16135 2415 16165 2435
rect 16185 2415 16215 2435
rect 16235 2415 16265 2435
rect 16285 2415 16315 2435
rect 16335 2415 16365 2435
rect 16385 2415 16415 2435
rect 16435 2415 16465 2435
rect 16485 2415 16515 2435
rect 16535 2415 16565 2435
rect 16585 2415 16615 2435
rect 16635 2415 16665 2435
rect 16685 2415 16715 2435
rect 16735 2415 16765 2435
rect 16785 2415 16815 2435
rect 16835 2415 16865 2435
rect 16885 2415 16915 2435
rect 16935 2415 16965 2435
rect 16985 2415 17015 2435
rect 17035 2415 17065 2435
rect 17085 2415 17115 2435
rect 17135 2415 17165 2435
rect 17185 2415 17215 2435
rect 17235 2415 17265 2435
rect 17285 2415 17315 2435
rect 17335 2415 17365 2435
rect 17385 2415 17415 2435
rect 17435 2415 17465 2435
rect 17485 2415 17515 2435
rect 17535 2415 17565 2435
rect 17585 2415 17615 2435
rect 17635 2415 17665 2435
rect 17685 2415 17715 2435
rect 17735 2415 17765 2435
rect 17785 2415 17815 2435
rect 17835 2415 17865 2435
rect 17885 2415 17915 2435
rect 17935 2415 17965 2435
rect 17985 2415 18015 2435
rect 18035 2415 18065 2435
rect 18085 2415 18115 2435
rect 18135 2415 18165 2435
rect 18185 2415 18215 2435
rect 18235 2415 18265 2435
rect 18285 2415 18315 2435
rect 18335 2415 18365 2435
rect 18385 2415 18415 2435
rect 18435 2415 18465 2435
rect 18485 2415 18515 2435
rect 18535 2415 18565 2435
rect 18585 2415 18615 2435
rect 18635 2415 18665 2435
rect 18685 2415 18715 2435
rect 18735 2415 18765 2435
rect 18785 2415 18815 2435
rect 18835 2415 18865 2435
rect 18885 2415 18915 2435
rect 18935 2415 18965 2435
rect 18985 2415 19015 2435
rect 19035 2415 19065 2435
rect 19085 2415 19115 2435
rect 19135 2415 19165 2435
rect 19185 2415 19215 2435
rect 19235 2415 19265 2435
rect 19285 2415 19315 2435
rect 19335 2415 19365 2435
rect 19385 2415 19415 2435
rect 19435 2415 19465 2435
rect 19485 2415 19515 2435
rect 19535 2415 19565 2435
rect 19585 2415 19615 2435
rect 19635 2415 19665 2435
rect 19685 2415 19715 2435
rect 19735 2415 19765 2435
rect 19785 2415 19815 2435
rect 19835 2415 19865 2435
rect 19885 2415 19915 2435
rect 19935 2415 19965 2435
rect 19985 2415 20015 2435
rect 20035 2415 20065 2435
rect 20085 2415 20115 2435
rect 20135 2415 20165 2435
rect 20185 2415 20215 2435
rect 20235 2415 20265 2435
rect 20285 2415 20315 2435
rect 20335 2415 20365 2435
rect 20385 2415 20400 2435
rect -900 2400 20400 2415
rect -900 2035 20400 2050
rect -900 2015 -885 2035
rect -865 2015 -835 2035
rect -815 2015 -785 2035
rect -765 2015 -735 2035
rect -715 2015 -685 2035
rect -665 2015 -635 2035
rect -615 2015 -585 2035
rect -565 2015 -535 2035
rect -515 2015 -485 2035
rect -465 2015 -435 2035
rect -415 2015 -385 2035
rect -365 2015 -335 2035
rect -315 2015 -285 2035
rect -265 2015 -235 2035
rect -215 2015 -185 2035
rect -165 2015 -135 2035
rect -115 2015 -85 2035
rect -65 2015 -35 2035
rect -15 2015 15 2035
rect 35 2015 65 2035
rect 85 2015 115 2035
rect 135 2015 165 2035
rect 185 2015 215 2035
rect 235 2015 265 2035
rect 285 2015 315 2035
rect 335 2015 365 2035
rect 385 2015 415 2035
rect 435 2015 465 2035
rect 485 2015 515 2035
rect 535 2015 565 2035
rect 585 2015 615 2035
rect 635 2015 665 2035
rect 685 2015 715 2035
rect 735 2015 765 2035
rect 785 2015 815 2035
rect 835 2015 865 2035
rect 885 2015 915 2035
rect 935 2015 965 2035
rect 985 2015 1015 2035
rect 1035 2015 1065 2035
rect 1085 2015 1115 2035
rect 1135 2015 1165 2035
rect 1185 2015 1215 2035
rect 1235 2015 1265 2035
rect 1285 2015 1315 2035
rect 1335 2015 1365 2035
rect 1385 2015 1415 2035
rect 1435 2015 1465 2035
rect 1485 2015 1515 2035
rect 1535 2015 1565 2035
rect 1585 2015 1615 2035
rect 1635 2015 1665 2035
rect 1685 2015 1715 2035
rect 1735 2015 1765 2035
rect 1785 2015 1815 2035
rect 1835 2015 1865 2035
rect 1885 2015 1915 2035
rect 1935 2015 1965 2035
rect 1985 2015 2015 2035
rect 2035 2015 2065 2035
rect 2085 2015 2115 2035
rect 2135 2015 2165 2035
rect 2185 2015 2215 2035
rect 2235 2015 2265 2035
rect 2285 2015 2315 2035
rect 2335 2015 2365 2035
rect 2385 2015 2415 2035
rect 2435 2015 2465 2035
rect 2485 2015 2515 2035
rect 2535 2015 2565 2035
rect 2585 2015 2615 2035
rect 2635 2015 2665 2035
rect 2685 2015 2715 2035
rect 2735 2015 2765 2035
rect 2785 2015 2815 2035
rect 2835 2015 2865 2035
rect 2885 2015 2915 2035
rect 2935 2015 2965 2035
rect 2985 2015 3015 2035
rect 3035 2015 3065 2035
rect 3085 2015 3115 2035
rect 3135 2015 3165 2035
rect 3185 2015 3215 2035
rect 3235 2015 3265 2035
rect 3285 2015 3315 2035
rect 3335 2015 3365 2035
rect 3385 2015 3415 2035
rect 3435 2015 3465 2035
rect 3485 2015 3515 2035
rect 3535 2015 3565 2035
rect 3585 2015 3615 2035
rect 3635 2015 3665 2035
rect 3685 2015 3715 2035
rect 3735 2015 3765 2035
rect 3785 2015 3815 2035
rect 3835 2015 3865 2035
rect 3885 2015 3915 2035
rect 3935 2015 3965 2035
rect 3985 2015 4015 2035
rect 4035 2015 4065 2035
rect 4085 2015 4115 2035
rect 4135 2015 4165 2035
rect 4185 2015 4215 2035
rect 4235 2015 4265 2035
rect 4285 2015 4315 2035
rect 4335 2015 4365 2035
rect 4385 2015 4415 2035
rect 4435 2015 4465 2035
rect 4485 2015 4515 2035
rect 4535 2015 4565 2035
rect 4585 2015 4615 2035
rect 4635 2015 4665 2035
rect 4685 2015 4715 2035
rect 4735 2015 4765 2035
rect 4785 2015 4815 2035
rect 4835 2015 4865 2035
rect 4885 2015 4915 2035
rect 4935 2015 4965 2035
rect 4985 2015 5015 2035
rect 5035 2015 5065 2035
rect 5085 2015 5115 2035
rect 5135 2015 5165 2035
rect 5185 2015 5215 2035
rect 5235 2015 5265 2035
rect 5285 2015 5315 2035
rect 5335 2015 5365 2035
rect 5385 2015 5415 2035
rect 5435 2015 5465 2035
rect 5485 2015 5515 2035
rect 5535 2015 5565 2035
rect 5585 2015 5615 2035
rect 5635 2015 5665 2035
rect 5685 2015 5715 2035
rect 5735 2015 5765 2035
rect 5785 2015 5815 2035
rect 5835 2015 5865 2035
rect 5885 2015 5915 2035
rect 5935 2015 5965 2035
rect 5985 2015 6015 2035
rect 6035 2015 6065 2035
rect 6085 2015 6115 2035
rect 6135 2015 6165 2035
rect 6185 2015 6215 2035
rect 6235 2015 6265 2035
rect 6285 2015 6315 2035
rect 6335 2015 6365 2035
rect 6385 2015 6415 2035
rect 6435 2015 6465 2035
rect 6485 2015 6515 2035
rect 6535 2015 6565 2035
rect 6585 2015 6615 2035
rect 6635 2015 6665 2035
rect 6685 2015 6715 2035
rect 6735 2015 6765 2035
rect 6785 2015 6815 2035
rect 6835 2015 6865 2035
rect 6885 2015 6915 2035
rect 6935 2015 6965 2035
rect 6985 2015 7015 2035
rect 7035 2015 7065 2035
rect 7085 2015 7115 2035
rect 7135 2015 7165 2035
rect 7185 2015 7215 2035
rect 7235 2015 7265 2035
rect 7285 2015 7315 2035
rect 7335 2015 7365 2035
rect 7385 2015 7415 2035
rect 7435 2015 7465 2035
rect 7485 2015 7515 2035
rect 7535 2015 7565 2035
rect 7585 2015 7615 2035
rect 7635 2015 7665 2035
rect 7685 2015 7715 2035
rect 7735 2015 7765 2035
rect 7785 2015 7815 2035
rect 7835 2015 7865 2035
rect 7885 2015 7915 2035
rect 7935 2015 7965 2035
rect 7985 2015 8015 2035
rect 8035 2015 8065 2035
rect 8085 2015 8115 2035
rect 8135 2015 8165 2035
rect 8185 2015 8215 2035
rect 8235 2015 8265 2035
rect 8285 2015 8315 2035
rect 8335 2015 8365 2035
rect 8385 2015 8415 2035
rect 8435 2015 8465 2035
rect 8485 2015 8515 2035
rect 8535 2015 8565 2035
rect 8585 2015 8615 2035
rect 8635 2015 8665 2035
rect 8685 2015 8715 2035
rect 8735 2015 8765 2035
rect 8785 2015 8815 2035
rect 8835 2015 8865 2035
rect 8885 2015 8915 2035
rect 8935 2015 8965 2035
rect 8985 2015 9015 2035
rect 9035 2015 9065 2035
rect 9085 2015 9115 2035
rect 9135 2015 9165 2035
rect 9185 2015 9215 2035
rect 9235 2015 9265 2035
rect 9285 2015 9315 2035
rect 9335 2015 9365 2035
rect 9385 2015 9415 2035
rect 9435 2015 9465 2035
rect 9485 2015 9515 2035
rect 9535 2015 9565 2035
rect 9585 2015 9615 2035
rect 9635 2015 9665 2035
rect 9685 2015 9715 2035
rect 9735 2015 9765 2035
rect 9785 2015 9815 2035
rect 9835 2015 9865 2035
rect 9885 2015 9915 2035
rect 9935 2015 9965 2035
rect 9985 2015 10015 2035
rect 10035 2015 10065 2035
rect 10085 2015 10115 2035
rect 10135 2015 10165 2035
rect 10185 2015 10215 2035
rect 10235 2015 10265 2035
rect 10285 2015 10315 2035
rect 10335 2015 10365 2035
rect 10385 2015 10415 2035
rect 10435 2015 10465 2035
rect 10485 2015 10515 2035
rect 10535 2015 10565 2035
rect 10585 2015 10615 2035
rect 10635 2015 10665 2035
rect 10685 2015 10715 2035
rect 10735 2015 10765 2035
rect 10785 2015 10815 2035
rect 10835 2015 10865 2035
rect 10885 2015 10915 2035
rect 10935 2015 10965 2035
rect 10985 2015 11015 2035
rect 11035 2015 11065 2035
rect 11085 2015 11115 2035
rect 11135 2015 11165 2035
rect 11185 2015 11215 2035
rect 11235 2015 11265 2035
rect 11285 2015 11315 2035
rect 11335 2015 11365 2035
rect 11385 2015 11415 2035
rect 11435 2015 11465 2035
rect 11485 2015 11515 2035
rect 11535 2015 11565 2035
rect 11585 2015 11615 2035
rect 11635 2015 11665 2035
rect 11685 2015 11715 2035
rect 11735 2015 11765 2035
rect 11785 2015 11815 2035
rect 11835 2015 11865 2035
rect 11885 2015 11915 2035
rect 11935 2015 11965 2035
rect 11985 2015 12015 2035
rect 12035 2015 12065 2035
rect 12085 2015 12115 2035
rect 12135 2015 12165 2035
rect 12185 2015 12215 2035
rect 12235 2015 12265 2035
rect 12285 2015 12315 2035
rect 12335 2015 12365 2035
rect 12385 2015 12415 2035
rect 12435 2015 12465 2035
rect 12485 2015 12515 2035
rect 12535 2015 12565 2035
rect 12585 2015 12615 2035
rect 12635 2015 12665 2035
rect 12685 2015 12715 2035
rect 12735 2015 12765 2035
rect 12785 2015 12815 2035
rect 12835 2015 12865 2035
rect 12885 2015 12915 2035
rect 12935 2015 12965 2035
rect 12985 2015 13015 2035
rect 13035 2015 13065 2035
rect 13085 2015 13115 2035
rect 13135 2015 13165 2035
rect 13185 2015 13215 2035
rect 13235 2015 13265 2035
rect 13285 2015 13315 2035
rect 13335 2015 13365 2035
rect 13385 2015 13415 2035
rect 13435 2015 13465 2035
rect 13485 2015 13515 2035
rect 13535 2015 13565 2035
rect 13585 2015 13615 2035
rect 13635 2015 13665 2035
rect 13685 2015 13715 2035
rect 13735 2015 13765 2035
rect 13785 2015 13815 2035
rect 13835 2015 13865 2035
rect 13885 2015 13915 2035
rect 13935 2015 13965 2035
rect 13985 2015 14015 2035
rect 14035 2015 14065 2035
rect 14085 2015 14115 2035
rect 14135 2015 14165 2035
rect 14185 2015 14215 2035
rect 14235 2015 14265 2035
rect 14285 2015 14315 2035
rect 14335 2015 14365 2035
rect 14385 2015 14415 2035
rect 14435 2015 14465 2035
rect 14485 2015 14515 2035
rect 14535 2015 14565 2035
rect 14585 2015 14615 2035
rect 14635 2015 14665 2035
rect 14685 2015 14715 2035
rect 14735 2015 14765 2035
rect 14785 2015 14815 2035
rect 14835 2015 14865 2035
rect 14885 2015 14915 2035
rect 14935 2015 14965 2035
rect 14985 2015 15015 2035
rect 15035 2015 15065 2035
rect 15085 2015 15115 2035
rect 15135 2015 15165 2035
rect 15185 2015 15215 2035
rect 15235 2015 15265 2035
rect 15285 2015 15315 2035
rect 15335 2015 15365 2035
rect 15385 2015 15415 2035
rect 15435 2015 15465 2035
rect 15485 2015 15515 2035
rect 15535 2015 15565 2035
rect 15585 2015 15615 2035
rect 15635 2015 15665 2035
rect 15685 2015 15715 2035
rect 15735 2015 15765 2035
rect 15785 2015 15815 2035
rect 15835 2015 15865 2035
rect 15885 2015 15915 2035
rect 15935 2015 15965 2035
rect 15985 2015 16015 2035
rect 16035 2015 16065 2035
rect 16085 2015 16115 2035
rect 16135 2015 16165 2035
rect 16185 2015 16215 2035
rect 16235 2015 16265 2035
rect 16285 2015 16315 2035
rect 16335 2015 16365 2035
rect 16385 2015 16415 2035
rect 16435 2015 16465 2035
rect 16485 2015 16515 2035
rect 16535 2015 16565 2035
rect 16585 2015 16615 2035
rect 16635 2015 16665 2035
rect 16685 2015 16715 2035
rect 16735 2015 16765 2035
rect 16785 2015 16815 2035
rect 16835 2015 16865 2035
rect 16885 2015 16915 2035
rect 16935 2015 16965 2035
rect 16985 2015 17015 2035
rect 17035 2015 17065 2035
rect 17085 2015 17115 2035
rect 17135 2015 17165 2035
rect 17185 2015 17215 2035
rect 17235 2015 17265 2035
rect 17285 2015 17315 2035
rect 17335 2015 17365 2035
rect 17385 2015 17415 2035
rect 17435 2015 17465 2035
rect 17485 2015 17515 2035
rect 17535 2015 17565 2035
rect 17585 2015 17615 2035
rect 17635 2015 17665 2035
rect 17685 2015 17715 2035
rect 17735 2015 17765 2035
rect 17785 2015 17815 2035
rect 17835 2015 17865 2035
rect 17885 2015 17915 2035
rect 17935 2015 17965 2035
rect 17985 2015 18015 2035
rect 18035 2015 18065 2035
rect 18085 2015 18115 2035
rect 18135 2015 18165 2035
rect 18185 2015 18215 2035
rect 18235 2015 18265 2035
rect 18285 2015 18315 2035
rect 18335 2015 18365 2035
rect 18385 2015 18415 2035
rect 18435 2015 18465 2035
rect 18485 2015 18515 2035
rect 18535 2015 18565 2035
rect 18585 2015 18615 2035
rect 18635 2015 18665 2035
rect 18685 2015 18715 2035
rect 18735 2015 18765 2035
rect 18785 2015 18815 2035
rect 18835 2015 18865 2035
rect 18885 2015 18915 2035
rect 18935 2015 18965 2035
rect 18985 2015 19015 2035
rect 19035 2015 19065 2035
rect 19085 2015 19115 2035
rect 19135 2015 19165 2035
rect 19185 2015 19215 2035
rect 19235 2015 19265 2035
rect 19285 2015 19315 2035
rect 19335 2015 19365 2035
rect 19385 2015 19415 2035
rect 19435 2015 19465 2035
rect 19485 2015 19515 2035
rect 19535 2015 19565 2035
rect 19585 2015 19615 2035
rect 19635 2015 19665 2035
rect 19685 2015 19715 2035
rect 19735 2015 19765 2035
rect 19785 2015 19815 2035
rect 19835 2015 19865 2035
rect 19885 2015 19915 2035
rect 19935 2015 19965 2035
rect 19985 2015 20015 2035
rect 20035 2015 20065 2035
rect 20085 2015 20115 2035
rect 20135 2015 20165 2035
rect 20185 2015 20215 2035
rect 20235 2015 20265 2035
rect 20285 2015 20315 2035
rect 20335 2015 20365 2035
rect 20385 2015 20400 2035
rect -900 2000 20400 2015
rect -650 1685 20400 1700
rect -650 1665 -635 1685
rect -615 1665 -585 1685
rect -565 1665 -535 1685
rect -515 1665 -485 1685
rect -465 1665 -435 1685
rect -415 1665 -385 1685
rect -365 1665 -335 1685
rect -315 1665 -285 1685
rect -265 1665 -235 1685
rect -215 1665 -185 1685
rect -165 1665 -135 1685
rect -115 1665 -85 1685
rect -65 1665 -35 1685
rect -15 1665 15 1685
rect 35 1665 65 1685
rect 85 1665 115 1685
rect 135 1665 165 1685
rect 185 1665 215 1685
rect 235 1665 265 1685
rect 285 1665 315 1685
rect 335 1665 365 1685
rect 385 1665 415 1685
rect 435 1665 465 1685
rect 485 1665 515 1685
rect 535 1665 565 1685
rect 585 1665 615 1685
rect 635 1665 665 1685
rect 685 1665 715 1685
rect 735 1665 765 1685
rect 785 1665 815 1685
rect 835 1665 865 1685
rect 885 1665 915 1685
rect 935 1665 965 1685
rect 985 1665 1015 1685
rect 1035 1665 1065 1685
rect 1085 1665 1115 1685
rect 1135 1665 1165 1685
rect 1185 1665 1215 1685
rect 1235 1665 1265 1685
rect 1285 1665 1315 1685
rect 1335 1665 1365 1685
rect 1385 1665 1415 1685
rect 1435 1665 1465 1685
rect 1485 1665 1515 1685
rect 1535 1665 1565 1685
rect 1585 1665 1615 1685
rect 1635 1665 1665 1685
rect 1685 1665 1715 1685
rect 1735 1665 1765 1685
rect 1785 1665 1815 1685
rect 1835 1665 1865 1685
rect 1885 1665 1915 1685
rect 1935 1665 1965 1685
rect 1985 1665 2015 1685
rect 2035 1665 2065 1685
rect 2085 1665 2115 1685
rect 2135 1665 2165 1685
rect 2185 1665 2215 1685
rect 2235 1665 2265 1685
rect 2285 1665 2315 1685
rect 2335 1665 2365 1685
rect 2385 1665 2415 1685
rect 2435 1665 2465 1685
rect 2485 1665 2515 1685
rect 2535 1665 2565 1685
rect 2585 1665 2615 1685
rect 2635 1665 2665 1685
rect 2685 1665 2715 1685
rect 2735 1665 2765 1685
rect 2785 1665 2815 1685
rect 2835 1665 2865 1685
rect 2885 1665 2915 1685
rect 2935 1665 2965 1685
rect 2985 1665 3015 1685
rect 3035 1665 3065 1685
rect 3085 1665 3115 1685
rect 3135 1665 3165 1685
rect 3185 1665 3215 1685
rect 3235 1665 3265 1685
rect 3285 1665 3315 1685
rect 3335 1665 3365 1685
rect 3385 1665 3415 1685
rect 3435 1665 3465 1685
rect 3485 1665 3515 1685
rect 3535 1665 3565 1685
rect 3585 1665 3615 1685
rect 3635 1665 3665 1685
rect 3685 1665 3715 1685
rect 3735 1665 3765 1685
rect 3785 1665 3815 1685
rect 3835 1665 3865 1685
rect 3885 1665 3915 1685
rect 3935 1665 3965 1685
rect 3985 1665 4015 1685
rect 4035 1665 4065 1685
rect 4085 1665 4115 1685
rect 4135 1665 4165 1685
rect 4185 1665 4215 1685
rect 4235 1665 4265 1685
rect 4285 1665 4315 1685
rect 4335 1665 4365 1685
rect 4385 1665 4415 1685
rect 4435 1665 4465 1685
rect 4485 1665 4515 1685
rect 4535 1665 4565 1685
rect 4585 1665 4615 1685
rect 4635 1665 4665 1685
rect 4685 1665 4715 1685
rect 4735 1665 4765 1685
rect 4785 1665 4815 1685
rect 4835 1665 4865 1685
rect 4885 1665 4915 1685
rect 4935 1665 4965 1685
rect 4985 1665 5015 1685
rect 5035 1665 5065 1685
rect 5085 1665 5115 1685
rect 5135 1665 5165 1685
rect 5185 1665 5215 1685
rect 5235 1665 5265 1685
rect 5285 1665 5315 1685
rect 5335 1665 5365 1685
rect 5385 1665 5415 1685
rect 5435 1665 5465 1685
rect 5485 1665 5515 1685
rect 5535 1665 5565 1685
rect 5585 1665 5615 1685
rect 5635 1665 5665 1685
rect 5685 1665 5715 1685
rect 5735 1665 5765 1685
rect 5785 1665 5815 1685
rect 5835 1665 5865 1685
rect 5885 1665 5915 1685
rect 5935 1665 5965 1685
rect 5985 1665 6015 1685
rect 6035 1665 6065 1685
rect 6085 1665 6115 1685
rect 6135 1665 6165 1685
rect 6185 1665 6215 1685
rect 6235 1665 6265 1685
rect 6285 1665 6315 1685
rect 6335 1665 6365 1685
rect 6385 1665 6415 1685
rect 6435 1665 6465 1685
rect 6485 1665 6515 1685
rect 6535 1665 6565 1685
rect 6585 1665 6615 1685
rect 6635 1665 6665 1685
rect 6685 1665 6715 1685
rect 6735 1665 6765 1685
rect 6785 1665 6815 1685
rect 6835 1665 6865 1685
rect 6885 1665 6915 1685
rect 6935 1665 6965 1685
rect 6985 1665 7015 1685
rect 7035 1665 7065 1685
rect 7085 1665 7115 1685
rect 7135 1665 7165 1685
rect 7185 1665 7215 1685
rect 7235 1665 7265 1685
rect 7285 1665 7315 1685
rect 7335 1665 7365 1685
rect 7385 1665 7415 1685
rect 7435 1665 7465 1685
rect 7485 1665 7515 1685
rect 7535 1665 7565 1685
rect 7585 1665 7615 1685
rect 7635 1665 7665 1685
rect 7685 1665 7715 1685
rect 7735 1665 7765 1685
rect 7785 1665 7815 1685
rect 7835 1665 7865 1685
rect 7885 1665 7915 1685
rect 7935 1665 7965 1685
rect 7985 1665 8015 1685
rect 8035 1665 8065 1685
rect 8085 1665 8115 1685
rect 8135 1665 8165 1685
rect 8185 1665 8215 1685
rect 8235 1665 8265 1685
rect 8285 1665 8315 1685
rect 8335 1665 8365 1685
rect 8385 1665 8415 1685
rect 8435 1665 8465 1685
rect 8485 1665 8515 1685
rect 8535 1665 8565 1685
rect 8585 1665 8615 1685
rect 8635 1665 8665 1685
rect 8685 1665 8715 1685
rect 8735 1665 8765 1685
rect 8785 1665 8815 1685
rect 8835 1665 8865 1685
rect 8885 1665 8915 1685
rect 8935 1665 8965 1685
rect 8985 1665 9015 1685
rect 9035 1665 9065 1685
rect 9085 1665 9115 1685
rect 9135 1665 9165 1685
rect 9185 1665 9215 1685
rect 9235 1665 9265 1685
rect 9285 1665 9315 1685
rect 9335 1665 9365 1685
rect 9385 1665 9415 1685
rect 9435 1665 9465 1685
rect 9485 1665 9515 1685
rect 9535 1665 9565 1685
rect 9585 1665 9615 1685
rect 9635 1665 9665 1685
rect 9685 1665 9715 1685
rect 9735 1665 9765 1685
rect 9785 1665 9815 1685
rect 9835 1665 9865 1685
rect 9885 1665 9915 1685
rect 9935 1665 9965 1685
rect 9985 1665 10015 1685
rect 10035 1665 10065 1685
rect 10085 1665 10115 1685
rect 10135 1665 10165 1685
rect 10185 1665 10215 1685
rect 10235 1665 10265 1685
rect 10285 1665 10315 1685
rect 10335 1665 10365 1685
rect 10385 1665 10415 1685
rect 10435 1665 10465 1685
rect 10485 1665 10515 1685
rect 10535 1665 10565 1685
rect 10585 1665 10615 1685
rect 10635 1665 10665 1685
rect 10685 1665 10715 1685
rect 10735 1665 10765 1685
rect 10785 1665 10815 1685
rect 10835 1665 10865 1685
rect 10885 1665 10915 1685
rect 10935 1665 10965 1685
rect 10985 1665 11015 1685
rect 11035 1665 11065 1685
rect 11085 1665 11115 1685
rect 11135 1665 11165 1685
rect 11185 1665 11215 1685
rect 11235 1665 11265 1685
rect 11285 1665 11315 1685
rect 11335 1665 11365 1685
rect 11385 1665 11415 1685
rect 11435 1665 11465 1685
rect 11485 1665 11515 1685
rect 11535 1665 11565 1685
rect 11585 1665 11615 1685
rect 11635 1665 11665 1685
rect 11685 1665 11715 1685
rect 11735 1665 11765 1685
rect 11785 1665 11815 1685
rect 11835 1665 11865 1685
rect 11885 1665 11915 1685
rect 11935 1665 11965 1685
rect 11985 1665 12015 1685
rect 12035 1665 12065 1685
rect 12085 1665 12115 1685
rect 12135 1665 12165 1685
rect 12185 1665 12215 1685
rect 12235 1665 12265 1685
rect 12285 1665 12315 1685
rect 12335 1665 12365 1685
rect 12385 1665 12415 1685
rect 12435 1665 12465 1685
rect 12485 1665 12515 1685
rect 12535 1665 12565 1685
rect 12585 1665 12615 1685
rect 12635 1665 12665 1685
rect 12685 1665 12715 1685
rect 12735 1665 12765 1685
rect 12785 1665 12815 1685
rect 12835 1665 12865 1685
rect 12885 1665 12915 1685
rect 12935 1665 12965 1685
rect 12985 1665 13015 1685
rect 13035 1665 13065 1685
rect 13085 1665 13115 1685
rect 13135 1665 13165 1685
rect 13185 1665 13215 1685
rect 13235 1665 13265 1685
rect 13285 1665 13315 1685
rect 13335 1665 13365 1685
rect 13385 1665 13415 1685
rect 13435 1665 13465 1685
rect 13485 1665 13515 1685
rect 13535 1665 13565 1685
rect 13585 1665 13615 1685
rect 13635 1665 13665 1685
rect 13685 1665 13715 1685
rect 13735 1665 13765 1685
rect 13785 1665 13815 1685
rect 13835 1665 13865 1685
rect 13885 1665 13915 1685
rect 13935 1665 13965 1685
rect 13985 1665 14015 1685
rect 14035 1665 14065 1685
rect 14085 1665 14115 1685
rect 14135 1665 14165 1685
rect 14185 1665 14215 1685
rect 14235 1665 14265 1685
rect 14285 1665 14315 1685
rect 14335 1665 14365 1685
rect 14385 1665 14415 1685
rect 14435 1665 14465 1685
rect 14485 1665 14515 1685
rect 14535 1665 14565 1685
rect 14585 1665 14615 1685
rect 14635 1665 14665 1685
rect 14685 1665 14715 1685
rect 14735 1665 14765 1685
rect 14785 1665 14815 1685
rect 14835 1665 14865 1685
rect 14885 1665 14915 1685
rect 14935 1665 14965 1685
rect 14985 1665 15015 1685
rect 15035 1665 15065 1685
rect 15085 1665 15115 1685
rect 15135 1665 15165 1685
rect 15185 1665 15215 1685
rect 15235 1665 15265 1685
rect 15285 1665 15315 1685
rect 15335 1665 15365 1685
rect 15385 1665 15415 1685
rect 15435 1665 15465 1685
rect 15485 1665 15515 1685
rect 15535 1665 15565 1685
rect 15585 1665 15615 1685
rect 15635 1665 15665 1685
rect 15685 1665 15715 1685
rect 15735 1665 15765 1685
rect 15785 1665 15815 1685
rect 15835 1665 15865 1685
rect 15885 1665 15915 1685
rect 15935 1665 15965 1685
rect 15985 1665 16015 1685
rect 16035 1665 16065 1685
rect 16085 1665 16115 1685
rect 16135 1665 16165 1685
rect 16185 1665 16215 1685
rect 16235 1665 16265 1685
rect 16285 1665 16315 1685
rect 16335 1665 16365 1685
rect 16385 1665 16415 1685
rect 16435 1665 16465 1685
rect 16485 1665 16515 1685
rect 16535 1665 16565 1685
rect 16585 1665 16615 1685
rect 16635 1665 16665 1685
rect 16685 1665 16715 1685
rect 16735 1665 16765 1685
rect 16785 1665 16815 1685
rect 16835 1665 16865 1685
rect 16885 1665 16915 1685
rect 16935 1665 16965 1685
rect 16985 1665 17015 1685
rect 17035 1665 17065 1685
rect 17085 1665 17115 1685
rect 17135 1665 17165 1685
rect 17185 1665 17215 1685
rect 17235 1665 17265 1685
rect 17285 1665 17315 1685
rect 17335 1665 17365 1685
rect 17385 1665 17415 1685
rect 17435 1665 17465 1685
rect 17485 1665 17515 1685
rect 17535 1665 17565 1685
rect 17585 1665 17615 1685
rect 17635 1665 17665 1685
rect 17685 1665 17715 1685
rect 17735 1665 17765 1685
rect 17785 1665 17815 1685
rect 17835 1665 17865 1685
rect 17885 1665 17915 1685
rect 17935 1665 17965 1685
rect 17985 1665 18015 1685
rect 18035 1665 18065 1685
rect 18085 1665 18115 1685
rect 18135 1665 18165 1685
rect 18185 1665 18215 1685
rect 18235 1665 18265 1685
rect 18285 1665 18315 1685
rect 18335 1665 18365 1685
rect 18385 1665 18415 1685
rect 18435 1665 18465 1685
rect 18485 1665 18515 1685
rect 18535 1665 18565 1685
rect 18585 1665 18615 1685
rect 18635 1665 18665 1685
rect 18685 1665 18715 1685
rect 18735 1665 18765 1685
rect 18785 1665 18815 1685
rect 18835 1665 18865 1685
rect 18885 1665 18915 1685
rect 18935 1665 18965 1685
rect 18985 1665 19015 1685
rect 19035 1665 19065 1685
rect 19085 1665 19115 1685
rect 19135 1665 19165 1685
rect 19185 1665 19215 1685
rect 19235 1665 19265 1685
rect 19285 1665 19315 1685
rect 19335 1665 19365 1685
rect 19385 1665 19415 1685
rect 19435 1665 19465 1685
rect 19485 1665 19515 1685
rect 19535 1665 19565 1685
rect 19585 1665 19615 1685
rect 19635 1665 19665 1685
rect 19685 1665 19715 1685
rect 19735 1665 19765 1685
rect 19785 1665 19815 1685
rect 19835 1665 19865 1685
rect 19885 1665 19915 1685
rect 19935 1665 19965 1685
rect 19985 1665 20015 1685
rect 20035 1665 20065 1685
rect 20085 1665 20115 1685
rect 20135 1665 20165 1685
rect 20185 1665 20215 1685
rect 20235 1665 20265 1685
rect 20285 1665 20315 1685
rect 20335 1665 20365 1685
rect 20385 1665 20400 1685
rect -650 1650 20400 1665
rect -650 -15 20400 0
rect -650 -35 -635 -15
rect -615 -35 -585 -15
rect -565 -35 -535 -15
rect -515 -35 -485 -15
rect -465 -35 -435 -15
rect -415 -35 -385 -15
rect -365 -35 -335 -15
rect -315 -35 -285 -15
rect -265 -35 -235 -15
rect -215 -35 -185 -15
rect -165 -35 -135 -15
rect -115 -35 -85 -15
rect -65 -35 -35 -15
rect -15 -35 15 -15
rect 35 -35 65 -15
rect 85 -35 115 -15
rect 135 -35 165 -15
rect 185 -35 215 -15
rect 235 -35 265 -15
rect 285 -35 315 -15
rect 335 -35 365 -15
rect 385 -35 415 -15
rect 435 -35 465 -15
rect 485 -35 515 -15
rect 535 -35 565 -15
rect 585 -35 615 -15
rect 635 -35 665 -15
rect 685 -35 715 -15
rect 735 -35 765 -15
rect 785 -35 815 -15
rect 835 -35 865 -15
rect 885 -35 915 -15
rect 935 -35 965 -15
rect 985 -35 1015 -15
rect 1035 -35 1065 -15
rect 1085 -35 1115 -15
rect 1135 -35 1165 -15
rect 1185 -35 1215 -15
rect 1235 -35 1265 -15
rect 1285 -35 1315 -15
rect 1335 -35 1365 -15
rect 1385 -35 1415 -15
rect 1435 -35 1465 -15
rect 1485 -35 1515 -15
rect 1535 -35 1565 -15
rect 1585 -35 1615 -15
rect 1635 -35 1665 -15
rect 1685 -35 1715 -15
rect 1735 -35 1765 -15
rect 1785 -35 1815 -15
rect 1835 -35 1865 -15
rect 1885 -35 1915 -15
rect 1935 -35 1965 -15
rect 1985 -35 2015 -15
rect 2035 -35 2065 -15
rect 2085 -35 2115 -15
rect 2135 -35 2165 -15
rect 2185 -35 2215 -15
rect 2235 -35 2265 -15
rect 2285 -35 2315 -15
rect 2335 -35 2365 -15
rect 2385 -35 2415 -15
rect 2435 -35 2465 -15
rect 2485 -35 2515 -15
rect 2535 -35 2565 -15
rect 2585 -35 2615 -15
rect 2635 -35 2665 -15
rect 2685 -35 2715 -15
rect 2735 -35 2765 -15
rect 2785 -35 2815 -15
rect 2835 -35 2865 -15
rect 2885 -35 2915 -15
rect 2935 -35 2965 -15
rect 2985 -35 3015 -15
rect 3035 -35 3065 -15
rect 3085 -35 3115 -15
rect 3135 -35 3165 -15
rect 3185 -35 3215 -15
rect 3235 -35 3265 -15
rect 3285 -35 3315 -15
rect 3335 -35 3365 -15
rect 3385 -35 3415 -15
rect 3435 -35 3465 -15
rect 3485 -35 3515 -15
rect 3535 -35 3565 -15
rect 3585 -35 3615 -15
rect 3635 -35 3665 -15
rect 3685 -35 3715 -15
rect 3735 -35 3765 -15
rect 3785 -35 3815 -15
rect 3835 -35 3865 -15
rect 3885 -35 3915 -15
rect 3935 -35 3965 -15
rect 3985 -35 4015 -15
rect 4035 -35 4065 -15
rect 4085 -35 4115 -15
rect 4135 -35 4165 -15
rect 4185 -35 4215 -15
rect 4235 -35 4265 -15
rect 4285 -35 4315 -15
rect 4335 -35 4365 -15
rect 4385 -35 4415 -15
rect 4435 -35 4465 -15
rect 4485 -35 4515 -15
rect 4535 -35 4565 -15
rect 4585 -35 4615 -15
rect 4635 -35 4665 -15
rect 4685 -35 4715 -15
rect 4735 -35 4765 -15
rect 4785 -35 4815 -15
rect 4835 -35 4865 -15
rect 4885 -35 4915 -15
rect 4935 -35 4965 -15
rect 4985 -35 5015 -15
rect 5035 -35 5065 -15
rect 5085 -35 5115 -15
rect 5135 -35 5165 -15
rect 5185 -35 5215 -15
rect 5235 -35 5265 -15
rect 5285 -35 5315 -15
rect 5335 -35 5365 -15
rect 5385 -35 5415 -15
rect 5435 -35 5465 -15
rect 5485 -35 5515 -15
rect 5535 -35 5565 -15
rect 5585 -35 5615 -15
rect 5635 -35 5665 -15
rect 5685 -35 5715 -15
rect 5735 -35 5765 -15
rect 5785 -35 5815 -15
rect 5835 -35 5865 -15
rect 5885 -35 5915 -15
rect 5935 -35 5965 -15
rect 5985 -35 6015 -15
rect 6035 -35 6065 -15
rect 6085 -35 6115 -15
rect 6135 -35 6165 -15
rect 6185 -35 6215 -15
rect 6235 -35 6265 -15
rect 6285 -35 6315 -15
rect 6335 -35 6365 -15
rect 6385 -35 6415 -15
rect 6435 -35 6465 -15
rect 6485 -35 6515 -15
rect 6535 -35 6565 -15
rect 6585 -35 6615 -15
rect 6635 -35 6665 -15
rect 6685 -35 6715 -15
rect 6735 -35 6765 -15
rect 6785 -35 6815 -15
rect 6835 -35 6865 -15
rect 6885 -35 6915 -15
rect 6935 -35 6965 -15
rect 6985 -35 7015 -15
rect 7035 -35 7065 -15
rect 7085 -35 7115 -15
rect 7135 -35 7165 -15
rect 7185 -35 7215 -15
rect 7235 -35 7265 -15
rect 7285 -35 7315 -15
rect 7335 -35 7365 -15
rect 7385 -35 7415 -15
rect 7435 -35 7465 -15
rect 7485 -35 7515 -15
rect 7535 -35 7565 -15
rect 7585 -35 7615 -15
rect 7635 -35 7665 -15
rect 7685 -35 7715 -15
rect 7735 -35 7765 -15
rect 7785 -35 7815 -15
rect 7835 -35 7865 -15
rect 7885 -35 7915 -15
rect 7935 -35 7965 -15
rect 7985 -35 8015 -15
rect 8035 -35 8065 -15
rect 8085 -35 8115 -15
rect 8135 -35 8165 -15
rect 8185 -35 8215 -15
rect 8235 -35 8265 -15
rect 8285 -35 8315 -15
rect 8335 -35 8365 -15
rect 8385 -35 8415 -15
rect 8435 -35 8465 -15
rect 8485 -35 8515 -15
rect 8535 -35 8565 -15
rect 8585 -35 8615 -15
rect 8635 -35 8665 -15
rect 8685 -35 8715 -15
rect 8735 -35 8765 -15
rect 8785 -35 8815 -15
rect 8835 -35 8865 -15
rect 8885 -35 8915 -15
rect 8935 -35 8965 -15
rect 8985 -35 9015 -15
rect 9035 -35 9065 -15
rect 9085 -35 9115 -15
rect 9135 -35 9165 -15
rect 9185 -35 9215 -15
rect 9235 -35 9265 -15
rect 9285 -35 9315 -15
rect 9335 -35 9365 -15
rect 9385 -35 9415 -15
rect 9435 -35 9465 -15
rect 9485 -35 9515 -15
rect 9535 -35 9565 -15
rect 9585 -35 9615 -15
rect 9635 -35 9665 -15
rect 9685 -35 9715 -15
rect 9735 -35 9765 -15
rect 9785 -35 9815 -15
rect 9835 -35 9865 -15
rect 9885 -35 9915 -15
rect 9935 -35 9965 -15
rect 9985 -35 10015 -15
rect 10035 -35 10065 -15
rect 10085 -35 10115 -15
rect 10135 -35 10165 -15
rect 10185 -35 10215 -15
rect 10235 -35 10265 -15
rect 10285 -35 10315 -15
rect 10335 -35 10365 -15
rect 10385 -35 10415 -15
rect 10435 -35 10465 -15
rect 10485 -35 10515 -15
rect 10535 -35 10565 -15
rect 10585 -35 10615 -15
rect 10635 -35 10665 -15
rect 10685 -35 10715 -15
rect 10735 -35 10765 -15
rect 10785 -35 10815 -15
rect 10835 -35 10865 -15
rect 10885 -35 10915 -15
rect 10935 -35 10965 -15
rect 10985 -35 11015 -15
rect 11035 -35 11065 -15
rect 11085 -35 11115 -15
rect 11135 -35 11165 -15
rect 11185 -35 11215 -15
rect 11235 -35 11265 -15
rect 11285 -35 11315 -15
rect 11335 -35 11365 -15
rect 11385 -35 11415 -15
rect 11435 -35 11465 -15
rect 11485 -35 11515 -15
rect 11535 -35 11565 -15
rect 11585 -35 11615 -15
rect 11635 -35 11665 -15
rect 11685 -35 11715 -15
rect 11735 -35 11765 -15
rect 11785 -35 11815 -15
rect 11835 -35 11865 -15
rect 11885 -35 11915 -15
rect 11935 -35 11965 -15
rect 11985 -35 12015 -15
rect 12035 -35 12065 -15
rect 12085 -35 12115 -15
rect 12135 -35 12165 -15
rect 12185 -35 12215 -15
rect 12235 -35 12265 -15
rect 12285 -35 12315 -15
rect 12335 -35 12365 -15
rect 12385 -35 12415 -15
rect 12435 -35 12465 -15
rect 12485 -35 12515 -15
rect 12535 -35 12565 -15
rect 12585 -35 12615 -15
rect 12635 -35 12665 -15
rect 12685 -35 12715 -15
rect 12735 -35 12765 -15
rect 12785 -35 12815 -15
rect 12835 -35 12865 -15
rect 12885 -35 12915 -15
rect 12935 -35 12965 -15
rect 12985 -35 13015 -15
rect 13035 -35 13065 -15
rect 13085 -35 13115 -15
rect 13135 -35 13165 -15
rect 13185 -35 13215 -15
rect 13235 -35 13265 -15
rect 13285 -35 13315 -15
rect 13335 -35 13365 -15
rect 13385 -35 13415 -15
rect 13435 -35 13465 -15
rect 13485 -35 13515 -15
rect 13535 -35 13565 -15
rect 13585 -35 13615 -15
rect 13635 -35 13665 -15
rect 13685 -35 13715 -15
rect 13735 -35 13765 -15
rect 13785 -35 13815 -15
rect 13835 -35 13865 -15
rect 13885 -35 13915 -15
rect 13935 -35 13965 -15
rect 13985 -35 14015 -15
rect 14035 -35 14065 -15
rect 14085 -35 14115 -15
rect 14135 -35 14165 -15
rect 14185 -35 14215 -15
rect 14235 -35 14265 -15
rect 14285 -35 14315 -15
rect 14335 -35 14365 -15
rect 14385 -35 14415 -15
rect 14435 -35 14465 -15
rect 14485 -35 14515 -15
rect 14535 -35 14565 -15
rect 14585 -35 14615 -15
rect 14635 -35 14665 -15
rect 14685 -35 14715 -15
rect 14735 -35 14765 -15
rect 14785 -35 14815 -15
rect 14835 -35 14865 -15
rect 14885 -35 14915 -15
rect 14935 -35 14965 -15
rect 14985 -35 15015 -15
rect 15035 -35 15065 -15
rect 15085 -35 15115 -15
rect 15135 -35 15165 -15
rect 15185 -35 15215 -15
rect 15235 -35 15265 -15
rect 15285 -35 15315 -15
rect 15335 -35 15365 -15
rect 15385 -35 15415 -15
rect 15435 -35 15465 -15
rect 15485 -35 15515 -15
rect 15535 -35 15565 -15
rect 15585 -35 15615 -15
rect 15635 -35 15665 -15
rect 15685 -35 15715 -15
rect 15735 -35 15765 -15
rect 15785 -35 15815 -15
rect 15835 -35 15865 -15
rect 15885 -35 15915 -15
rect 15935 -35 15965 -15
rect 15985 -35 16015 -15
rect 16035 -35 16065 -15
rect 16085 -35 16115 -15
rect 16135 -35 16165 -15
rect 16185 -35 16215 -15
rect 16235 -35 16265 -15
rect 16285 -35 16315 -15
rect 16335 -35 16365 -15
rect 16385 -35 16415 -15
rect 16435 -35 16465 -15
rect 16485 -35 16515 -15
rect 16535 -35 16565 -15
rect 16585 -35 16615 -15
rect 16635 -35 16665 -15
rect 16685 -35 16715 -15
rect 16735 -35 16765 -15
rect 16785 -35 16815 -15
rect 16835 -35 16865 -15
rect 16885 -35 16915 -15
rect 16935 -35 16965 -15
rect 16985 -35 17015 -15
rect 17035 -35 17065 -15
rect 17085 -35 17115 -15
rect 17135 -35 17165 -15
rect 17185 -35 17215 -15
rect 17235 -35 17265 -15
rect 17285 -35 17315 -15
rect 17335 -35 17365 -15
rect 17385 -35 17415 -15
rect 17435 -35 17465 -15
rect 17485 -35 17515 -15
rect 17535 -35 17565 -15
rect 17585 -35 17615 -15
rect 17635 -35 17665 -15
rect 17685 -35 17715 -15
rect 17735 -35 17765 -15
rect 17785 -35 17815 -15
rect 17835 -35 17865 -15
rect 17885 -35 17915 -15
rect 17935 -35 17965 -15
rect 17985 -35 18015 -15
rect 18035 -35 18065 -15
rect 18085 -35 18115 -15
rect 18135 -35 18165 -15
rect 18185 -35 18215 -15
rect 18235 -35 18265 -15
rect 18285 -35 18315 -15
rect 18335 -35 18365 -15
rect 18385 -35 18415 -15
rect 18435 -35 18465 -15
rect 18485 -35 18515 -15
rect 18535 -35 18565 -15
rect 18585 -35 18615 -15
rect 18635 -35 18665 -15
rect 18685 -35 18715 -15
rect 18735 -35 18765 -15
rect 18785 -35 18815 -15
rect 18835 -35 18865 -15
rect 18885 -35 18915 -15
rect 18935 -35 18965 -15
rect 18985 -35 19015 -15
rect 19035 -35 19065 -15
rect 19085 -35 19115 -15
rect 19135 -35 19165 -15
rect 19185 -35 19215 -15
rect 19235 -35 19265 -15
rect 19285 -35 19315 -15
rect 19335 -35 19365 -15
rect 19385 -35 19415 -15
rect 19435 -35 19465 -15
rect 19485 -35 19515 -15
rect 19535 -35 19565 -15
rect 19585 -35 19615 -15
rect 19635 -35 19665 -15
rect 19685 -35 19715 -15
rect 19735 -35 19765 -15
rect 19785 -35 19815 -15
rect 19835 -35 19865 -15
rect 19885 -35 19915 -15
rect 19935 -35 19965 -15
rect 19985 -35 20015 -15
rect 20035 -35 20065 -15
rect 20085 -35 20115 -15
rect 20135 -35 20165 -15
rect 20185 -35 20215 -15
rect 20235 -35 20265 -15
rect 20285 -35 20315 -15
rect 20335 -35 20365 -15
rect 20385 -35 20400 -15
rect -650 -50 20400 -35
rect -650 -1715 20400 -1700
rect -650 -1735 -635 -1715
rect -615 -1735 -585 -1715
rect -565 -1735 -535 -1715
rect -515 -1735 -485 -1715
rect -465 -1735 -435 -1715
rect -415 -1735 -385 -1715
rect -365 -1735 -335 -1715
rect -315 -1735 -285 -1715
rect -265 -1735 -235 -1715
rect -215 -1735 -185 -1715
rect -165 -1735 -135 -1715
rect -115 -1735 -85 -1715
rect -65 -1735 -35 -1715
rect -15 -1735 15 -1715
rect 35 -1735 65 -1715
rect 85 -1735 115 -1715
rect 135 -1735 165 -1715
rect 185 -1735 215 -1715
rect 235 -1735 265 -1715
rect 285 -1735 315 -1715
rect 335 -1735 365 -1715
rect 385 -1735 415 -1715
rect 435 -1735 465 -1715
rect 485 -1735 515 -1715
rect 535 -1735 565 -1715
rect 585 -1735 615 -1715
rect 635 -1735 665 -1715
rect 685 -1735 715 -1715
rect 735 -1735 765 -1715
rect 785 -1735 815 -1715
rect 835 -1735 865 -1715
rect 885 -1735 915 -1715
rect 935 -1735 965 -1715
rect 985 -1735 1015 -1715
rect 1035 -1735 1065 -1715
rect 1085 -1735 1115 -1715
rect 1135 -1735 1165 -1715
rect 1185 -1735 1215 -1715
rect 1235 -1735 1265 -1715
rect 1285 -1735 1315 -1715
rect 1335 -1735 1365 -1715
rect 1385 -1735 1415 -1715
rect 1435 -1735 1465 -1715
rect 1485 -1735 1515 -1715
rect 1535 -1735 1565 -1715
rect 1585 -1735 1615 -1715
rect 1635 -1735 1665 -1715
rect 1685 -1735 1715 -1715
rect 1735 -1735 1765 -1715
rect 1785 -1735 1815 -1715
rect 1835 -1735 1865 -1715
rect 1885 -1735 1915 -1715
rect 1935 -1735 1965 -1715
rect 1985 -1735 2015 -1715
rect 2035 -1735 2065 -1715
rect 2085 -1735 2115 -1715
rect 2135 -1735 2165 -1715
rect 2185 -1735 2215 -1715
rect 2235 -1735 2265 -1715
rect 2285 -1735 2315 -1715
rect 2335 -1735 2365 -1715
rect 2385 -1735 2415 -1715
rect 2435 -1735 2465 -1715
rect 2485 -1735 2515 -1715
rect 2535 -1735 2565 -1715
rect 2585 -1735 2615 -1715
rect 2635 -1735 2665 -1715
rect 2685 -1735 2715 -1715
rect 2735 -1735 2765 -1715
rect 2785 -1735 2815 -1715
rect 2835 -1735 2865 -1715
rect 2885 -1735 2915 -1715
rect 2935 -1735 2965 -1715
rect 2985 -1735 3015 -1715
rect 3035 -1735 3065 -1715
rect 3085 -1735 3115 -1715
rect 3135 -1735 3165 -1715
rect 3185 -1735 3215 -1715
rect 3235 -1735 3265 -1715
rect 3285 -1735 3315 -1715
rect 3335 -1735 3365 -1715
rect 3385 -1735 3415 -1715
rect 3435 -1735 3465 -1715
rect 3485 -1735 3515 -1715
rect 3535 -1735 3565 -1715
rect 3585 -1735 3615 -1715
rect 3635 -1735 3665 -1715
rect 3685 -1735 3715 -1715
rect 3735 -1735 3765 -1715
rect 3785 -1735 3815 -1715
rect 3835 -1735 3865 -1715
rect 3885 -1735 3915 -1715
rect 3935 -1735 3965 -1715
rect 3985 -1735 4015 -1715
rect 4035 -1735 4065 -1715
rect 4085 -1735 4115 -1715
rect 4135 -1735 4165 -1715
rect 4185 -1735 4215 -1715
rect 4235 -1735 4265 -1715
rect 4285 -1735 4315 -1715
rect 4335 -1735 4365 -1715
rect 4385 -1735 4415 -1715
rect 4435 -1735 4465 -1715
rect 4485 -1735 4515 -1715
rect 4535 -1735 4565 -1715
rect 4585 -1735 4615 -1715
rect 4635 -1735 4665 -1715
rect 4685 -1735 4715 -1715
rect 4735 -1735 4765 -1715
rect 4785 -1735 4815 -1715
rect 4835 -1735 4865 -1715
rect 4885 -1735 4915 -1715
rect 4935 -1735 4965 -1715
rect 4985 -1735 5015 -1715
rect 5035 -1735 5065 -1715
rect 5085 -1735 5115 -1715
rect 5135 -1735 5165 -1715
rect 5185 -1735 5215 -1715
rect 5235 -1735 5265 -1715
rect 5285 -1735 5315 -1715
rect 5335 -1735 5365 -1715
rect 5385 -1735 5415 -1715
rect 5435 -1735 5465 -1715
rect 5485 -1735 5515 -1715
rect 5535 -1735 5565 -1715
rect 5585 -1735 5615 -1715
rect 5635 -1735 5665 -1715
rect 5685 -1735 5715 -1715
rect 5735 -1735 5765 -1715
rect 5785 -1735 5815 -1715
rect 5835 -1735 5865 -1715
rect 5885 -1735 5915 -1715
rect 5935 -1735 5965 -1715
rect 5985 -1735 6015 -1715
rect 6035 -1735 6065 -1715
rect 6085 -1735 6115 -1715
rect 6135 -1735 6165 -1715
rect 6185 -1735 6215 -1715
rect 6235 -1735 6265 -1715
rect 6285 -1735 6315 -1715
rect 6335 -1735 6365 -1715
rect 6385 -1735 6415 -1715
rect 6435 -1735 6465 -1715
rect 6485 -1735 6515 -1715
rect 6535 -1735 6565 -1715
rect 6585 -1735 6615 -1715
rect 6635 -1735 6665 -1715
rect 6685 -1735 6715 -1715
rect 6735 -1735 6765 -1715
rect 6785 -1735 6815 -1715
rect 6835 -1735 6865 -1715
rect 6885 -1735 6915 -1715
rect 6935 -1735 6965 -1715
rect 6985 -1735 7015 -1715
rect 7035 -1735 7065 -1715
rect 7085 -1735 7115 -1715
rect 7135 -1735 7165 -1715
rect 7185 -1735 7215 -1715
rect 7235 -1735 7265 -1715
rect 7285 -1735 7315 -1715
rect 7335 -1735 7365 -1715
rect 7385 -1735 7415 -1715
rect 7435 -1735 7465 -1715
rect 7485 -1735 7515 -1715
rect 7535 -1735 7565 -1715
rect 7585 -1735 7615 -1715
rect 7635 -1735 7665 -1715
rect 7685 -1735 7715 -1715
rect 7735 -1735 7765 -1715
rect 7785 -1735 7815 -1715
rect 7835 -1735 7865 -1715
rect 7885 -1735 7915 -1715
rect 7935 -1735 7965 -1715
rect 7985 -1735 8015 -1715
rect 8035 -1735 8065 -1715
rect 8085 -1735 8115 -1715
rect 8135 -1735 8165 -1715
rect 8185 -1735 8215 -1715
rect 8235 -1735 8265 -1715
rect 8285 -1735 8315 -1715
rect 8335 -1735 8365 -1715
rect 8385 -1735 8415 -1715
rect 8435 -1735 8465 -1715
rect 8485 -1735 8515 -1715
rect 8535 -1735 8565 -1715
rect 8585 -1735 8615 -1715
rect 8635 -1735 8665 -1715
rect 8685 -1735 8715 -1715
rect 8735 -1735 8765 -1715
rect 8785 -1735 8815 -1715
rect 8835 -1735 8865 -1715
rect 8885 -1735 8915 -1715
rect 8935 -1735 8965 -1715
rect 8985 -1735 9015 -1715
rect 9035 -1735 9065 -1715
rect 9085 -1735 9115 -1715
rect 9135 -1735 9165 -1715
rect 9185 -1735 9215 -1715
rect 9235 -1735 9265 -1715
rect 9285 -1735 9315 -1715
rect 9335 -1735 9365 -1715
rect 9385 -1735 9415 -1715
rect 9435 -1735 9465 -1715
rect 9485 -1735 9515 -1715
rect 9535 -1735 9565 -1715
rect 9585 -1735 9615 -1715
rect 9635 -1735 9665 -1715
rect 9685 -1735 9715 -1715
rect 9735 -1735 9765 -1715
rect 9785 -1735 9815 -1715
rect 9835 -1735 9865 -1715
rect 9885 -1735 9915 -1715
rect 9935 -1735 9965 -1715
rect 9985 -1735 10015 -1715
rect 10035 -1735 10065 -1715
rect 10085 -1735 10115 -1715
rect 10135 -1735 10165 -1715
rect 10185 -1735 10215 -1715
rect 10235 -1735 10265 -1715
rect 10285 -1735 10315 -1715
rect 10335 -1735 10365 -1715
rect 10385 -1735 10415 -1715
rect 10435 -1735 10465 -1715
rect 10485 -1735 10515 -1715
rect 10535 -1735 10565 -1715
rect 10585 -1735 10615 -1715
rect 10635 -1735 10665 -1715
rect 10685 -1735 10715 -1715
rect 10735 -1735 10765 -1715
rect 10785 -1735 10815 -1715
rect 10835 -1735 10865 -1715
rect 10885 -1735 10915 -1715
rect 10935 -1735 10965 -1715
rect 10985 -1735 11015 -1715
rect 11035 -1735 11065 -1715
rect 11085 -1735 11115 -1715
rect 11135 -1735 11165 -1715
rect 11185 -1735 11215 -1715
rect 11235 -1735 11265 -1715
rect 11285 -1735 11315 -1715
rect 11335 -1735 11365 -1715
rect 11385 -1735 11415 -1715
rect 11435 -1735 11465 -1715
rect 11485 -1735 11515 -1715
rect 11535 -1735 11565 -1715
rect 11585 -1735 11615 -1715
rect 11635 -1735 11665 -1715
rect 11685 -1735 11715 -1715
rect 11735 -1735 11765 -1715
rect 11785 -1735 11815 -1715
rect 11835 -1735 11865 -1715
rect 11885 -1735 11915 -1715
rect 11935 -1735 11965 -1715
rect 11985 -1735 12015 -1715
rect 12035 -1735 12065 -1715
rect 12085 -1735 12115 -1715
rect 12135 -1735 12165 -1715
rect 12185 -1735 12215 -1715
rect 12235 -1735 12265 -1715
rect 12285 -1735 12315 -1715
rect 12335 -1735 12365 -1715
rect 12385 -1735 12415 -1715
rect 12435 -1735 12465 -1715
rect 12485 -1735 12515 -1715
rect 12535 -1735 12565 -1715
rect 12585 -1735 12615 -1715
rect 12635 -1735 12665 -1715
rect 12685 -1735 12715 -1715
rect 12735 -1735 12765 -1715
rect 12785 -1735 12815 -1715
rect 12835 -1735 12865 -1715
rect 12885 -1735 12915 -1715
rect 12935 -1735 12965 -1715
rect 12985 -1735 13015 -1715
rect 13035 -1735 13065 -1715
rect 13085 -1735 13115 -1715
rect 13135 -1735 13165 -1715
rect 13185 -1735 13215 -1715
rect 13235 -1735 13265 -1715
rect 13285 -1735 13315 -1715
rect 13335 -1735 13365 -1715
rect 13385 -1735 13415 -1715
rect 13435 -1735 13465 -1715
rect 13485 -1735 13515 -1715
rect 13535 -1735 13565 -1715
rect 13585 -1735 13615 -1715
rect 13635 -1735 13665 -1715
rect 13685 -1735 13715 -1715
rect 13735 -1735 13765 -1715
rect 13785 -1735 13815 -1715
rect 13835 -1735 13865 -1715
rect 13885 -1735 13915 -1715
rect 13935 -1735 13965 -1715
rect 13985 -1735 14015 -1715
rect 14035 -1735 14065 -1715
rect 14085 -1735 14115 -1715
rect 14135 -1735 14165 -1715
rect 14185 -1735 14215 -1715
rect 14235 -1735 14265 -1715
rect 14285 -1735 14315 -1715
rect 14335 -1735 14365 -1715
rect 14385 -1735 14415 -1715
rect 14435 -1735 14465 -1715
rect 14485 -1735 14515 -1715
rect 14535 -1735 14565 -1715
rect 14585 -1735 14615 -1715
rect 14635 -1735 14665 -1715
rect 14685 -1735 14715 -1715
rect 14735 -1735 14765 -1715
rect 14785 -1735 14815 -1715
rect 14835 -1735 14865 -1715
rect 14885 -1735 14915 -1715
rect 14935 -1735 14965 -1715
rect 14985 -1735 15015 -1715
rect 15035 -1735 15065 -1715
rect 15085 -1735 15115 -1715
rect 15135 -1735 15165 -1715
rect 15185 -1735 15215 -1715
rect 15235 -1735 15265 -1715
rect 15285 -1735 15315 -1715
rect 15335 -1735 15365 -1715
rect 15385 -1735 15415 -1715
rect 15435 -1735 15465 -1715
rect 15485 -1735 15515 -1715
rect 15535 -1735 15565 -1715
rect 15585 -1735 15615 -1715
rect 15635 -1735 15665 -1715
rect 15685 -1735 15715 -1715
rect 15735 -1735 15765 -1715
rect 15785 -1735 15815 -1715
rect 15835 -1735 15865 -1715
rect 15885 -1735 15915 -1715
rect 15935 -1735 15965 -1715
rect 15985 -1735 16015 -1715
rect 16035 -1735 16065 -1715
rect 16085 -1735 16115 -1715
rect 16135 -1735 16165 -1715
rect 16185 -1735 16215 -1715
rect 16235 -1735 16265 -1715
rect 16285 -1735 16315 -1715
rect 16335 -1735 16365 -1715
rect 16385 -1735 16415 -1715
rect 16435 -1735 16465 -1715
rect 16485 -1735 16515 -1715
rect 16535 -1735 16565 -1715
rect 16585 -1735 16615 -1715
rect 16635 -1735 16665 -1715
rect 16685 -1735 16715 -1715
rect 16735 -1735 16765 -1715
rect 16785 -1735 16815 -1715
rect 16835 -1735 16865 -1715
rect 16885 -1735 16915 -1715
rect 16935 -1735 16965 -1715
rect 16985 -1735 17015 -1715
rect 17035 -1735 17065 -1715
rect 17085 -1735 17115 -1715
rect 17135 -1735 17165 -1715
rect 17185 -1735 17215 -1715
rect 17235 -1735 17265 -1715
rect 17285 -1735 17315 -1715
rect 17335 -1735 17365 -1715
rect 17385 -1735 17415 -1715
rect 17435 -1735 17465 -1715
rect 17485 -1735 17515 -1715
rect 17535 -1735 17565 -1715
rect 17585 -1735 17615 -1715
rect 17635 -1735 17665 -1715
rect 17685 -1735 17715 -1715
rect 17735 -1735 17765 -1715
rect 17785 -1735 17815 -1715
rect 17835 -1735 17865 -1715
rect 17885 -1735 17915 -1715
rect 17935 -1735 17965 -1715
rect 17985 -1735 18015 -1715
rect 18035 -1735 18065 -1715
rect 18085 -1735 18115 -1715
rect 18135 -1735 18165 -1715
rect 18185 -1735 18215 -1715
rect 18235 -1735 18265 -1715
rect 18285 -1735 18315 -1715
rect 18335 -1735 18365 -1715
rect 18385 -1735 18415 -1715
rect 18435 -1735 18465 -1715
rect 18485 -1735 18515 -1715
rect 18535 -1735 18565 -1715
rect 18585 -1735 18615 -1715
rect 18635 -1735 18665 -1715
rect 18685 -1735 18715 -1715
rect 18735 -1735 18765 -1715
rect 18785 -1735 18815 -1715
rect 18835 -1735 18865 -1715
rect 18885 -1735 18915 -1715
rect 18935 -1735 18965 -1715
rect 18985 -1735 19015 -1715
rect 19035 -1735 19065 -1715
rect 19085 -1735 19115 -1715
rect 19135 -1735 19165 -1715
rect 19185 -1735 19215 -1715
rect 19235 -1735 19265 -1715
rect 19285 -1735 19315 -1715
rect 19335 -1735 19365 -1715
rect 19385 -1735 19415 -1715
rect 19435 -1735 19465 -1715
rect 19485 -1735 19515 -1715
rect 19535 -1735 19565 -1715
rect 19585 -1735 19615 -1715
rect 19635 -1735 19665 -1715
rect 19685 -1735 19715 -1715
rect 19735 -1735 19765 -1715
rect 19785 -1735 19815 -1715
rect 19835 -1735 19865 -1715
rect 19885 -1735 19915 -1715
rect 19935 -1735 19965 -1715
rect 19985 -1735 20015 -1715
rect 20035 -1735 20065 -1715
rect 20085 -1735 20115 -1715
rect 20135 -1735 20165 -1715
rect 20185 -1735 20215 -1715
rect 20235 -1735 20265 -1715
rect 20285 -1735 20315 -1715
rect 20335 -1735 20365 -1715
rect 20385 -1735 20400 -1715
rect -650 -1750 20400 -1735
<< mvnsubdiff >>
rect -650 5185 20400 5200
rect -650 5165 -635 5185
rect -615 5165 -585 5185
rect -565 5165 -535 5185
rect -515 5165 -485 5185
rect -465 5165 -435 5185
rect -415 5165 -385 5185
rect -365 5165 -335 5185
rect -315 5165 -285 5185
rect -265 5165 -235 5185
rect -215 5165 -185 5185
rect -165 5165 -135 5185
rect -115 5165 -85 5185
rect -65 5165 -35 5185
rect -15 5165 15 5185
rect 35 5165 65 5185
rect 85 5165 115 5185
rect 135 5165 165 5185
rect 185 5165 215 5185
rect 235 5165 265 5185
rect 285 5165 315 5185
rect 335 5165 365 5185
rect 385 5165 415 5185
rect 435 5165 465 5185
rect 485 5165 515 5185
rect 535 5165 565 5185
rect 585 5165 615 5185
rect 635 5165 665 5185
rect 685 5165 715 5185
rect 735 5165 765 5185
rect 785 5165 815 5185
rect 835 5165 865 5185
rect 885 5165 915 5185
rect 935 5165 965 5185
rect 985 5165 1015 5185
rect 1035 5165 1065 5185
rect 1085 5165 1115 5185
rect 1135 5165 1165 5185
rect 1185 5165 1215 5185
rect 1235 5165 1265 5185
rect 1285 5165 1315 5185
rect 1335 5165 1365 5185
rect 1385 5165 1415 5185
rect 1435 5165 1465 5185
rect 1485 5165 1515 5185
rect 1535 5165 1565 5185
rect 1585 5165 1615 5185
rect 1635 5165 1665 5185
rect 1685 5165 1715 5185
rect 1735 5165 1765 5185
rect 1785 5165 1815 5185
rect 1835 5165 1865 5185
rect 1885 5165 1915 5185
rect 1935 5165 1965 5185
rect 1985 5165 2015 5185
rect 2035 5165 2065 5185
rect 2085 5165 2115 5185
rect 2135 5165 2165 5185
rect 2185 5165 2215 5185
rect 2235 5165 2265 5185
rect 2285 5165 2315 5185
rect 2335 5165 2365 5185
rect 2385 5165 2415 5185
rect 2435 5165 2465 5185
rect 2485 5165 2515 5185
rect 2535 5165 2565 5185
rect 2585 5165 2615 5185
rect 2635 5165 2665 5185
rect 2685 5165 2715 5185
rect 2735 5165 2765 5185
rect 2785 5165 2815 5185
rect 2835 5165 2865 5185
rect 2885 5165 2915 5185
rect 2935 5165 2965 5185
rect 2985 5165 3015 5185
rect 3035 5165 3065 5185
rect 3085 5165 3115 5185
rect 3135 5165 3165 5185
rect 3185 5165 3215 5185
rect 3235 5165 3265 5185
rect 3285 5165 3315 5185
rect 3335 5165 3365 5185
rect 3385 5165 3415 5185
rect 3435 5165 3465 5185
rect 3485 5165 3515 5185
rect 3535 5165 3565 5185
rect 3585 5165 3615 5185
rect 3635 5165 3665 5185
rect 3685 5165 3715 5185
rect 3735 5165 3765 5185
rect 3785 5165 3815 5185
rect 3835 5165 3865 5185
rect 3885 5165 3915 5185
rect 3935 5165 3965 5185
rect 3985 5165 4015 5185
rect 4035 5165 4065 5185
rect 4085 5165 4115 5185
rect 4135 5165 4165 5185
rect 4185 5165 4215 5185
rect 4235 5165 4265 5185
rect 4285 5165 4315 5185
rect 4335 5165 4365 5185
rect 4385 5165 4415 5185
rect 4435 5165 4465 5185
rect 4485 5165 4515 5185
rect 4535 5165 4565 5185
rect 4585 5165 4615 5185
rect 4635 5165 4665 5185
rect 4685 5165 4715 5185
rect 4735 5165 4765 5185
rect 4785 5165 4815 5185
rect 4835 5165 4865 5185
rect 4885 5165 4915 5185
rect 4935 5165 4965 5185
rect 4985 5165 5015 5185
rect 5035 5165 5065 5185
rect 5085 5165 5115 5185
rect 5135 5165 5165 5185
rect 5185 5165 5215 5185
rect 5235 5165 5265 5185
rect 5285 5165 5315 5185
rect 5335 5165 5365 5185
rect 5385 5165 5415 5185
rect 5435 5165 5465 5185
rect 5485 5165 5515 5185
rect 5535 5165 5565 5185
rect 5585 5165 5615 5185
rect 5635 5165 5665 5185
rect 5685 5165 5715 5185
rect 5735 5165 5765 5185
rect 5785 5165 5815 5185
rect 5835 5165 5865 5185
rect 5885 5165 5915 5185
rect 5935 5165 5965 5185
rect 5985 5165 6015 5185
rect 6035 5165 6065 5185
rect 6085 5165 6115 5185
rect 6135 5165 6165 5185
rect 6185 5165 6215 5185
rect 6235 5165 6265 5185
rect 6285 5165 6315 5185
rect 6335 5165 6365 5185
rect 6385 5165 6415 5185
rect 6435 5165 6465 5185
rect 6485 5165 6515 5185
rect 6535 5165 6565 5185
rect 6585 5165 6615 5185
rect 6635 5165 6665 5185
rect 6685 5165 6715 5185
rect 6735 5165 6765 5185
rect 6785 5165 6815 5185
rect 6835 5165 6865 5185
rect 6885 5165 6915 5185
rect 6935 5165 6965 5185
rect 6985 5165 7015 5185
rect 7035 5165 7065 5185
rect 7085 5165 7115 5185
rect 7135 5165 7165 5185
rect 7185 5165 7215 5185
rect 7235 5165 7265 5185
rect 7285 5165 7315 5185
rect 7335 5165 7365 5185
rect 7385 5165 7415 5185
rect 7435 5165 7465 5185
rect 7485 5165 7515 5185
rect 7535 5165 7565 5185
rect 7585 5165 7615 5185
rect 7635 5165 7665 5185
rect 7685 5165 7715 5185
rect 7735 5165 7765 5185
rect 7785 5165 7815 5185
rect 7835 5165 7865 5185
rect 7885 5165 7915 5185
rect 7935 5165 7965 5185
rect 7985 5165 8015 5185
rect 8035 5165 8065 5185
rect 8085 5165 8115 5185
rect 8135 5165 8165 5185
rect 8185 5165 8215 5185
rect 8235 5165 8265 5185
rect 8285 5165 8315 5185
rect 8335 5165 8365 5185
rect 8385 5165 8415 5185
rect 8435 5165 8465 5185
rect 8485 5165 8515 5185
rect 8535 5165 8565 5185
rect 8585 5165 8615 5185
rect 8635 5165 8665 5185
rect 8685 5165 8715 5185
rect 8735 5165 8765 5185
rect 8785 5165 8815 5185
rect 8835 5165 8865 5185
rect 8885 5165 8915 5185
rect 8935 5165 8965 5185
rect 8985 5165 9015 5185
rect 9035 5165 9065 5185
rect 9085 5165 9115 5185
rect 9135 5165 9165 5185
rect 9185 5165 9215 5185
rect 9235 5165 9265 5185
rect 9285 5165 9315 5185
rect 9335 5165 9365 5185
rect 9385 5165 9415 5185
rect 9435 5165 9465 5185
rect 9485 5165 9515 5185
rect 9535 5165 9565 5185
rect 9585 5165 9615 5185
rect 9635 5165 9665 5185
rect 9685 5165 9715 5185
rect 9735 5165 9765 5185
rect 9785 5165 9815 5185
rect 9835 5165 9865 5185
rect 9885 5165 9915 5185
rect 9935 5165 9965 5185
rect 9985 5165 10015 5185
rect 10035 5165 10065 5185
rect 10085 5165 10115 5185
rect 10135 5165 10165 5185
rect 10185 5165 10215 5185
rect 10235 5165 10265 5185
rect 10285 5165 10315 5185
rect 10335 5165 10365 5185
rect 10385 5165 10415 5185
rect 10435 5165 10465 5185
rect 10485 5165 10515 5185
rect 10535 5165 10565 5185
rect 10585 5165 10615 5185
rect 10635 5165 10665 5185
rect 10685 5165 10715 5185
rect 10735 5165 10765 5185
rect 10785 5165 10815 5185
rect 10835 5165 10865 5185
rect 10885 5165 10915 5185
rect 10935 5165 10965 5185
rect 10985 5165 11015 5185
rect 11035 5165 11065 5185
rect 11085 5165 11115 5185
rect 11135 5165 11165 5185
rect 11185 5165 11215 5185
rect 11235 5165 11265 5185
rect 11285 5165 11315 5185
rect 11335 5165 11365 5185
rect 11385 5165 11415 5185
rect 11435 5165 11465 5185
rect 11485 5165 11515 5185
rect 11535 5165 11565 5185
rect 11585 5165 11615 5185
rect 11635 5165 11665 5185
rect 11685 5165 11715 5185
rect 11735 5165 11765 5185
rect 11785 5165 11815 5185
rect 11835 5165 11865 5185
rect 11885 5165 11915 5185
rect 11935 5165 11965 5185
rect 11985 5165 12015 5185
rect 12035 5165 12065 5185
rect 12085 5165 12115 5185
rect 12135 5165 12165 5185
rect 12185 5165 12215 5185
rect 12235 5165 12265 5185
rect 12285 5165 12315 5185
rect 12335 5165 12365 5185
rect 12385 5165 12415 5185
rect 12435 5165 12465 5185
rect 12485 5165 12515 5185
rect 12535 5165 12565 5185
rect 12585 5165 12615 5185
rect 12635 5165 12665 5185
rect 12685 5165 12715 5185
rect 12735 5165 12765 5185
rect 12785 5165 12815 5185
rect 12835 5165 12865 5185
rect 12885 5165 12915 5185
rect 12935 5165 12965 5185
rect 12985 5165 13015 5185
rect 13035 5165 13065 5185
rect 13085 5165 13115 5185
rect 13135 5165 13165 5185
rect 13185 5165 13215 5185
rect 13235 5165 13265 5185
rect 13285 5165 13315 5185
rect 13335 5165 13365 5185
rect 13385 5165 13415 5185
rect 13435 5165 13465 5185
rect 13485 5165 13515 5185
rect 13535 5165 13565 5185
rect 13585 5165 13615 5185
rect 13635 5165 13665 5185
rect 13685 5165 13715 5185
rect 13735 5165 13765 5185
rect 13785 5165 13815 5185
rect 13835 5165 13865 5185
rect 13885 5165 13915 5185
rect 13935 5165 13965 5185
rect 13985 5165 14015 5185
rect 14035 5165 14065 5185
rect 14085 5165 14115 5185
rect 14135 5165 14165 5185
rect 14185 5165 14215 5185
rect 14235 5165 14265 5185
rect 14285 5165 14315 5185
rect 14335 5165 14365 5185
rect 14385 5165 14415 5185
rect 14435 5165 14465 5185
rect 14485 5165 14515 5185
rect 14535 5165 14565 5185
rect 14585 5165 14615 5185
rect 14635 5165 14665 5185
rect 14685 5165 14715 5185
rect 14735 5165 14765 5185
rect 14785 5165 14815 5185
rect 14835 5165 14865 5185
rect 14885 5165 14915 5185
rect 14935 5165 14965 5185
rect 14985 5165 15015 5185
rect 15035 5165 15065 5185
rect 15085 5165 15115 5185
rect 15135 5165 15165 5185
rect 15185 5165 15215 5185
rect 15235 5165 15265 5185
rect 15285 5165 15315 5185
rect 15335 5165 15365 5185
rect 15385 5165 15415 5185
rect 15435 5165 15465 5185
rect 15485 5165 15515 5185
rect 15535 5165 15565 5185
rect 15585 5165 15615 5185
rect 15635 5165 15665 5185
rect 15685 5165 15715 5185
rect 15735 5165 15765 5185
rect 15785 5165 15815 5185
rect 15835 5165 15865 5185
rect 15885 5165 15915 5185
rect 15935 5165 15965 5185
rect 15985 5165 16015 5185
rect 16035 5165 16065 5185
rect 16085 5165 16115 5185
rect 16135 5165 16165 5185
rect 16185 5165 16215 5185
rect 16235 5165 16265 5185
rect 16285 5165 16315 5185
rect 16335 5165 16365 5185
rect 16385 5165 16415 5185
rect 16435 5165 16465 5185
rect 16485 5165 16515 5185
rect 16535 5165 16565 5185
rect 16585 5165 16615 5185
rect 16635 5165 16665 5185
rect 16685 5165 16715 5185
rect 16735 5165 16765 5185
rect 16785 5165 16815 5185
rect 16835 5165 16865 5185
rect 16885 5165 16915 5185
rect 16935 5165 16965 5185
rect 16985 5165 17015 5185
rect 17035 5165 17065 5185
rect 17085 5165 17115 5185
rect 17135 5165 17165 5185
rect 17185 5165 17215 5185
rect 17235 5165 17265 5185
rect 17285 5165 17315 5185
rect 17335 5165 17365 5185
rect 17385 5165 17415 5185
rect 17435 5165 17465 5185
rect 17485 5165 17515 5185
rect 17535 5165 17565 5185
rect 17585 5165 17615 5185
rect 17635 5165 17665 5185
rect 17685 5165 17715 5185
rect 17735 5165 17765 5185
rect 17785 5165 17815 5185
rect 17835 5165 17865 5185
rect 17885 5165 17915 5185
rect 17935 5165 17965 5185
rect 17985 5165 18015 5185
rect 18035 5165 18065 5185
rect 18085 5165 18115 5185
rect 18135 5165 18165 5185
rect 18185 5165 18215 5185
rect 18235 5165 18265 5185
rect 18285 5165 18315 5185
rect 18335 5165 18365 5185
rect 18385 5165 18415 5185
rect 18435 5165 18465 5185
rect 18485 5165 18515 5185
rect 18535 5165 18565 5185
rect 18585 5165 18615 5185
rect 18635 5165 18665 5185
rect 18685 5165 18715 5185
rect 18735 5165 18765 5185
rect 18785 5165 18815 5185
rect 18835 5165 18865 5185
rect 18885 5165 18915 5185
rect 18935 5165 18965 5185
rect 18985 5165 19015 5185
rect 19035 5165 19065 5185
rect 19085 5165 19115 5185
rect 19135 5165 19165 5185
rect 19185 5165 19215 5185
rect 19235 5165 19265 5185
rect 19285 5165 19315 5185
rect 19335 5165 19365 5185
rect 19385 5165 19415 5185
rect 19435 5165 19465 5185
rect 19485 5165 19515 5185
rect 19535 5165 19565 5185
rect 19585 5165 19615 5185
rect 19635 5165 19665 5185
rect 19685 5165 19715 5185
rect 19735 5165 19765 5185
rect 19785 5165 19815 5185
rect 19835 5165 19865 5185
rect 19885 5165 19915 5185
rect 19935 5165 19965 5185
rect 19985 5165 20015 5185
rect 20035 5165 20065 5185
rect 20085 5165 20115 5185
rect 20135 5165 20165 5185
rect 20185 5165 20215 5185
rect 20235 5165 20265 5185
rect 20285 5165 20315 5185
rect 20335 5165 20365 5185
rect 20385 5165 20400 5185
rect -650 5150 20400 5165
rect -650 3885 20400 3900
rect -650 3865 -635 3885
rect -615 3865 -585 3885
rect -565 3865 -535 3885
rect -515 3865 -485 3885
rect -465 3865 -435 3885
rect -415 3865 -385 3885
rect -365 3865 -335 3885
rect -315 3865 -285 3885
rect -265 3865 -235 3885
rect -215 3865 -185 3885
rect -165 3865 -135 3885
rect -115 3865 -85 3885
rect -65 3865 -35 3885
rect -15 3865 15 3885
rect 35 3865 65 3885
rect 85 3865 115 3885
rect 135 3865 165 3885
rect 185 3865 215 3885
rect 235 3865 265 3885
rect 285 3865 315 3885
rect 335 3865 365 3885
rect 385 3865 415 3885
rect 435 3865 465 3885
rect 485 3865 515 3885
rect 535 3865 565 3885
rect 585 3865 615 3885
rect 635 3865 665 3885
rect 685 3865 715 3885
rect 735 3865 765 3885
rect 785 3865 815 3885
rect 835 3865 865 3885
rect 885 3865 915 3885
rect 935 3865 965 3885
rect 985 3865 1015 3885
rect 1035 3865 1065 3885
rect 1085 3865 1115 3885
rect 1135 3865 1165 3885
rect 1185 3865 1215 3885
rect 1235 3865 1265 3885
rect 1285 3865 1315 3885
rect 1335 3865 1365 3885
rect 1385 3865 1415 3885
rect 1435 3865 1465 3885
rect 1485 3865 1515 3885
rect 1535 3865 1565 3885
rect 1585 3865 1615 3885
rect 1635 3865 1665 3885
rect 1685 3865 1715 3885
rect 1735 3865 1765 3885
rect 1785 3865 1815 3885
rect 1835 3865 1865 3885
rect 1885 3865 1915 3885
rect 1935 3865 1965 3885
rect 1985 3865 2015 3885
rect 2035 3865 2065 3885
rect 2085 3865 2115 3885
rect 2135 3865 2165 3885
rect 2185 3865 2215 3885
rect 2235 3865 2265 3885
rect 2285 3865 2315 3885
rect 2335 3865 2365 3885
rect 2385 3865 2415 3885
rect 2435 3865 2465 3885
rect 2485 3865 2515 3885
rect 2535 3865 2565 3885
rect 2585 3865 2615 3885
rect 2635 3865 2665 3885
rect 2685 3865 2715 3885
rect 2735 3865 2765 3885
rect 2785 3865 2815 3885
rect 2835 3865 2865 3885
rect 2885 3865 2915 3885
rect 2935 3865 2965 3885
rect 2985 3865 3015 3885
rect 3035 3865 3065 3885
rect 3085 3865 3115 3885
rect 3135 3865 3165 3885
rect 3185 3865 3215 3885
rect 3235 3865 3265 3885
rect 3285 3865 3315 3885
rect 3335 3865 3365 3885
rect 3385 3865 3415 3885
rect 3435 3865 3465 3885
rect 3485 3865 3515 3885
rect 3535 3865 3565 3885
rect 3585 3865 3615 3885
rect 3635 3865 3665 3885
rect 3685 3865 3715 3885
rect 3735 3865 3765 3885
rect 3785 3865 3815 3885
rect 3835 3865 3865 3885
rect 3885 3865 3915 3885
rect 3935 3865 3965 3885
rect 3985 3865 4015 3885
rect 4035 3865 4065 3885
rect 4085 3865 4115 3885
rect 4135 3865 4165 3885
rect 4185 3865 4215 3885
rect 4235 3865 4265 3885
rect 4285 3865 4315 3885
rect 4335 3865 4365 3885
rect 4385 3865 4415 3885
rect 4435 3865 4465 3885
rect 4485 3865 4515 3885
rect 4535 3865 4565 3885
rect 4585 3865 4615 3885
rect 4635 3865 4665 3885
rect 4685 3865 4715 3885
rect 4735 3865 4765 3885
rect 4785 3865 4815 3885
rect 4835 3865 4865 3885
rect 4885 3865 4915 3885
rect 4935 3865 4965 3885
rect 4985 3865 5015 3885
rect 5035 3865 5065 3885
rect 5085 3865 5115 3885
rect 5135 3865 5165 3885
rect 5185 3865 5215 3885
rect 5235 3865 5265 3885
rect 5285 3865 5315 3885
rect 5335 3865 5365 3885
rect 5385 3865 5415 3885
rect 5435 3865 5465 3885
rect 5485 3865 5515 3885
rect 5535 3865 5565 3885
rect 5585 3865 5615 3885
rect 5635 3865 5665 3885
rect 5685 3865 5715 3885
rect 5735 3865 5765 3885
rect 5785 3865 5815 3885
rect 5835 3865 5865 3885
rect 5885 3865 5915 3885
rect 5935 3865 5965 3885
rect 5985 3865 6015 3885
rect 6035 3865 6065 3885
rect 6085 3865 6115 3885
rect 6135 3865 6165 3885
rect 6185 3865 6215 3885
rect 6235 3865 6265 3885
rect 6285 3865 6315 3885
rect 6335 3865 6365 3885
rect 6385 3865 6415 3885
rect 6435 3865 6465 3885
rect 6485 3865 6515 3885
rect 6535 3865 6565 3885
rect 6585 3865 6615 3885
rect 6635 3865 6665 3885
rect 6685 3865 6715 3885
rect 6735 3865 6765 3885
rect 6785 3865 6815 3885
rect 6835 3865 6865 3885
rect 6885 3865 6915 3885
rect 6935 3865 6965 3885
rect 6985 3865 7015 3885
rect 7035 3865 7065 3885
rect 7085 3865 7115 3885
rect 7135 3865 7165 3885
rect 7185 3865 7215 3885
rect 7235 3865 7265 3885
rect 7285 3865 7315 3885
rect 7335 3865 7365 3885
rect 7385 3865 7415 3885
rect 7435 3865 7465 3885
rect 7485 3865 7515 3885
rect 7535 3865 7565 3885
rect 7585 3865 7615 3885
rect 7635 3865 7665 3885
rect 7685 3865 7715 3885
rect 7735 3865 7765 3885
rect 7785 3865 7815 3885
rect 7835 3865 7865 3885
rect 7885 3865 7915 3885
rect 7935 3865 7965 3885
rect 7985 3865 8015 3885
rect 8035 3865 8065 3885
rect 8085 3865 8115 3885
rect 8135 3865 8165 3885
rect 8185 3865 8215 3885
rect 8235 3865 8265 3885
rect 8285 3865 8315 3885
rect 8335 3865 8365 3885
rect 8385 3865 8415 3885
rect 8435 3865 8465 3885
rect 8485 3865 8515 3885
rect 8535 3865 8565 3885
rect 8585 3865 8615 3885
rect 8635 3865 8665 3885
rect 8685 3865 8715 3885
rect 8735 3865 8765 3885
rect 8785 3865 8815 3885
rect 8835 3865 8865 3885
rect 8885 3865 8915 3885
rect 8935 3865 8965 3885
rect 8985 3865 9015 3885
rect 9035 3865 9065 3885
rect 9085 3865 9115 3885
rect 9135 3865 9165 3885
rect 9185 3865 9215 3885
rect 9235 3865 9265 3885
rect 9285 3865 9315 3885
rect 9335 3865 9365 3885
rect 9385 3865 9415 3885
rect 9435 3865 9465 3885
rect 9485 3865 9515 3885
rect 9535 3865 9565 3885
rect 9585 3865 9615 3885
rect 9635 3865 9665 3885
rect 9685 3865 9715 3885
rect 9735 3865 9765 3885
rect 9785 3865 9815 3885
rect 9835 3865 9865 3885
rect 9885 3865 9915 3885
rect 9935 3865 9965 3885
rect 9985 3865 10015 3885
rect 10035 3865 10065 3885
rect 10085 3865 10115 3885
rect 10135 3865 10165 3885
rect 10185 3865 10215 3885
rect 10235 3865 10265 3885
rect 10285 3865 10315 3885
rect 10335 3865 10365 3885
rect 10385 3865 10415 3885
rect 10435 3865 10465 3885
rect 10485 3865 10515 3885
rect 10535 3865 10565 3885
rect 10585 3865 10615 3885
rect 10635 3865 10665 3885
rect 10685 3865 10715 3885
rect 10735 3865 10765 3885
rect 10785 3865 10815 3885
rect 10835 3865 10865 3885
rect 10885 3865 10915 3885
rect 10935 3865 10965 3885
rect 10985 3865 11015 3885
rect 11035 3865 11065 3885
rect 11085 3865 11115 3885
rect 11135 3865 11165 3885
rect 11185 3865 11215 3885
rect 11235 3865 11265 3885
rect 11285 3865 11315 3885
rect 11335 3865 11365 3885
rect 11385 3865 11415 3885
rect 11435 3865 11465 3885
rect 11485 3865 11515 3885
rect 11535 3865 11565 3885
rect 11585 3865 11615 3885
rect 11635 3865 11665 3885
rect 11685 3865 11715 3885
rect 11735 3865 11765 3885
rect 11785 3865 11815 3885
rect 11835 3865 11865 3885
rect 11885 3865 11915 3885
rect 11935 3865 11965 3885
rect 11985 3865 12015 3885
rect 12035 3865 12065 3885
rect 12085 3865 12115 3885
rect 12135 3865 12165 3885
rect 12185 3865 12215 3885
rect 12235 3865 12265 3885
rect 12285 3865 12315 3885
rect 12335 3865 12365 3885
rect 12385 3865 12415 3885
rect 12435 3865 12465 3885
rect 12485 3865 12515 3885
rect 12535 3865 12565 3885
rect 12585 3865 12615 3885
rect 12635 3865 12665 3885
rect 12685 3865 12715 3885
rect 12735 3865 12765 3885
rect 12785 3865 12815 3885
rect 12835 3865 12865 3885
rect 12885 3865 12915 3885
rect 12935 3865 12965 3885
rect 12985 3865 13015 3885
rect 13035 3865 13065 3885
rect 13085 3865 13115 3885
rect 13135 3865 13165 3885
rect 13185 3865 13215 3885
rect 13235 3865 13265 3885
rect 13285 3865 13315 3885
rect 13335 3865 13365 3885
rect 13385 3865 13415 3885
rect 13435 3865 13465 3885
rect 13485 3865 13515 3885
rect 13535 3865 13565 3885
rect 13585 3865 13615 3885
rect 13635 3865 13665 3885
rect 13685 3865 13715 3885
rect 13735 3865 13765 3885
rect 13785 3865 13815 3885
rect 13835 3865 13865 3885
rect 13885 3865 13915 3885
rect 13935 3865 13965 3885
rect 13985 3865 14015 3885
rect 14035 3865 14065 3885
rect 14085 3865 14115 3885
rect 14135 3865 14165 3885
rect 14185 3865 14215 3885
rect 14235 3865 14265 3885
rect 14285 3865 14315 3885
rect 14335 3865 14365 3885
rect 14385 3865 14415 3885
rect 14435 3865 14465 3885
rect 14485 3865 14515 3885
rect 14535 3865 14565 3885
rect 14585 3865 14615 3885
rect 14635 3865 14665 3885
rect 14685 3865 14715 3885
rect 14735 3865 14765 3885
rect 14785 3865 14815 3885
rect 14835 3865 14865 3885
rect 14885 3865 14915 3885
rect 14935 3865 14965 3885
rect 14985 3865 15015 3885
rect 15035 3865 15065 3885
rect 15085 3865 15115 3885
rect 15135 3865 15165 3885
rect 15185 3865 15215 3885
rect 15235 3865 15265 3885
rect 15285 3865 15315 3885
rect 15335 3865 15365 3885
rect 15385 3865 15415 3885
rect 15435 3865 15465 3885
rect 15485 3865 15515 3885
rect 15535 3865 15565 3885
rect 15585 3865 15615 3885
rect 15635 3865 15665 3885
rect 15685 3865 15715 3885
rect 15735 3865 15765 3885
rect 15785 3865 15815 3885
rect 15835 3865 15865 3885
rect 15885 3865 15915 3885
rect 15935 3865 15965 3885
rect 15985 3865 16015 3885
rect 16035 3865 16065 3885
rect 16085 3865 16115 3885
rect 16135 3865 16165 3885
rect 16185 3865 16215 3885
rect 16235 3865 16265 3885
rect 16285 3865 16315 3885
rect 16335 3865 16365 3885
rect 16385 3865 16415 3885
rect 16435 3865 16465 3885
rect 16485 3865 16515 3885
rect 16535 3865 16565 3885
rect 16585 3865 16615 3885
rect 16635 3865 16665 3885
rect 16685 3865 16715 3885
rect 16735 3865 16765 3885
rect 16785 3865 16815 3885
rect 16835 3865 16865 3885
rect 16885 3865 16915 3885
rect 16935 3865 16965 3885
rect 16985 3865 17015 3885
rect 17035 3865 17065 3885
rect 17085 3865 17115 3885
rect 17135 3865 17165 3885
rect 17185 3865 17215 3885
rect 17235 3865 17265 3885
rect 17285 3865 17315 3885
rect 17335 3865 17365 3885
rect 17385 3865 17415 3885
rect 17435 3865 17465 3885
rect 17485 3865 17515 3885
rect 17535 3865 17565 3885
rect 17585 3865 17615 3885
rect 17635 3865 17665 3885
rect 17685 3865 17715 3885
rect 17735 3865 17765 3885
rect 17785 3865 17815 3885
rect 17835 3865 17865 3885
rect 17885 3865 17915 3885
rect 17935 3865 17965 3885
rect 17985 3865 18015 3885
rect 18035 3865 18065 3885
rect 18085 3865 18115 3885
rect 18135 3865 18165 3885
rect 18185 3865 18215 3885
rect 18235 3865 18265 3885
rect 18285 3865 18315 3885
rect 18335 3865 18365 3885
rect 18385 3865 18415 3885
rect 18435 3865 18465 3885
rect 18485 3865 18515 3885
rect 18535 3865 18565 3885
rect 18585 3865 18615 3885
rect 18635 3865 18665 3885
rect 18685 3865 18715 3885
rect 18735 3865 18765 3885
rect 18785 3865 18815 3885
rect 18835 3865 18865 3885
rect 18885 3865 18915 3885
rect 18935 3865 18965 3885
rect 18985 3865 19015 3885
rect 19035 3865 19065 3885
rect 19085 3865 19115 3885
rect 19135 3865 19165 3885
rect 19185 3865 19215 3885
rect 19235 3865 19265 3885
rect 19285 3865 19315 3885
rect 19335 3865 19365 3885
rect 19385 3865 19415 3885
rect 19435 3865 19465 3885
rect 19485 3865 19515 3885
rect 19535 3865 19565 3885
rect 19585 3865 19615 3885
rect 19635 3865 19665 3885
rect 19685 3865 19715 3885
rect 19735 3865 19765 3885
rect 19785 3865 19815 3885
rect 19835 3865 19865 3885
rect 19885 3865 19915 3885
rect 19935 3865 19965 3885
rect 19985 3865 20015 3885
rect 20035 3865 20065 3885
rect 20085 3865 20115 3885
rect 20135 3865 20165 3885
rect 20185 3865 20215 3885
rect 20235 3865 20265 3885
rect 20285 3865 20315 3885
rect 20335 3865 20365 3885
rect 20385 3865 20400 3885
rect -650 3850 20400 3865
rect -650 2585 20400 2600
rect -650 2565 -635 2585
rect -615 2565 -585 2585
rect -565 2565 -535 2585
rect -515 2565 -485 2585
rect -465 2565 -435 2585
rect -415 2565 -385 2585
rect -365 2565 -335 2585
rect -315 2565 -285 2585
rect -265 2565 -235 2585
rect -215 2565 -185 2585
rect -165 2565 -135 2585
rect -115 2565 -85 2585
rect -65 2565 -35 2585
rect -15 2565 15 2585
rect 35 2565 65 2585
rect 85 2565 115 2585
rect 135 2565 165 2585
rect 185 2565 215 2585
rect 235 2565 265 2585
rect 285 2565 315 2585
rect 335 2565 365 2585
rect 385 2565 415 2585
rect 435 2565 465 2585
rect 485 2565 515 2585
rect 535 2565 565 2585
rect 585 2565 615 2585
rect 635 2565 665 2585
rect 685 2565 715 2585
rect 735 2565 765 2585
rect 785 2565 815 2585
rect 835 2565 865 2585
rect 885 2565 915 2585
rect 935 2565 965 2585
rect 985 2565 1015 2585
rect 1035 2565 1065 2585
rect 1085 2565 1115 2585
rect 1135 2565 1165 2585
rect 1185 2565 1215 2585
rect 1235 2565 1265 2585
rect 1285 2565 1315 2585
rect 1335 2565 1365 2585
rect 1385 2565 1415 2585
rect 1435 2565 1465 2585
rect 1485 2565 1515 2585
rect 1535 2565 1565 2585
rect 1585 2565 1615 2585
rect 1635 2565 1665 2585
rect 1685 2565 1715 2585
rect 1735 2565 1765 2585
rect 1785 2565 1815 2585
rect 1835 2565 1865 2585
rect 1885 2565 1915 2585
rect 1935 2565 1965 2585
rect 1985 2565 2015 2585
rect 2035 2565 2065 2585
rect 2085 2565 2115 2585
rect 2135 2565 2165 2585
rect 2185 2565 2215 2585
rect 2235 2565 2265 2585
rect 2285 2565 2315 2585
rect 2335 2565 2365 2585
rect 2385 2565 2415 2585
rect 2435 2565 2465 2585
rect 2485 2565 2515 2585
rect 2535 2565 2565 2585
rect 2585 2565 2615 2585
rect 2635 2565 2665 2585
rect 2685 2565 2715 2585
rect 2735 2565 2765 2585
rect 2785 2565 2815 2585
rect 2835 2565 2865 2585
rect 2885 2565 2915 2585
rect 2935 2565 2965 2585
rect 2985 2565 3015 2585
rect 3035 2565 3065 2585
rect 3085 2565 3115 2585
rect 3135 2565 3165 2585
rect 3185 2565 3215 2585
rect 3235 2565 3265 2585
rect 3285 2565 3315 2585
rect 3335 2565 3365 2585
rect 3385 2565 3415 2585
rect 3435 2565 3465 2585
rect 3485 2565 3515 2585
rect 3535 2565 3565 2585
rect 3585 2565 3615 2585
rect 3635 2565 3665 2585
rect 3685 2565 3715 2585
rect 3735 2565 3765 2585
rect 3785 2565 3815 2585
rect 3835 2565 3865 2585
rect 3885 2565 3915 2585
rect 3935 2565 3965 2585
rect 3985 2565 4015 2585
rect 4035 2565 4065 2585
rect 4085 2565 4115 2585
rect 4135 2565 4165 2585
rect 4185 2565 4215 2585
rect 4235 2565 4265 2585
rect 4285 2565 4315 2585
rect 4335 2565 4365 2585
rect 4385 2565 4415 2585
rect 4435 2565 4465 2585
rect 4485 2565 4515 2585
rect 4535 2565 4565 2585
rect 4585 2565 4615 2585
rect 4635 2565 4665 2585
rect 4685 2565 4715 2585
rect 4735 2565 4765 2585
rect 4785 2565 4815 2585
rect 4835 2565 4865 2585
rect 4885 2565 4915 2585
rect 4935 2565 4965 2585
rect 4985 2565 5015 2585
rect 5035 2565 5065 2585
rect 5085 2565 5115 2585
rect 5135 2565 5165 2585
rect 5185 2565 5215 2585
rect 5235 2565 5265 2585
rect 5285 2565 5315 2585
rect 5335 2565 5365 2585
rect 5385 2565 5415 2585
rect 5435 2565 5465 2585
rect 5485 2565 5515 2585
rect 5535 2565 5565 2585
rect 5585 2565 5615 2585
rect 5635 2565 5665 2585
rect 5685 2565 5715 2585
rect 5735 2565 5765 2585
rect 5785 2565 5815 2585
rect 5835 2565 5865 2585
rect 5885 2565 5915 2585
rect 5935 2565 5965 2585
rect 5985 2565 6015 2585
rect 6035 2565 6065 2585
rect 6085 2565 6115 2585
rect 6135 2565 6165 2585
rect 6185 2565 6215 2585
rect 6235 2565 6265 2585
rect 6285 2565 6315 2585
rect 6335 2565 6365 2585
rect 6385 2565 6415 2585
rect 6435 2565 6465 2585
rect 6485 2565 6515 2585
rect 6535 2565 6565 2585
rect 6585 2565 6615 2585
rect 6635 2565 6665 2585
rect 6685 2565 6715 2585
rect 6735 2565 6765 2585
rect 6785 2565 6815 2585
rect 6835 2565 6865 2585
rect 6885 2565 6915 2585
rect 6935 2565 6965 2585
rect 6985 2565 7015 2585
rect 7035 2565 7065 2585
rect 7085 2565 7115 2585
rect 7135 2565 7165 2585
rect 7185 2565 7215 2585
rect 7235 2565 7265 2585
rect 7285 2565 7315 2585
rect 7335 2565 7365 2585
rect 7385 2565 7415 2585
rect 7435 2565 7465 2585
rect 7485 2565 7515 2585
rect 7535 2565 7565 2585
rect 7585 2565 7615 2585
rect 7635 2565 7665 2585
rect 7685 2565 7715 2585
rect 7735 2565 7765 2585
rect 7785 2565 7815 2585
rect 7835 2565 7865 2585
rect 7885 2565 7915 2585
rect 7935 2565 7965 2585
rect 7985 2565 8015 2585
rect 8035 2565 8065 2585
rect 8085 2565 8115 2585
rect 8135 2565 8165 2585
rect 8185 2565 8215 2585
rect 8235 2565 8265 2585
rect 8285 2565 8315 2585
rect 8335 2565 8365 2585
rect 8385 2565 8415 2585
rect 8435 2565 8465 2585
rect 8485 2565 8515 2585
rect 8535 2565 8565 2585
rect 8585 2565 8615 2585
rect 8635 2565 8665 2585
rect 8685 2565 8715 2585
rect 8735 2565 8765 2585
rect 8785 2565 8815 2585
rect 8835 2565 8865 2585
rect 8885 2565 8915 2585
rect 8935 2565 8965 2585
rect 8985 2565 9015 2585
rect 9035 2565 9065 2585
rect 9085 2565 9115 2585
rect 9135 2565 9165 2585
rect 9185 2565 9215 2585
rect 9235 2565 9265 2585
rect 9285 2565 9315 2585
rect 9335 2565 9365 2585
rect 9385 2565 9415 2585
rect 9435 2565 9465 2585
rect 9485 2565 9515 2585
rect 9535 2565 9565 2585
rect 9585 2565 9615 2585
rect 9635 2565 9665 2585
rect 9685 2565 9715 2585
rect 9735 2565 9765 2585
rect 9785 2565 9815 2585
rect 9835 2565 9865 2585
rect 9885 2565 9915 2585
rect 9935 2565 9965 2585
rect 9985 2565 10015 2585
rect 10035 2565 10065 2585
rect 10085 2565 10115 2585
rect 10135 2565 10165 2585
rect 10185 2565 10215 2585
rect 10235 2565 10265 2585
rect 10285 2565 10315 2585
rect 10335 2565 10365 2585
rect 10385 2565 10415 2585
rect 10435 2565 10465 2585
rect 10485 2565 10515 2585
rect 10535 2565 10565 2585
rect 10585 2565 10615 2585
rect 10635 2565 10665 2585
rect 10685 2565 10715 2585
rect 10735 2565 10765 2585
rect 10785 2565 10815 2585
rect 10835 2565 10865 2585
rect 10885 2565 10915 2585
rect 10935 2565 10965 2585
rect 10985 2565 11015 2585
rect 11035 2565 11065 2585
rect 11085 2565 11115 2585
rect 11135 2565 11165 2585
rect 11185 2565 11215 2585
rect 11235 2565 11265 2585
rect 11285 2565 11315 2585
rect 11335 2565 11365 2585
rect 11385 2565 11415 2585
rect 11435 2565 11465 2585
rect 11485 2565 11515 2585
rect 11535 2565 11565 2585
rect 11585 2565 11615 2585
rect 11635 2565 11665 2585
rect 11685 2565 11715 2585
rect 11735 2565 11765 2585
rect 11785 2565 11815 2585
rect 11835 2565 11865 2585
rect 11885 2565 11915 2585
rect 11935 2565 11965 2585
rect 11985 2565 12015 2585
rect 12035 2565 12065 2585
rect 12085 2565 12115 2585
rect 12135 2565 12165 2585
rect 12185 2565 12215 2585
rect 12235 2565 12265 2585
rect 12285 2565 12315 2585
rect 12335 2565 12365 2585
rect 12385 2565 12415 2585
rect 12435 2565 12465 2585
rect 12485 2565 12515 2585
rect 12535 2565 12565 2585
rect 12585 2565 12615 2585
rect 12635 2565 12665 2585
rect 12685 2565 12715 2585
rect 12735 2565 12765 2585
rect 12785 2565 12815 2585
rect 12835 2565 12865 2585
rect 12885 2565 12915 2585
rect 12935 2565 12965 2585
rect 12985 2565 13015 2585
rect 13035 2565 13065 2585
rect 13085 2565 13115 2585
rect 13135 2565 13165 2585
rect 13185 2565 13215 2585
rect 13235 2565 13265 2585
rect 13285 2565 13315 2585
rect 13335 2565 13365 2585
rect 13385 2565 13415 2585
rect 13435 2565 13465 2585
rect 13485 2565 13515 2585
rect 13535 2565 13565 2585
rect 13585 2565 13615 2585
rect 13635 2565 13665 2585
rect 13685 2565 13715 2585
rect 13735 2565 13765 2585
rect 13785 2565 13815 2585
rect 13835 2565 13865 2585
rect 13885 2565 13915 2585
rect 13935 2565 13965 2585
rect 13985 2565 14015 2585
rect 14035 2565 14065 2585
rect 14085 2565 14115 2585
rect 14135 2565 14165 2585
rect 14185 2565 14215 2585
rect 14235 2565 14265 2585
rect 14285 2565 14315 2585
rect 14335 2565 14365 2585
rect 14385 2565 14415 2585
rect 14435 2565 14465 2585
rect 14485 2565 14515 2585
rect 14535 2565 14565 2585
rect 14585 2565 14615 2585
rect 14635 2565 14665 2585
rect 14685 2565 14715 2585
rect 14735 2565 14765 2585
rect 14785 2565 14815 2585
rect 14835 2565 14865 2585
rect 14885 2565 14915 2585
rect 14935 2565 14965 2585
rect 14985 2565 15015 2585
rect 15035 2565 15065 2585
rect 15085 2565 15115 2585
rect 15135 2565 15165 2585
rect 15185 2565 15215 2585
rect 15235 2565 15265 2585
rect 15285 2565 15315 2585
rect 15335 2565 15365 2585
rect 15385 2565 15415 2585
rect 15435 2565 15465 2585
rect 15485 2565 15515 2585
rect 15535 2565 15565 2585
rect 15585 2565 15615 2585
rect 15635 2565 15665 2585
rect 15685 2565 15715 2585
rect 15735 2565 15765 2585
rect 15785 2565 15815 2585
rect 15835 2565 15865 2585
rect 15885 2565 15915 2585
rect 15935 2565 15965 2585
rect 15985 2565 16015 2585
rect 16035 2565 16065 2585
rect 16085 2565 16115 2585
rect 16135 2565 16165 2585
rect 16185 2565 16215 2585
rect 16235 2565 16265 2585
rect 16285 2565 16315 2585
rect 16335 2565 16365 2585
rect 16385 2565 16415 2585
rect 16435 2565 16465 2585
rect 16485 2565 16515 2585
rect 16535 2565 16565 2585
rect 16585 2565 16615 2585
rect 16635 2565 16665 2585
rect 16685 2565 16715 2585
rect 16735 2565 16765 2585
rect 16785 2565 16815 2585
rect 16835 2565 16865 2585
rect 16885 2565 16915 2585
rect 16935 2565 16965 2585
rect 16985 2565 17015 2585
rect 17035 2565 17065 2585
rect 17085 2565 17115 2585
rect 17135 2565 17165 2585
rect 17185 2565 17215 2585
rect 17235 2565 17265 2585
rect 17285 2565 17315 2585
rect 17335 2565 17365 2585
rect 17385 2565 17415 2585
rect 17435 2565 17465 2585
rect 17485 2565 17515 2585
rect 17535 2565 17565 2585
rect 17585 2565 17615 2585
rect 17635 2565 17665 2585
rect 17685 2565 17715 2585
rect 17735 2565 17765 2585
rect 17785 2565 17815 2585
rect 17835 2565 17865 2585
rect 17885 2565 17915 2585
rect 17935 2565 17965 2585
rect 17985 2565 18015 2585
rect 18035 2565 18065 2585
rect 18085 2565 18115 2585
rect 18135 2565 18165 2585
rect 18185 2565 18215 2585
rect 18235 2565 18265 2585
rect 18285 2565 18315 2585
rect 18335 2565 18365 2585
rect 18385 2565 18415 2585
rect 18435 2565 18465 2585
rect 18485 2565 18515 2585
rect 18535 2565 18565 2585
rect 18585 2565 18615 2585
rect 18635 2565 18665 2585
rect 18685 2565 18715 2585
rect 18735 2565 18765 2585
rect 18785 2565 18815 2585
rect 18835 2565 18865 2585
rect 18885 2565 18915 2585
rect 18935 2565 18965 2585
rect 18985 2565 19015 2585
rect 19035 2565 19065 2585
rect 19085 2565 19115 2585
rect 19135 2565 19165 2585
rect 19185 2565 19215 2585
rect 19235 2565 19265 2585
rect 19285 2565 19315 2585
rect 19335 2565 19365 2585
rect 19385 2565 19415 2585
rect 19435 2565 19465 2585
rect 19485 2565 19515 2585
rect 19535 2565 19565 2585
rect 19585 2565 19615 2585
rect 19635 2565 19665 2585
rect 19685 2565 19715 2585
rect 19735 2565 19765 2585
rect 19785 2565 19815 2585
rect 19835 2565 19865 2585
rect 19885 2565 19915 2585
rect 19935 2565 19965 2585
rect 19985 2565 20015 2585
rect 20035 2565 20065 2585
rect 20085 2565 20115 2585
rect 20135 2565 20165 2585
rect 20185 2565 20215 2585
rect 20235 2565 20265 2585
rect 20285 2565 20315 2585
rect 20335 2565 20365 2585
rect 20385 2565 20400 2585
rect -650 2550 20400 2565
rect -650 1835 20400 1850
rect -650 1815 -635 1835
rect -615 1815 -585 1835
rect -565 1815 -535 1835
rect -515 1815 -485 1835
rect -465 1815 -435 1835
rect -415 1815 -385 1835
rect -365 1815 -335 1835
rect -315 1815 -285 1835
rect -265 1815 -235 1835
rect -215 1815 -185 1835
rect -165 1815 -135 1835
rect -115 1815 -85 1835
rect -65 1815 -35 1835
rect -15 1815 15 1835
rect 35 1815 65 1835
rect 85 1815 115 1835
rect 135 1815 165 1835
rect 185 1815 215 1835
rect 235 1815 265 1835
rect 285 1815 315 1835
rect 335 1815 365 1835
rect 385 1815 415 1835
rect 435 1815 465 1835
rect 485 1815 515 1835
rect 535 1815 565 1835
rect 585 1815 615 1835
rect 635 1815 665 1835
rect 685 1815 715 1835
rect 735 1815 765 1835
rect 785 1815 815 1835
rect 835 1815 865 1835
rect 885 1815 915 1835
rect 935 1815 965 1835
rect 985 1815 1015 1835
rect 1035 1815 1065 1835
rect 1085 1815 1115 1835
rect 1135 1815 1165 1835
rect 1185 1815 1215 1835
rect 1235 1815 1265 1835
rect 1285 1815 1315 1835
rect 1335 1815 1365 1835
rect 1385 1815 1415 1835
rect 1435 1815 1465 1835
rect 1485 1815 1515 1835
rect 1535 1815 1565 1835
rect 1585 1815 1615 1835
rect 1635 1815 1665 1835
rect 1685 1815 1715 1835
rect 1735 1815 1765 1835
rect 1785 1815 1815 1835
rect 1835 1815 1865 1835
rect 1885 1815 1915 1835
rect 1935 1815 1965 1835
rect 1985 1815 2015 1835
rect 2035 1815 2065 1835
rect 2085 1815 2115 1835
rect 2135 1815 2165 1835
rect 2185 1815 2215 1835
rect 2235 1815 2265 1835
rect 2285 1815 2315 1835
rect 2335 1815 2365 1835
rect 2385 1815 2415 1835
rect 2435 1815 2465 1835
rect 2485 1815 2515 1835
rect 2535 1815 2565 1835
rect 2585 1815 2615 1835
rect 2635 1815 2665 1835
rect 2685 1815 2715 1835
rect 2735 1815 2765 1835
rect 2785 1815 2815 1835
rect 2835 1815 2865 1835
rect 2885 1815 2915 1835
rect 2935 1815 2965 1835
rect 2985 1815 3015 1835
rect 3035 1815 3065 1835
rect 3085 1815 3115 1835
rect 3135 1815 3165 1835
rect 3185 1815 3215 1835
rect 3235 1815 3265 1835
rect 3285 1815 3315 1835
rect 3335 1815 3365 1835
rect 3385 1815 3415 1835
rect 3435 1815 3465 1835
rect 3485 1815 3515 1835
rect 3535 1815 3565 1835
rect 3585 1815 3615 1835
rect 3635 1815 3665 1835
rect 3685 1815 3715 1835
rect 3735 1815 3765 1835
rect 3785 1815 3815 1835
rect 3835 1815 3865 1835
rect 3885 1815 3915 1835
rect 3935 1815 3965 1835
rect 3985 1815 4015 1835
rect 4035 1815 4065 1835
rect 4085 1815 4115 1835
rect 4135 1815 4165 1835
rect 4185 1815 4215 1835
rect 4235 1815 4265 1835
rect 4285 1815 4315 1835
rect 4335 1815 4365 1835
rect 4385 1815 4415 1835
rect 4435 1815 4465 1835
rect 4485 1815 4515 1835
rect 4535 1815 4565 1835
rect 4585 1815 4615 1835
rect 4635 1815 4665 1835
rect 4685 1815 4715 1835
rect 4735 1815 4765 1835
rect 4785 1815 4815 1835
rect 4835 1815 4865 1835
rect 4885 1815 4915 1835
rect 4935 1815 4965 1835
rect 4985 1815 5015 1835
rect 5035 1815 5065 1835
rect 5085 1815 5115 1835
rect 5135 1815 5165 1835
rect 5185 1815 5215 1835
rect 5235 1815 5265 1835
rect 5285 1815 5315 1835
rect 5335 1815 5365 1835
rect 5385 1815 5415 1835
rect 5435 1815 5465 1835
rect 5485 1815 5515 1835
rect 5535 1815 5565 1835
rect 5585 1815 5615 1835
rect 5635 1815 5665 1835
rect 5685 1815 5715 1835
rect 5735 1815 5765 1835
rect 5785 1815 5815 1835
rect 5835 1815 5865 1835
rect 5885 1815 5915 1835
rect 5935 1815 5965 1835
rect 5985 1815 6015 1835
rect 6035 1815 6065 1835
rect 6085 1815 6115 1835
rect 6135 1815 6165 1835
rect 6185 1815 6215 1835
rect 6235 1815 6265 1835
rect 6285 1815 6315 1835
rect 6335 1815 6365 1835
rect 6385 1815 6415 1835
rect 6435 1815 6465 1835
rect 6485 1815 6515 1835
rect 6535 1815 6565 1835
rect 6585 1815 6615 1835
rect 6635 1815 6665 1835
rect 6685 1815 6715 1835
rect 6735 1815 6765 1835
rect 6785 1815 6815 1835
rect 6835 1815 6865 1835
rect 6885 1815 6915 1835
rect 6935 1815 6965 1835
rect 6985 1815 7015 1835
rect 7035 1815 7065 1835
rect 7085 1815 7115 1835
rect 7135 1815 7165 1835
rect 7185 1815 7215 1835
rect 7235 1815 7265 1835
rect 7285 1815 7315 1835
rect 7335 1815 7365 1835
rect 7385 1815 7415 1835
rect 7435 1815 7465 1835
rect 7485 1815 7515 1835
rect 7535 1815 7565 1835
rect 7585 1815 7615 1835
rect 7635 1815 7665 1835
rect 7685 1815 7715 1835
rect 7735 1815 7765 1835
rect 7785 1815 7815 1835
rect 7835 1815 7865 1835
rect 7885 1815 7915 1835
rect 7935 1815 7965 1835
rect 7985 1815 8015 1835
rect 8035 1815 8065 1835
rect 8085 1815 8115 1835
rect 8135 1815 8165 1835
rect 8185 1815 8215 1835
rect 8235 1815 8265 1835
rect 8285 1815 8315 1835
rect 8335 1815 8365 1835
rect 8385 1815 8415 1835
rect 8435 1815 8465 1835
rect 8485 1815 8515 1835
rect 8535 1815 8565 1835
rect 8585 1815 8615 1835
rect 8635 1815 8665 1835
rect 8685 1815 8715 1835
rect 8735 1815 8765 1835
rect 8785 1815 8815 1835
rect 8835 1815 8865 1835
rect 8885 1815 8915 1835
rect 8935 1815 8965 1835
rect 8985 1815 9015 1835
rect 9035 1815 9065 1835
rect 9085 1815 9115 1835
rect 9135 1815 9165 1835
rect 9185 1815 9215 1835
rect 9235 1815 9265 1835
rect 9285 1815 9315 1835
rect 9335 1815 9365 1835
rect 9385 1815 9415 1835
rect 9435 1815 9465 1835
rect 9485 1815 9515 1835
rect 9535 1815 9565 1835
rect 9585 1815 9615 1835
rect 9635 1815 9665 1835
rect 9685 1815 9715 1835
rect 9735 1815 9765 1835
rect 9785 1815 9815 1835
rect 9835 1815 9865 1835
rect 9885 1815 9915 1835
rect 9935 1815 9965 1835
rect 9985 1815 10015 1835
rect 10035 1815 10065 1835
rect 10085 1815 10115 1835
rect 10135 1815 10165 1835
rect 10185 1815 10215 1835
rect 10235 1815 10265 1835
rect 10285 1815 10315 1835
rect 10335 1815 10365 1835
rect 10385 1815 10415 1835
rect 10435 1815 10465 1835
rect 10485 1815 10515 1835
rect 10535 1815 10565 1835
rect 10585 1815 10615 1835
rect 10635 1815 10665 1835
rect 10685 1815 10715 1835
rect 10735 1815 10765 1835
rect 10785 1815 10815 1835
rect 10835 1815 10865 1835
rect 10885 1815 10915 1835
rect 10935 1815 10965 1835
rect 10985 1815 11015 1835
rect 11035 1815 11065 1835
rect 11085 1815 11115 1835
rect 11135 1815 11165 1835
rect 11185 1815 11215 1835
rect 11235 1815 11265 1835
rect 11285 1815 11315 1835
rect 11335 1815 11365 1835
rect 11385 1815 11415 1835
rect 11435 1815 11465 1835
rect 11485 1815 11515 1835
rect 11535 1815 11565 1835
rect 11585 1815 11615 1835
rect 11635 1815 11665 1835
rect 11685 1815 11715 1835
rect 11735 1815 11765 1835
rect 11785 1815 11815 1835
rect 11835 1815 11865 1835
rect 11885 1815 11915 1835
rect 11935 1815 11965 1835
rect 11985 1815 12015 1835
rect 12035 1815 12065 1835
rect 12085 1815 12115 1835
rect 12135 1815 12165 1835
rect 12185 1815 12215 1835
rect 12235 1815 12265 1835
rect 12285 1815 12315 1835
rect 12335 1815 12365 1835
rect 12385 1815 12415 1835
rect 12435 1815 12465 1835
rect 12485 1815 12515 1835
rect 12535 1815 12565 1835
rect 12585 1815 12615 1835
rect 12635 1815 12665 1835
rect 12685 1815 12715 1835
rect 12735 1815 12765 1835
rect 12785 1815 12815 1835
rect 12835 1815 12865 1835
rect 12885 1815 12915 1835
rect 12935 1815 12965 1835
rect 12985 1815 13015 1835
rect 13035 1815 13065 1835
rect 13085 1815 13115 1835
rect 13135 1815 13165 1835
rect 13185 1815 13215 1835
rect 13235 1815 13265 1835
rect 13285 1815 13315 1835
rect 13335 1815 13365 1835
rect 13385 1815 13415 1835
rect 13435 1815 13465 1835
rect 13485 1815 13515 1835
rect 13535 1815 13565 1835
rect 13585 1815 13615 1835
rect 13635 1815 13665 1835
rect 13685 1815 13715 1835
rect 13735 1815 13765 1835
rect 13785 1815 13815 1835
rect 13835 1815 13865 1835
rect 13885 1815 13915 1835
rect 13935 1815 13965 1835
rect 13985 1815 14015 1835
rect 14035 1815 14065 1835
rect 14085 1815 14115 1835
rect 14135 1815 14165 1835
rect 14185 1815 14215 1835
rect 14235 1815 14265 1835
rect 14285 1815 14315 1835
rect 14335 1815 14365 1835
rect 14385 1815 14415 1835
rect 14435 1815 14465 1835
rect 14485 1815 14515 1835
rect 14535 1815 14565 1835
rect 14585 1815 14615 1835
rect 14635 1815 14665 1835
rect 14685 1815 14715 1835
rect 14735 1815 14765 1835
rect 14785 1815 14815 1835
rect 14835 1815 14865 1835
rect 14885 1815 14915 1835
rect 14935 1815 14965 1835
rect 14985 1815 15015 1835
rect 15035 1815 15065 1835
rect 15085 1815 15115 1835
rect 15135 1815 15165 1835
rect 15185 1815 15215 1835
rect 15235 1815 15265 1835
rect 15285 1815 15315 1835
rect 15335 1815 15365 1835
rect 15385 1815 15415 1835
rect 15435 1815 15465 1835
rect 15485 1815 15515 1835
rect 15535 1815 15565 1835
rect 15585 1815 15615 1835
rect 15635 1815 15665 1835
rect 15685 1815 15715 1835
rect 15735 1815 15765 1835
rect 15785 1815 15815 1835
rect 15835 1815 15865 1835
rect 15885 1815 15915 1835
rect 15935 1815 15965 1835
rect 15985 1815 16015 1835
rect 16035 1815 16065 1835
rect 16085 1815 16115 1835
rect 16135 1815 16165 1835
rect 16185 1815 16215 1835
rect 16235 1815 16265 1835
rect 16285 1815 16315 1835
rect 16335 1815 16365 1835
rect 16385 1815 16415 1835
rect 16435 1815 16465 1835
rect 16485 1815 16515 1835
rect 16535 1815 16565 1835
rect 16585 1815 16615 1835
rect 16635 1815 16665 1835
rect 16685 1815 16715 1835
rect 16735 1815 16765 1835
rect 16785 1815 16815 1835
rect 16835 1815 16865 1835
rect 16885 1815 16915 1835
rect 16935 1815 16965 1835
rect 16985 1815 17015 1835
rect 17035 1815 17065 1835
rect 17085 1815 17115 1835
rect 17135 1815 17165 1835
rect 17185 1815 17215 1835
rect 17235 1815 17265 1835
rect 17285 1815 17315 1835
rect 17335 1815 17365 1835
rect 17385 1815 17415 1835
rect 17435 1815 17465 1835
rect 17485 1815 17515 1835
rect 17535 1815 17565 1835
rect 17585 1815 17615 1835
rect 17635 1815 17665 1835
rect 17685 1815 17715 1835
rect 17735 1815 17765 1835
rect 17785 1815 17815 1835
rect 17835 1815 17865 1835
rect 17885 1815 17915 1835
rect 17935 1815 17965 1835
rect 17985 1815 18015 1835
rect 18035 1815 18065 1835
rect 18085 1815 18115 1835
rect 18135 1815 18165 1835
rect 18185 1815 18215 1835
rect 18235 1815 18265 1835
rect 18285 1815 18315 1835
rect 18335 1815 18365 1835
rect 18385 1815 18415 1835
rect 18435 1815 18465 1835
rect 18485 1815 18515 1835
rect 18535 1815 18565 1835
rect 18585 1815 18615 1835
rect 18635 1815 18665 1835
rect 18685 1815 18715 1835
rect 18735 1815 18765 1835
rect 18785 1815 18815 1835
rect 18835 1815 18865 1835
rect 18885 1815 18915 1835
rect 18935 1815 18965 1835
rect 18985 1815 19015 1835
rect 19035 1815 19065 1835
rect 19085 1815 19115 1835
rect 19135 1815 19165 1835
rect 19185 1815 19215 1835
rect 19235 1815 19265 1835
rect 19285 1815 19315 1835
rect 19335 1815 19365 1835
rect 19385 1815 19415 1835
rect 19435 1815 19465 1835
rect 19485 1815 19515 1835
rect 19535 1815 19565 1835
rect 19585 1815 19615 1835
rect 19635 1815 19665 1835
rect 19685 1815 19715 1835
rect 19735 1815 19765 1835
rect 19785 1815 19815 1835
rect 19835 1815 19865 1835
rect 19885 1815 19915 1835
rect 19935 1815 19965 1835
rect 19985 1815 20015 1835
rect 20035 1815 20065 1835
rect 20085 1815 20115 1835
rect 20135 1815 20165 1835
rect 20185 1815 20215 1835
rect 20235 1815 20265 1835
rect 20285 1815 20315 1835
rect 20335 1815 20365 1835
rect 20385 1815 20400 1835
rect -650 1800 20400 1815
rect -650 -1865 20400 -1850
rect -650 -1885 -635 -1865
rect -615 -1885 -585 -1865
rect -565 -1885 -535 -1865
rect -515 -1885 -485 -1865
rect -465 -1885 -435 -1865
rect -415 -1885 -385 -1865
rect -365 -1885 -335 -1865
rect -315 -1885 -285 -1865
rect -265 -1885 -235 -1865
rect -215 -1885 -185 -1865
rect -165 -1885 -135 -1865
rect -115 -1885 -85 -1865
rect -65 -1885 -35 -1865
rect -15 -1885 15 -1865
rect 35 -1885 65 -1865
rect 85 -1885 115 -1865
rect 135 -1885 165 -1865
rect 185 -1885 215 -1865
rect 235 -1885 265 -1865
rect 285 -1885 315 -1865
rect 335 -1885 365 -1865
rect 385 -1885 415 -1865
rect 435 -1885 465 -1865
rect 485 -1885 515 -1865
rect 535 -1885 565 -1865
rect 585 -1885 615 -1865
rect 635 -1885 665 -1865
rect 685 -1885 715 -1865
rect 735 -1885 765 -1865
rect 785 -1885 815 -1865
rect 835 -1885 865 -1865
rect 885 -1885 915 -1865
rect 935 -1885 965 -1865
rect 985 -1885 1015 -1865
rect 1035 -1885 1065 -1865
rect 1085 -1885 1115 -1865
rect 1135 -1885 1165 -1865
rect 1185 -1885 1215 -1865
rect 1235 -1885 1265 -1865
rect 1285 -1885 1315 -1865
rect 1335 -1885 1365 -1865
rect 1385 -1885 1415 -1865
rect 1435 -1885 1465 -1865
rect 1485 -1885 1515 -1865
rect 1535 -1885 1565 -1865
rect 1585 -1885 1615 -1865
rect 1635 -1885 1665 -1865
rect 1685 -1885 1715 -1865
rect 1735 -1885 1765 -1865
rect 1785 -1885 1815 -1865
rect 1835 -1885 1865 -1865
rect 1885 -1885 1915 -1865
rect 1935 -1885 1965 -1865
rect 1985 -1885 2015 -1865
rect 2035 -1885 2065 -1865
rect 2085 -1885 2115 -1865
rect 2135 -1885 2165 -1865
rect 2185 -1885 2215 -1865
rect 2235 -1885 2265 -1865
rect 2285 -1885 2315 -1865
rect 2335 -1885 2365 -1865
rect 2385 -1885 2415 -1865
rect 2435 -1885 2465 -1865
rect 2485 -1885 2515 -1865
rect 2535 -1885 2565 -1865
rect 2585 -1885 2615 -1865
rect 2635 -1885 2665 -1865
rect 2685 -1885 2715 -1865
rect 2735 -1885 2765 -1865
rect 2785 -1885 2815 -1865
rect 2835 -1885 2865 -1865
rect 2885 -1885 2915 -1865
rect 2935 -1885 2965 -1865
rect 2985 -1885 3015 -1865
rect 3035 -1885 3065 -1865
rect 3085 -1885 3115 -1865
rect 3135 -1885 3165 -1865
rect 3185 -1885 3215 -1865
rect 3235 -1885 3265 -1865
rect 3285 -1885 3315 -1865
rect 3335 -1885 3365 -1865
rect 3385 -1885 3415 -1865
rect 3435 -1885 3465 -1865
rect 3485 -1885 3515 -1865
rect 3535 -1885 3565 -1865
rect 3585 -1885 3615 -1865
rect 3635 -1885 3665 -1865
rect 3685 -1885 3715 -1865
rect 3735 -1885 3765 -1865
rect 3785 -1885 3815 -1865
rect 3835 -1885 3865 -1865
rect 3885 -1885 3915 -1865
rect 3935 -1885 3965 -1865
rect 3985 -1885 4015 -1865
rect 4035 -1885 4065 -1865
rect 4085 -1885 4115 -1865
rect 4135 -1885 4165 -1865
rect 4185 -1885 4215 -1865
rect 4235 -1885 4265 -1865
rect 4285 -1885 4315 -1865
rect 4335 -1885 4365 -1865
rect 4385 -1885 4415 -1865
rect 4435 -1885 4465 -1865
rect 4485 -1885 4515 -1865
rect 4535 -1885 4565 -1865
rect 4585 -1885 4615 -1865
rect 4635 -1885 4665 -1865
rect 4685 -1885 4715 -1865
rect 4735 -1885 4765 -1865
rect 4785 -1885 4815 -1865
rect 4835 -1885 4865 -1865
rect 4885 -1885 4915 -1865
rect 4935 -1885 4965 -1865
rect 4985 -1885 5015 -1865
rect 5035 -1885 5065 -1865
rect 5085 -1885 5115 -1865
rect 5135 -1885 5165 -1865
rect 5185 -1885 5215 -1865
rect 5235 -1885 5265 -1865
rect 5285 -1885 5315 -1865
rect 5335 -1885 5365 -1865
rect 5385 -1885 5415 -1865
rect 5435 -1885 5465 -1865
rect 5485 -1885 5515 -1865
rect 5535 -1885 5565 -1865
rect 5585 -1885 5615 -1865
rect 5635 -1885 5665 -1865
rect 5685 -1885 5715 -1865
rect 5735 -1885 5765 -1865
rect 5785 -1885 5815 -1865
rect 5835 -1885 5865 -1865
rect 5885 -1885 5915 -1865
rect 5935 -1885 5965 -1865
rect 5985 -1885 6015 -1865
rect 6035 -1885 6065 -1865
rect 6085 -1885 6115 -1865
rect 6135 -1885 6165 -1865
rect 6185 -1885 6215 -1865
rect 6235 -1885 6265 -1865
rect 6285 -1885 6315 -1865
rect 6335 -1885 6365 -1865
rect 6385 -1885 6415 -1865
rect 6435 -1885 6465 -1865
rect 6485 -1885 6515 -1865
rect 6535 -1885 6565 -1865
rect 6585 -1885 6615 -1865
rect 6635 -1885 6665 -1865
rect 6685 -1885 6715 -1865
rect 6735 -1885 6765 -1865
rect 6785 -1885 6815 -1865
rect 6835 -1885 6865 -1865
rect 6885 -1885 6915 -1865
rect 6935 -1885 6965 -1865
rect 6985 -1885 7015 -1865
rect 7035 -1885 7065 -1865
rect 7085 -1885 7115 -1865
rect 7135 -1885 7165 -1865
rect 7185 -1885 7215 -1865
rect 7235 -1885 7265 -1865
rect 7285 -1885 7315 -1865
rect 7335 -1885 7365 -1865
rect 7385 -1885 7415 -1865
rect 7435 -1885 7465 -1865
rect 7485 -1885 7515 -1865
rect 7535 -1885 7565 -1865
rect 7585 -1885 7615 -1865
rect 7635 -1885 7665 -1865
rect 7685 -1885 7715 -1865
rect 7735 -1885 7765 -1865
rect 7785 -1885 7815 -1865
rect 7835 -1885 7865 -1865
rect 7885 -1885 7915 -1865
rect 7935 -1885 7965 -1865
rect 7985 -1885 8015 -1865
rect 8035 -1885 8065 -1865
rect 8085 -1885 8115 -1865
rect 8135 -1885 8165 -1865
rect 8185 -1885 8215 -1865
rect 8235 -1885 8265 -1865
rect 8285 -1885 8315 -1865
rect 8335 -1885 8365 -1865
rect 8385 -1885 8415 -1865
rect 8435 -1885 8465 -1865
rect 8485 -1885 8515 -1865
rect 8535 -1885 8565 -1865
rect 8585 -1885 8615 -1865
rect 8635 -1885 8665 -1865
rect 8685 -1885 8715 -1865
rect 8735 -1885 8765 -1865
rect 8785 -1885 8815 -1865
rect 8835 -1885 8865 -1865
rect 8885 -1885 8915 -1865
rect 8935 -1885 8965 -1865
rect 8985 -1885 9015 -1865
rect 9035 -1885 9065 -1865
rect 9085 -1885 9115 -1865
rect 9135 -1885 9165 -1865
rect 9185 -1885 9215 -1865
rect 9235 -1885 9265 -1865
rect 9285 -1885 9315 -1865
rect 9335 -1885 9365 -1865
rect 9385 -1885 9415 -1865
rect 9435 -1885 9465 -1865
rect 9485 -1885 9515 -1865
rect 9535 -1885 9565 -1865
rect 9585 -1885 9615 -1865
rect 9635 -1885 9665 -1865
rect 9685 -1885 9715 -1865
rect 9735 -1885 9765 -1865
rect 9785 -1885 9815 -1865
rect 9835 -1885 9865 -1865
rect 9885 -1885 9915 -1865
rect 9935 -1885 9965 -1865
rect 9985 -1885 10015 -1865
rect 10035 -1885 10065 -1865
rect 10085 -1885 10115 -1865
rect 10135 -1885 10165 -1865
rect 10185 -1885 10215 -1865
rect 10235 -1885 10265 -1865
rect 10285 -1885 10315 -1865
rect 10335 -1885 10365 -1865
rect 10385 -1885 10415 -1865
rect 10435 -1885 10465 -1865
rect 10485 -1885 10515 -1865
rect 10535 -1885 10565 -1865
rect 10585 -1885 10615 -1865
rect 10635 -1885 10665 -1865
rect 10685 -1885 10715 -1865
rect 10735 -1885 10765 -1865
rect 10785 -1885 10815 -1865
rect 10835 -1885 10865 -1865
rect 10885 -1885 10915 -1865
rect 10935 -1885 10965 -1865
rect 10985 -1885 11015 -1865
rect 11035 -1885 11065 -1865
rect 11085 -1885 11115 -1865
rect 11135 -1885 11165 -1865
rect 11185 -1885 11215 -1865
rect 11235 -1885 11265 -1865
rect 11285 -1885 11315 -1865
rect 11335 -1885 11365 -1865
rect 11385 -1885 11415 -1865
rect 11435 -1885 11465 -1865
rect 11485 -1885 11515 -1865
rect 11535 -1885 11565 -1865
rect 11585 -1885 11615 -1865
rect 11635 -1885 11665 -1865
rect 11685 -1885 11715 -1865
rect 11735 -1885 11765 -1865
rect 11785 -1885 11815 -1865
rect 11835 -1885 11865 -1865
rect 11885 -1885 11915 -1865
rect 11935 -1885 11965 -1865
rect 11985 -1885 12015 -1865
rect 12035 -1885 12065 -1865
rect 12085 -1885 12115 -1865
rect 12135 -1885 12165 -1865
rect 12185 -1885 12215 -1865
rect 12235 -1885 12265 -1865
rect 12285 -1885 12315 -1865
rect 12335 -1885 12365 -1865
rect 12385 -1885 12415 -1865
rect 12435 -1885 12465 -1865
rect 12485 -1885 12515 -1865
rect 12535 -1885 12565 -1865
rect 12585 -1885 12615 -1865
rect 12635 -1885 12665 -1865
rect 12685 -1885 12715 -1865
rect 12735 -1885 12765 -1865
rect 12785 -1885 12815 -1865
rect 12835 -1885 12865 -1865
rect 12885 -1885 12915 -1865
rect 12935 -1885 12965 -1865
rect 12985 -1885 13015 -1865
rect 13035 -1885 13065 -1865
rect 13085 -1885 13115 -1865
rect 13135 -1885 13165 -1865
rect 13185 -1885 13215 -1865
rect 13235 -1885 13265 -1865
rect 13285 -1885 13315 -1865
rect 13335 -1885 13365 -1865
rect 13385 -1885 13415 -1865
rect 13435 -1885 13465 -1865
rect 13485 -1885 13515 -1865
rect 13535 -1885 13565 -1865
rect 13585 -1885 13615 -1865
rect 13635 -1885 13665 -1865
rect 13685 -1885 13715 -1865
rect 13735 -1885 13765 -1865
rect 13785 -1885 13815 -1865
rect 13835 -1885 13865 -1865
rect 13885 -1885 13915 -1865
rect 13935 -1885 13965 -1865
rect 13985 -1885 14015 -1865
rect 14035 -1885 14065 -1865
rect 14085 -1885 14115 -1865
rect 14135 -1885 14165 -1865
rect 14185 -1885 14215 -1865
rect 14235 -1885 14265 -1865
rect 14285 -1885 14315 -1865
rect 14335 -1885 14365 -1865
rect 14385 -1885 14415 -1865
rect 14435 -1885 14465 -1865
rect 14485 -1885 14515 -1865
rect 14535 -1885 14565 -1865
rect 14585 -1885 14615 -1865
rect 14635 -1885 14665 -1865
rect 14685 -1885 14715 -1865
rect 14735 -1885 14765 -1865
rect 14785 -1885 14815 -1865
rect 14835 -1885 14865 -1865
rect 14885 -1885 14915 -1865
rect 14935 -1885 14965 -1865
rect 14985 -1885 15015 -1865
rect 15035 -1885 15065 -1865
rect 15085 -1885 15115 -1865
rect 15135 -1885 15165 -1865
rect 15185 -1885 15215 -1865
rect 15235 -1885 15265 -1865
rect 15285 -1885 15315 -1865
rect 15335 -1885 15365 -1865
rect 15385 -1885 15415 -1865
rect 15435 -1885 15465 -1865
rect 15485 -1885 15515 -1865
rect 15535 -1885 15565 -1865
rect 15585 -1885 15615 -1865
rect 15635 -1885 15665 -1865
rect 15685 -1885 15715 -1865
rect 15735 -1885 15765 -1865
rect 15785 -1885 15815 -1865
rect 15835 -1885 15865 -1865
rect 15885 -1885 15915 -1865
rect 15935 -1885 15965 -1865
rect 15985 -1885 16015 -1865
rect 16035 -1885 16065 -1865
rect 16085 -1885 16115 -1865
rect 16135 -1885 16165 -1865
rect 16185 -1885 16215 -1865
rect 16235 -1885 16265 -1865
rect 16285 -1885 16315 -1865
rect 16335 -1885 16365 -1865
rect 16385 -1885 16415 -1865
rect 16435 -1885 16465 -1865
rect 16485 -1885 16515 -1865
rect 16535 -1885 16565 -1865
rect 16585 -1885 16615 -1865
rect 16635 -1885 16665 -1865
rect 16685 -1885 16715 -1865
rect 16735 -1885 16765 -1865
rect 16785 -1885 16815 -1865
rect 16835 -1885 16865 -1865
rect 16885 -1885 16915 -1865
rect 16935 -1885 16965 -1865
rect 16985 -1885 17015 -1865
rect 17035 -1885 17065 -1865
rect 17085 -1885 17115 -1865
rect 17135 -1885 17165 -1865
rect 17185 -1885 17215 -1865
rect 17235 -1885 17265 -1865
rect 17285 -1885 17315 -1865
rect 17335 -1885 17365 -1865
rect 17385 -1885 17415 -1865
rect 17435 -1885 17465 -1865
rect 17485 -1885 17515 -1865
rect 17535 -1885 17565 -1865
rect 17585 -1885 17615 -1865
rect 17635 -1885 17665 -1865
rect 17685 -1885 17715 -1865
rect 17735 -1885 17765 -1865
rect 17785 -1885 17815 -1865
rect 17835 -1885 17865 -1865
rect 17885 -1885 17915 -1865
rect 17935 -1885 17965 -1865
rect 17985 -1885 18015 -1865
rect 18035 -1885 18065 -1865
rect 18085 -1885 18115 -1865
rect 18135 -1885 18165 -1865
rect 18185 -1885 18215 -1865
rect 18235 -1885 18265 -1865
rect 18285 -1885 18315 -1865
rect 18335 -1885 18365 -1865
rect 18385 -1885 18415 -1865
rect 18435 -1885 18465 -1865
rect 18485 -1885 18515 -1865
rect 18535 -1885 18565 -1865
rect 18585 -1885 18615 -1865
rect 18635 -1885 18665 -1865
rect 18685 -1885 18715 -1865
rect 18735 -1885 18765 -1865
rect 18785 -1885 18815 -1865
rect 18835 -1885 18865 -1865
rect 18885 -1885 18915 -1865
rect 18935 -1885 18965 -1865
rect 18985 -1885 19015 -1865
rect 19035 -1885 19065 -1865
rect 19085 -1885 19115 -1865
rect 19135 -1885 19165 -1865
rect 19185 -1885 19215 -1865
rect 19235 -1885 19265 -1865
rect 19285 -1885 19315 -1865
rect 19335 -1885 19365 -1865
rect 19385 -1885 19415 -1865
rect 19435 -1885 19465 -1865
rect 19485 -1885 19515 -1865
rect 19535 -1885 19565 -1865
rect 19585 -1885 19615 -1865
rect 19635 -1885 19665 -1865
rect 19685 -1885 19715 -1865
rect 19735 -1885 19765 -1865
rect 19785 -1885 19815 -1865
rect 19835 -1885 19865 -1865
rect 19885 -1885 19915 -1865
rect 19935 -1885 19965 -1865
rect 19985 -1885 20015 -1865
rect 20035 -1885 20065 -1865
rect 20085 -1885 20115 -1865
rect 20135 -1885 20165 -1865
rect 20185 -1885 20215 -1865
rect 20235 -1885 20265 -1865
rect 20285 -1885 20315 -1865
rect 20335 -1885 20365 -1865
rect 20385 -1885 20400 -1865
rect -650 -1900 20400 -1885
<< mvpsubdiffcont >>
rect -885 2415 -865 2435
rect -835 2415 -815 2435
rect -785 2415 -765 2435
rect -735 2415 -715 2435
rect -685 2415 -665 2435
rect -635 2415 -615 2435
rect -585 2415 -565 2435
rect -535 2415 -515 2435
rect -485 2415 -465 2435
rect -435 2415 -415 2435
rect -385 2415 -365 2435
rect -335 2415 -315 2435
rect -285 2415 -265 2435
rect -235 2415 -215 2435
rect -185 2415 -165 2435
rect -135 2415 -115 2435
rect -85 2415 -65 2435
rect -35 2415 -15 2435
rect 15 2415 35 2435
rect 65 2415 85 2435
rect 115 2415 135 2435
rect 165 2415 185 2435
rect 215 2415 235 2435
rect 265 2415 285 2435
rect 315 2415 335 2435
rect 365 2415 385 2435
rect 415 2415 435 2435
rect 465 2415 485 2435
rect 515 2415 535 2435
rect 565 2415 585 2435
rect 615 2415 635 2435
rect 665 2415 685 2435
rect 715 2415 735 2435
rect 765 2415 785 2435
rect 815 2415 835 2435
rect 865 2415 885 2435
rect 915 2415 935 2435
rect 965 2415 985 2435
rect 1015 2415 1035 2435
rect 1065 2415 1085 2435
rect 1115 2415 1135 2435
rect 1165 2415 1185 2435
rect 1215 2415 1235 2435
rect 1265 2415 1285 2435
rect 1315 2415 1335 2435
rect 1365 2415 1385 2435
rect 1415 2415 1435 2435
rect 1465 2415 1485 2435
rect 1515 2415 1535 2435
rect 1565 2415 1585 2435
rect 1615 2415 1635 2435
rect 1665 2415 1685 2435
rect 1715 2415 1735 2435
rect 1765 2415 1785 2435
rect 1815 2415 1835 2435
rect 1865 2415 1885 2435
rect 1915 2415 1935 2435
rect 1965 2415 1985 2435
rect 2015 2415 2035 2435
rect 2065 2415 2085 2435
rect 2115 2415 2135 2435
rect 2165 2415 2185 2435
rect 2215 2415 2235 2435
rect 2265 2415 2285 2435
rect 2315 2415 2335 2435
rect 2365 2415 2385 2435
rect 2415 2415 2435 2435
rect 2465 2415 2485 2435
rect 2515 2415 2535 2435
rect 2565 2415 2585 2435
rect 2615 2415 2635 2435
rect 2665 2415 2685 2435
rect 2715 2415 2735 2435
rect 2765 2415 2785 2435
rect 2815 2415 2835 2435
rect 2865 2415 2885 2435
rect 2915 2415 2935 2435
rect 2965 2415 2985 2435
rect 3015 2415 3035 2435
rect 3065 2415 3085 2435
rect 3115 2415 3135 2435
rect 3165 2415 3185 2435
rect 3215 2415 3235 2435
rect 3265 2415 3285 2435
rect 3315 2415 3335 2435
rect 3365 2415 3385 2435
rect 3415 2415 3435 2435
rect 3465 2415 3485 2435
rect 3515 2415 3535 2435
rect 3565 2415 3585 2435
rect 3615 2415 3635 2435
rect 3665 2415 3685 2435
rect 3715 2415 3735 2435
rect 3765 2415 3785 2435
rect 3815 2415 3835 2435
rect 3865 2415 3885 2435
rect 3915 2415 3935 2435
rect 3965 2415 3985 2435
rect 4015 2415 4035 2435
rect 4065 2415 4085 2435
rect 4115 2415 4135 2435
rect 4165 2415 4185 2435
rect 4215 2415 4235 2435
rect 4265 2415 4285 2435
rect 4315 2415 4335 2435
rect 4365 2415 4385 2435
rect 4415 2415 4435 2435
rect 4465 2415 4485 2435
rect 4515 2415 4535 2435
rect 4565 2415 4585 2435
rect 4615 2415 4635 2435
rect 4665 2415 4685 2435
rect 4715 2415 4735 2435
rect 4765 2415 4785 2435
rect 4815 2415 4835 2435
rect 4865 2415 4885 2435
rect 4915 2415 4935 2435
rect 4965 2415 4985 2435
rect 5015 2415 5035 2435
rect 5065 2415 5085 2435
rect 5115 2415 5135 2435
rect 5165 2415 5185 2435
rect 5215 2415 5235 2435
rect 5265 2415 5285 2435
rect 5315 2415 5335 2435
rect 5365 2415 5385 2435
rect 5415 2415 5435 2435
rect 5465 2415 5485 2435
rect 5515 2415 5535 2435
rect 5565 2415 5585 2435
rect 5615 2415 5635 2435
rect 5665 2415 5685 2435
rect 5715 2415 5735 2435
rect 5765 2415 5785 2435
rect 5815 2415 5835 2435
rect 5865 2415 5885 2435
rect 5915 2415 5935 2435
rect 5965 2415 5985 2435
rect 6015 2415 6035 2435
rect 6065 2415 6085 2435
rect 6115 2415 6135 2435
rect 6165 2415 6185 2435
rect 6215 2415 6235 2435
rect 6265 2415 6285 2435
rect 6315 2415 6335 2435
rect 6365 2415 6385 2435
rect 6415 2415 6435 2435
rect 6465 2415 6485 2435
rect 6515 2415 6535 2435
rect 6565 2415 6585 2435
rect 6615 2415 6635 2435
rect 6665 2415 6685 2435
rect 6715 2415 6735 2435
rect 6765 2415 6785 2435
rect 6815 2415 6835 2435
rect 6865 2415 6885 2435
rect 6915 2415 6935 2435
rect 6965 2415 6985 2435
rect 7015 2415 7035 2435
rect 7065 2415 7085 2435
rect 7115 2415 7135 2435
rect 7165 2415 7185 2435
rect 7215 2415 7235 2435
rect 7265 2415 7285 2435
rect 7315 2415 7335 2435
rect 7365 2415 7385 2435
rect 7415 2415 7435 2435
rect 7465 2415 7485 2435
rect 7515 2415 7535 2435
rect 7565 2415 7585 2435
rect 7615 2415 7635 2435
rect 7665 2415 7685 2435
rect 7715 2415 7735 2435
rect 7765 2415 7785 2435
rect 7815 2415 7835 2435
rect 7865 2415 7885 2435
rect 7915 2415 7935 2435
rect 7965 2415 7985 2435
rect 8015 2415 8035 2435
rect 8065 2415 8085 2435
rect 8115 2415 8135 2435
rect 8165 2415 8185 2435
rect 8215 2415 8235 2435
rect 8265 2415 8285 2435
rect 8315 2415 8335 2435
rect 8365 2415 8385 2435
rect 8415 2415 8435 2435
rect 8465 2415 8485 2435
rect 8515 2415 8535 2435
rect 8565 2415 8585 2435
rect 8615 2415 8635 2435
rect 8665 2415 8685 2435
rect 8715 2415 8735 2435
rect 8765 2415 8785 2435
rect 8815 2415 8835 2435
rect 8865 2415 8885 2435
rect 8915 2415 8935 2435
rect 8965 2415 8985 2435
rect 9015 2415 9035 2435
rect 9065 2415 9085 2435
rect 9115 2415 9135 2435
rect 9165 2415 9185 2435
rect 9215 2415 9235 2435
rect 9265 2415 9285 2435
rect 9315 2415 9335 2435
rect 9365 2415 9385 2435
rect 9415 2415 9435 2435
rect 9465 2415 9485 2435
rect 9515 2415 9535 2435
rect 9565 2415 9585 2435
rect 9615 2415 9635 2435
rect 9665 2415 9685 2435
rect 9715 2415 9735 2435
rect 9765 2415 9785 2435
rect 9815 2415 9835 2435
rect 9865 2415 9885 2435
rect 9915 2415 9935 2435
rect 9965 2415 9985 2435
rect 10015 2415 10035 2435
rect 10065 2415 10085 2435
rect 10115 2415 10135 2435
rect 10165 2415 10185 2435
rect 10215 2415 10235 2435
rect 10265 2415 10285 2435
rect 10315 2415 10335 2435
rect 10365 2415 10385 2435
rect 10415 2415 10435 2435
rect 10465 2415 10485 2435
rect 10515 2415 10535 2435
rect 10565 2415 10585 2435
rect 10615 2415 10635 2435
rect 10665 2415 10685 2435
rect 10715 2415 10735 2435
rect 10765 2415 10785 2435
rect 10815 2415 10835 2435
rect 10865 2415 10885 2435
rect 10915 2415 10935 2435
rect 10965 2415 10985 2435
rect 11015 2415 11035 2435
rect 11065 2415 11085 2435
rect 11115 2415 11135 2435
rect 11165 2415 11185 2435
rect 11215 2415 11235 2435
rect 11265 2415 11285 2435
rect 11315 2415 11335 2435
rect 11365 2415 11385 2435
rect 11415 2415 11435 2435
rect 11465 2415 11485 2435
rect 11515 2415 11535 2435
rect 11565 2415 11585 2435
rect 11615 2415 11635 2435
rect 11665 2415 11685 2435
rect 11715 2415 11735 2435
rect 11765 2415 11785 2435
rect 11815 2415 11835 2435
rect 11865 2415 11885 2435
rect 11915 2415 11935 2435
rect 11965 2415 11985 2435
rect 12015 2415 12035 2435
rect 12065 2415 12085 2435
rect 12115 2415 12135 2435
rect 12165 2415 12185 2435
rect 12215 2415 12235 2435
rect 12265 2415 12285 2435
rect 12315 2415 12335 2435
rect 12365 2415 12385 2435
rect 12415 2415 12435 2435
rect 12465 2415 12485 2435
rect 12515 2415 12535 2435
rect 12565 2415 12585 2435
rect 12615 2415 12635 2435
rect 12665 2415 12685 2435
rect 12715 2415 12735 2435
rect 12765 2415 12785 2435
rect 12815 2415 12835 2435
rect 12865 2415 12885 2435
rect 12915 2415 12935 2435
rect 12965 2415 12985 2435
rect 13015 2415 13035 2435
rect 13065 2415 13085 2435
rect 13115 2415 13135 2435
rect 13165 2415 13185 2435
rect 13215 2415 13235 2435
rect 13265 2415 13285 2435
rect 13315 2415 13335 2435
rect 13365 2415 13385 2435
rect 13415 2415 13435 2435
rect 13465 2415 13485 2435
rect 13515 2415 13535 2435
rect 13565 2415 13585 2435
rect 13615 2415 13635 2435
rect 13665 2415 13685 2435
rect 13715 2415 13735 2435
rect 13765 2415 13785 2435
rect 13815 2415 13835 2435
rect 13865 2415 13885 2435
rect 13915 2415 13935 2435
rect 13965 2415 13985 2435
rect 14015 2415 14035 2435
rect 14065 2415 14085 2435
rect 14115 2415 14135 2435
rect 14165 2415 14185 2435
rect 14215 2415 14235 2435
rect 14265 2415 14285 2435
rect 14315 2415 14335 2435
rect 14365 2415 14385 2435
rect 14415 2415 14435 2435
rect 14465 2415 14485 2435
rect 14515 2415 14535 2435
rect 14565 2415 14585 2435
rect 14615 2415 14635 2435
rect 14665 2415 14685 2435
rect 14715 2415 14735 2435
rect 14765 2415 14785 2435
rect 14815 2415 14835 2435
rect 14865 2415 14885 2435
rect 14915 2415 14935 2435
rect 14965 2415 14985 2435
rect 15015 2415 15035 2435
rect 15065 2415 15085 2435
rect 15115 2415 15135 2435
rect 15165 2415 15185 2435
rect 15215 2415 15235 2435
rect 15265 2415 15285 2435
rect 15315 2415 15335 2435
rect 15365 2415 15385 2435
rect 15415 2415 15435 2435
rect 15465 2415 15485 2435
rect 15515 2415 15535 2435
rect 15565 2415 15585 2435
rect 15615 2415 15635 2435
rect 15665 2415 15685 2435
rect 15715 2415 15735 2435
rect 15765 2415 15785 2435
rect 15815 2415 15835 2435
rect 15865 2415 15885 2435
rect 15915 2415 15935 2435
rect 15965 2415 15985 2435
rect 16015 2415 16035 2435
rect 16065 2415 16085 2435
rect 16115 2415 16135 2435
rect 16165 2415 16185 2435
rect 16215 2415 16235 2435
rect 16265 2415 16285 2435
rect 16315 2415 16335 2435
rect 16365 2415 16385 2435
rect 16415 2415 16435 2435
rect 16465 2415 16485 2435
rect 16515 2415 16535 2435
rect 16565 2415 16585 2435
rect 16615 2415 16635 2435
rect 16665 2415 16685 2435
rect 16715 2415 16735 2435
rect 16765 2415 16785 2435
rect 16815 2415 16835 2435
rect 16865 2415 16885 2435
rect 16915 2415 16935 2435
rect 16965 2415 16985 2435
rect 17015 2415 17035 2435
rect 17065 2415 17085 2435
rect 17115 2415 17135 2435
rect 17165 2415 17185 2435
rect 17215 2415 17235 2435
rect 17265 2415 17285 2435
rect 17315 2415 17335 2435
rect 17365 2415 17385 2435
rect 17415 2415 17435 2435
rect 17465 2415 17485 2435
rect 17515 2415 17535 2435
rect 17565 2415 17585 2435
rect 17615 2415 17635 2435
rect 17665 2415 17685 2435
rect 17715 2415 17735 2435
rect 17765 2415 17785 2435
rect 17815 2415 17835 2435
rect 17865 2415 17885 2435
rect 17915 2415 17935 2435
rect 17965 2415 17985 2435
rect 18015 2415 18035 2435
rect 18065 2415 18085 2435
rect 18115 2415 18135 2435
rect 18165 2415 18185 2435
rect 18215 2415 18235 2435
rect 18265 2415 18285 2435
rect 18315 2415 18335 2435
rect 18365 2415 18385 2435
rect 18415 2415 18435 2435
rect 18465 2415 18485 2435
rect 18515 2415 18535 2435
rect 18565 2415 18585 2435
rect 18615 2415 18635 2435
rect 18665 2415 18685 2435
rect 18715 2415 18735 2435
rect 18765 2415 18785 2435
rect 18815 2415 18835 2435
rect 18865 2415 18885 2435
rect 18915 2415 18935 2435
rect 18965 2415 18985 2435
rect 19015 2415 19035 2435
rect 19065 2415 19085 2435
rect 19115 2415 19135 2435
rect 19165 2415 19185 2435
rect 19215 2415 19235 2435
rect 19265 2415 19285 2435
rect 19315 2415 19335 2435
rect 19365 2415 19385 2435
rect 19415 2415 19435 2435
rect 19465 2415 19485 2435
rect 19515 2415 19535 2435
rect 19565 2415 19585 2435
rect 19615 2415 19635 2435
rect 19665 2415 19685 2435
rect 19715 2415 19735 2435
rect 19765 2415 19785 2435
rect 19815 2415 19835 2435
rect 19865 2415 19885 2435
rect 19915 2415 19935 2435
rect 19965 2415 19985 2435
rect 20015 2415 20035 2435
rect 20065 2415 20085 2435
rect 20115 2415 20135 2435
rect 20165 2415 20185 2435
rect 20215 2415 20235 2435
rect 20265 2415 20285 2435
rect 20315 2415 20335 2435
rect 20365 2415 20385 2435
rect -885 2015 -865 2035
rect -835 2015 -815 2035
rect -785 2015 -765 2035
rect -735 2015 -715 2035
rect -685 2015 -665 2035
rect -635 2015 -615 2035
rect -585 2015 -565 2035
rect -535 2015 -515 2035
rect -485 2015 -465 2035
rect -435 2015 -415 2035
rect -385 2015 -365 2035
rect -335 2015 -315 2035
rect -285 2015 -265 2035
rect -235 2015 -215 2035
rect -185 2015 -165 2035
rect -135 2015 -115 2035
rect -85 2015 -65 2035
rect -35 2015 -15 2035
rect 15 2015 35 2035
rect 65 2015 85 2035
rect 115 2015 135 2035
rect 165 2015 185 2035
rect 215 2015 235 2035
rect 265 2015 285 2035
rect 315 2015 335 2035
rect 365 2015 385 2035
rect 415 2015 435 2035
rect 465 2015 485 2035
rect 515 2015 535 2035
rect 565 2015 585 2035
rect 615 2015 635 2035
rect 665 2015 685 2035
rect 715 2015 735 2035
rect 765 2015 785 2035
rect 815 2015 835 2035
rect 865 2015 885 2035
rect 915 2015 935 2035
rect 965 2015 985 2035
rect 1015 2015 1035 2035
rect 1065 2015 1085 2035
rect 1115 2015 1135 2035
rect 1165 2015 1185 2035
rect 1215 2015 1235 2035
rect 1265 2015 1285 2035
rect 1315 2015 1335 2035
rect 1365 2015 1385 2035
rect 1415 2015 1435 2035
rect 1465 2015 1485 2035
rect 1515 2015 1535 2035
rect 1565 2015 1585 2035
rect 1615 2015 1635 2035
rect 1665 2015 1685 2035
rect 1715 2015 1735 2035
rect 1765 2015 1785 2035
rect 1815 2015 1835 2035
rect 1865 2015 1885 2035
rect 1915 2015 1935 2035
rect 1965 2015 1985 2035
rect 2015 2015 2035 2035
rect 2065 2015 2085 2035
rect 2115 2015 2135 2035
rect 2165 2015 2185 2035
rect 2215 2015 2235 2035
rect 2265 2015 2285 2035
rect 2315 2015 2335 2035
rect 2365 2015 2385 2035
rect 2415 2015 2435 2035
rect 2465 2015 2485 2035
rect 2515 2015 2535 2035
rect 2565 2015 2585 2035
rect 2615 2015 2635 2035
rect 2665 2015 2685 2035
rect 2715 2015 2735 2035
rect 2765 2015 2785 2035
rect 2815 2015 2835 2035
rect 2865 2015 2885 2035
rect 2915 2015 2935 2035
rect 2965 2015 2985 2035
rect 3015 2015 3035 2035
rect 3065 2015 3085 2035
rect 3115 2015 3135 2035
rect 3165 2015 3185 2035
rect 3215 2015 3235 2035
rect 3265 2015 3285 2035
rect 3315 2015 3335 2035
rect 3365 2015 3385 2035
rect 3415 2015 3435 2035
rect 3465 2015 3485 2035
rect 3515 2015 3535 2035
rect 3565 2015 3585 2035
rect 3615 2015 3635 2035
rect 3665 2015 3685 2035
rect 3715 2015 3735 2035
rect 3765 2015 3785 2035
rect 3815 2015 3835 2035
rect 3865 2015 3885 2035
rect 3915 2015 3935 2035
rect 3965 2015 3985 2035
rect 4015 2015 4035 2035
rect 4065 2015 4085 2035
rect 4115 2015 4135 2035
rect 4165 2015 4185 2035
rect 4215 2015 4235 2035
rect 4265 2015 4285 2035
rect 4315 2015 4335 2035
rect 4365 2015 4385 2035
rect 4415 2015 4435 2035
rect 4465 2015 4485 2035
rect 4515 2015 4535 2035
rect 4565 2015 4585 2035
rect 4615 2015 4635 2035
rect 4665 2015 4685 2035
rect 4715 2015 4735 2035
rect 4765 2015 4785 2035
rect 4815 2015 4835 2035
rect 4865 2015 4885 2035
rect 4915 2015 4935 2035
rect 4965 2015 4985 2035
rect 5015 2015 5035 2035
rect 5065 2015 5085 2035
rect 5115 2015 5135 2035
rect 5165 2015 5185 2035
rect 5215 2015 5235 2035
rect 5265 2015 5285 2035
rect 5315 2015 5335 2035
rect 5365 2015 5385 2035
rect 5415 2015 5435 2035
rect 5465 2015 5485 2035
rect 5515 2015 5535 2035
rect 5565 2015 5585 2035
rect 5615 2015 5635 2035
rect 5665 2015 5685 2035
rect 5715 2015 5735 2035
rect 5765 2015 5785 2035
rect 5815 2015 5835 2035
rect 5865 2015 5885 2035
rect 5915 2015 5935 2035
rect 5965 2015 5985 2035
rect 6015 2015 6035 2035
rect 6065 2015 6085 2035
rect 6115 2015 6135 2035
rect 6165 2015 6185 2035
rect 6215 2015 6235 2035
rect 6265 2015 6285 2035
rect 6315 2015 6335 2035
rect 6365 2015 6385 2035
rect 6415 2015 6435 2035
rect 6465 2015 6485 2035
rect 6515 2015 6535 2035
rect 6565 2015 6585 2035
rect 6615 2015 6635 2035
rect 6665 2015 6685 2035
rect 6715 2015 6735 2035
rect 6765 2015 6785 2035
rect 6815 2015 6835 2035
rect 6865 2015 6885 2035
rect 6915 2015 6935 2035
rect 6965 2015 6985 2035
rect 7015 2015 7035 2035
rect 7065 2015 7085 2035
rect 7115 2015 7135 2035
rect 7165 2015 7185 2035
rect 7215 2015 7235 2035
rect 7265 2015 7285 2035
rect 7315 2015 7335 2035
rect 7365 2015 7385 2035
rect 7415 2015 7435 2035
rect 7465 2015 7485 2035
rect 7515 2015 7535 2035
rect 7565 2015 7585 2035
rect 7615 2015 7635 2035
rect 7665 2015 7685 2035
rect 7715 2015 7735 2035
rect 7765 2015 7785 2035
rect 7815 2015 7835 2035
rect 7865 2015 7885 2035
rect 7915 2015 7935 2035
rect 7965 2015 7985 2035
rect 8015 2015 8035 2035
rect 8065 2015 8085 2035
rect 8115 2015 8135 2035
rect 8165 2015 8185 2035
rect 8215 2015 8235 2035
rect 8265 2015 8285 2035
rect 8315 2015 8335 2035
rect 8365 2015 8385 2035
rect 8415 2015 8435 2035
rect 8465 2015 8485 2035
rect 8515 2015 8535 2035
rect 8565 2015 8585 2035
rect 8615 2015 8635 2035
rect 8665 2015 8685 2035
rect 8715 2015 8735 2035
rect 8765 2015 8785 2035
rect 8815 2015 8835 2035
rect 8865 2015 8885 2035
rect 8915 2015 8935 2035
rect 8965 2015 8985 2035
rect 9015 2015 9035 2035
rect 9065 2015 9085 2035
rect 9115 2015 9135 2035
rect 9165 2015 9185 2035
rect 9215 2015 9235 2035
rect 9265 2015 9285 2035
rect 9315 2015 9335 2035
rect 9365 2015 9385 2035
rect 9415 2015 9435 2035
rect 9465 2015 9485 2035
rect 9515 2015 9535 2035
rect 9565 2015 9585 2035
rect 9615 2015 9635 2035
rect 9665 2015 9685 2035
rect 9715 2015 9735 2035
rect 9765 2015 9785 2035
rect 9815 2015 9835 2035
rect 9865 2015 9885 2035
rect 9915 2015 9935 2035
rect 9965 2015 9985 2035
rect 10015 2015 10035 2035
rect 10065 2015 10085 2035
rect 10115 2015 10135 2035
rect 10165 2015 10185 2035
rect 10215 2015 10235 2035
rect 10265 2015 10285 2035
rect 10315 2015 10335 2035
rect 10365 2015 10385 2035
rect 10415 2015 10435 2035
rect 10465 2015 10485 2035
rect 10515 2015 10535 2035
rect 10565 2015 10585 2035
rect 10615 2015 10635 2035
rect 10665 2015 10685 2035
rect 10715 2015 10735 2035
rect 10765 2015 10785 2035
rect 10815 2015 10835 2035
rect 10865 2015 10885 2035
rect 10915 2015 10935 2035
rect 10965 2015 10985 2035
rect 11015 2015 11035 2035
rect 11065 2015 11085 2035
rect 11115 2015 11135 2035
rect 11165 2015 11185 2035
rect 11215 2015 11235 2035
rect 11265 2015 11285 2035
rect 11315 2015 11335 2035
rect 11365 2015 11385 2035
rect 11415 2015 11435 2035
rect 11465 2015 11485 2035
rect 11515 2015 11535 2035
rect 11565 2015 11585 2035
rect 11615 2015 11635 2035
rect 11665 2015 11685 2035
rect 11715 2015 11735 2035
rect 11765 2015 11785 2035
rect 11815 2015 11835 2035
rect 11865 2015 11885 2035
rect 11915 2015 11935 2035
rect 11965 2015 11985 2035
rect 12015 2015 12035 2035
rect 12065 2015 12085 2035
rect 12115 2015 12135 2035
rect 12165 2015 12185 2035
rect 12215 2015 12235 2035
rect 12265 2015 12285 2035
rect 12315 2015 12335 2035
rect 12365 2015 12385 2035
rect 12415 2015 12435 2035
rect 12465 2015 12485 2035
rect 12515 2015 12535 2035
rect 12565 2015 12585 2035
rect 12615 2015 12635 2035
rect 12665 2015 12685 2035
rect 12715 2015 12735 2035
rect 12765 2015 12785 2035
rect 12815 2015 12835 2035
rect 12865 2015 12885 2035
rect 12915 2015 12935 2035
rect 12965 2015 12985 2035
rect 13015 2015 13035 2035
rect 13065 2015 13085 2035
rect 13115 2015 13135 2035
rect 13165 2015 13185 2035
rect 13215 2015 13235 2035
rect 13265 2015 13285 2035
rect 13315 2015 13335 2035
rect 13365 2015 13385 2035
rect 13415 2015 13435 2035
rect 13465 2015 13485 2035
rect 13515 2015 13535 2035
rect 13565 2015 13585 2035
rect 13615 2015 13635 2035
rect 13665 2015 13685 2035
rect 13715 2015 13735 2035
rect 13765 2015 13785 2035
rect 13815 2015 13835 2035
rect 13865 2015 13885 2035
rect 13915 2015 13935 2035
rect 13965 2015 13985 2035
rect 14015 2015 14035 2035
rect 14065 2015 14085 2035
rect 14115 2015 14135 2035
rect 14165 2015 14185 2035
rect 14215 2015 14235 2035
rect 14265 2015 14285 2035
rect 14315 2015 14335 2035
rect 14365 2015 14385 2035
rect 14415 2015 14435 2035
rect 14465 2015 14485 2035
rect 14515 2015 14535 2035
rect 14565 2015 14585 2035
rect 14615 2015 14635 2035
rect 14665 2015 14685 2035
rect 14715 2015 14735 2035
rect 14765 2015 14785 2035
rect 14815 2015 14835 2035
rect 14865 2015 14885 2035
rect 14915 2015 14935 2035
rect 14965 2015 14985 2035
rect 15015 2015 15035 2035
rect 15065 2015 15085 2035
rect 15115 2015 15135 2035
rect 15165 2015 15185 2035
rect 15215 2015 15235 2035
rect 15265 2015 15285 2035
rect 15315 2015 15335 2035
rect 15365 2015 15385 2035
rect 15415 2015 15435 2035
rect 15465 2015 15485 2035
rect 15515 2015 15535 2035
rect 15565 2015 15585 2035
rect 15615 2015 15635 2035
rect 15665 2015 15685 2035
rect 15715 2015 15735 2035
rect 15765 2015 15785 2035
rect 15815 2015 15835 2035
rect 15865 2015 15885 2035
rect 15915 2015 15935 2035
rect 15965 2015 15985 2035
rect 16015 2015 16035 2035
rect 16065 2015 16085 2035
rect 16115 2015 16135 2035
rect 16165 2015 16185 2035
rect 16215 2015 16235 2035
rect 16265 2015 16285 2035
rect 16315 2015 16335 2035
rect 16365 2015 16385 2035
rect 16415 2015 16435 2035
rect 16465 2015 16485 2035
rect 16515 2015 16535 2035
rect 16565 2015 16585 2035
rect 16615 2015 16635 2035
rect 16665 2015 16685 2035
rect 16715 2015 16735 2035
rect 16765 2015 16785 2035
rect 16815 2015 16835 2035
rect 16865 2015 16885 2035
rect 16915 2015 16935 2035
rect 16965 2015 16985 2035
rect 17015 2015 17035 2035
rect 17065 2015 17085 2035
rect 17115 2015 17135 2035
rect 17165 2015 17185 2035
rect 17215 2015 17235 2035
rect 17265 2015 17285 2035
rect 17315 2015 17335 2035
rect 17365 2015 17385 2035
rect 17415 2015 17435 2035
rect 17465 2015 17485 2035
rect 17515 2015 17535 2035
rect 17565 2015 17585 2035
rect 17615 2015 17635 2035
rect 17665 2015 17685 2035
rect 17715 2015 17735 2035
rect 17765 2015 17785 2035
rect 17815 2015 17835 2035
rect 17865 2015 17885 2035
rect 17915 2015 17935 2035
rect 17965 2015 17985 2035
rect 18015 2015 18035 2035
rect 18065 2015 18085 2035
rect 18115 2015 18135 2035
rect 18165 2015 18185 2035
rect 18215 2015 18235 2035
rect 18265 2015 18285 2035
rect 18315 2015 18335 2035
rect 18365 2015 18385 2035
rect 18415 2015 18435 2035
rect 18465 2015 18485 2035
rect 18515 2015 18535 2035
rect 18565 2015 18585 2035
rect 18615 2015 18635 2035
rect 18665 2015 18685 2035
rect 18715 2015 18735 2035
rect 18765 2015 18785 2035
rect 18815 2015 18835 2035
rect 18865 2015 18885 2035
rect 18915 2015 18935 2035
rect 18965 2015 18985 2035
rect 19015 2015 19035 2035
rect 19065 2015 19085 2035
rect 19115 2015 19135 2035
rect 19165 2015 19185 2035
rect 19215 2015 19235 2035
rect 19265 2015 19285 2035
rect 19315 2015 19335 2035
rect 19365 2015 19385 2035
rect 19415 2015 19435 2035
rect 19465 2015 19485 2035
rect 19515 2015 19535 2035
rect 19565 2015 19585 2035
rect 19615 2015 19635 2035
rect 19665 2015 19685 2035
rect 19715 2015 19735 2035
rect 19765 2015 19785 2035
rect 19815 2015 19835 2035
rect 19865 2015 19885 2035
rect 19915 2015 19935 2035
rect 19965 2015 19985 2035
rect 20015 2015 20035 2035
rect 20065 2015 20085 2035
rect 20115 2015 20135 2035
rect 20165 2015 20185 2035
rect 20215 2015 20235 2035
rect 20265 2015 20285 2035
rect 20315 2015 20335 2035
rect 20365 2015 20385 2035
rect -635 1665 -615 1685
rect -585 1665 -565 1685
rect -535 1665 -515 1685
rect -485 1665 -465 1685
rect -435 1665 -415 1685
rect -385 1665 -365 1685
rect -335 1665 -315 1685
rect -285 1665 -265 1685
rect -235 1665 -215 1685
rect -185 1665 -165 1685
rect -135 1665 -115 1685
rect -85 1665 -65 1685
rect -35 1665 -15 1685
rect 15 1665 35 1685
rect 65 1665 85 1685
rect 115 1665 135 1685
rect 165 1665 185 1685
rect 215 1665 235 1685
rect 265 1665 285 1685
rect 315 1665 335 1685
rect 365 1665 385 1685
rect 415 1665 435 1685
rect 465 1665 485 1685
rect 515 1665 535 1685
rect 565 1665 585 1685
rect 615 1665 635 1685
rect 665 1665 685 1685
rect 715 1665 735 1685
rect 765 1665 785 1685
rect 815 1665 835 1685
rect 865 1665 885 1685
rect 915 1665 935 1685
rect 965 1665 985 1685
rect 1015 1665 1035 1685
rect 1065 1665 1085 1685
rect 1115 1665 1135 1685
rect 1165 1665 1185 1685
rect 1215 1665 1235 1685
rect 1265 1665 1285 1685
rect 1315 1665 1335 1685
rect 1365 1665 1385 1685
rect 1415 1665 1435 1685
rect 1465 1665 1485 1685
rect 1515 1665 1535 1685
rect 1565 1665 1585 1685
rect 1615 1665 1635 1685
rect 1665 1665 1685 1685
rect 1715 1665 1735 1685
rect 1765 1665 1785 1685
rect 1815 1665 1835 1685
rect 1865 1665 1885 1685
rect 1915 1665 1935 1685
rect 1965 1665 1985 1685
rect 2015 1665 2035 1685
rect 2065 1665 2085 1685
rect 2115 1665 2135 1685
rect 2165 1665 2185 1685
rect 2215 1665 2235 1685
rect 2265 1665 2285 1685
rect 2315 1665 2335 1685
rect 2365 1665 2385 1685
rect 2415 1665 2435 1685
rect 2465 1665 2485 1685
rect 2515 1665 2535 1685
rect 2565 1665 2585 1685
rect 2615 1665 2635 1685
rect 2665 1665 2685 1685
rect 2715 1665 2735 1685
rect 2765 1665 2785 1685
rect 2815 1665 2835 1685
rect 2865 1665 2885 1685
rect 2915 1665 2935 1685
rect 2965 1665 2985 1685
rect 3015 1665 3035 1685
rect 3065 1665 3085 1685
rect 3115 1665 3135 1685
rect 3165 1665 3185 1685
rect 3215 1665 3235 1685
rect 3265 1665 3285 1685
rect 3315 1665 3335 1685
rect 3365 1665 3385 1685
rect 3415 1665 3435 1685
rect 3465 1665 3485 1685
rect 3515 1665 3535 1685
rect 3565 1665 3585 1685
rect 3615 1665 3635 1685
rect 3665 1665 3685 1685
rect 3715 1665 3735 1685
rect 3765 1665 3785 1685
rect 3815 1665 3835 1685
rect 3865 1665 3885 1685
rect 3915 1665 3935 1685
rect 3965 1665 3985 1685
rect 4015 1665 4035 1685
rect 4065 1665 4085 1685
rect 4115 1665 4135 1685
rect 4165 1665 4185 1685
rect 4215 1665 4235 1685
rect 4265 1665 4285 1685
rect 4315 1665 4335 1685
rect 4365 1665 4385 1685
rect 4415 1665 4435 1685
rect 4465 1665 4485 1685
rect 4515 1665 4535 1685
rect 4565 1665 4585 1685
rect 4615 1665 4635 1685
rect 4665 1665 4685 1685
rect 4715 1665 4735 1685
rect 4765 1665 4785 1685
rect 4815 1665 4835 1685
rect 4865 1665 4885 1685
rect 4915 1665 4935 1685
rect 4965 1665 4985 1685
rect 5015 1665 5035 1685
rect 5065 1665 5085 1685
rect 5115 1665 5135 1685
rect 5165 1665 5185 1685
rect 5215 1665 5235 1685
rect 5265 1665 5285 1685
rect 5315 1665 5335 1685
rect 5365 1665 5385 1685
rect 5415 1665 5435 1685
rect 5465 1665 5485 1685
rect 5515 1665 5535 1685
rect 5565 1665 5585 1685
rect 5615 1665 5635 1685
rect 5665 1665 5685 1685
rect 5715 1665 5735 1685
rect 5765 1665 5785 1685
rect 5815 1665 5835 1685
rect 5865 1665 5885 1685
rect 5915 1665 5935 1685
rect 5965 1665 5985 1685
rect 6015 1665 6035 1685
rect 6065 1665 6085 1685
rect 6115 1665 6135 1685
rect 6165 1665 6185 1685
rect 6215 1665 6235 1685
rect 6265 1665 6285 1685
rect 6315 1665 6335 1685
rect 6365 1665 6385 1685
rect 6415 1665 6435 1685
rect 6465 1665 6485 1685
rect 6515 1665 6535 1685
rect 6565 1665 6585 1685
rect 6615 1665 6635 1685
rect 6665 1665 6685 1685
rect 6715 1665 6735 1685
rect 6765 1665 6785 1685
rect 6815 1665 6835 1685
rect 6865 1665 6885 1685
rect 6915 1665 6935 1685
rect 6965 1665 6985 1685
rect 7015 1665 7035 1685
rect 7065 1665 7085 1685
rect 7115 1665 7135 1685
rect 7165 1665 7185 1685
rect 7215 1665 7235 1685
rect 7265 1665 7285 1685
rect 7315 1665 7335 1685
rect 7365 1665 7385 1685
rect 7415 1665 7435 1685
rect 7465 1665 7485 1685
rect 7515 1665 7535 1685
rect 7565 1665 7585 1685
rect 7615 1665 7635 1685
rect 7665 1665 7685 1685
rect 7715 1665 7735 1685
rect 7765 1665 7785 1685
rect 7815 1665 7835 1685
rect 7865 1665 7885 1685
rect 7915 1665 7935 1685
rect 7965 1665 7985 1685
rect 8015 1665 8035 1685
rect 8065 1665 8085 1685
rect 8115 1665 8135 1685
rect 8165 1665 8185 1685
rect 8215 1665 8235 1685
rect 8265 1665 8285 1685
rect 8315 1665 8335 1685
rect 8365 1665 8385 1685
rect 8415 1665 8435 1685
rect 8465 1665 8485 1685
rect 8515 1665 8535 1685
rect 8565 1665 8585 1685
rect 8615 1665 8635 1685
rect 8665 1665 8685 1685
rect 8715 1665 8735 1685
rect 8765 1665 8785 1685
rect 8815 1665 8835 1685
rect 8865 1665 8885 1685
rect 8915 1665 8935 1685
rect 8965 1665 8985 1685
rect 9015 1665 9035 1685
rect 9065 1665 9085 1685
rect 9115 1665 9135 1685
rect 9165 1665 9185 1685
rect 9215 1665 9235 1685
rect 9265 1665 9285 1685
rect 9315 1665 9335 1685
rect 9365 1665 9385 1685
rect 9415 1665 9435 1685
rect 9465 1665 9485 1685
rect 9515 1665 9535 1685
rect 9565 1665 9585 1685
rect 9615 1665 9635 1685
rect 9665 1665 9685 1685
rect 9715 1665 9735 1685
rect 9765 1665 9785 1685
rect 9815 1665 9835 1685
rect 9865 1665 9885 1685
rect 9915 1665 9935 1685
rect 9965 1665 9985 1685
rect 10015 1665 10035 1685
rect 10065 1665 10085 1685
rect 10115 1665 10135 1685
rect 10165 1665 10185 1685
rect 10215 1665 10235 1685
rect 10265 1665 10285 1685
rect 10315 1665 10335 1685
rect 10365 1665 10385 1685
rect 10415 1665 10435 1685
rect 10465 1665 10485 1685
rect 10515 1665 10535 1685
rect 10565 1665 10585 1685
rect 10615 1665 10635 1685
rect 10665 1665 10685 1685
rect 10715 1665 10735 1685
rect 10765 1665 10785 1685
rect 10815 1665 10835 1685
rect 10865 1665 10885 1685
rect 10915 1665 10935 1685
rect 10965 1665 10985 1685
rect 11015 1665 11035 1685
rect 11065 1665 11085 1685
rect 11115 1665 11135 1685
rect 11165 1665 11185 1685
rect 11215 1665 11235 1685
rect 11265 1665 11285 1685
rect 11315 1665 11335 1685
rect 11365 1665 11385 1685
rect 11415 1665 11435 1685
rect 11465 1665 11485 1685
rect 11515 1665 11535 1685
rect 11565 1665 11585 1685
rect 11615 1665 11635 1685
rect 11665 1665 11685 1685
rect 11715 1665 11735 1685
rect 11765 1665 11785 1685
rect 11815 1665 11835 1685
rect 11865 1665 11885 1685
rect 11915 1665 11935 1685
rect 11965 1665 11985 1685
rect 12015 1665 12035 1685
rect 12065 1665 12085 1685
rect 12115 1665 12135 1685
rect 12165 1665 12185 1685
rect 12215 1665 12235 1685
rect 12265 1665 12285 1685
rect 12315 1665 12335 1685
rect 12365 1665 12385 1685
rect 12415 1665 12435 1685
rect 12465 1665 12485 1685
rect 12515 1665 12535 1685
rect 12565 1665 12585 1685
rect 12615 1665 12635 1685
rect 12665 1665 12685 1685
rect 12715 1665 12735 1685
rect 12765 1665 12785 1685
rect 12815 1665 12835 1685
rect 12865 1665 12885 1685
rect 12915 1665 12935 1685
rect 12965 1665 12985 1685
rect 13015 1665 13035 1685
rect 13065 1665 13085 1685
rect 13115 1665 13135 1685
rect 13165 1665 13185 1685
rect 13215 1665 13235 1685
rect 13265 1665 13285 1685
rect 13315 1665 13335 1685
rect 13365 1665 13385 1685
rect 13415 1665 13435 1685
rect 13465 1665 13485 1685
rect 13515 1665 13535 1685
rect 13565 1665 13585 1685
rect 13615 1665 13635 1685
rect 13665 1665 13685 1685
rect 13715 1665 13735 1685
rect 13765 1665 13785 1685
rect 13815 1665 13835 1685
rect 13865 1665 13885 1685
rect 13915 1665 13935 1685
rect 13965 1665 13985 1685
rect 14015 1665 14035 1685
rect 14065 1665 14085 1685
rect 14115 1665 14135 1685
rect 14165 1665 14185 1685
rect 14215 1665 14235 1685
rect 14265 1665 14285 1685
rect 14315 1665 14335 1685
rect 14365 1665 14385 1685
rect 14415 1665 14435 1685
rect 14465 1665 14485 1685
rect 14515 1665 14535 1685
rect 14565 1665 14585 1685
rect 14615 1665 14635 1685
rect 14665 1665 14685 1685
rect 14715 1665 14735 1685
rect 14765 1665 14785 1685
rect 14815 1665 14835 1685
rect 14865 1665 14885 1685
rect 14915 1665 14935 1685
rect 14965 1665 14985 1685
rect 15015 1665 15035 1685
rect 15065 1665 15085 1685
rect 15115 1665 15135 1685
rect 15165 1665 15185 1685
rect 15215 1665 15235 1685
rect 15265 1665 15285 1685
rect 15315 1665 15335 1685
rect 15365 1665 15385 1685
rect 15415 1665 15435 1685
rect 15465 1665 15485 1685
rect 15515 1665 15535 1685
rect 15565 1665 15585 1685
rect 15615 1665 15635 1685
rect 15665 1665 15685 1685
rect 15715 1665 15735 1685
rect 15765 1665 15785 1685
rect 15815 1665 15835 1685
rect 15865 1665 15885 1685
rect 15915 1665 15935 1685
rect 15965 1665 15985 1685
rect 16015 1665 16035 1685
rect 16065 1665 16085 1685
rect 16115 1665 16135 1685
rect 16165 1665 16185 1685
rect 16215 1665 16235 1685
rect 16265 1665 16285 1685
rect 16315 1665 16335 1685
rect 16365 1665 16385 1685
rect 16415 1665 16435 1685
rect 16465 1665 16485 1685
rect 16515 1665 16535 1685
rect 16565 1665 16585 1685
rect 16615 1665 16635 1685
rect 16665 1665 16685 1685
rect 16715 1665 16735 1685
rect 16765 1665 16785 1685
rect 16815 1665 16835 1685
rect 16865 1665 16885 1685
rect 16915 1665 16935 1685
rect 16965 1665 16985 1685
rect 17015 1665 17035 1685
rect 17065 1665 17085 1685
rect 17115 1665 17135 1685
rect 17165 1665 17185 1685
rect 17215 1665 17235 1685
rect 17265 1665 17285 1685
rect 17315 1665 17335 1685
rect 17365 1665 17385 1685
rect 17415 1665 17435 1685
rect 17465 1665 17485 1685
rect 17515 1665 17535 1685
rect 17565 1665 17585 1685
rect 17615 1665 17635 1685
rect 17665 1665 17685 1685
rect 17715 1665 17735 1685
rect 17765 1665 17785 1685
rect 17815 1665 17835 1685
rect 17865 1665 17885 1685
rect 17915 1665 17935 1685
rect 17965 1665 17985 1685
rect 18015 1665 18035 1685
rect 18065 1665 18085 1685
rect 18115 1665 18135 1685
rect 18165 1665 18185 1685
rect 18215 1665 18235 1685
rect 18265 1665 18285 1685
rect 18315 1665 18335 1685
rect 18365 1665 18385 1685
rect 18415 1665 18435 1685
rect 18465 1665 18485 1685
rect 18515 1665 18535 1685
rect 18565 1665 18585 1685
rect 18615 1665 18635 1685
rect 18665 1665 18685 1685
rect 18715 1665 18735 1685
rect 18765 1665 18785 1685
rect 18815 1665 18835 1685
rect 18865 1665 18885 1685
rect 18915 1665 18935 1685
rect 18965 1665 18985 1685
rect 19015 1665 19035 1685
rect 19065 1665 19085 1685
rect 19115 1665 19135 1685
rect 19165 1665 19185 1685
rect 19215 1665 19235 1685
rect 19265 1665 19285 1685
rect 19315 1665 19335 1685
rect 19365 1665 19385 1685
rect 19415 1665 19435 1685
rect 19465 1665 19485 1685
rect 19515 1665 19535 1685
rect 19565 1665 19585 1685
rect 19615 1665 19635 1685
rect 19665 1665 19685 1685
rect 19715 1665 19735 1685
rect 19765 1665 19785 1685
rect 19815 1665 19835 1685
rect 19865 1665 19885 1685
rect 19915 1665 19935 1685
rect 19965 1665 19985 1685
rect 20015 1665 20035 1685
rect 20065 1665 20085 1685
rect 20115 1665 20135 1685
rect 20165 1665 20185 1685
rect 20215 1665 20235 1685
rect 20265 1665 20285 1685
rect 20315 1665 20335 1685
rect 20365 1665 20385 1685
rect -635 -35 -615 -15
rect -585 -35 -565 -15
rect -535 -35 -515 -15
rect -485 -35 -465 -15
rect -435 -35 -415 -15
rect -385 -35 -365 -15
rect -335 -35 -315 -15
rect -285 -35 -265 -15
rect -235 -35 -215 -15
rect -185 -35 -165 -15
rect -135 -35 -115 -15
rect -85 -35 -65 -15
rect -35 -35 -15 -15
rect 15 -35 35 -15
rect 65 -35 85 -15
rect 115 -35 135 -15
rect 165 -35 185 -15
rect 215 -35 235 -15
rect 265 -35 285 -15
rect 315 -35 335 -15
rect 365 -35 385 -15
rect 415 -35 435 -15
rect 465 -35 485 -15
rect 515 -35 535 -15
rect 565 -35 585 -15
rect 615 -35 635 -15
rect 665 -35 685 -15
rect 715 -35 735 -15
rect 765 -35 785 -15
rect 815 -35 835 -15
rect 865 -35 885 -15
rect 915 -35 935 -15
rect 965 -35 985 -15
rect 1015 -35 1035 -15
rect 1065 -35 1085 -15
rect 1115 -35 1135 -15
rect 1165 -35 1185 -15
rect 1215 -35 1235 -15
rect 1265 -35 1285 -15
rect 1315 -35 1335 -15
rect 1365 -35 1385 -15
rect 1415 -35 1435 -15
rect 1465 -35 1485 -15
rect 1515 -35 1535 -15
rect 1565 -35 1585 -15
rect 1615 -35 1635 -15
rect 1665 -35 1685 -15
rect 1715 -35 1735 -15
rect 1765 -35 1785 -15
rect 1815 -35 1835 -15
rect 1865 -35 1885 -15
rect 1915 -35 1935 -15
rect 1965 -35 1985 -15
rect 2015 -35 2035 -15
rect 2065 -35 2085 -15
rect 2115 -35 2135 -15
rect 2165 -35 2185 -15
rect 2215 -35 2235 -15
rect 2265 -35 2285 -15
rect 2315 -35 2335 -15
rect 2365 -35 2385 -15
rect 2415 -35 2435 -15
rect 2465 -35 2485 -15
rect 2515 -35 2535 -15
rect 2565 -35 2585 -15
rect 2615 -35 2635 -15
rect 2665 -35 2685 -15
rect 2715 -35 2735 -15
rect 2765 -35 2785 -15
rect 2815 -35 2835 -15
rect 2865 -35 2885 -15
rect 2915 -35 2935 -15
rect 2965 -35 2985 -15
rect 3015 -35 3035 -15
rect 3065 -35 3085 -15
rect 3115 -35 3135 -15
rect 3165 -35 3185 -15
rect 3215 -35 3235 -15
rect 3265 -35 3285 -15
rect 3315 -35 3335 -15
rect 3365 -35 3385 -15
rect 3415 -35 3435 -15
rect 3465 -35 3485 -15
rect 3515 -35 3535 -15
rect 3565 -35 3585 -15
rect 3615 -35 3635 -15
rect 3665 -35 3685 -15
rect 3715 -35 3735 -15
rect 3765 -35 3785 -15
rect 3815 -35 3835 -15
rect 3865 -35 3885 -15
rect 3915 -35 3935 -15
rect 3965 -35 3985 -15
rect 4015 -35 4035 -15
rect 4065 -35 4085 -15
rect 4115 -35 4135 -15
rect 4165 -35 4185 -15
rect 4215 -35 4235 -15
rect 4265 -35 4285 -15
rect 4315 -35 4335 -15
rect 4365 -35 4385 -15
rect 4415 -35 4435 -15
rect 4465 -35 4485 -15
rect 4515 -35 4535 -15
rect 4565 -35 4585 -15
rect 4615 -35 4635 -15
rect 4665 -35 4685 -15
rect 4715 -35 4735 -15
rect 4765 -35 4785 -15
rect 4815 -35 4835 -15
rect 4865 -35 4885 -15
rect 4915 -35 4935 -15
rect 4965 -35 4985 -15
rect 5015 -35 5035 -15
rect 5065 -35 5085 -15
rect 5115 -35 5135 -15
rect 5165 -35 5185 -15
rect 5215 -35 5235 -15
rect 5265 -35 5285 -15
rect 5315 -35 5335 -15
rect 5365 -35 5385 -15
rect 5415 -35 5435 -15
rect 5465 -35 5485 -15
rect 5515 -35 5535 -15
rect 5565 -35 5585 -15
rect 5615 -35 5635 -15
rect 5665 -35 5685 -15
rect 5715 -35 5735 -15
rect 5765 -35 5785 -15
rect 5815 -35 5835 -15
rect 5865 -35 5885 -15
rect 5915 -35 5935 -15
rect 5965 -35 5985 -15
rect 6015 -35 6035 -15
rect 6065 -35 6085 -15
rect 6115 -35 6135 -15
rect 6165 -35 6185 -15
rect 6215 -35 6235 -15
rect 6265 -35 6285 -15
rect 6315 -35 6335 -15
rect 6365 -35 6385 -15
rect 6415 -35 6435 -15
rect 6465 -35 6485 -15
rect 6515 -35 6535 -15
rect 6565 -35 6585 -15
rect 6615 -35 6635 -15
rect 6665 -35 6685 -15
rect 6715 -35 6735 -15
rect 6765 -35 6785 -15
rect 6815 -35 6835 -15
rect 6865 -35 6885 -15
rect 6915 -35 6935 -15
rect 6965 -35 6985 -15
rect 7015 -35 7035 -15
rect 7065 -35 7085 -15
rect 7115 -35 7135 -15
rect 7165 -35 7185 -15
rect 7215 -35 7235 -15
rect 7265 -35 7285 -15
rect 7315 -35 7335 -15
rect 7365 -35 7385 -15
rect 7415 -35 7435 -15
rect 7465 -35 7485 -15
rect 7515 -35 7535 -15
rect 7565 -35 7585 -15
rect 7615 -35 7635 -15
rect 7665 -35 7685 -15
rect 7715 -35 7735 -15
rect 7765 -35 7785 -15
rect 7815 -35 7835 -15
rect 7865 -35 7885 -15
rect 7915 -35 7935 -15
rect 7965 -35 7985 -15
rect 8015 -35 8035 -15
rect 8065 -35 8085 -15
rect 8115 -35 8135 -15
rect 8165 -35 8185 -15
rect 8215 -35 8235 -15
rect 8265 -35 8285 -15
rect 8315 -35 8335 -15
rect 8365 -35 8385 -15
rect 8415 -35 8435 -15
rect 8465 -35 8485 -15
rect 8515 -35 8535 -15
rect 8565 -35 8585 -15
rect 8615 -35 8635 -15
rect 8665 -35 8685 -15
rect 8715 -35 8735 -15
rect 8765 -35 8785 -15
rect 8815 -35 8835 -15
rect 8865 -35 8885 -15
rect 8915 -35 8935 -15
rect 8965 -35 8985 -15
rect 9015 -35 9035 -15
rect 9065 -35 9085 -15
rect 9115 -35 9135 -15
rect 9165 -35 9185 -15
rect 9215 -35 9235 -15
rect 9265 -35 9285 -15
rect 9315 -35 9335 -15
rect 9365 -35 9385 -15
rect 9415 -35 9435 -15
rect 9465 -35 9485 -15
rect 9515 -35 9535 -15
rect 9565 -35 9585 -15
rect 9615 -35 9635 -15
rect 9665 -35 9685 -15
rect 9715 -35 9735 -15
rect 9765 -35 9785 -15
rect 9815 -35 9835 -15
rect 9865 -35 9885 -15
rect 9915 -35 9935 -15
rect 9965 -35 9985 -15
rect 10015 -35 10035 -15
rect 10065 -35 10085 -15
rect 10115 -35 10135 -15
rect 10165 -35 10185 -15
rect 10215 -35 10235 -15
rect 10265 -35 10285 -15
rect 10315 -35 10335 -15
rect 10365 -35 10385 -15
rect 10415 -35 10435 -15
rect 10465 -35 10485 -15
rect 10515 -35 10535 -15
rect 10565 -35 10585 -15
rect 10615 -35 10635 -15
rect 10665 -35 10685 -15
rect 10715 -35 10735 -15
rect 10765 -35 10785 -15
rect 10815 -35 10835 -15
rect 10865 -35 10885 -15
rect 10915 -35 10935 -15
rect 10965 -35 10985 -15
rect 11015 -35 11035 -15
rect 11065 -35 11085 -15
rect 11115 -35 11135 -15
rect 11165 -35 11185 -15
rect 11215 -35 11235 -15
rect 11265 -35 11285 -15
rect 11315 -35 11335 -15
rect 11365 -35 11385 -15
rect 11415 -35 11435 -15
rect 11465 -35 11485 -15
rect 11515 -35 11535 -15
rect 11565 -35 11585 -15
rect 11615 -35 11635 -15
rect 11665 -35 11685 -15
rect 11715 -35 11735 -15
rect 11765 -35 11785 -15
rect 11815 -35 11835 -15
rect 11865 -35 11885 -15
rect 11915 -35 11935 -15
rect 11965 -35 11985 -15
rect 12015 -35 12035 -15
rect 12065 -35 12085 -15
rect 12115 -35 12135 -15
rect 12165 -35 12185 -15
rect 12215 -35 12235 -15
rect 12265 -35 12285 -15
rect 12315 -35 12335 -15
rect 12365 -35 12385 -15
rect 12415 -35 12435 -15
rect 12465 -35 12485 -15
rect 12515 -35 12535 -15
rect 12565 -35 12585 -15
rect 12615 -35 12635 -15
rect 12665 -35 12685 -15
rect 12715 -35 12735 -15
rect 12765 -35 12785 -15
rect 12815 -35 12835 -15
rect 12865 -35 12885 -15
rect 12915 -35 12935 -15
rect 12965 -35 12985 -15
rect 13015 -35 13035 -15
rect 13065 -35 13085 -15
rect 13115 -35 13135 -15
rect 13165 -35 13185 -15
rect 13215 -35 13235 -15
rect 13265 -35 13285 -15
rect 13315 -35 13335 -15
rect 13365 -35 13385 -15
rect 13415 -35 13435 -15
rect 13465 -35 13485 -15
rect 13515 -35 13535 -15
rect 13565 -35 13585 -15
rect 13615 -35 13635 -15
rect 13665 -35 13685 -15
rect 13715 -35 13735 -15
rect 13765 -35 13785 -15
rect 13815 -35 13835 -15
rect 13865 -35 13885 -15
rect 13915 -35 13935 -15
rect 13965 -35 13985 -15
rect 14015 -35 14035 -15
rect 14065 -35 14085 -15
rect 14115 -35 14135 -15
rect 14165 -35 14185 -15
rect 14215 -35 14235 -15
rect 14265 -35 14285 -15
rect 14315 -35 14335 -15
rect 14365 -35 14385 -15
rect 14415 -35 14435 -15
rect 14465 -35 14485 -15
rect 14515 -35 14535 -15
rect 14565 -35 14585 -15
rect 14615 -35 14635 -15
rect 14665 -35 14685 -15
rect 14715 -35 14735 -15
rect 14765 -35 14785 -15
rect 14815 -35 14835 -15
rect 14865 -35 14885 -15
rect 14915 -35 14935 -15
rect 14965 -35 14985 -15
rect 15015 -35 15035 -15
rect 15065 -35 15085 -15
rect 15115 -35 15135 -15
rect 15165 -35 15185 -15
rect 15215 -35 15235 -15
rect 15265 -35 15285 -15
rect 15315 -35 15335 -15
rect 15365 -35 15385 -15
rect 15415 -35 15435 -15
rect 15465 -35 15485 -15
rect 15515 -35 15535 -15
rect 15565 -35 15585 -15
rect 15615 -35 15635 -15
rect 15665 -35 15685 -15
rect 15715 -35 15735 -15
rect 15765 -35 15785 -15
rect 15815 -35 15835 -15
rect 15865 -35 15885 -15
rect 15915 -35 15935 -15
rect 15965 -35 15985 -15
rect 16015 -35 16035 -15
rect 16065 -35 16085 -15
rect 16115 -35 16135 -15
rect 16165 -35 16185 -15
rect 16215 -35 16235 -15
rect 16265 -35 16285 -15
rect 16315 -35 16335 -15
rect 16365 -35 16385 -15
rect 16415 -35 16435 -15
rect 16465 -35 16485 -15
rect 16515 -35 16535 -15
rect 16565 -35 16585 -15
rect 16615 -35 16635 -15
rect 16665 -35 16685 -15
rect 16715 -35 16735 -15
rect 16765 -35 16785 -15
rect 16815 -35 16835 -15
rect 16865 -35 16885 -15
rect 16915 -35 16935 -15
rect 16965 -35 16985 -15
rect 17015 -35 17035 -15
rect 17065 -35 17085 -15
rect 17115 -35 17135 -15
rect 17165 -35 17185 -15
rect 17215 -35 17235 -15
rect 17265 -35 17285 -15
rect 17315 -35 17335 -15
rect 17365 -35 17385 -15
rect 17415 -35 17435 -15
rect 17465 -35 17485 -15
rect 17515 -35 17535 -15
rect 17565 -35 17585 -15
rect 17615 -35 17635 -15
rect 17665 -35 17685 -15
rect 17715 -35 17735 -15
rect 17765 -35 17785 -15
rect 17815 -35 17835 -15
rect 17865 -35 17885 -15
rect 17915 -35 17935 -15
rect 17965 -35 17985 -15
rect 18015 -35 18035 -15
rect 18065 -35 18085 -15
rect 18115 -35 18135 -15
rect 18165 -35 18185 -15
rect 18215 -35 18235 -15
rect 18265 -35 18285 -15
rect 18315 -35 18335 -15
rect 18365 -35 18385 -15
rect 18415 -35 18435 -15
rect 18465 -35 18485 -15
rect 18515 -35 18535 -15
rect 18565 -35 18585 -15
rect 18615 -35 18635 -15
rect 18665 -35 18685 -15
rect 18715 -35 18735 -15
rect 18765 -35 18785 -15
rect 18815 -35 18835 -15
rect 18865 -35 18885 -15
rect 18915 -35 18935 -15
rect 18965 -35 18985 -15
rect 19015 -35 19035 -15
rect 19065 -35 19085 -15
rect 19115 -35 19135 -15
rect 19165 -35 19185 -15
rect 19215 -35 19235 -15
rect 19265 -35 19285 -15
rect 19315 -35 19335 -15
rect 19365 -35 19385 -15
rect 19415 -35 19435 -15
rect 19465 -35 19485 -15
rect 19515 -35 19535 -15
rect 19565 -35 19585 -15
rect 19615 -35 19635 -15
rect 19665 -35 19685 -15
rect 19715 -35 19735 -15
rect 19765 -35 19785 -15
rect 19815 -35 19835 -15
rect 19865 -35 19885 -15
rect 19915 -35 19935 -15
rect 19965 -35 19985 -15
rect 20015 -35 20035 -15
rect 20065 -35 20085 -15
rect 20115 -35 20135 -15
rect 20165 -35 20185 -15
rect 20215 -35 20235 -15
rect 20265 -35 20285 -15
rect 20315 -35 20335 -15
rect 20365 -35 20385 -15
rect -635 -1735 -615 -1715
rect -585 -1735 -565 -1715
rect -535 -1735 -515 -1715
rect -485 -1735 -465 -1715
rect -435 -1735 -415 -1715
rect -385 -1735 -365 -1715
rect -335 -1735 -315 -1715
rect -285 -1735 -265 -1715
rect -235 -1735 -215 -1715
rect -185 -1735 -165 -1715
rect -135 -1735 -115 -1715
rect -85 -1735 -65 -1715
rect -35 -1735 -15 -1715
rect 15 -1735 35 -1715
rect 65 -1735 85 -1715
rect 115 -1735 135 -1715
rect 165 -1735 185 -1715
rect 215 -1735 235 -1715
rect 265 -1735 285 -1715
rect 315 -1735 335 -1715
rect 365 -1735 385 -1715
rect 415 -1735 435 -1715
rect 465 -1735 485 -1715
rect 515 -1735 535 -1715
rect 565 -1735 585 -1715
rect 615 -1735 635 -1715
rect 665 -1735 685 -1715
rect 715 -1735 735 -1715
rect 765 -1735 785 -1715
rect 815 -1735 835 -1715
rect 865 -1735 885 -1715
rect 915 -1735 935 -1715
rect 965 -1735 985 -1715
rect 1015 -1735 1035 -1715
rect 1065 -1735 1085 -1715
rect 1115 -1735 1135 -1715
rect 1165 -1735 1185 -1715
rect 1215 -1735 1235 -1715
rect 1265 -1735 1285 -1715
rect 1315 -1735 1335 -1715
rect 1365 -1735 1385 -1715
rect 1415 -1735 1435 -1715
rect 1465 -1735 1485 -1715
rect 1515 -1735 1535 -1715
rect 1565 -1735 1585 -1715
rect 1615 -1735 1635 -1715
rect 1665 -1735 1685 -1715
rect 1715 -1735 1735 -1715
rect 1765 -1735 1785 -1715
rect 1815 -1735 1835 -1715
rect 1865 -1735 1885 -1715
rect 1915 -1735 1935 -1715
rect 1965 -1735 1985 -1715
rect 2015 -1735 2035 -1715
rect 2065 -1735 2085 -1715
rect 2115 -1735 2135 -1715
rect 2165 -1735 2185 -1715
rect 2215 -1735 2235 -1715
rect 2265 -1735 2285 -1715
rect 2315 -1735 2335 -1715
rect 2365 -1735 2385 -1715
rect 2415 -1735 2435 -1715
rect 2465 -1735 2485 -1715
rect 2515 -1735 2535 -1715
rect 2565 -1735 2585 -1715
rect 2615 -1735 2635 -1715
rect 2665 -1735 2685 -1715
rect 2715 -1735 2735 -1715
rect 2765 -1735 2785 -1715
rect 2815 -1735 2835 -1715
rect 2865 -1735 2885 -1715
rect 2915 -1735 2935 -1715
rect 2965 -1735 2985 -1715
rect 3015 -1735 3035 -1715
rect 3065 -1735 3085 -1715
rect 3115 -1735 3135 -1715
rect 3165 -1735 3185 -1715
rect 3215 -1735 3235 -1715
rect 3265 -1735 3285 -1715
rect 3315 -1735 3335 -1715
rect 3365 -1735 3385 -1715
rect 3415 -1735 3435 -1715
rect 3465 -1735 3485 -1715
rect 3515 -1735 3535 -1715
rect 3565 -1735 3585 -1715
rect 3615 -1735 3635 -1715
rect 3665 -1735 3685 -1715
rect 3715 -1735 3735 -1715
rect 3765 -1735 3785 -1715
rect 3815 -1735 3835 -1715
rect 3865 -1735 3885 -1715
rect 3915 -1735 3935 -1715
rect 3965 -1735 3985 -1715
rect 4015 -1735 4035 -1715
rect 4065 -1735 4085 -1715
rect 4115 -1735 4135 -1715
rect 4165 -1735 4185 -1715
rect 4215 -1735 4235 -1715
rect 4265 -1735 4285 -1715
rect 4315 -1735 4335 -1715
rect 4365 -1735 4385 -1715
rect 4415 -1735 4435 -1715
rect 4465 -1735 4485 -1715
rect 4515 -1735 4535 -1715
rect 4565 -1735 4585 -1715
rect 4615 -1735 4635 -1715
rect 4665 -1735 4685 -1715
rect 4715 -1735 4735 -1715
rect 4765 -1735 4785 -1715
rect 4815 -1735 4835 -1715
rect 4865 -1735 4885 -1715
rect 4915 -1735 4935 -1715
rect 4965 -1735 4985 -1715
rect 5015 -1735 5035 -1715
rect 5065 -1735 5085 -1715
rect 5115 -1735 5135 -1715
rect 5165 -1735 5185 -1715
rect 5215 -1735 5235 -1715
rect 5265 -1735 5285 -1715
rect 5315 -1735 5335 -1715
rect 5365 -1735 5385 -1715
rect 5415 -1735 5435 -1715
rect 5465 -1735 5485 -1715
rect 5515 -1735 5535 -1715
rect 5565 -1735 5585 -1715
rect 5615 -1735 5635 -1715
rect 5665 -1735 5685 -1715
rect 5715 -1735 5735 -1715
rect 5765 -1735 5785 -1715
rect 5815 -1735 5835 -1715
rect 5865 -1735 5885 -1715
rect 5915 -1735 5935 -1715
rect 5965 -1735 5985 -1715
rect 6015 -1735 6035 -1715
rect 6065 -1735 6085 -1715
rect 6115 -1735 6135 -1715
rect 6165 -1735 6185 -1715
rect 6215 -1735 6235 -1715
rect 6265 -1735 6285 -1715
rect 6315 -1735 6335 -1715
rect 6365 -1735 6385 -1715
rect 6415 -1735 6435 -1715
rect 6465 -1735 6485 -1715
rect 6515 -1735 6535 -1715
rect 6565 -1735 6585 -1715
rect 6615 -1735 6635 -1715
rect 6665 -1735 6685 -1715
rect 6715 -1735 6735 -1715
rect 6765 -1735 6785 -1715
rect 6815 -1735 6835 -1715
rect 6865 -1735 6885 -1715
rect 6915 -1735 6935 -1715
rect 6965 -1735 6985 -1715
rect 7015 -1735 7035 -1715
rect 7065 -1735 7085 -1715
rect 7115 -1735 7135 -1715
rect 7165 -1735 7185 -1715
rect 7215 -1735 7235 -1715
rect 7265 -1735 7285 -1715
rect 7315 -1735 7335 -1715
rect 7365 -1735 7385 -1715
rect 7415 -1735 7435 -1715
rect 7465 -1735 7485 -1715
rect 7515 -1735 7535 -1715
rect 7565 -1735 7585 -1715
rect 7615 -1735 7635 -1715
rect 7665 -1735 7685 -1715
rect 7715 -1735 7735 -1715
rect 7765 -1735 7785 -1715
rect 7815 -1735 7835 -1715
rect 7865 -1735 7885 -1715
rect 7915 -1735 7935 -1715
rect 7965 -1735 7985 -1715
rect 8015 -1735 8035 -1715
rect 8065 -1735 8085 -1715
rect 8115 -1735 8135 -1715
rect 8165 -1735 8185 -1715
rect 8215 -1735 8235 -1715
rect 8265 -1735 8285 -1715
rect 8315 -1735 8335 -1715
rect 8365 -1735 8385 -1715
rect 8415 -1735 8435 -1715
rect 8465 -1735 8485 -1715
rect 8515 -1735 8535 -1715
rect 8565 -1735 8585 -1715
rect 8615 -1735 8635 -1715
rect 8665 -1735 8685 -1715
rect 8715 -1735 8735 -1715
rect 8765 -1735 8785 -1715
rect 8815 -1735 8835 -1715
rect 8865 -1735 8885 -1715
rect 8915 -1735 8935 -1715
rect 8965 -1735 8985 -1715
rect 9015 -1735 9035 -1715
rect 9065 -1735 9085 -1715
rect 9115 -1735 9135 -1715
rect 9165 -1735 9185 -1715
rect 9215 -1735 9235 -1715
rect 9265 -1735 9285 -1715
rect 9315 -1735 9335 -1715
rect 9365 -1735 9385 -1715
rect 9415 -1735 9435 -1715
rect 9465 -1735 9485 -1715
rect 9515 -1735 9535 -1715
rect 9565 -1735 9585 -1715
rect 9615 -1735 9635 -1715
rect 9665 -1735 9685 -1715
rect 9715 -1735 9735 -1715
rect 9765 -1735 9785 -1715
rect 9815 -1735 9835 -1715
rect 9865 -1735 9885 -1715
rect 9915 -1735 9935 -1715
rect 9965 -1735 9985 -1715
rect 10015 -1735 10035 -1715
rect 10065 -1735 10085 -1715
rect 10115 -1735 10135 -1715
rect 10165 -1735 10185 -1715
rect 10215 -1735 10235 -1715
rect 10265 -1735 10285 -1715
rect 10315 -1735 10335 -1715
rect 10365 -1735 10385 -1715
rect 10415 -1735 10435 -1715
rect 10465 -1735 10485 -1715
rect 10515 -1735 10535 -1715
rect 10565 -1735 10585 -1715
rect 10615 -1735 10635 -1715
rect 10665 -1735 10685 -1715
rect 10715 -1735 10735 -1715
rect 10765 -1735 10785 -1715
rect 10815 -1735 10835 -1715
rect 10865 -1735 10885 -1715
rect 10915 -1735 10935 -1715
rect 10965 -1735 10985 -1715
rect 11015 -1735 11035 -1715
rect 11065 -1735 11085 -1715
rect 11115 -1735 11135 -1715
rect 11165 -1735 11185 -1715
rect 11215 -1735 11235 -1715
rect 11265 -1735 11285 -1715
rect 11315 -1735 11335 -1715
rect 11365 -1735 11385 -1715
rect 11415 -1735 11435 -1715
rect 11465 -1735 11485 -1715
rect 11515 -1735 11535 -1715
rect 11565 -1735 11585 -1715
rect 11615 -1735 11635 -1715
rect 11665 -1735 11685 -1715
rect 11715 -1735 11735 -1715
rect 11765 -1735 11785 -1715
rect 11815 -1735 11835 -1715
rect 11865 -1735 11885 -1715
rect 11915 -1735 11935 -1715
rect 11965 -1735 11985 -1715
rect 12015 -1735 12035 -1715
rect 12065 -1735 12085 -1715
rect 12115 -1735 12135 -1715
rect 12165 -1735 12185 -1715
rect 12215 -1735 12235 -1715
rect 12265 -1735 12285 -1715
rect 12315 -1735 12335 -1715
rect 12365 -1735 12385 -1715
rect 12415 -1735 12435 -1715
rect 12465 -1735 12485 -1715
rect 12515 -1735 12535 -1715
rect 12565 -1735 12585 -1715
rect 12615 -1735 12635 -1715
rect 12665 -1735 12685 -1715
rect 12715 -1735 12735 -1715
rect 12765 -1735 12785 -1715
rect 12815 -1735 12835 -1715
rect 12865 -1735 12885 -1715
rect 12915 -1735 12935 -1715
rect 12965 -1735 12985 -1715
rect 13015 -1735 13035 -1715
rect 13065 -1735 13085 -1715
rect 13115 -1735 13135 -1715
rect 13165 -1735 13185 -1715
rect 13215 -1735 13235 -1715
rect 13265 -1735 13285 -1715
rect 13315 -1735 13335 -1715
rect 13365 -1735 13385 -1715
rect 13415 -1735 13435 -1715
rect 13465 -1735 13485 -1715
rect 13515 -1735 13535 -1715
rect 13565 -1735 13585 -1715
rect 13615 -1735 13635 -1715
rect 13665 -1735 13685 -1715
rect 13715 -1735 13735 -1715
rect 13765 -1735 13785 -1715
rect 13815 -1735 13835 -1715
rect 13865 -1735 13885 -1715
rect 13915 -1735 13935 -1715
rect 13965 -1735 13985 -1715
rect 14015 -1735 14035 -1715
rect 14065 -1735 14085 -1715
rect 14115 -1735 14135 -1715
rect 14165 -1735 14185 -1715
rect 14215 -1735 14235 -1715
rect 14265 -1735 14285 -1715
rect 14315 -1735 14335 -1715
rect 14365 -1735 14385 -1715
rect 14415 -1735 14435 -1715
rect 14465 -1735 14485 -1715
rect 14515 -1735 14535 -1715
rect 14565 -1735 14585 -1715
rect 14615 -1735 14635 -1715
rect 14665 -1735 14685 -1715
rect 14715 -1735 14735 -1715
rect 14765 -1735 14785 -1715
rect 14815 -1735 14835 -1715
rect 14865 -1735 14885 -1715
rect 14915 -1735 14935 -1715
rect 14965 -1735 14985 -1715
rect 15015 -1735 15035 -1715
rect 15065 -1735 15085 -1715
rect 15115 -1735 15135 -1715
rect 15165 -1735 15185 -1715
rect 15215 -1735 15235 -1715
rect 15265 -1735 15285 -1715
rect 15315 -1735 15335 -1715
rect 15365 -1735 15385 -1715
rect 15415 -1735 15435 -1715
rect 15465 -1735 15485 -1715
rect 15515 -1735 15535 -1715
rect 15565 -1735 15585 -1715
rect 15615 -1735 15635 -1715
rect 15665 -1735 15685 -1715
rect 15715 -1735 15735 -1715
rect 15765 -1735 15785 -1715
rect 15815 -1735 15835 -1715
rect 15865 -1735 15885 -1715
rect 15915 -1735 15935 -1715
rect 15965 -1735 15985 -1715
rect 16015 -1735 16035 -1715
rect 16065 -1735 16085 -1715
rect 16115 -1735 16135 -1715
rect 16165 -1735 16185 -1715
rect 16215 -1735 16235 -1715
rect 16265 -1735 16285 -1715
rect 16315 -1735 16335 -1715
rect 16365 -1735 16385 -1715
rect 16415 -1735 16435 -1715
rect 16465 -1735 16485 -1715
rect 16515 -1735 16535 -1715
rect 16565 -1735 16585 -1715
rect 16615 -1735 16635 -1715
rect 16665 -1735 16685 -1715
rect 16715 -1735 16735 -1715
rect 16765 -1735 16785 -1715
rect 16815 -1735 16835 -1715
rect 16865 -1735 16885 -1715
rect 16915 -1735 16935 -1715
rect 16965 -1735 16985 -1715
rect 17015 -1735 17035 -1715
rect 17065 -1735 17085 -1715
rect 17115 -1735 17135 -1715
rect 17165 -1735 17185 -1715
rect 17215 -1735 17235 -1715
rect 17265 -1735 17285 -1715
rect 17315 -1735 17335 -1715
rect 17365 -1735 17385 -1715
rect 17415 -1735 17435 -1715
rect 17465 -1735 17485 -1715
rect 17515 -1735 17535 -1715
rect 17565 -1735 17585 -1715
rect 17615 -1735 17635 -1715
rect 17665 -1735 17685 -1715
rect 17715 -1735 17735 -1715
rect 17765 -1735 17785 -1715
rect 17815 -1735 17835 -1715
rect 17865 -1735 17885 -1715
rect 17915 -1735 17935 -1715
rect 17965 -1735 17985 -1715
rect 18015 -1735 18035 -1715
rect 18065 -1735 18085 -1715
rect 18115 -1735 18135 -1715
rect 18165 -1735 18185 -1715
rect 18215 -1735 18235 -1715
rect 18265 -1735 18285 -1715
rect 18315 -1735 18335 -1715
rect 18365 -1735 18385 -1715
rect 18415 -1735 18435 -1715
rect 18465 -1735 18485 -1715
rect 18515 -1735 18535 -1715
rect 18565 -1735 18585 -1715
rect 18615 -1735 18635 -1715
rect 18665 -1735 18685 -1715
rect 18715 -1735 18735 -1715
rect 18765 -1735 18785 -1715
rect 18815 -1735 18835 -1715
rect 18865 -1735 18885 -1715
rect 18915 -1735 18935 -1715
rect 18965 -1735 18985 -1715
rect 19015 -1735 19035 -1715
rect 19065 -1735 19085 -1715
rect 19115 -1735 19135 -1715
rect 19165 -1735 19185 -1715
rect 19215 -1735 19235 -1715
rect 19265 -1735 19285 -1715
rect 19315 -1735 19335 -1715
rect 19365 -1735 19385 -1715
rect 19415 -1735 19435 -1715
rect 19465 -1735 19485 -1715
rect 19515 -1735 19535 -1715
rect 19565 -1735 19585 -1715
rect 19615 -1735 19635 -1715
rect 19665 -1735 19685 -1715
rect 19715 -1735 19735 -1715
rect 19765 -1735 19785 -1715
rect 19815 -1735 19835 -1715
rect 19865 -1735 19885 -1715
rect 19915 -1735 19935 -1715
rect 19965 -1735 19985 -1715
rect 20015 -1735 20035 -1715
rect 20065 -1735 20085 -1715
rect 20115 -1735 20135 -1715
rect 20165 -1735 20185 -1715
rect 20215 -1735 20235 -1715
rect 20265 -1735 20285 -1715
rect 20315 -1735 20335 -1715
rect 20365 -1735 20385 -1715
<< mvnsubdiffcont >>
rect -635 5165 -615 5185
rect -585 5165 -565 5185
rect -535 5165 -515 5185
rect -485 5165 -465 5185
rect -435 5165 -415 5185
rect -385 5165 -365 5185
rect -335 5165 -315 5185
rect -285 5165 -265 5185
rect -235 5165 -215 5185
rect -185 5165 -165 5185
rect -135 5165 -115 5185
rect -85 5165 -65 5185
rect -35 5165 -15 5185
rect 15 5165 35 5185
rect 65 5165 85 5185
rect 115 5165 135 5185
rect 165 5165 185 5185
rect 215 5165 235 5185
rect 265 5165 285 5185
rect 315 5165 335 5185
rect 365 5165 385 5185
rect 415 5165 435 5185
rect 465 5165 485 5185
rect 515 5165 535 5185
rect 565 5165 585 5185
rect 615 5165 635 5185
rect 665 5165 685 5185
rect 715 5165 735 5185
rect 765 5165 785 5185
rect 815 5165 835 5185
rect 865 5165 885 5185
rect 915 5165 935 5185
rect 965 5165 985 5185
rect 1015 5165 1035 5185
rect 1065 5165 1085 5185
rect 1115 5165 1135 5185
rect 1165 5165 1185 5185
rect 1215 5165 1235 5185
rect 1265 5165 1285 5185
rect 1315 5165 1335 5185
rect 1365 5165 1385 5185
rect 1415 5165 1435 5185
rect 1465 5165 1485 5185
rect 1515 5165 1535 5185
rect 1565 5165 1585 5185
rect 1615 5165 1635 5185
rect 1665 5165 1685 5185
rect 1715 5165 1735 5185
rect 1765 5165 1785 5185
rect 1815 5165 1835 5185
rect 1865 5165 1885 5185
rect 1915 5165 1935 5185
rect 1965 5165 1985 5185
rect 2015 5165 2035 5185
rect 2065 5165 2085 5185
rect 2115 5165 2135 5185
rect 2165 5165 2185 5185
rect 2215 5165 2235 5185
rect 2265 5165 2285 5185
rect 2315 5165 2335 5185
rect 2365 5165 2385 5185
rect 2415 5165 2435 5185
rect 2465 5165 2485 5185
rect 2515 5165 2535 5185
rect 2565 5165 2585 5185
rect 2615 5165 2635 5185
rect 2665 5165 2685 5185
rect 2715 5165 2735 5185
rect 2765 5165 2785 5185
rect 2815 5165 2835 5185
rect 2865 5165 2885 5185
rect 2915 5165 2935 5185
rect 2965 5165 2985 5185
rect 3015 5165 3035 5185
rect 3065 5165 3085 5185
rect 3115 5165 3135 5185
rect 3165 5165 3185 5185
rect 3215 5165 3235 5185
rect 3265 5165 3285 5185
rect 3315 5165 3335 5185
rect 3365 5165 3385 5185
rect 3415 5165 3435 5185
rect 3465 5165 3485 5185
rect 3515 5165 3535 5185
rect 3565 5165 3585 5185
rect 3615 5165 3635 5185
rect 3665 5165 3685 5185
rect 3715 5165 3735 5185
rect 3765 5165 3785 5185
rect 3815 5165 3835 5185
rect 3865 5165 3885 5185
rect 3915 5165 3935 5185
rect 3965 5165 3985 5185
rect 4015 5165 4035 5185
rect 4065 5165 4085 5185
rect 4115 5165 4135 5185
rect 4165 5165 4185 5185
rect 4215 5165 4235 5185
rect 4265 5165 4285 5185
rect 4315 5165 4335 5185
rect 4365 5165 4385 5185
rect 4415 5165 4435 5185
rect 4465 5165 4485 5185
rect 4515 5165 4535 5185
rect 4565 5165 4585 5185
rect 4615 5165 4635 5185
rect 4665 5165 4685 5185
rect 4715 5165 4735 5185
rect 4765 5165 4785 5185
rect 4815 5165 4835 5185
rect 4865 5165 4885 5185
rect 4915 5165 4935 5185
rect 4965 5165 4985 5185
rect 5015 5165 5035 5185
rect 5065 5165 5085 5185
rect 5115 5165 5135 5185
rect 5165 5165 5185 5185
rect 5215 5165 5235 5185
rect 5265 5165 5285 5185
rect 5315 5165 5335 5185
rect 5365 5165 5385 5185
rect 5415 5165 5435 5185
rect 5465 5165 5485 5185
rect 5515 5165 5535 5185
rect 5565 5165 5585 5185
rect 5615 5165 5635 5185
rect 5665 5165 5685 5185
rect 5715 5165 5735 5185
rect 5765 5165 5785 5185
rect 5815 5165 5835 5185
rect 5865 5165 5885 5185
rect 5915 5165 5935 5185
rect 5965 5165 5985 5185
rect 6015 5165 6035 5185
rect 6065 5165 6085 5185
rect 6115 5165 6135 5185
rect 6165 5165 6185 5185
rect 6215 5165 6235 5185
rect 6265 5165 6285 5185
rect 6315 5165 6335 5185
rect 6365 5165 6385 5185
rect 6415 5165 6435 5185
rect 6465 5165 6485 5185
rect 6515 5165 6535 5185
rect 6565 5165 6585 5185
rect 6615 5165 6635 5185
rect 6665 5165 6685 5185
rect 6715 5165 6735 5185
rect 6765 5165 6785 5185
rect 6815 5165 6835 5185
rect 6865 5165 6885 5185
rect 6915 5165 6935 5185
rect 6965 5165 6985 5185
rect 7015 5165 7035 5185
rect 7065 5165 7085 5185
rect 7115 5165 7135 5185
rect 7165 5165 7185 5185
rect 7215 5165 7235 5185
rect 7265 5165 7285 5185
rect 7315 5165 7335 5185
rect 7365 5165 7385 5185
rect 7415 5165 7435 5185
rect 7465 5165 7485 5185
rect 7515 5165 7535 5185
rect 7565 5165 7585 5185
rect 7615 5165 7635 5185
rect 7665 5165 7685 5185
rect 7715 5165 7735 5185
rect 7765 5165 7785 5185
rect 7815 5165 7835 5185
rect 7865 5165 7885 5185
rect 7915 5165 7935 5185
rect 7965 5165 7985 5185
rect 8015 5165 8035 5185
rect 8065 5165 8085 5185
rect 8115 5165 8135 5185
rect 8165 5165 8185 5185
rect 8215 5165 8235 5185
rect 8265 5165 8285 5185
rect 8315 5165 8335 5185
rect 8365 5165 8385 5185
rect 8415 5165 8435 5185
rect 8465 5165 8485 5185
rect 8515 5165 8535 5185
rect 8565 5165 8585 5185
rect 8615 5165 8635 5185
rect 8665 5165 8685 5185
rect 8715 5165 8735 5185
rect 8765 5165 8785 5185
rect 8815 5165 8835 5185
rect 8865 5165 8885 5185
rect 8915 5165 8935 5185
rect 8965 5165 8985 5185
rect 9015 5165 9035 5185
rect 9065 5165 9085 5185
rect 9115 5165 9135 5185
rect 9165 5165 9185 5185
rect 9215 5165 9235 5185
rect 9265 5165 9285 5185
rect 9315 5165 9335 5185
rect 9365 5165 9385 5185
rect 9415 5165 9435 5185
rect 9465 5165 9485 5185
rect 9515 5165 9535 5185
rect 9565 5165 9585 5185
rect 9615 5165 9635 5185
rect 9665 5165 9685 5185
rect 9715 5165 9735 5185
rect 9765 5165 9785 5185
rect 9815 5165 9835 5185
rect 9865 5165 9885 5185
rect 9915 5165 9935 5185
rect 9965 5165 9985 5185
rect 10015 5165 10035 5185
rect 10065 5165 10085 5185
rect 10115 5165 10135 5185
rect 10165 5165 10185 5185
rect 10215 5165 10235 5185
rect 10265 5165 10285 5185
rect 10315 5165 10335 5185
rect 10365 5165 10385 5185
rect 10415 5165 10435 5185
rect 10465 5165 10485 5185
rect 10515 5165 10535 5185
rect 10565 5165 10585 5185
rect 10615 5165 10635 5185
rect 10665 5165 10685 5185
rect 10715 5165 10735 5185
rect 10765 5165 10785 5185
rect 10815 5165 10835 5185
rect 10865 5165 10885 5185
rect 10915 5165 10935 5185
rect 10965 5165 10985 5185
rect 11015 5165 11035 5185
rect 11065 5165 11085 5185
rect 11115 5165 11135 5185
rect 11165 5165 11185 5185
rect 11215 5165 11235 5185
rect 11265 5165 11285 5185
rect 11315 5165 11335 5185
rect 11365 5165 11385 5185
rect 11415 5165 11435 5185
rect 11465 5165 11485 5185
rect 11515 5165 11535 5185
rect 11565 5165 11585 5185
rect 11615 5165 11635 5185
rect 11665 5165 11685 5185
rect 11715 5165 11735 5185
rect 11765 5165 11785 5185
rect 11815 5165 11835 5185
rect 11865 5165 11885 5185
rect 11915 5165 11935 5185
rect 11965 5165 11985 5185
rect 12015 5165 12035 5185
rect 12065 5165 12085 5185
rect 12115 5165 12135 5185
rect 12165 5165 12185 5185
rect 12215 5165 12235 5185
rect 12265 5165 12285 5185
rect 12315 5165 12335 5185
rect 12365 5165 12385 5185
rect 12415 5165 12435 5185
rect 12465 5165 12485 5185
rect 12515 5165 12535 5185
rect 12565 5165 12585 5185
rect 12615 5165 12635 5185
rect 12665 5165 12685 5185
rect 12715 5165 12735 5185
rect 12765 5165 12785 5185
rect 12815 5165 12835 5185
rect 12865 5165 12885 5185
rect 12915 5165 12935 5185
rect 12965 5165 12985 5185
rect 13015 5165 13035 5185
rect 13065 5165 13085 5185
rect 13115 5165 13135 5185
rect 13165 5165 13185 5185
rect 13215 5165 13235 5185
rect 13265 5165 13285 5185
rect 13315 5165 13335 5185
rect 13365 5165 13385 5185
rect 13415 5165 13435 5185
rect 13465 5165 13485 5185
rect 13515 5165 13535 5185
rect 13565 5165 13585 5185
rect 13615 5165 13635 5185
rect 13665 5165 13685 5185
rect 13715 5165 13735 5185
rect 13765 5165 13785 5185
rect 13815 5165 13835 5185
rect 13865 5165 13885 5185
rect 13915 5165 13935 5185
rect 13965 5165 13985 5185
rect 14015 5165 14035 5185
rect 14065 5165 14085 5185
rect 14115 5165 14135 5185
rect 14165 5165 14185 5185
rect 14215 5165 14235 5185
rect 14265 5165 14285 5185
rect 14315 5165 14335 5185
rect 14365 5165 14385 5185
rect 14415 5165 14435 5185
rect 14465 5165 14485 5185
rect 14515 5165 14535 5185
rect 14565 5165 14585 5185
rect 14615 5165 14635 5185
rect 14665 5165 14685 5185
rect 14715 5165 14735 5185
rect 14765 5165 14785 5185
rect 14815 5165 14835 5185
rect 14865 5165 14885 5185
rect 14915 5165 14935 5185
rect 14965 5165 14985 5185
rect 15015 5165 15035 5185
rect 15065 5165 15085 5185
rect 15115 5165 15135 5185
rect 15165 5165 15185 5185
rect 15215 5165 15235 5185
rect 15265 5165 15285 5185
rect 15315 5165 15335 5185
rect 15365 5165 15385 5185
rect 15415 5165 15435 5185
rect 15465 5165 15485 5185
rect 15515 5165 15535 5185
rect 15565 5165 15585 5185
rect 15615 5165 15635 5185
rect 15665 5165 15685 5185
rect 15715 5165 15735 5185
rect 15765 5165 15785 5185
rect 15815 5165 15835 5185
rect 15865 5165 15885 5185
rect 15915 5165 15935 5185
rect 15965 5165 15985 5185
rect 16015 5165 16035 5185
rect 16065 5165 16085 5185
rect 16115 5165 16135 5185
rect 16165 5165 16185 5185
rect 16215 5165 16235 5185
rect 16265 5165 16285 5185
rect 16315 5165 16335 5185
rect 16365 5165 16385 5185
rect 16415 5165 16435 5185
rect 16465 5165 16485 5185
rect 16515 5165 16535 5185
rect 16565 5165 16585 5185
rect 16615 5165 16635 5185
rect 16665 5165 16685 5185
rect 16715 5165 16735 5185
rect 16765 5165 16785 5185
rect 16815 5165 16835 5185
rect 16865 5165 16885 5185
rect 16915 5165 16935 5185
rect 16965 5165 16985 5185
rect 17015 5165 17035 5185
rect 17065 5165 17085 5185
rect 17115 5165 17135 5185
rect 17165 5165 17185 5185
rect 17215 5165 17235 5185
rect 17265 5165 17285 5185
rect 17315 5165 17335 5185
rect 17365 5165 17385 5185
rect 17415 5165 17435 5185
rect 17465 5165 17485 5185
rect 17515 5165 17535 5185
rect 17565 5165 17585 5185
rect 17615 5165 17635 5185
rect 17665 5165 17685 5185
rect 17715 5165 17735 5185
rect 17765 5165 17785 5185
rect 17815 5165 17835 5185
rect 17865 5165 17885 5185
rect 17915 5165 17935 5185
rect 17965 5165 17985 5185
rect 18015 5165 18035 5185
rect 18065 5165 18085 5185
rect 18115 5165 18135 5185
rect 18165 5165 18185 5185
rect 18215 5165 18235 5185
rect 18265 5165 18285 5185
rect 18315 5165 18335 5185
rect 18365 5165 18385 5185
rect 18415 5165 18435 5185
rect 18465 5165 18485 5185
rect 18515 5165 18535 5185
rect 18565 5165 18585 5185
rect 18615 5165 18635 5185
rect 18665 5165 18685 5185
rect 18715 5165 18735 5185
rect 18765 5165 18785 5185
rect 18815 5165 18835 5185
rect 18865 5165 18885 5185
rect 18915 5165 18935 5185
rect 18965 5165 18985 5185
rect 19015 5165 19035 5185
rect 19065 5165 19085 5185
rect 19115 5165 19135 5185
rect 19165 5165 19185 5185
rect 19215 5165 19235 5185
rect 19265 5165 19285 5185
rect 19315 5165 19335 5185
rect 19365 5165 19385 5185
rect 19415 5165 19435 5185
rect 19465 5165 19485 5185
rect 19515 5165 19535 5185
rect 19565 5165 19585 5185
rect 19615 5165 19635 5185
rect 19665 5165 19685 5185
rect 19715 5165 19735 5185
rect 19765 5165 19785 5185
rect 19815 5165 19835 5185
rect 19865 5165 19885 5185
rect 19915 5165 19935 5185
rect 19965 5165 19985 5185
rect 20015 5165 20035 5185
rect 20065 5165 20085 5185
rect 20115 5165 20135 5185
rect 20165 5165 20185 5185
rect 20215 5165 20235 5185
rect 20265 5165 20285 5185
rect 20315 5165 20335 5185
rect 20365 5165 20385 5185
rect -635 3865 -615 3885
rect -585 3865 -565 3885
rect -535 3865 -515 3885
rect -485 3865 -465 3885
rect -435 3865 -415 3885
rect -385 3865 -365 3885
rect -335 3865 -315 3885
rect -285 3865 -265 3885
rect -235 3865 -215 3885
rect -185 3865 -165 3885
rect -135 3865 -115 3885
rect -85 3865 -65 3885
rect -35 3865 -15 3885
rect 15 3865 35 3885
rect 65 3865 85 3885
rect 115 3865 135 3885
rect 165 3865 185 3885
rect 215 3865 235 3885
rect 265 3865 285 3885
rect 315 3865 335 3885
rect 365 3865 385 3885
rect 415 3865 435 3885
rect 465 3865 485 3885
rect 515 3865 535 3885
rect 565 3865 585 3885
rect 615 3865 635 3885
rect 665 3865 685 3885
rect 715 3865 735 3885
rect 765 3865 785 3885
rect 815 3865 835 3885
rect 865 3865 885 3885
rect 915 3865 935 3885
rect 965 3865 985 3885
rect 1015 3865 1035 3885
rect 1065 3865 1085 3885
rect 1115 3865 1135 3885
rect 1165 3865 1185 3885
rect 1215 3865 1235 3885
rect 1265 3865 1285 3885
rect 1315 3865 1335 3885
rect 1365 3865 1385 3885
rect 1415 3865 1435 3885
rect 1465 3865 1485 3885
rect 1515 3865 1535 3885
rect 1565 3865 1585 3885
rect 1615 3865 1635 3885
rect 1665 3865 1685 3885
rect 1715 3865 1735 3885
rect 1765 3865 1785 3885
rect 1815 3865 1835 3885
rect 1865 3865 1885 3885
rect 1915 3865 1935 3885
rect 1965 3865 1985 3885
rect 2015 3865 2035 3885
rect 2065 3865 2085 3885
rect 2115 3865 2135 3885
rect 2165 3865 2185 3885
rect 2215 3865 2235 3885
rect 2265 3865 2285 3885
rect 2315 3865 2335 3885
rect 2365 3865 2385 3885
rect 2415 3865 2435 3885
rect 2465 3865 2485 3885
rect 2515 3865 2535 3885
rect 2565 3865 2585 3885
rect 2615 3865 2635 3885
rect 2665 3865 2685 3885
rect 2715 3865 2735 3885
rect 2765 3865 2785 3885
rect 2815 3865 2835 3885
rect 2865 3865 2885 3885
rect 2915 3865 2935 3885
rect 2965 3865 2985 3885
rect 3015 3865 3035 3885
rect 3065 3865 3085 3885
rect 3115 3865 3135 3885
rect 3165 3865 3185 3885
rect 3215 3865 3235 3885
rect 3265 3865 3285 3885
rect 3315 3865 3335 3885
rect 3365 3865 3385 3885
rect 3415 3865 3435 3885
rect 3465 3865 3485 3885
rect 3515 3865 3535 3885
rect 3565 3865 3585 3885
rect 3615 3865 3635 3885
rect 3665 3865 3685 3885
rect 3715 3865 3735 3885
rect 3765 3865 3785 3885
rect 3815 3865 3835 3885
rect 3865 3865 3885 3885
rect 3915 3865 3935 3885
rect 3965 3865 3985 3885
rect 4015 3865 4035 3885
rect 4065 3865 4085 3885
rect 4115 3865 4135 3885
rect 4165 3865 4185 3885
rect 4215 3865 4235 3885
rect 4265 3865 4285 3885
rect 4315 3865 4335 3885
rect 4365 3865 4385 3885
rect 4415 3865 4435 3885
rect 4465 3865 4485 3885
rect 4515 3865 4535 3885
rect 4565 3865 4585 3885
rect 4615 3865 4635 3885
rect 4665 3865 4685 3885
rect 4715 3865 4735 3885
rect 4765 3865 4785 3885
rect 4815 3865 4835 3885
rect 4865 3865 4885 3885
rect 4915 3865 4935 3885
rect 4965 3865 4985 3885
rect 5015 3865 5035 3885
rect 5065 3865 5085 3885
rect 5115 3865 5135 3885
rect 5165 3865 5185 3885
rect 5215 3865 5235 3885
rect 5265 3865 5285 3885
rect 5315 3865 5335 3885
rect 5365 3865 5385 3885
rect 5415 3865 5435 3885
rect 5465 3865 5485 3885
rect 5515 3865 5535 3885
rect 5565 3865 5585 3885
rect 5615 3865 5635 3885
rect 5665 3865 5685 3885
rect 5715 3865 5735 3885
rect 5765 3865 5785 3885
rect 5815 3865 5835 3885
rect 5865 3865 5885 3885
rect 5915 3865 5935 3885
rect 5965 3865 5985 3885
rect 6015 3865 6035 3885
rect 6065 3865 6085 3885
rect 6115 3865 6135 3885
rect 6165 3865 6185 3885
rect 6215 3865 6235 3885
rect 6265 3865 6285 3885
rect 6315 3865 6335 3885
rect 6365 3865 6385 3885
rect 6415 3865 6435 3885
rect 6465 3865 6485 3885
rect 6515 3865 6535 3885
rect 6565 3865 6585 3885
rect 6615 3865 6635 3885
rect 6665 3865 6685 3885
rect 6715 3865 6735 3885
rect 6765 3865 6785 3885
rect 6815 3865 6835 3885
rect 6865 3865 6885 3885
rect 6915 3865 6935 3885
rect 6965 3865 6985 3885
rect 7015 3865 7035 3885
rect 7065 3865 7085 3885
rect 7115 3865 7135 3885
rect 7165 3865 7185 3885
rect 7215 3865 7235 3885
rect 7265 3865 7285 3885
rect 7315 3865 7335 3885
rect 7365 3865 7385 3885
rect 7415 3865 7435 3885
rect 7465 3865 7485 3885
rect 7515 3865 7535 3885
rect 7565 3865 7585 3885
rect 7615 3865 7635 3885
rect 7665 3865 7685 3885
rect 7715 3865 7735 3885
rect 7765 3865 7785 3885
rect 7815 3865 7835 3885
rect 7865 3865 7885 3885
rect 7915 3865 7935 3885
rect 7965 3865 7985 3885
rect 8015 3865 8035 3885
rect 8065 3865 8085 3885
rect 8115 3865 8135 3885
rect 8165 3865 8185 3885
rect 8215 3865 8235 3885
rect 8265 3865 8285 3885
rect 8315 3865 8335 3885
rect 8365 3865 8385 3885
rect 8415 3865 8435 3885
rect 8465 3865 8485 3885
rect 8515 3865 8535 3885
rect 8565 3865 8585 3885
rect 8615 3865 8635 3885
rect 8665 3865 8685 3885
rect 8715 3865 8735 3885
rect 8765 3865 8785 3885
rect 8815 3865 8835 3885
rect 8865 3865 8885 3885
rect 8915 3865 8935 3885
rect 8965 3865 8985 3885
rect 9015 3865 9035 3885
rect 9065 3865 9085 3885
rect 9115 3865 9135 3885
rect 9165 3865 9185 3885
rect 9215 3865 9235 3885
rect 9265 3865 9285 3885
rect 9315 3865 9335 3885
rect 9365 3865 9385 3885
rect 9415 3865 9435 3885
rect 9465 3865 9485 3885
rect 9515 3865 9535 3885
rect 9565 3865 9585 3885
rect 9615 3865 9635 3885
rect 9665 3865 9685 3885
rect 9715 3865 9735 3885
rect 9765 3865 9785 3885
rect 9815 3865 9835 3885
rect 9865 3865 9885 3885
rect 9915 3865 9935 3885
rect 9965 3865 9985 3885
rect 10015 3865 10035 3885
rect 10065 3865 10085 3885
rect 10115 3865 10135 3885
rect 10165 3865 10185 3885
rect 10215 3865 10235 3885
rect 10265 3865 10285 3885
rect 10315 3865 10335 3885
rect 10365 3865 10385 3885
rect 10415 3865 10435 3885
rect 10465 3865 10485 3885
rect 10515 3865 10535 3885
rect 10565 3865 10585 3885
rect 10615 3865 10635 3885
rect 10665 3865 10685 3885
rect 10715 3865 10735 3885
rect 10765 3865 10785 3885
rect 10815 3865 10835 3885
rect 10865 3865 10885 3885
rect 10915 3865 10935 3885
rect 10965 3865 10985 3885
rect 11015 3865 11035 3885
rect 11065 3865 11085 3885
rect 11115 3865 11135 3885
rect 11165 3865 11185 3885
rect 11215 3865 11235 3885
rect 11265 3865 11285 3885
rect 11315 3865 11335 3885
rect 11365 3865 11385 3885
rect 11415 3865 11435 3885
rect 11465 3865 11485 3885
rect 11515 3865 11535 3885
rect 11565 3865 11585 3885
rect 11615 3865 11635 3885
rect 11665 3865 11685 3885
rect 11715 3865 11735 3885
rect 11765 3865 11785 3885
rect 11815 3865 11835 3885
rect 11865 3865 11885 3885
rect 11915 3865 11935 3885
rect 11965 3865 11985 3885
rect 12015 3865 12035 3885
rect 12065 3865 12085 3885
rect 12115 3865 12135 3885
rect 12165 3865 12185 3885
rect 12215 3865 12235 3885
rect 12265 3865 12285 3885
rect 12315 3865 12335 3885
rect 12365 3865 12385 3885
rect 12415 3865 12435 3885
rect 12465 3865 12485 3885
rect 12515 3865 12535 3885
rect 12565 3865 12585 3885
rect 12615 3865 12635 3885
rect 12665 3865 12685 3885
rect 12715 3865 12735 3885
rect 12765 3865 12785 3885
rect 12815 3865 12835 3885
rect 12865 3865 12885 3885
rect 12915 3865 12935 3885
rect 12965 3865 12985 3885
rect 13015 3865 13035 3885
rect 13065 3865 13085 3885
rect 13115 3865 13135 3885
rect 13165 3865 13185 3885
rect 13215 3865 13235 3885
rect 13265 3865 13285 3885
rect 13315 3865 13335 3885
rect 13365 3865 13385 3885
rect 13415 3865 13435 3885
rect 13465 3865 13485 3885
rect 13515 3865 13535 3885
rect 13565 3865 13585 3885
rect 13615 3865 13635 3885
rect 13665 3865 13685 3885
rect 13715 3865 13735 3885
rect 13765 3865 13785 3885
rect 13815 3865 13835 3885
rect 13865 3865 13885 3885
rect 13915 3865 13935 3885
rect 13965 3865 13985 3885
rect 14015 3865 14035 3885
rect 14065 3865 14085 3885
rect 14115 3865 14135 3885
rect 14165 3865 14185 3885
rect 14215 3865 14235 3885
rect 14265 3865 14285 3885
rect 14315 3865 14335 3885
rect 14365 3865 14385 3885
rect 14415 3865 14435 3885
rect 14465 3865 14485 3885
rect 14515 3865 14535 3885
rect 14565 3865 14585 3885
rect 14615 3865 14635 3885
rect 14665 3865 14685 3885
rect 14715 3865 14735 3885
rect 14765 3865 14785 3885
rect 14815 3865 14835 3885
rect 14865 3865 14885 3885
rect 14915 3865 14935 3885
rect 14965 3865 14985 3885
rect 15015 3865 15035 3885
rect 15065 3865 15085 3885
rect 15115 3865 15135 3885
rect 15165 3865 15185 3885
rect 15215 3865 15235 3885
rect 15265 3865 15285 3885
rect 15315 3865 15335 3885
rect 15365 3865 15385 3885
rect 15415 3865 15435 3885
rect 15465 3865 15485 3885
rect 15515 3865 15535 3885
rect 15565 3865 15585 3885
rect 15615 3865 15635 3885
rect 15665 3865 15685 3885
rect 15715 3865 15735 3885
rect 15765 3865 15785 3885
rect 15815 3865 15835 3885
rect 15865 3865 15885 3885
rect 15915 3865 15935 3885
rect 15965 3865 15985 3885
rect 16015 3865 16035 3885
rect 16065 3865 16085 3885
rect 16115 3865 16135 3885
rect 16165 3865 16185 3885
rect 16215 3865 16235 3885
rect 16265 3865 16285 3885
rect 16315 3865 16335 3885
rect 16365 3865 16385 3885
rect 16415 3865 16435 3885
rect 16465 3865 16485 3885
rect 16515 3865 16535 3885
rect 16565 3865 16585 3885
rect 16615 3865 16635 3885
rect 16665 3865 16685 3885
rect 16715 3865 16735 3885
rect 16765 3865 16785 3885
rect 16815 3865 16835 3885
rect 16865 3865 16885 3885
rect 16915 3865 16935 3885
rect 16965 3865 16985 3885
rect 17015 3865 17035 3885
rect 17065 3865 17085 3885
rect 17115 3865 17135 3885
rect 17165 3865 17185 3885
rect 17215 3865 17235 3885
rect 17265 3865 17285 3885
rect 17315 3865 17335 3885
rect 17365 3865 17385 3885
rect 17415 3865 17435 3885
rect 17465 3865 17485 3885
rect 17515 3865 17535 3885
rect 17565 3865 17585 3885
rect 17615 3865 17635 3885
rect 17665 3865 17685 3885
rect 17715 3865 17735 3885
rect 17765 3865 17785 3885
rect 17815 3865 17835 3885
rect 17865 3865 17885 3885
rect 17915 3865 17935 3885
rect 17965 3865 17985 3885
rect 18015 3865 18035 3885
rect 18065 3865 18085 3885
rect 18115 3865 18135 3885
rect 18165 3865 18185 3885
rect 18215 3865 18235 3885
rect 18265 3865 18285 3885
rect 18315 3865 18335 3885
rect 18365 3865 18385 3885
rect 18415 3865 18435 3885
rect 18465 3865 18485 3885
rect 18515 3865 18535 3885
rect 18565 3865 18585 3885
rect 18615 3865 18635 3885
rect 18665 3865 18685 3885
rect 18715 3865 18735 3885
rect 18765 3865 18785 3885
rect 18815 3865 18835 3885
rect 18865 3865 18885 3885
rect 18915 3865 18935 3885
rect 18965 3865 18985 3885
rect 19015 3865 19035 3885
rect 19065 3865 19085 3885
rect 19115 3865 19135 3885
rect 19165 3865 19185 3885
rect 19215 3865 19235 3885
rect 19265 3865 19285 3885
rect 19315 3865 19335 3885
rect 19365 3865 19385 3885
rect 19415 3865 19435 3885
rect 19465 3865 19485 3885
rect 19515 3865 19535 3885
rect 19565 3865 19585 3885
rect 19615 3865 19635 3885
rect 19665 3865 19685 3885
rect 19715 3865 19735 3885
rect 19765 3865 19785 3885
rect 19815 3865 19835 3885
rect 19865 3865 19885 3885
rect 19915 3865 19935 3885
rect 19965 3865 19985 3885
rect 20015 3865 20035 3885
rect 20065 3865 20085 3885
rect 20115 3865 20135 3885
rect 20165 3865 20185 3885
rect 20215 3865 20235 3885
rect 20265 3865 20285 3885
rect 20315 3865 20335 3885
rect 20365 3865 20385 3885
rect -635 2565 -615 2585
rect -585 2565 -565 2585
rect -535 2565 -515 2585
rect -485 2565 -465 2585
rect -435 2565 -415 2585
rect -385 2565 -365 2585
rect -335 2565 -315 2585
rect -285 2565 -265 2585
rect -235 2565 -215 2585
rect -185 2565 -165 2585
rect -135 2565 -115 2585
rect -85 2565 -65 2585
rect -35 2565 -15 2585
rect 15 2565 35 2585
rect 65 2565 85 2585
rect 115 2565 135 2585
rect 165 2565 185 2585
rect 215 2565 235 2585
rect 265 2565 285 2585
rect 315 2565 335 2585
rect 365 2565 385 2585
rect 415 2565 435 2585
rect 465 2565 485 2585
rect 515 2565 535 2585
rect 565 2565 585 2585
rect 615 2565 635 2585
rect 665 2565 685 2585
rect 715 2565 735 2585
rect 765 2565 785 2585
rect 815 2565 835 2585
rect 865 2565 885 2585
rect 915 2565 935 2585
rect 965 2565 985 2585
rect 1015 2565 1035 2585
rect 1065 2565 1085 2585
rect 1115 2565 1135 2585
rect 1165 2565 1185 2585
rect 1215 2565 1235 2585
rect 1265 2565 1285 2585
rect 1315 2565 1335 2585
rect 1365 2565 1385 2585
rect 1415 2565 1435 2585
rect 1465 2565 1485 2585
rect 1515 2565 1535 2585
rect 1565 2565 1585 2585
rect 1615 2565 1635 2585
rect 1665 2565 1685 2585
rect 1715 2565 1735 2585
rect 1765 2565 1785 2585
rect 1815 2565 1835 2585
rect 1865 2565 1885 2585
rect 1915 2565 1935 2585
rect 1965 2565 1985 2585
rect 2015 2565 2035 2585
rect 2065 2565 2085 2585
rect 2115 2565 2135 2585
rect 2165 2565 2185 2585
rect 2215 2565 2235 2585
rect 2265 2565 2285 2585
rect 2315 2565 2335 2585
rect 2365 2565 2385 2585
rect 2415 2565 2435 2585
rect 2465 2565 2485 2585
rect 2515 2565 2535 2585
rect 2565 2565 2585 2585
rect 2615 2565 2635 2585
rect 2665 2565 2685 2585
rect 2715 2565 2735 2585
rect 2765 2565 2785 2585
rect 2815 2565 2835 2585
rect 2865 2565 2885 2585
rect 2915 2565 2935 2585
rect 2965 2565 2985 2585
rect 3015 2565 3035 2585
rect 3065 2565 3085 2585
rect 3115 2565 3135 2585
rect 3165 2565 3185 2585
rect 3215 2565 3235 2585
rect 3265 2565 3285 2585
rect 3315 2565 3335 2585
rect 3365 2565 3385 2585
rect 3415 2565 3435 2585
rect 3465 2565 3485 2585
rect 3515 2565 3535 2585
rect 3565 2565 3585 2585
rect 3615 2565 3635 2585
rect 3665 2565 3685 2585
rect 3715 2565 3735 2585
rect 3765 2565 3785 2585
rect 3815 2565 3835 2585
rect 3865 2565 3885 2585
rect 3915 2565 3935 2585
rect 3965 2565 3985 2585
rect 4015 2565 4035 2585
rect 4065 2565 4085 2585
rect 4115 2565 4135 2585
rect 4165 2565 4185 2585
rect 4215 2565 4235 2585
rect 4265 2565 4285 2585
rect 4315 2565 4335 2585
rect 4365 2565 4385 2585
rect 4415 2565 4435 2585
rect 4465 2565 4485 2585
rect 4515 2565 4535 2585
rect 4565 2565 4585 2585
rect 4615 2565 4635 2585
rect 4665 2565 4685 2585
rect 4715 2565 4735 2585
rect 4765 2565 4785 2585
rect 4815 2565 4835 2585
rect 4865 2565 4885 2585
rect 4915 2565 4935 2585
rect 4965 2565 4985 2585
rect 5015 2565 5035 2585
rect 5065 2565 5085 2585
rect 5115 2565 5135 2585
rect 5165 2565 5185 2585
rect 5215 2565 5235 2585
rect 5265 2565 5285 2585
rect 5315 2565 5335 2585
rect 5365 2565 5385 2585
rect 5415 2565 5435 2585
rect 5465 2565 5485 2585
rect 5515 2565 5535 2585
rect 5565 2565 5585 2585
rect 5615 2565 5635 2585
rect 5665 2565 5685 2585
rect 5715 2565 5735 2585
rect 5765 2565 5785 2585
rect 5815 2565 5835 2585
rect 5865 2565 5885 2585
rect 5915 2565 5935 2585
rect 5965 2565 5985 2585
rect 6015 2565 6035 2585
rect 6065 2565 6085 2585
rect 6115 2565 6135 2585
rect 6165 2565 6185 2585
rect 6215 2565 6235 2585
rect 6265 2565 6285 2585
rect 6315 2565 6335 2585
rect 6365 2565 6385 2585
rect 6415 2565 6435 2585
rect 6465 2565 6485 2585
rect 6515 2565 6535 2585
rect 6565 2565 6585 2585
rect 6615 2565 6635 2585
rect 6665 2565 6685 2585
rect 6715 2565 6735 2585
rect 6765 2565 6785 2585
rect 6815 2565 6835 2585
rect 6865 2565 6885 2585
rect 6915 2565 6935 2585
rect 6965 2565 6985 2585
rect 7015 2565 7035 2585
rect 7065 2565 7085 2585
rect 7115 2565 7135 2585
rect 7165 2565 7185 2585
rect 7215 2565 7235 2585
rect 7265 2565 7285 2585
rect 7315 2565 7335 2585
rect 7365 2565 7385 2585
rect 7415 2565 7435 2585
rect 7465 2565 7485 2585
rect 7515 2565 7535 2585
rect 7565 2565 7585 2585
rect 7615 2565 7635 2585
rect 7665 2565 7685 2585
rect 7715 2565 7735 2585
rect 7765 2565 7785 2585
rect 7815 2565 7835 2585
rect 7865 2565 7885 2585
rect 7915 2565 7935 2585
rect 7965 2565 7985 2585
rect 8015 2565 8035 2585
rect 8065 2565 8085 2585
rect 8115 2565 8135 2585
rect 8165 2565 8185 2585
rect 8215 2565 8235 2585
rect 8265 2565 8285 2585
rect 8315 2565 8335 2585
rect 8365 2565 8385 2585
rect 8415 2565 8435 2585
rect 8465 2565 8485 2585
rect 8515 2565 8535 2585
rect 8565 2565 8585 2585
rect 8615 2565 8635 2585
rect 8665 2565 8685 2585
rect 8715 2565 8735 2585
rect 8765 2565 8785 2585
rect 8815 2565 8835 2585
rect 8865 2565 8885 2585
rect 8915 2565 8935 2585
rect 8965 2565 8985 2585
rect 9015 2565 9035 2585
rect 9065 2565 9085 2585
rect 9115 2565 9135 2585
rect 9165 2565 9185 2585
rect 9215 2565 9235 2585
rect 9265 2565 9285 2585
rect 9315 2565 9335 2585
rect 9365 2565 9385 2585
rect 9415 2565 9435 2585
rect 9465 2565 9485 2585
rect 9515 2565 9535 2585
rect 9565 2565 9585 2585
rect 9615 2565 9635 2585
rect 9665 2565 9685 2585
rect 9715 2565 9735 2585
rect 9765 2565 9785 2585
rect 9815 2565 9835 2585
rect 9865 2565 9885 2585
rect 9915 2565 9935 2585
rect 9965 2565 9985 2585
rect 10015 2565 10035 2585
rect 10065 2565 10085 2585
rect 10115 2565 10135 2585
rect 10165 2565 10185 2585
rect 10215 2565 10235 2585
rect 10265 2565 10285 2585
rect 10315 2565 10335 2585
rect 10365 2565 10385 2585
rect 10415 2565 10435 2585
rect 10465 2565 10485 2585
rect 10515 2565 10535 2585
rect 10565 2565 10585 2585
rect 10615 2565 10635 2585
rect 10665 2565 10685 2585
rect 10715 2565 10735 2585
rect 10765 2565 10785 2585
rect 10815 2565 10835 2585
rect 10865 2565 10885 2585
rect 10915 2565 10935 2585
rect 10965 2565 10985 2585
rect 11015 2565 11035 2585
rect 11065 2565 11085 2585
rect 11115 2565 11135 2585
rect 11165 2565 11185 2585
rect 11215 2565 11235 2585
rect 11265 2565 11285 2585
rect 11315 2565 11335 2585
rect 11365 2565 11385 2585
rect 11415 2565 11435 2585
rect 11465 2565 11485 2585
rect 11515 2565 11535 2585
rect 11565 2565 11585 2585
rect 11615 2565 11635 2585
rect 11665 2565 11685 2585
rect 11715 2565 11735 2585
rect 11765 2565 11785 2585
rect 11815 2565 11835 2585
rect 11865 2565 11885 2585
rect 11915 2565 11935 2585
rect 11965 2565 11985 2585
rect 12015 2565 12035 2585
rect 12065 2565 12085 2585
rect 12115 2565 12135 2585
rect 12165 2565 12185 2585
rect 12215 2565 12235 2585
rect 12265 2565 12285 2585
rect 12315 2565 12335 2585
rect 12365 2565 12385 2585
rect 12415 2565 12435 2585
rect 12465 2565 12485 2585
rect 12515 2565 12535 2585
rect 12565 2565 12585 2585
rect 12615 2565 12635 2585
rect 12665 2565 12685 2585
rect 12715 2565 12735 2585
rect 12765 2565 12785 2585
rect 12815 2565 12835 2585
rect 12865 2565 12885 2585
rect 12915 2565 12935 2585
rect 12965 2565 12985 2585
rect 13015 2565 13035 2585
rect 13065 2565 13085 2585
rect 13115 2565 13135 2585
rect 13165 2565 13185 2585
rect 13215 2565 13235 2585
rect 13265 2565 13285 2585
rect 13315 2565 13335 2585
rect 13365 2565 13385 2585
rect 13415 2565 13435 2585
rect 13465 2565 13485 2585
rect 13515 2565 13535 2585
rect 13565 2565 13585 2585
rect 13615 2565 13635 2585
rect 13665 2565 13685 2585
rect 13715 2565 13735 2585
rect 13765 2565 13785 2585
rect 13815 2565 13835 2585
rect 13865 2565 13885 2585
rect 13915 2565 13935 2585
rect 13965 2565 13985 2585
rect 14015 2565 14035 2585
rect 14065 2565 14085 2585
rect 14115 2565 14135 2585
rect 14165 2565 14185 2585
rect 14215 2565 14235 2585
rect 14265 2565 14285 2585
rect 14315 2565 14335 2585
rect 14365 2565 14385 2585
rect 14415 2565 14435 2585
rect 14465 2565 14485 2585
rect 14515 2565 14535 2585
rect 14565 2565 14585 2585
rect 14615 2565 14635 2585
rect 14665 2565 14685 2585
rect 14715 2565 14735 2585
rect 14765 2565 14785 2585
rect 14815 2565 14835 2585
rect 14865 2565 14885 2585
rect 14915 2565 14935 2585
rect 14965 2565 14985 2585
rect 15015 2565 15035 2585
rect 15065 2565 15085 2585
rect 15115 2565 15135 2585
rect 15165 2565 15185 2585
rect 15215 2565 15235 2585
rect 15265 2565 15285 2585
rect 15315 2565 15335 2585
rect 15365 2565 15385 2585
rect 15415 2565 15435 2585
rect 15465 2565 15485 2585
rect 15515 2565 15535 2585
rect 15565 2565 15585 2585
rect 15615 2565 15635 2585
rect 15665 2565 15685 2585
rect 15715 2565 15735 2585
rect 15765 2565 15785 2585
rect 15815 2565 15835 2585
rect 15865 2565 15885 2585
rect 15915 2565 15935 2585
rect 15965 2565 15985 2585
rect 16015 2565 16035 2585
rect 16065 2565 16085 2585
rect 16115 2565 16135 2585
rect 16165 2565 16185 2585
rect 16215 2565 16235 2585
rect 16265 2565 16285 2585
rect 16315 2565 16335 2585
rect 16365 2565 16385 2585
rect 16415 2565 16435 2585
rect 16465 2565 16485 2585
rect 16515 2565 16535 2585
rect 16565 2565 16585 2585
rect 16615 2565 16635 2585
rect 16665 2565 16685 2585
rect 16715 2565 16735 2585
rect 16765 2565 16785 2585
rect 16815 2565 16835 2585
rect 16865 2565 16885 2585
rect 16915 2565 16935 2585
rect 16965 2565 16985 2585
rect 17015 2565 17035 2585
rect 17065 2565 17085 2585
rect 17115 2565 17135 2585
rect 17165 2565 17185 2585
rect 17215 2565 17235 2585
rect 17265 2565 17285 2585
rect 17315 2565 17335 2585
rect 17365 2565 17385 2585
rect 17415 2565 17435 2585
rect 17465 2565 17485 2585
rect 17515 2565 17535 2585
rect 17565 2565 17585 2585
rect 17615 2565 17635 2585
rect 17665 2565 17685 2585
rect 17715 2565 17735 2585
rect 17765 2565 17785 2585
rect 17815 2565 17835 2585
rect 17865 2565 17885 2585
rect 17915 2565 17935 2585
rect 17965 2565 17985 2585
rect 18015 2565 18035 2585
rect 18065 2565 18085 2585
rect 18115 2565 18135 2585
rect 18165 2565 18185 2585
rect 18215 2565 18235 2585
rect 18265 2565 18285 2585
rect 18315 2565 18335 2585
rect 18365 2565 18385 2585
rect 18415 2565 18435 2585
rect 18465 2565 18485 2585
rect 18515 2565 18535 2585
rect 18565 2565 18585 2585
rect 18615 2565 18635 2585
rect 18665 2565 18685 2585
rect 18715 2565 18735 2585
rect 18765 2565 18785 2585
rect 18815 2565 18835 2585
rect 18865 2565 18885 2585
rect 18915 2565 18935 2585
rect 18965 2565 18985 2585
rect 19015 2565 19035 2585
rect 19065 2565 19085 2585
rect 19115 2565 19135 2585
rect 19165 2565 19185 2585
rect 19215 2565 19235 2585
rect 19265 2565 19285 2585
rect 19315 2565 19335 2585
rect 19365 2565 19385 2585
rect 19415 2565 19435 2585
rect 19465 2565 19485 2585
rect 19515 2565 19535 2585
rect 19565 2565 19585 2585
rect 19615 2565 19635 2585
rect 19665 2565 19685 2585
rect 19715 2565 19735 2585
rect 19765 2565 19785 2585
rect 19815 2565 19835 2585
rect 19865 2565 19885 2585
rect 19915 2565 19935 2585
rect 19965 2565 19985 2585
rect 20015 2565 20035 2585
rect 20065 2565 20085 2585
rect 20115 2565 20135 2585
rect 20165 2565 20185 2585
rect 20215 2565 20235 2585
rect 20265 2565 20285 2585
rect 20315 2565 20335 2585
rect 20365 2565 20385 2585
rect -635 1815 -615 1835
rect -585 1815 -565 1835
rect -535 1815 -515 1835
rect -485 1815 -465 1835
rect -435 1815 -415 1835
rect -385 1815 -365 1835
rect -335 1815 -315 1835
rect -285 1815 -265 1835
rect -235 1815 -215 1835
rect -185 1815 -165 1835
rect -135 1815 -115 1835
rect -85 1815 -65 1835
rect -35 1815 -15 1835
rect 15 1815 35 1835
rect 65 1815 85 1835
rect 115 1815 135 1835
rect 165 1815 185 1835
rect 215 1815 235 1835
rect 265 1815 285 1835
rect 315 1815 335 1835
rect 365 1815 385 1835
rect 415 1815 435 1835
rect 465 1815 485 1835
rect 515 1815 535 1835
rect 565 1815 585 1835
rect 615 1815 635 1835
rect 665 1815 685 1835
rect 715 1815 735 1835
rect 765 1815 785 1835
rect 815 1815 835 1835
rect 865 1815 885 1835
rect 915 1815 935 1835
rect 965 1815 985 1835
rect 1015 1815 1035 1835
rect 1065 1815 1085 1835
rect 1115 1815 1135 1835
rect 1165 1815 1185 1835
rect 1215 1815 1235 1835
rect 1265 1815 1285 1835
rect 1315 1815 1335 1835
rect 1365 1815 1385 1835
rect 1415 1815 1435 1835
rect 1465 1815 1485 1835
rect 1515 1815 1535 1835
rect 1565 1815 1585 1835
rect 1615 1815 1635 1835
rect 1665 1815 1685 1835
rect 1715 1815 1735 1835
rect 1765 1815 1785 1835
rect 1815 1815 1835 1835
rect 1865 1815 1885 1835
rect 1915 1815 1935 1835
rect 1965 1815 1985 1835
rect 2015 1815 2035 1835
rect 2065 1815 2085 1835
rect 2115 1815 2135 1835
rect 2165 1815 2185 1835
rect 2215 1815 2235 1835
rect 2265 1815 2285 1835
rect 2315 1815 2335 1835
rect 2365 1815 2385 1835
rect 2415 1815 2435 1835
rect 2465 1815 2485 1835
rect 2515 1815 2535 1835
rect 2565 1815 2585 1835
rect 2615 1815 2635 1835
rect 2665 1815 2685 1835
rect 2715 1815 2735 1835
rect 2765 1815 2785 1835
rect 2815 1815 2835 1835
rect 2865 1815 2885 1835
rect 2915 1815 2935 1835
rect 2965 1815 2985 1835
rect 3015 1815 3035 1835
rect 3065 1815 3085 1835
rect 3115 1815 3135 1835
rect 3165 1815 3185 1835
rect 3215 1815 3235 1835
rect 3265 1815 3285 1835
rect 3315 1815 3335 1835
rect 3365 1815 3385 1835
rect 3415 1815 3435 1835
rect 3465 1815 3485 1835
rect 3515 1815 3535 1835
rect 3565 1815 3585 1835
rect 3615 1815 3635 1835
rect 3665 1815 3685 1835
rect 3715 1815 3735 1835
rect 3765 1815 3785 1835
rect 3815 1815 3835 1835
rect 3865 1815 3885 1835
rect 3915 1815 3935 1835
rect 3965 1815 3985 1835
rect 4015 1815 4035 1835
rect 4065 1815 4085 1835
rect 4115 1815 4135 1835
rect 4165 1815 4185 1835
rect 4215 1815 4235 1835
rect 4265 1815 4285 1835
rect 4315 1815 4335 1835
rect 4365 1815 4385 1835
rect 4415 1815 4435 1835
rect 4465 1815 4485 1835
rect 4515 1815 4535 1835
rect 4565 1815 4585 1835
rect 4615 1815 4635 1835
rect 4665 1815 4685 1835
rect 4715 1815 4735 1835
rect 4765 1815 4785 1835
rect 4815 1815 4835 1835
rect 4865 1815 4885 1835
rect 4915 1815 4935 1835
rect 4965 1815 4985 1835
rect 5015 1815 5035 1835
rect 5065 1815 5085 1835
rect 5115 1815 5135 1835
rect 5165 1815 5185 1835
rect 5215 1815 5235 1835
rect 5265 1815 5285 1835
rect 5315 1815 5335 1835
rect 5365 1815 5385 1835
rect 5415 1815 5435 1835
rect 5465 1815 5485 1835
rect 5515 1815 5535 1835
rect 5565 1815 5585 1835
rect 5615 1815 5635 1835
rect 5665 1815 5685 1835
rect 5715 1815 5735 1835
rect 5765 1815 5785 1835
rect 5815 1815 5835 1835
rect 5865 1815 5885 1835
rect 5915 1815 5935 1835
rect 5965 1815 5985 1835
rect 6015 1815 6035 1835
rect 6065 1815 6085 1835
rect 6115 1815 6135 1835
rect 6165 1815 6185 1835
rect 6215 1815 6235 1835
rect 6265 1815 6285 1835
rect 6315 1815 6335 1835
rect 6365 1815 6385 1835
rect 6415 1815 6435 1835
rect 6465 1815 6485 1835
rect 6515 1815 6535 1835
rect 6565 1815 6585 1835
rect 6615 1815 6635 1835
rect 6665 1815 6685 1835
rect 6715 1815 6735 1835
rect 6765 1815 6785 1835
rect 6815 1815 6835 1835
rect 6865 1815 6885 1835
rect 6915 1815 6935 1835
rect 6965 1815 6985 1835
rect 7015 1815 7035 1835
rect 7065 1815 7085 1835
rect 7115 1815 7135 1835
rect 7165 1815 7185 1835
rect 7215 1815 7235 1835
rect 7265 1815 7285 1835
rect 7315 1815 7335 1835
rect 7365 1815 7385 1835
rect 7415 1815 7435 1835
rect 7465 1815 7485 1835
rect 7515 1815 7535 1835
rect 7565 1815 7585 1835
rect 7615 1815 7635 1835
rect 7665 1815 7685 1835
rect 7715 1815 7735 1835
rect 7765 1815 7785 1835
rect 7815 1815 7835 1835
rect 7865 1815 7885 1835
rect 7915 1815 7935 1835
rect 7965 1815 7985 1835
rect 8015 1815 8035 1835
rect 8065 1815 8085 1835
rect 8115 1815 8135 1835
rect 8165 1815 8185 1835
rect 8215 1815 8235 1835
rect 8265 1815 8285 1835
rect 8315 1815 8335 1835
rect 8365 1815 8385 1835
rect 8415 1815 8435 1835
rect 8465 1815 8485 1835
rect 8515 1815 8535 1835
rect 8565 1815 8585 1835
rect 8615 1815 8635 1835
rect 8665 1815 8685 1835
rect 8715 1815 8735 1835
rect 8765 1815 8785 1835
rect 8815 1815 8835 1835
rect 8865 1815 8885 1835
rect 8915 1815 8935 1835
rect 8965 1815 8985 1835
rect 9015 1815 9035 1835
rect 9065 1815 9085 1835
rect 9115 1815 9135 1835
rect 9165 1815 9185 1835
rect 9215 1815 9235 1835
rect 9265 1815 9285 1835
rect 9315 1815 9335 1835
rect 9365 1815 9385 1835
rect 9415 1815 9435 1835
rect 9465 1815 9485 1835
rect 9515 1815 9535 1835
rect 9565 1815 9585 1835
rect 9615 1815 9635 1835
rect 9665 1815 9685 1835
rect 9715 1815 9735 1835
rect 9765 1815 9785 1835
rect 9815 1815 9835 1835
rect 9865 1815 9885 1835
rect 9915 1815 9935 1835
rect 9965 1815 9985 1835
rect 10015 1815 10035 1835
rect 10065 1815 10085 1835
rect 10115 1815 10135 1835
rect 10165 1815 10185 1835
rect 10215 1815 10235 1835
rect 10265 1815 10285 1835
rect 10315 1815 10335 1835
rect 10365 1815 10385 1835
rect 10415 1815 10435 1835
rect 10465 1815 10485 1835
rect 10515 1815 10535 1835
rect 10565 1815 10585 1835
rect 10615 1815 10635 1835
rect 10665 1815 10685 1835
rect 10715 1815 10735 1835
rect 10765 1815 10785 1835
rect 10815 1815 10835 1835
rect 10865 1815 10885 1835
rect 10915 1815 10935 1835
rect 10965 1815 10985 1835
rect 11015 1815 11035 1835
rect 11065 1815 11085 1835
rect 11115 1815 11135 1835
rect 11165 1815 11185 1835
rect 11215 1815 11235 1835
rect 11265 1815 11285 1835
rect 11315 1815 11335 1835
rect 11365 1815 11385 1835
rect 11415 1815 11435 1835
rect 11465 1815 11485 1835
rect 11515 1815 11535 1835
rect 11565 1815 11585 1835
rect 11615 1815 11635 1835
rect 11665 1815 11685 1835
rect 11715 1815 11735 1835
rect 11765 1815 11785 1835
rect 11815 1815 11835 1835
rect 11865 1815 11885 1835
rect 11915 1815 11935 1835
rect 11965 1815 11985 1835
rect 12015 1815 12035 1835
rect 12065 1815 12085 1835
rect 12115 1815 12135 1835
rect 12165 1815 12185 1835
rect 12215 1815 12235 1835
rect 12265 1815 12285 1835
rect 12315 1815 12335 1835
rect 12365 1815 12385 1835
rect 12415 1815 12435 1835
rect 12465 1815 12485 1835
rect 12515 1815 12535 1835
rect 12565 1815 12585 1835
rect 12615 1815 12635 1835
rect 12665 1815 12685 1835
rect 12715 1815 12735 1835
rect 12765 1815 12785 1835
rect 12815 1815 12835 1835
rect 12865 1815 12885 1835
rect 12915 1815 12935 1835
rect 12965 1815 12985 1835
rect 13015 1815 13035 1835
rect 13065 1815 13085 1835
rect 13115 1815 13135 1835
rect 13165 1815 13185 1835
rect 13215 1815 13235 1835
rect 13265 1815 13285 1835
rect 13315 1815 13335 1835
rect 13365 1815 13385 1835
rect 13415 1815 13435 1835
rect 13465 1815 13485 1835
rect 13515 1815 13535 1835
rect 13565 1815 13585 1835
rect 13615 1815 13635 1835
rect 13665 1815 13685 1835
rect 13715 1815 13735 1835
rect 13765 1815 13785 1835
rect 13815 1815 13835 1835
rect 13865 1815 13885 1835
rect 13915 1815 13935 1835
rect 13965 1815 13985 1835
rect 14015 1815 14035 1835
rect 14065 1815 14085 1835
rect 14115 1815 14135 1835
rect 14165 1815 14185 1835
rect 14215 1815 14235 1835
rect 14265 1815 14285 1835
rect 14315 1815 14335 1835
rect 14365 1815 14385 1835
rect 14415 1815 14435 1835
rect 14465 1815 14485 1835
rect 14515 1815 14535 1835
rect 14565 1815 14585 1835
rect 14615 1815 14635 1835
rect 14665 1815 14685 1835
rect 14715 1815 14735 1835
rect 14765 1815 14785 1835
rect 14815 1815 14835 1835
rect 14865 1815 14885 1835
rect 14915 1815 14935 1835
rect 14965 1815 14985 1835
rect 15015 1815 15035 1835
rect 15065 1815 15085 1835
rect 15115 1815 15135 1835
rect 15165 1815 15185 1835
rect 15215 1815 15235 1835
rect 15265 1815 15285 1835
rect 15315 1815 15335 1835
rect 15365 1815 15385 1835
rect 15415 1815 15435 1835
rect 15465 1815 15485 1835
rect 15515 1815 15535 1835
rect 15565 1815 15585 1835
rect 15615 1815 15635 1835
rect 15665 1815 15685 1835
rect 15715 1815 15735 1835
rect 15765 1815 15785 1835
rect 15815 1815 15835 1835
rect 15865 1815 15885 1835
rect 15915 1815 15935 1835
rect 15965 1815 15985 1835
rect 16015 1815 16035 1835
rect 16065 1815 16085 1835
rect 16115 1815 16135 1835
rect 16165 1815 16185 1835
rect 16215 1815 16235 1835
rect 16265 1815 16285 1835
rect 16315 1815 16335 1835
rect 16365 1815 16385 1835
rect 16415 1815 16435 1835
rect 16465 1815 16485 1835
rect 16515 1815 16535 1835
rect 16565 1815 16585 1835
rect 16615 1815 16635 1835
rect 16665 1815 16685 1835
rect 16715 1815 16735 1835
rect 16765 1815 16785 1835
rect 16815 1815 16835 1835
rect 16865 1815 16885 1835
rect 16915 1815 16935 1835
rect 16965 1815 16985 1835
rect 17015 1815 17035 1835
rect 17065 1815 17085 1835
rect 17115 1815 17135 1835
rect 17165 1815 17185 1835
rect 17215 1815 17235 1835
rect 17265 1815 17285 1835
rect 17315 1815 17335 1835
rect 17365 1815 17385 1835
rect 17415 1815 17435 1835
rect 17465 1815 17485 1835
rect 17515 1815 17535 1835
rect 17565 1815 17585 1835
rect 17615 1815 17635 1835
rect 17665 1815 17685 1835
rect 17715 1815 17735 1835
rect 17765 1815 17785 1835
rect 17815 1815 17835 1835
rect 17865 1815 17885 1835
rect 17915 1815 17935 1835
rect 17965 1815 17985 1835
rect 18015 1815 18035 1835
rect 18065 1815 18085 1835
rect 18115 1815 18135 1835
rect 18165 1815 18185 1835
rect 18215 1815 18235 1835
rect 18265 1815 18285 1835
rect 18315 1815 18335 1835
rect 18365 1815 18385 1835
rect 18415 1815 18435 1835
rect 18465 1815 18485 1835
rect 18515 1815 18535 1835
rect 18565 1815 18585 1835
rect 18615 1815 18635 1835
rect 18665 1815 18685 1835
rect 18715 1815 18735 1835
rect 18765 1815 18785 1835
rect 18815 1815 18835 1835
rect 18865 1815 18885 1835
rect 18915 1815 18935 1835
rect 18965 1815 18985 1835
rect 19015 1815 19035 1835
rect 19065 1815 19085 1835
rect 19115 1815 19135 1835
rect 19165 1815 19185 1835
rect 19215 1815 19235 1835
rect 19265 1815 19285 1835
rect 19315 1815 19335 1835
rect 19365 1815 19385 1835
rect 19415 1815 19435 1835
rect 19465 1815 19485 1835
rect 19515 1815 19535 1835
rect 19565 1815 19585 1835
rect 19615 1815 19635 1835
rect 19665 1815 19685 1835
rect 19715 1815 19735 1835
rect 19765 1815 19785 1835
rect 19815 1815 19835 1835
rect 19865 1815 19885 1835
rect 19915 1815 19935 1835
rect 19965 1815 19985 1835
rect 20015 1815 20035 1835
rect 20065 1815 20085 1835
rect 20115 1815 20135 1835
rect 20165 1815 20185 1835
rect 20215 1815 20235 1835
rect 20265 1815 20285 1835
rect 20315 1815 20335 1835
rect 20365 1815 20385 1835
rect -635 -1885 -615 -1865
rect -585 -1885 -565 -1865
rect -535 -1885 -515 -1865
rect -485 -1885 -465 -1865
rect -435 -1885 -415 -1865
rect -385 -1885 -365 -1865
rect -335 -1885 -315 -1865
rect -285 -1885 -265 -1865
rect -235 -1885 -215 -1865
rect -185 -1885 -165 -1865
rect -135 -1885 -115 -1865
rect -85 -1885 -65 -1865
rect -35 -1885 -15 -1865
rect 15 -1885 35 -1865
rect 65 -1885 85 -1865
rect 115 -1885 135 -1865
rect 165 -1885 185 -1865
rect 215 -1885 235 -1865
rect 265 -1885 285 -1865
rect 315 -1885 335 -1865
rect 365 -1885 385 -1865
rect 415 -1885 435 -1865
rect 465 -1885 485 -1865
rect 515 -1885 535 -1865
rect 565 -1885 585 -1865
rect 615 -1885 635 -1865
rect 665 -1885 685 -1865
rect 715 -1885 735 -1865
rect 765 -1885 785 -1865
rect 815 -1885 835 -1865
rect 865 -1885 885 -1865
rect 915 -1885 935 -1865
rect 965 -1885 985 -1865
rect 1015 -1885 1035 -1865
rect 1065 -1885 1085 -1865
rect 1115 -1885 1135 -1865
rect 1165 -1885 1185 -1865
rect 1215 -1885 1235 -1865
rect 1265 -1885 1285 -1865
rect 1315 -1885 1335 -1865
rect 1365 -1885 1385 -1865
rect 1415 -1885 1435 -1865
rect 1465 -1885 1485 -1865
rect 1515 -1885 1535 -1865
rect 1565 -1885 1585 -1865
rect 1615 -1885 1635 -1865
rect 1665 -1885 1685 -1865
rect 1715 -1885 1735 -1865
rect 1765 -1885 1785 -1865
rect 1815 -1885 1835 -1865
rect 1865 -1885 1885 -1865
rect 1915 -1885 1935 -1865
rect 1965 -1885 1985 -1865
rect 2015 -1885 2035 -1865
rect 2065 -1885 2085 -1865
rect 2115 -1885 2135 -1865
rect 2165 -1885 2185 -1865
rect 2215 -1885 2235 -1865
rect 2265 -1885 2285 -1865
rect 2315 -1885 2335 -1865
rect 2365 -1885 2385 -1865
rect 2415 -1885 2435 -1865
rect 2465 -1885 2485 -1865
rect 2515 -1885 2535 -1865
rect 2565 -1885 2585 -1865
rect 2615 -1885 2635 -1865
rect 2665 -1885 2685 -1865
rect 2715 -1885 2735 -1865
rect 2765 -1885 2785 -1865
rect 2815 -1885 2835 -1865
rect 2865 -1885 2885 -1865
rect 2915 -1885 2935 -1865
rect 2965 -1885 2985 -1865
rect 3015 -1885 3035 -1865
rect 3065 -1885 3085 -1865
rect 3115 -1885 3135 -1865
rect 3165 -1885 3185 -1865
rect 3215 -1885 3235 -1865
rect 3265 -1885 3285 -1865
rect 3315 -1885 3335 -1865
rect 3365 -1885 3385 -1865
rect 3415 -1885 3435 -1865
rect 3465 -1885 3485 -1865
rect 3515 -1885 3535 -1865
rect 3565 -1885 3585 -1865
rect 3615 -1885 3635 -1865
rect 3665 -1885 3685 -1865
rect 3715 -1885 3735 -1865
rect 3765 -1885 3785 -1865
rect 3815 -1885 3835 -1865
rect 3865 -1885 3885 -1865
rect 3915 -1885 3935 -1865
rect 3965 -1885 3985 -1865
rect 4015 -1885 4035 -1865
rect 4065 -1885 4085 -1865
rect 4115 -1885 4135 -1865
rect 4165 -1885 4185 -1865
rect 4215 -1885 4235 -1865
rect 4265 -1885 4285 -1865
rect 4315 -1885 4335 -1865
rect 4365 -1885 4385 -1865
rect 4415 -1885 4435 -1865
rect 4465 -1885 4485 -1865
rect 4515 -1885 4535 -1865
rect 4565 -1885 4585 -1865
rect 4615 -1885 4635 -1865
rect 4665 -1885 4685 -1865
rect 4715 -1885 4735 -1865
rect 4765 -1885 4785 -1865
rect 4815 -1885 4835 -1865
rect 4865 -1885 4885 -1865
rect 4915 -1885 4935 -1865
rect 4965 -1885 4985 -1865
rect 5015 -1885 5035 -1865
rect 5065 -1885 5085 -1865
rect 5115 -1885 5135 -1865
rect 5165 -1885 5185 -1865
rect 5215 -1885 5235 -1865
rect 5265 -1885 5285 -1865
rect 5315 -1885 5335 -1865
rect 5365 -1885 5385 -1865
rect 5415 -1885 5435 -1865
rect 5465 -1885 5485 -1865
rect 5515 -1885 5535 -1865
rect 5565 -1885 5585 -1865
rect 5615 -1885 5635 -1865
rect 5665 -1885 5685 -1865
rect 5715 -1885 5735 -1865
rect 5765 -1885 5785 -1865
rect 5815 -1885 5835 -1865
rect 5865 -1885 5885 -1865
rect 5915 -1885 5935 -1865
rect 5965 -1885 5985 -1865
rect 6015 -1885 6035 -1865
rect 6065 -1885 6085 -1865
rect 6115 -1885 6135 -1865
rect 6165 -1885 6185 -1865
rect 6215 -1885 6235 -1865
rect 6265 -1885 6285 -1865
rect 6315 -1885 6335 -1865
rect 6365 -1885 6385 -1865
rect 6415 -1885 6435 -1865
rect 6465 -1885 6485 -1865
rect 6515 -1885 6535 -1865
rect 6565 -1885 6585 -1865
rect 6615 -1885 6635 -1865
rect 6665 -1885 6685 -1865
rect 6715 -1885 6735 -1865
rect 6765 -1885 6785 -1865
rect 6815 -1885 6835 -1865
rect 6865 -1885 6885 -1865
rect 6915 -1885 6935 -1865
rect 6965 -1885 6985 -1865
rect 7015 -1885 7035 -1865
rect 7065 -1885 7085 -1865
rect 7115 -1885 7135 -1865
rect 7165 -1885 7185 -1865
rect 7215 -1885 7235 -1865
rect 7265 -1885 7285 -1865
rect 7315 -1885 7335 -1865
rect 7365 -1885 7385 -1865
rect 7415 -1885 7435 -1865
rect 7465 -1885 7485 -1865
rect 7515 -1885 7535 -1865
rect 7565 -1885 7585 -1865
rect 7615 -1885 7635 -1865
rect 7665 -1885 7685 -1865
rect 7715 -1885 7735 -1865
rect 7765 -1885 7785 -1865
rect 7815 -1885 7835 -1865
rect 7865 -1885 7885 -1865
rect 7915 -1885 7935 -1865
rect 7965 -1885 7985 -1865
rect 8015 -1885 8035 -1865
rect 8065 -1885 8085 -1865
rect 8115 -1885 8135 -1865
rect 8165 -1885 8185 -1865
rect 8215 -1885 8235 -1865
rect 8265 -1885 8285 -1865
rect 8315 -1885 8335 -1865
rect 8365 -1885 8385 -1865
rect 8415 -1885 8435 -1865
rect 8465 -1885 8485 -1865
rect 8515 -1885 8535 -1865
rect 8565 -1885 8585 -1865
rect 8615 -1885 8635 -1865
rect 8665 -1885 8685 -1865
rect 8715 -1885 8735 -1865
rect 8765 -1885 8785 -1865
rect 8815 -1885 8835 -1865
rect 8865 -1885 8885 -1865
rect 8915 -1885 8935 -1865
rect 8965 -1885 8985 -1865
rect 9015 -1885 9035 -1865
rect 9065 -1885 9085 -1865
rect 9115 -1885 9135 -1865
rect 9165 -1885 9185 -1865
rect 9215 -1885 9235 -1865
rect 9265 -1885 9285 -1865
rect 9315 -1885 9335 -1865
rect 9365 -1885 9385 -1865
rect 9415 -1885 9435 -1865
rect 9465 -1885 9485 -1865
rect 9515 -1885 9535 -1865
rect 9565 -1885 9585 -1865
rect 9615 -1885 9635 -1865
rect 9665 -1885 9685 -1865
rect 9715 -1885 9735 -1865
rect 9765 -1885 9785 -1865
rect 9815 -1885 9835 -1865
rect 9865 -1885 9885 -1865
rect 9915 -1885 9935 -1865
rect 9965 -1885 9985 -1865
rect 10015 -1885 10035 -1865
rect 10065 -1885 10085 -1865
rect 10115 -1885 10135 -1865
rect 10165 -1885 10185 -1865
rect 10215 -1885 10235 -1865
rect 10265 -1885 10285 -1865
rect 10315 -1885 10335 -1865
rect 10365 -1885 10385 -1865
rect 10415 -1885 10435 -1865
rect 10465 -1885 10485 -1865
rect 10515 -1885 10535 -1865
rect 10565 -1885 10585 -1865
rect 10615 -1885 10635 -1865
rect 10665 -1885 10685 -1865
rect 10715 -1885 10735 -1865
rect 10765 -1885 10785 -1865
rect 10815 -1885 10835 -1865
rect 10865 -1885 10885 -1865
rect 10915 -1885 10935 -1865
rect 10965 -1885 10985 -1865
rect 11015 -1885 11035 -1865
rect 11065 -1885 11085 -1865
rect 11115 -1885 11135 -1865
rect 11165 -1885 11185 -1865
rect 11215 -1885 11235 -1865
rect 11265 -1885 11285 -1865
rect 11315 -1885 11335 -1865
rect 11365 -1885 11385 -1865
rect 11415 -1885 11435 -1865
rect 11465 -1885 11485 -1865
rect 11515 -1885 11535 -1865
rect 11565 -1885 11585 -1865
rect 11615 -1885 11635 -1865
rect 11665 -1885 11685 -1865
rect 11715 -1885 11735 -1865
rect 11765 -1885 11785 -1865
rect 11815 -1885 11835 -1865
rect 11865 -1885 11885 -1865
rect 11915 -1885 11935 -1865
rect 11965 -1885 11985 -1865
rect 12015 -1885 12035 -1865
rect 12065 -1885 12085 -1865
rect 12115 -1885 12135 -1865
rect 12165 -1885 12185 -1865
rect 12215 -1885 12235 -1865
rect 12265 -1885 12285 -1865
rect 12315 -1885 12335 -1865
rect 12365 -1885 12385 -1865
rect 12415 -1885 12435 -1865
rect 12465 -1885 12485 -1865
rect 12515 -1885 12535 -1865
rect 12565 -1885 12585 -1865
rect 12615 -1885 12635 -1865
rect 12665 -1885 12685 -1865
rect 12715 -1885 12735 -1865
rect 12765 -1885 12785 -1865
rect 12815 -1885 12835 -1865
rect 12865 -1885 12885 -1865
rect 12915 -1885 12935 -1865
rect 12965 -1885 12985 -1865
rect 13015 -1885 13035 -1865
rect 13065 -1885 13085 -1865
rect 13115 -1885 13135 -1865
rect 13165 -1885 13185 -1865
rect 13215 -1885 13235 -1865
rect 13265 -1885 13285 -1865
rect 13315 -1885 13335 -1865
rect 13365 -1885 13385 -1865
rect 13415 -1885 13435 -1865
rect 13465 -1885 13485 -1865
rect 13515 -1885 13535 -1865
rect 13565 -1885 13585 -1865
rect 13615 -1885 13635 -1865
rect 13665 -1885 13685 -1865
rect 13715 -1885 13735 -1865
rect 13765 -1885 13785 -1865
rect 13815 -1885 13835 -1865
rect 13865 -1885 13885 -1865
rect 13915 -1885 13935 -1865
rect 13965 -1885 13985 -1865
rect 14015 -1885 14035 -1865
rect 14065 -1885 14085 -1865
rect 14115 -1885 14135 -1865
rect 14165 -1885 14185 -1865
rect 14215 -1885 14235 -1865
rect 14265 -1885 14285 -1865
rect 14315 -1885 14335 -1865
rect 14365 -1885 14385 -1865
rect 14415 -1885 14435 -1865
rect 14465 -1885 14485 -1865
rect 14515 -1885 14535 -1865
rect 14565 -1885 14585 -1865
rect 14615 -1885 14635 -1865
rect 14665 -1885 14685 -1865
rect 14715 -1885 14735 -1865
rect 14765 -1885 14785 -1865
rect 14815 -1885 14835 -1865
rect 14865 -1885 14885 -1865
rect 14915 -1885 14935 -1865
rect 14965 -1885 14985 -1865
rect 15015 -1885 15035 -1865
rect 15065 -1885 15085 -1865
rect 15115 -1885 15135 -1865
rect 15165 -1885 15185 -1865
rect 15215 -1885 15235 -1865
rect 15265 -1885 15285 -1865
rect 15315 -1885 15335 -1865
rect 15365 -1885 15385 -1865
rect 15415 -1885 15435 -1865
rect 15465 -1885 15485 -1865
rect 15515 -1885 15535 -1865
rect 15565 -1885 15585 -1865
rect 15615 -1885 15635 -1865
rect 15665 -1885 15685 -1865
rect 15715 -1885 15735 -1865
rect 15765 -1885 15785 -1865
rect 15815 -1885 15835 -1865
rect 15865 -1885 15885 -1865
rect 15915 -1885 15935 -1865
rect 15965 -1885 15985 -1865
rect 16015 -1885 16035 -1865
rect 16065 -1885 16085 -1865
rect 16115 -1885 16135 -1865
rect 16165 -1885 16185 -1865
rect 16215 -1885 16235 -1865
rect 16265 -1885 16285 -1865
rect 16315 -1885 16335 -1865
rect 16365 -1885 16385 -1865
rect 16415 -1885 16435 -1865
rect 16465 -1885 16485 -1865
rect 16515 -1885 16535 -1865
rect 16565 -1885 16585 -1865
rect 16615 -1885 16635 -1865
rect 16665 -1885 16685 -1865
rect 16715 -1885 16735 -1865
rect 16765 -1885 16785 -1865
rect 16815 -1885 16835 -1865
rect 16865 -1885 16885 -1865
rect 16915 -1885 16935 -1865
rect 16965 -1885 16985 -1865
rect 17015 -1885 17035 -1865
rect 17065 -1885 17085 -1865
rect 17115 -1885 17135 -1865
rect 17165 -1885 17185 -1865
rect 17215 -1885 17235 -1865
rect 17265 -1885 17285 -1865
rect 17315 -1885 17335 -1865
rect 17365 -1885 17385 -1865
rect 17415 -1885 17435 -1865
rect 17465 -1885 17485 -1865
rect 17515 -1885 17535 -1865
rect 17565 -1885 17585 -1865
rect 17615 -1885 17635 -1865
rect 17665 -1885 17685 -1865
rect 17715 -1885 17735 -1865
rect 17765 -1885 17785 -1865
rect 17815 -1885 17835 -1865
rect 17865 -1885 17885 -1865
rect 17915 -1885 17935 -1865
rect 17965 -1885 17985 -1865
rect 18015 -1885 18035 -1865
rect 18065 -1885 18085 -1865
rect 18115 -1885 18135 -1865
rect 18165 -1885 18185 -1865
rect 18215 -1885 18235 -1865
rect 18265 -1885 18285 -1865
rect 18315 -1885 18335 -1865
rect 18365 -1885 18385 -1865
rect 18415 -1885 18435 -1865
rect 18465 -1885 18485 -1865
rect 18515 -1885 18535 -1865
rect 18565 -1885 18585 -1865
rect 18615 -1885 18635 -1865
rect 18665 -1885 18685 -1865
rect 18715 -1885 18735 -1865
rect 18765 -1885 18785 -1865
rect 18815 -1885 18835 -1865
rect 18865 -1885 18885 -1865
rect 18915 -1885 18935 -1865
rect 18965 -1885 18985 -1865
rect 19015 -1885 19035 -1865
rect 19065 -1885 19085 -1865
rect 19115 -1885 19135 -1865
rect 19165 -1885 19185 -1865
rect 19215 -1885 19235 -1865
rect 19265 -1885 19285 -1865
rect 19315 -1885 19335 -1865
rect 19365 -1885 19385 -1865
rect 19415 -1885 19435 -1865
rect 19465 -1885 19485 -1865
rect 19515 -1885 19535 -1865
rect 19565 -1885 19585 -1865
rect 19615 -1885 19635 -1865
rect 19665 -1885 19685 -1865
rect 19715 -1885 19735 -1865
rect 19765 -1885 19785 -1865
rect 19815 -1885 19835 -1865
rect 19865 -1885 19885 -1865
rect 19915 -1885 19935 -1865
rect 19965 -1885 19985 -1865
rect 20015 -1885 20035 -1865
rect 20065 -1885 20085 -1865
rect 20115 -1885 20135 -1865
rect 20165 -1885 20185 -1865
rect 20215 -1885 20235 -1865
rect 20265 -1885 20285 -1865
rect 20315 -1885 20335 -1865
rect 20365 -1885 20385 -1865
<< poly >>
rect -600 5100 -500 5115
rect -450 5100 -350 5115
rect -300 5100 -200 5115
rect -150 5100 -50 5115
rect 0 5100 100 5115
rect 150 5100 250 5115
rect 300 5100 400 5115
rect 450 5100 550 5115
rect 600 5100 700 5115
rect 750 5100 850 5115
rect 900 5100 1000 5115
rect 1050 5100 1150 5115
rect 1200 5100 1300 5115
rect 1350 5100 1450 5115
rect 1500 5100 1600 5115
rect 1650 5100 1750 5115
rect 1800 5100 1900 5115
rect 1950 5100 2050 5115
rect 2100 5100 2200 5115
rect 2250 5100 2350 5115
rect 2400 5100 2500 5115
rect 2550 5100 2650 5115
rect 2700 5100 2800 5115
rect 2850 5100 2950 5115
rect 3000 5100 3100 5115
rect 3150 5100 3250 5115
rect 3300 5100 3400 5115
rect 3450 5100 3550 5115
rect 3600 5100 3700 5115
rect 3750 5100 3850 5115
rect 3900 5100 4000 5115
rect 4050 5100 4150 5115
rect 4200 5100 4300 5115
rect 4350 5100 4450 5115
rect 4500 5100 4600 5115
rect 4650 5100 4750 5115
rect 4800 5100 4900 5115
rect 4950 5100 5050 5115
rect 5100 5100 5200 5115
rect 5250 5100 5350 5115
rect 5400 5100 5500 5115
rect 5550 5100 5650 5115
rect 5700 5100 5800 5115
rect 5850 5100 5950 5115
rect 6000 5100 6100 5115
rect 6150 5100 6250 5115
rect 6300 5100 6400 5115
rect 6450 5100 6550 5115
rect 6600 5100 6700 5115
rect 6750 5100 6850 5115
rect 6900 5100 7000 5115
rect 7050 5100 7150 5115
rect 7200 5100 7300 5115
rect 7350 5100 7450 5115
rect 7500 5100 7600 5115
rect 7650 5100 7750 5115
rect 7800 5100 7900 5115
rect 7950 5100 8050 5115
rect 8100 5100 8200 5115
rect 8250 5100 8350 5115
rect 8400 5100 8500 5115
rect 8550 5100 8650 5115
rect 8700 5100 8800 5115
rect 8850 5100 8950 5115
rect 9000 5100 9100 5115
rect 9150 5100 9250 5115
rect 9300 5100 9400 5115
rect 9450 5100 9550 5115
rect 9600 5100 9700 5115
rect 9750 5100 9850 5115
rect 9900 5100 10000 5115
rect 10050 5100 10150 5115
rect 10200 5100 10300 5115
rect 10350 5100 10450 5115
rect 10500 5100 10600 5115
rect 10650 5100 10750 5115
rect 10800 5100 10900 5115
rect 10950 5100 11050 5115
rect 11100 5100 11200 5115
rect 11250 5100 11350 5115
rect 11400 5100 11500 5115
rect 11550 5100 11650 5115
rect 11700 5100 11800 5115
rect 11850 5100 11950 5115
rect 12000 5100 12100 5115
rect 12150 5100 12250 5115
rect 12300 5100 12400 5115
rect 12450 5100 12550 5115
rect 12600 5100 12700 5115
rect 12750 5100 12850 5115
rect 12900 5100 13000 5115
rect 13050 5100 13150 5115
rect 13200 5100 13300 5115
rect 13350 5100 13450 5115
rect 13500 5100 13600 5115
rect 13650 5100 13750 5115
rect 13800 5100 13900 5115
rect 13950 5100 14050 5115
rect 14100 5100 14200 5115
rect 14250 5100 14350 5115
rect 14400 5100 14500 5115
rect 14550 5100 14650 5115
rect 14700 5100 14800 5115
rect 14850 5100 14950 5115
rect 15000 5100 15100 5115
rect 15150 5100 15250 5115
rect 15300 5100 15400 5115
rect 15450 5100 15550 5115
rect 15600 5100 15700 5115
rect 15750 5100 15850 5115
rect 15900 5100 16000 5115
rect 16050 5100 16150 5115
rect 16200 5100 16300 5115
rect 16350 5100 16450 5115
rect 16500 5100 16600 5115
rect 16650 5100 16750 5115
rect 16800 5100 16900 5115
rect 16950 5100 17050 5115
rect 17100 5100 17200 5115
rect 17250 5100 17350 5115
rect 17400 5100 17500 5115
rect 17550 5100 17650 5115
rect 17700 5100 17800 5115
rect 17850 5100 17950 5115
rect 18000 5100 18100 5115
rect 18150 5100 18250 5115
rect 18300 5100 18400 5115
rect 18450 5100 18550 5115
rect 18600 5100 18700 5115
rect 18750 5100 18850 5115
rect 18900 5100 19000 5115
rect 19050 5100 19150 5115
rect 19200 5100 19300 5115
rect 19350 5100 19450 5115
rect 19500 5100 19600 5115
rect 19650 5100 19750 5115
rect 19800 5100 19900 5115
rect 19950 5100 20050 5115
rect 20100 5100 20200 5115
rect 20250 5100 20350 5115
rect -600 4550 -500 4600
rect -450 4550 -350 4600
rect -600 4535 -350 4550
rect -600 4515 -585 4535
rect -565 4515 -535 4535
rect -515 4515 -485 4535
rect -465 4515 -435 4535
rect -415 4515 -385 4535
rect -365 4515 -350 4535
rect -600 4500 -350 4515
rect -600 4450 -500 4500
rect -450 4450 -350 4500
rect -300 4550 -200 4600
rect -150 4550 -50 4600
rect -300 4535 -50 4550
rect -300 4515 -285 4535
rect -265 4515 -235 4535
rect -215 4515 -185 4535
rect -165 4515 -135 4535
rect -115 4515 -85 4535
rect -65 4515 -50 4535
rect -300 4500 -50 4515
rect -300 4450 -200 4500
rect -150 4450 -50 4500
rect 0 4550 100 4600
rect 150 4550 250 4600
rect 0 4535 250 4550
rect 0 4515 15 4535
rect 35 4515 65 4535
rect 85 4515 115 4535
rect 135 4515 165 4535
rect 185 4515 215 4535
rect 235 4515 250 4535
rect 0 4500 250 4515
rect 0 4450 100 4500
rect 150 4450 250 4500
rect 300 4550 400 4600
rect 450 4550 550 4600
rect 300 4535 550 4550
rect 300 4515 315 4535
rect 335 4515 365 4535
rect 385 4515 415 4535
rect 435 4515 465 4535
rect 485 4515 515 4535
rect 535 4515 550 4535
rect 300 4500 550 4515
rect 300 4450 400 4500
rect 450 4450 550 4500
rect 600 4550 700 4600
rect 750 4550 850 4600
rect 600 4535 850 4550
rect 600 4515 615 4535
rect 635 4515 665 4535
rect 685 4515 715 4535
rect 735 4515 765 4535
rect 785 4515 815 4535
rect 835 4515 850 4535
rect 600 4500 850 4515
rect 600 4450 700 4500
rect 750 4450 850 4500
rect 900 4550 1000 4600
rect 1050 4550 1150 4600
rect 900 4535 1150 4550
rect 900 4515 915 4535
rect 935 4515 965 4535
rect 985 4515 1015 4535
rect 1035 4515 1065 4535
rect 1085 4515 1115 4535
rect 1135 4515 1150 4535
rect 900 4500 1150 4515
rect 900 4450 1000 4500
rect 1050 4450 1150 4500
rect 1200 4550 1300 4600
rect 1350 4550 1450 4600
rect 1200 4535 1450 4550
rect 1200 4515 1215 4535
rect 1235 4515 1265 4535
rect 1285 4515 1315 4535
rect 1335 4515 1365 4535
rect 1385 4515 1415 4535
rect 1435 4515 1450 4535
rect 1200 4500 1450 4515
rect 1200 4450 1300 4500
rect 1350 4450 1450 4500
rect 1500 4550 1600 4600
rect 1650 4550 1750 4600
rect 1500 4535 1750 4550
rect 1500 4515 1515 4535
rect 1535 4515 1565 4535
rect 1585 4515 1615 4535
rect 1635 4515 1665 4535
rect 1685 4515 1715 4535
rect 1735 4515 1750 4535
rect 1500 4500 1750 4515
rect 1500 4450 1600 4500
rect 1650 4450 1750 4500
rect 1800 4550 1900 4600
rect 1950 4550 2050 4600
rect 1800 4535 2050 4550
rect 1800 4515 1815 4535
rect 1835 4515 1865 4535
rect 1885 4515 1915 4535
rect 1935 4515 1965 4535
rect 1985 4515 2015 4535
rect 2035 4515 2050 4535
rect 1800 4500 2050 4515
rect 1800 4450 1900 4500
rect 1950 4450 2050 4500
rect 2100 4550 2200 4600
rect 2250 4550 2350 4600
rect 2100 4535 2350 4550
rect 2100 4515 2115 4535
rect 2135 4515 2165 4535
rect 2185 4515 2215 4535
rect 2235 4515 2265 4535
rect 2285 4515 2315 4535
rect 2335 4515 2350 4535
rect 2100 4500 2350 4515
rect 2100 4450 2200 4500
rect 2250 4450 2350 4500
rect 2400 4550 2500 4600
rect 2550 4550 2650 4600
rect 2400 4535 2650 4550
rect 2400 4515 2415 4535
rect 2435 4515 2465 4535
rect 2485 4515 2515 4535
rect 2535 4515 2565 4535
rect 2585 4515 2615 4535
rect 2635 4515 2650 4535
rect 2400 4500 2650 4515
rect 2400 4450 2500 4500
rect 2550 4450 2650 4500
rect 2700 4550 2800 4600
rect 2850 4550 2950 4600
rect 2700 4535 2950 4550
rect 2700 4515 2715 4535
rect 2735 4515 2765 4535
rect 2785 4515 2815 4535
rect 2835 4515 2865 4535
rect 2885 4515 2915 4535
rect 2935 4515 2950 4535
rect 2700 4500 2950 4515
rect 2700 4450 2800 4500
rect 2850 4450 2950 4500
rect 3000 4550 3100 4600
rect 3150 4550 3250 4600
rect 3000 4535 3250 4550
rect 3000 4515 3015 4535
rect 3035 4515 3065 4535
rect 3085 4515 3115 4535
rect 3135 4515 3165 4535
rect 3185 4515 3215 4535
rect 3235 4515 3250 4535
rect 3000 4500 3250 4515
rect 3000 4450 3100 4500
rect 3150 4450 3250 4500
rect 3300 4550 3400 4600
rect 3450 4550 3550 4600
rect 3300 4535 3550 4550
rect 3300 4515 3315 4535
rect 3335 4515 3365 4535
rect 3385 4515 3415 4535
rect 3435 4515 3465 4535
rect 3485 4515 3515 4535
rect 3535 4515 3550 4535
rect 3300 4500 3550 4515
rect 3300 4450 3400 4500
rect 3450 4450 3550 4500
rect 3600 4550 3700 4600
rect 3750 4550 3850 4600
rect 3600 4535 3850 4550
rect 3600 4515 3615 4535
rect 3635 4515 3665 4535
rect 3685 4515 3715 4535
rect 3735 4515 3765 4535
rect 3785 4515 3815 4535
rect 3835 4515 3850 4535
rect 3600 4500 3850 4515
rect 3600 4450 3700 4500
rect 3750 4450 3850 4500
rect 3900 4550 4000 4600
rect 4050 4550 4150 4600
rect 3900 4535 4150 4550
rect 3900 4515 3915 4535
rect 3935 4515 3965 4535
rect 3985 4515 4015 4535
rect 4035 4515 4065 4535
rect 4085 4515 4115 4535
rect 4135 4515 4150 4535
rect 3900 4500 4150 4515
rect 3900 4450 4000 4500
rect 4050 4450 4150 4500
rect 4200 4550 4300 4600
rect 4350 4550 4450 4600
rect 4200 4535 4450 4550
rect 4200 4515 4215 4535
rect 4235 4515 4265 4535
rect 4285 4515 4315 4535
rect 4335 4515 4365 4535
rect 4385 4515 4415 4535
rect 4435 4515 4450 4535
rect 4200 4500 4450 4515
rect 4200 4450 4300 4500
rect 4350 4450 4450 4500
rect 4500 4550 4600 4600
rect 4650 4550 4750 4600
rect 4500 4535 4750 4550
rect 4500 4515 4515 4535
rect 4535 4515 4565 4535
rect 4585 4515 4615 4535
rect 4635 4515 4665 4535
rect 4685 4515 4715 4535
rect 4735 4515 4750 4535
rect 4500 4500 4750 4515
rect 4500 4450 4600 4500
rect 4650 4450 4750 4500
rect 4800 4550 4900 4600
rect 4950 4550 5050 4600
rect 4800 4535 5050 4550
rect 4800 4515 4815 4535
rect 4835 4515 4865 4535
rect 4885 4515 4915 4535
rect 4935 4515 4965 4535
rect 4985 4515 5015 4535
rect 5035 4515 5050 4535
rect 4800 4500 5050 4515
rect 4800 4450 4900 4500
rect 4950 4450 5050 4500
rect 5100 4550 5200 4600
rect 5250 4550 5350 4600
rect 5100 4535 5350 4550
rect 5100 4515 5115 4535
rect 5135 4515 5165 4535
rect 5185 4515 5215 4535
rect 5235 4515 5265 4535
rect 5285 4515 5315 4535
rect 5335 4515 5350 4535
rect 5100 4500 5350 4515
rect 5100 4450 5200 4500
rect 5250 4450 5350 4500
rect 5400 4550 5500 4600
rect 5550 4550 5650 4600
rect 5400 4535 5650 4550
rect 5400 4515 5415 4535
rect 5435 4515 5465 4535
rect 5485 4515 5515 4535
rect 5535 4515 5565 4535
rect 5585 4515 5615 4535
rect 5635 4515 5650 4535
rect 5400 4500 5650 4515
rect 5400 4450 5500 4500
rect 5550 4450 5650 4500
rect 5700 4550 5800 4600
rect 5850 4550 5950 4600
rect 5700 4535 5950 4550
rect 5700 4515 5715 4535
rect 5735 4515 5765 4535
rect 5785 4515 5815 4535
rect 5835 4515 5865 4535
rect 5885 4515 5915 4535
rect 5935 4515 5950 4535
rect 5700 4500 5950 4515
rect 5700 4450 5800 4500
rect 5850 4450 5950 4500
rect 6000 4550 6100 4600
rect 6150 4550 6250 4600
rect 6000 4535 6250 4550
rect 6000 4515 6015 4535
rect 6035 4515 6065 4535
rect 6085 4515 6115 4535
rect 6135 4515 6165 4535
rect 6185 4515 6215 4535
rect 6235 4515 6250 4535
rect 6000 4500 6250 4515
rect 6000 4450 6100 4500
rect 6150 4450 6250 4500
rect 6300 4550 6400 4600
rect 6450 4550 6550 4600
rect 6300 4535 6550 4550
rect 6300 4515 6315 4535
rect 6335 4515 6365 4535
rect 6385 4515 6415 4535
rect 6435 4515 6465 4535
rect 6485 4515 6515 4535
rect 6535 4515 6550 4535
rect 6300 4500 6550 4515
rect 6300 4450 6400 4500
rect 6450 4450 6550 4500
rect 6600 4550 6700 4600
rect 6750 4550 6850 4600
rect 6600 4535 6850 4550
rect 6600 4515 6615 4535
rect 6635 4515 6665 4535
rect 6685 4515 6715 4535
rect 6735 4515 6765 4535
rect 6785 4515 6815 4535
rect 6835 4515 6850 4535
rect 6600 4500 6850 4515
rect 6600 4450 6700 4500
rect 6750 4450 6850 4500
rect 6900 4550 7000 4600
rect 7050 4550 7150 4600
rect 6900 4535 7150 4550
rect 6900 4515 6915 4535
rect 6935 4515 6965 4535
rect 6985 4515 7015 4535
rect 7035 4515 7065 4535
rect 7085 4515 7115 4535
rect 7135 4515 7150 4535
rect 6900 4500 7150 4515
rect 6900 4450 7000 4500
rect 7050 4450 7150 4500
rect 7200 4550 7300 4600
rect 7350 4550 7450 4600
rect 7200 4535 7450 4550
rect 7200 4515 7215 4535
rect 7235 4515 7265 4535
rect 7285 4515 7315 4535
rect 7335 4515 7365 4535
rect 7385 4515 7415 4535
rect 7435 4515 7450 4535
rect 7200 4500 7450 4515
rect 7200 4450 7300 4500
rect 7350 4450 7450 4500
rect 7500 4550 7600 4600
rect 7650 4550 7750 4600
rect 7500 4535 7750 4550
rect 7500 4515 7515 4535
rect 7535 4515 7565 4535
rect 7585 4515 7615 4535
rect 7635 4515 7665 4535
rect 7685 4515 7715 4535
rect 7735 4515 7750 4535
rect 7500 4500 7750 4515
rect 7500 4450 7600 4500
rect 7650 4450 7750 4500
rect 7800 4550 7900 4600
rect 7950 4550 8050 4600
rect 7800 4535 8050 4550
rect 7800 4515 7815 4535
rect 7835 4515 7865 4535
rect 7885 4515 7915 4535
rect 7935 4515 7965 4535
rect 7985 4515 8015 4535
rect 8035 4515 8050 4535
rect 7800 4500 8050 4515
rect 7800 4450 7900 4500
rect 7950 4450 8050 4500
rect 8100 4550 8200 4600
rect 8250 4550 8350 4600
rect 8100 4535 8350 4550
rect 8100 4515 8115 4535
rect 8135 4515 8165 4535
rect 8185 4515 8215 4535
rect 8235 4515 8265 4535
rect 8285 4515 8315 4535
rect 8335 4515 8350 4535
rect 8100 4500 8350 4515
rect 8100 4450 8200 4500
rect 8250 4450 8350 4500
rect 8400 4550 8500 4600
rect 8550 4550 8650 4600
rect 8400 4535 8650 4550
rect 8400 4515 8415 4535
rect 8435 4515 8465 4535
rect 8485 4515 8515 4535
rect 8535 4515 8565 4535
rect 8585 4515 8615 4535
rect 8635 4515 8650 4535
rect 8400 4500 8650 4515
rect 8400 4450 8500 4500
rect 8550 4450 8650 4500
rect 8700 4550 8800 4600
rect 8850 4550 8950 4600
rect 8700 4535 8950 4550
rect 8700 4515 8715 4535
rect 8735 4515 8765 4535
rect 8785 4515 8815 4535
rect 8835 4515 8865 4535
rect 8885 4515 8915 4535
rect 8935 4515 8950 4535
rect 8700 4500 8950 4515
rect 8700 4450 8800 4500
rect 8850 4450 8950 4500
rect 9000 4550 9100 4600
rect 9150 4550 9250 4600
rect 9000 4535 9250 4550
rect 9000 4515 9015 4535
rect 9035 4515 9065 4535
rect 9085 4515 9115 4535
rect 9135 4515 9165 4535
rect 9185 4515 9215 4535
rect 9235 4515 9250 4535
rect 9000 4500 9250 4515
rect 9000 4450 9100 4500
rect 9150 4450 9250 4500
rect 9300 4550 9400 4600
rect 9450 4550 9550 4600
rect 9300 4535 9550 4550
rect 9300 4515 9315 4535
rect 9335 4515 9365 4535
rect 9385 4515 9415 4535
rect 9435 4515 9465 4535
rect 9485 4515 9515 4535
rect 9535 4515 9550 4535
rect 9300 4500 9550 4515
rect 9300 4450 9400 4500
rect 9450 4450 9550 4500
rect 9600 4550 9700 4600
rect 9750 4550 9850 4600
rect 9600 4535 9850 4550
rect 9600 4515 9615 4535
rect 9635 4515 9665 4535
rect 9685 4515 9715 4535
rect 9735 4515 9765 4535
rect 9785 4515 9815 4535
rect 9835 4515 9850 4535
rect 9600 4500 9850 4515
rect 9600 4450 9700 4500
rect 9750 4450 9850 4500
rect 9900 4550 10000 4600
rect 10050 4550 10150 4600
rect 9900 4535 10150 4550
rect 9900 4515 9915 4535
rect 9935 4515 9965 4535
rect 9985 4515 10015 4535
rect 10035 4515 10065 4535
rect 10085 4515 10115 4535
rect 10135 4515 10150 4535
rect 9900 4500 10150 4515
rect 9900 4450 10000 4500
rect 10050 4450 10150 4500
rect 10200 4550 10300 4600
rect 10350 4550 10450 4600
rect 10200 4535 10450 4550
rect 10200 4515 10215 4535
rect 10235 4515 10265 4535
rect 10285 4515 10315 4535
rect 10335 4515 10365 4535
rect 10385 4515 10415 4535
rect 10435 4515 10450 4535
rect 10200 4500 10450 4515
rect 10200 4450 10300 4500
rect 10350 4450 10450 4500
rect 10500 4550 10600 4600
rect 10650 4550 10750 4600
rect 10500 4535 10750 4550
rect 10500 4515 10515 4535
rect 10535 4515 10565 4535
rect 10585 4515 10615 4535
rect 10635 4515 10665 4535
rect 10685 4515 10715 4535
rect 10735 4515 10750 4535
rect 10500 4500 10750 4515
rect 10500 4450 10600 4500
rect 10650 4450 10750 4500
rect 10800 4550 10900 4600
rect 10950 4550 11050 4600
rect 10800 4535 11050 4550
rect 10800 4515 10815 4535
rect 10835 4515 10865 4535
rect 10885 4515 10915 4535
rect 10935 4515 10965 4535
rect 10985 4515 11015 4535
rect 11035 4515 11050 4535
rect 10800 4500 11050 4515
rect 10800 4450 10900 4500
rect 10950 4450 11050 4500
rect 11100 4550 11200 4600
rect 11250 4550 11350 4600
rect 11100 4535 11350 4550
rect 11100 4515 11115 4535
rect 11135 4515 11165 4535
rect 11185 4515 11215 4535
rect 11235 4515 11265 4535
rect 11285 4515 11315 4535
rect 11335 4515 11350 4535
rect 11100 4500 11350 4515
rect 11100 4450 11200 4500
rect 11250 4450 11350 4500
rect 11400 4550 11500 4600
rect 11550 4550 11650 4600
rect 11400 4535 11650 4550
rect 11400 4515 11415 4535
rect 11435 4515 11465 4535
rect 11485 4515 11515 4535
rect 11535 4515 11565 4535
rect 11585 4515 11615 4535
rect 11635 4515 11650 4535
rect 11400 4500 11650 4515
rect 11400 4450 11500 4500
rect 11550 4450 11650 4500
rect 11700 4550 11800 4600
rect 11850 4550 11950 4600
rect 11700 4535 11950 4550
rect 11700 4515 11715 4535
rect 11735 4515 11765 4535
rect 11785 4515 11815 4535
rect 11835 4515 11865 4535
rect 11885 4515 11915 4535
rect 11935 4515 11950 4535
rect 11700 4500 11950 4515
rect 11700 4450 11800 4500
rect 11850 4450 11950 4500
rect 12000 4550 12100 4600
rect 12150 4550 12250 4600
rect 12000 4535 12250 4550
rect 12000 4515 12015 4535
rect 12035 4515 12065 4535
rect 12085 4515 12115 4535
rect 12135 4515 12165 4535
rect 12185 4515 12215 4535
rect 12235 4515 12250 4535
rect 12000 4500 12250 4515
rect 12000 4450 12100 4500
rect 12150 4450 12250 4500
rect 12300 4550 12400 4600
rect 12450 4550 12550 4600
rect 12300 4535 12550 4550
rect 12300 4515 12315 4535
rect 12335 4515 12365 4535
rect 12385 4515 12415 4535
rect 12435 4515 12465 4535
rect 12485 4515 12515 4535
rect 12535 4515 12550 4535
rect 12300 4500 12550 4515
rect 12300 4450 12400 4500
rect 12450 4450 12550 4500
rect 12600 4550 12700 4600
rect 12750 4550 12850 4600
rect 12600 4535 12850 4550
rect 12600 4515 12615 4535
rect 12635 4515 12665 4535
rect 12685 4515 12715 4535
rect 12735 4515 12765 4535
rect 12785 4515 12815 4535
rect 12835 4515 12850 4535
rect 12600 4500 12850 4515
rect 12600 4450 12700 4500
rect 12750 4450 12850 4500
rect 12900 4550 13000 4600
rect 13050 4550 13150 4600
rect 12900 4535 13150 4550
rect 12900 4515 12915 4535
rect 12935 4515 12965 4535
rect 12985 4515 13015 4535
rect 13035 4515 13065 4535
rect 13085 4515 13115 4535
rect 13135 4515 13150 4535
rect 12900 4500 13150 4515
rect 12900 4450 13000 4500
rect 13050 4450 13150 4500
rect 13200 4550 13300 4600
rect 13350 4550 13450 4600
rect 13200 4535 13450 4550
rect 13200 4515 13215 4535
rect 13235 4515 13265 4535
rect 13285 4515 13315 4535
rect 13335 4515 13365 4535
rect 13385 4515 13415 4535
rect 13435 4515 13450 4535
rect 13200 4500 13450 4515
rect 13200 4450 13300 4500
rect 13350 4450 13450 4500
rect 13500 4550 13600 4600
rect 13650 4550 13750 4600
rect 13500 4535 13750 4550
rect 13500 4515 13515 4535
rect 13535 4515 13565 4535
rect 13585 4515 13615 4535
rect 13635 4515 13665 4535
rect 13685 4515 13715 4535
rect 13735 4515 13750 4535
rect 13500 4500 13750 4515
rect 13500 4450 13600 4500
rect 13650 4450 13750 4500
rect 13800 4550 13900 4600
rect 13950 4550 14050 4600
rect 13800 4535 14050 4550
rect 13800 4515 13815 4535
rect 13835 4515 13865 4535
rect 13885 4515 13915 4535
rect 13935 4515 13965 4535
rect 13985 4515 14015 4535
rect 14035 4515 14050 4535
rect 13800 4500 14050 4515
rect 13800 4450 13900 4500
rect 13950 4450 14050 4500
rect 14100 4550 14200 4600
rect 14250 4550 14350 4600
rect 14100 4535 14350 4550
rect 14100 4515 14115 4535
rect 14135 4515 14165 4535
rect 14185 4515 14215 4535
rect 14235 4515 14265 4535
rect 14285 4515 14315 4535
rect 14335 4515 14350 4535
rect 14100 4500 14350 4515
rect 14100 4450 14200 4500
rect 14250 4450 14350 4500
rect 14400 4550 14500 4600
rect 14550 4550 14650 4600
rect 14400 4535 14650 4550
rect 14400 4515 14415 4535
rect 14435 4515 14465 4535
rect 14485 4515 14515 4535
rect 14535 4515 14565 4535
rect 14585 4515 14615 4535
rect 14635 4515 14650 4535
rect 14400 4500 14650 4515
rect 14400 4450 14500 4500
rect 14550 4450 14650 4500
rect 14700 4550 14800 4600
rect 14850 4550 14950 4600
rect 14700 4535 14950 4550
rect 14700 4515 14715 4535
rect 14735 4515 14765 4535
rect 14785 4515 14815 4535
rect 14835 4515 14865 4535
rect 14885 4515 14915 4535
rect 14935 4515 14950 4535
rect 14700 4500 14950 4515
rect 14700 4450 14800 4500
rect 14850 4450 14950 4500
rect 15000 4550 15100 4600
rect 15150 4550 15250 4600
rect 15000 4535 15250 4550
rect 15000 4515 15015 4535
rect 15035 4515 15065 4535
rect 15085 4515 15115 4535
rect 15135 4515 15165 4535
rect 15185 4515 15215 4535
rect 15235 4515 15250 4535
rect 15000 4500 15250 4515
rect 15000 4450 15100 4500
rect 15150 4450 15250 4500
rect 15300 4550 15400 4600
rect 15450 4550 15550 4600
rect 15300 4535 15550 4550
rect 15300 4515 15315 4535
rect 15335 4515 15365 4535
rect 15385 4515 15415 4535
rect 15435 4515 15465 4535
rect 15485 4515 15515 4535
rect 15535 4515 15550 4535
rect 15300 4500 15550 4515
rect 15300 4450 15400 4500
rect 15450 4450 15550 4500
rect 15600 4550 15700 4600
rect 15750 4550 15850 4600
rect 15600 4535 15850 4550
rect 15600 4515 15615 4535
rect 15635 4515 15665 4535
rect 15685 4515 15715 4535
rect 15735 4515 15765 4535
rect 15785 4515 15815 4535
rect 15835 4515 15850 4535
rect 15600 4500 15850 4515
rect 15600 4450 15700 4500
rect 15750 4450 15850 4500
rect 15900 4550 16000 4600
rect 16050 4550 16150 4600
rect 15900 4535 16150 4550
rect 15900 4515 15915 4535
rect 15935 4515 15965 4535
rect 15985 4515 16015 4535
rect 16035 4515 16065 4535
rect 16085 4515 16115 4535
rect 16135 4515 16150 4535
rect 15900 4500 16150 4515
rect 15900 4450 16000 4500
rect 16050 4450 16150 4500
rect 16200 4550 16300 4600
rect 16350 4550 16450 4600
rect 16200 4535 16450 4550
rect 16200 4515 16215 4535
rect 16235 4515 16265 4535
rect 16285 4515 16315 4535
rect 16335 4515 16365 4535
rect 16385 4515 16415 4535
rect 16435 4515 16450 4535
rect 16200 4500 16450 4515
rect 16200 4450 16300 4500
rect 16350 4450 16450 4500
rect 16500 4550 16600 4600
rect 16650 4550 16750 4600
rect 16500 4535 16750 4550
rect 16500 4515 16515 4535
rect 16535 4515 16565 4535
rect 16585 4515 16615 4535
rect 16635 4515 16665 4535
rect 16685 4515 16715 4535
rect 16735 4515 16750 4535
rect 16500 4500 16750 4515
rect 16500 4450 16600 4500
rect 16650 4450 16750 4500
rect 16800 4550 16900 4600
rect 16950 4550 17050 4600
rect 16800 4535 17050 4550
rect 16800 4515 16815 4535
rect 16835 4515 16865 4535
rect 16885 4515 16915 4535
rect 16935 4515 16965 4535
rect 16985 4515 17015 4535
rect 17035 4515 17050 4535
rect 16800 4500 17050 4515
rect 16800 4450 16900 4500
rect 16950 4450 17050 4500
rect 17100 4550 17200 4600
rect 17250 4550 17350 4600
rect 17100 4535 17350 4550
rect 17100 4515 17115 4535
rect 17135 4515 17165 4535
rect 17185 4515 17215 4535
rect 17235 4515 17265 4535
rect 17285 4515 17315 4535
rect 17335 4515 17350 4535
rect 17100 4500 17350 4515
rect 17100 4450 17200 4500
rect 17250 4450 17350 4500
rect 17400 4550 17500 4600
rect 17550 4550 17650 4600
rect 17400 4535 17650 4550
rect 17400 4515 17415 4535
rect 17435 4515 17465 4535
rect 17485 4515 17515 4535
rect 17535 4515 17565 4535
rect 17585 4515 17615 4535
rect 17635 4515 17650 4535
rect 17400 4500 17650 4515
rect 17400 4450 17500 4500
rect 17550 4450 17650 4500
rect 17700 4550 17800 4600
rect 17850 4550 17950 4600
rect 17700 4535 17950 4550
rect 17700 4515 17715 4535
rect 17735 4515 17765 4535
rect 17785 4515 17815 4535
rect 17835 4515 17865 4535
rect 17885 4515 17915 4535
rect 17935 4515 17950 4535
rect 17700 4500 17950 4515
rect 17700 4450 17800 4500
rect 17850 4450 17950 4500
rect 18000 4550 18100 4600
rect 18150 4550 18250 4600
rect 18000 4535 18250 4550
rect 18000 4515 18015 4535
rect 18035 4515 18065 4535
rect 18085 4515 18115 4535
rect 18135 4515 18165 4535
rect 18185 4515 18215 4535
rect 18235 4515 18250 4535
rect 18000 4500 18250 4515
rect 18000 4450 18100 4500
rect 18150 4450 18250 4500
rect 18300 4550 18400 4600
rect 18450 4550 18550 4600
rect 18300 4535 18550 4550
rect 18300 4515 18315 4535
rect 18335 4515 18365 4535
rect 18385 4515 18415 4535
rect 18435 4515 18465 4535
rect 18485 4515 18515 4535
rect 18535 4515 18550 4535
rect 18300 4500 18550 4515
rect 18300 4450 18400 4500
rect 18450 4450 18550 4500
rect 18600 4550 18700 4600
rect 18750 4550 18850 4600
rect 18600 4535 18850 4550
rect 18600 4515 18615 4535
rect 18635 4515 18665 4535
rect 18685 4515 18715 4535
rect 18735 4515 18765 4535
rect 18785 4515 18815 4535
rect 18835 4515 18850 4535
rect 18600 4500 18850 4515
rect 18600 4450 18700 4500
rect 18750 4450 18850 4500
rect 18900 4550 19000 4600
rect 19050 4550 19150 4600
rect 18900 4535 19150 4550
rect 18900 4515 18915 4535
rect 18935 4515 18965 4535
rect 18985 4515 19015 4535
rect 19035 4515 19065 4535
rect 19085 4515 19115 4535
rect 19135 4515 19150 4535
rect 18900 4500 19150 4515
rect 18900 4450 19000 4500
rect 19050 4450 19150 4500
rect 19200 4550 19300 4600
rect 19350 4550 19450 4600
rect 19200 4535 19450 4550
rect 19200 4515 19215 4535
rect 19235 4515 19265 4535
rect 19285 4515 19315 4535
rect 19335 4515 19365 4535
rect 19385 4515 19415 4535
rect 19435 4515 19450 4535
rect 19200 4500 19450 4515
rect 19200 4450 19300 4500
rect 19350 4450 19450 4500
rect 19500 4550 19600 4600
rect 19650 4550 19750 4600
rect 19500 4535 19750 4550
rect 19500 4515 19515 4535
rect 19535 4515 19565 4535
rect 19585 4515 19615 4535
rect 19635 4515 19665 4535
rect 19685 4515 19715 4535
rect 19735 4515 19750 4535
rect 19500 4500 19750 4515
rect 19500 4450 19600 4500
rect 19650 4450 19750 4500
rect 19800 4550 19900 4600
rect 19950 4550 20050 4600
rect 19800 4535 20050 4550
rect 19800 4515 19815 4535
rect 19835 4515 19865 4535
rect 19885 4515 19915 4535
rect 19935 4515 19965 4535
rect 19985 4515 20015 4535
rect 20035 4515 20050 4535
rect 19800 4500 20050 4515
rect 19800 4450 19900 4500
rect 19950 4450 20050 4500
rect 20100 4550 20200 4600
rect 20250 4550 20350 4600
rect 20100 4535 20350 4550
rect 20100 4515 20115 4535
rect 20135 4515 20165 4535
rect 20185 4515 20215 4535
rect 20235 4515 20265 4535
rect 20285 4515 20315 4535
rect 20335 4515 20350 4535
rect 20100 4500 20350 4515
rect 20100 4450 20200 4500
rect 20250 4450 20350 4500
rect -600 3935 -500 3950
rect -450 3935 -350 3950
rect -300 3935 -200 3950
rect -150 3935 -50 3950
rect 0 3935 100 3950
rect 150 3935 250 3950
rect 300 3935 400 3950
rect 450 3935 550 3950
rect 600 3935 700 3950
rect 750 3935 850 3950
rect 900 3935 1000 3950
rect 1050 3935 1150 3950
rect 1200 3935 1300 3950
rect 1350 3935 1450 3950
rect 1500 3935 1600 3950
rect 1650 3935 1750 3950
rect 1800 3935 1900 3950
rect 1950 3935 2050 3950
rect 2100 3935 2200 3950
rect 2250 3935 2350 3950
rect 2400 3935 2500 3950
rect 2550 3935 2650 3950
rect 2700 3935 2800 3950
rect 2850 3935 2950 3950
rect 3000 3935 3100 3950
rect 3150 3935 3250 3950
rect 3300 3935 3400 3950
rect 3450 3935 3550 3950
rect 3600 3935 3700 3950
rect 3750 3935 3850 3950
rect 3900 3935 4000 3950
rect 4050 3935 4150 3950
rect 4200 3935 4300 3950
rect 4350 3935 4450 3950
rect 4500 3935 4600 3950
rect 4650 3935 4750 3950
rect 4800 3935 4900 3950
rect 4950 3935 5050 3950
rect 5100 3935 5200 3950
rect 5250 3935 5350 3950
rect 5400 3935 5500 3950
rect 5550 3935 5650 3950
rect 5700 3935 5800 3950
rect 5850 3935 5950 3950
rect 6000 3935 6100 3950
rect 6150 3935 6250 3950
rect 6300 3935 6400 3950
rect 6450 3935 6550 3950
rect 6600 3935 6700 3950
rect 6750 3935 6850 3950
rect 6900 3935 7000 3950
rect 7050 3935 7150 3950
rect 7200 3935 7300 3950
rect 7350 3935 7450 3950
rect 7500 3935 7600 3950
rect 7650 3935 7750 3950
rect 7800 3935 7900 3950
rect 7950 3935 8050 3950
rect 8100 3935 8200 3950
rect 8250 3935 8350 3950
rect 8400 3935 8500 3950
rect 8550 3935 8650 3950
rect 8700 3935 8800 3950
rect 8850 3935 8950 3950
rect 9000 3935 9100 3950
rect 9150 3935 9250 3950
rect 9300 3935 9400 3950
rect 9450 3935 9550 3950
rect 9600 3935 9700 3950
rect 9750 3935 9850 3950
rect 9900 3935 10000 3950
rect 10050 3935 10150 3950
rect 10200 3935 10300 3950
rect 10350 3935 10450 3950
rect 10500 3935 10600 3950
rect 10650 3935 10750 3950
rect 10800 3935 10900 3950
rect 10950 3935 11050 3950
rect 11100 3935 11200 3950
rect 11250 3935 11350 3950
rect 11400 3935 11500 3950
rect 11550 3935 11650 3950
rect 11700 3935 11800 3950
rect 11850 3935 11950 3950
rect 12000 3935 12100 3950
rect 12150 3935 12250 3950
rect 12300 3935 12400 3950
rect 12450 3935 12550 3950
rect 12600 3935 12700 3950
rect 12750 3935 12850 3950
rect 12900 3935 13000 3950
rect 13050 3935 13150 3950
rect 13200 3935 13300 3950
rect 13350 3935 13450 3950
rect 13500 3935 13600 3950
rect 13650 3935 13750 3950
rect 13800 3935 13900 3950
rect 13950 3935 14050 3950
rect 14100 3935 14200 3950
rect 14250 3935 14350 3950
rect 14400 3935 14500 3950
rect 14550 3935 14650 3950
rect 14700 3935 14800 3950
rect 14850 3935 14950 3950
rect 15000 3935 15100 3950
rect 15150 3935 15250 3950
rect 15300 3935 15400 3950
rect 15450 3935 15550 3950
rect 15600 3935 15700 3950
rect 15750 3935 15850 3950
rect 15900 3935 16000 3950
rect 16050 3935 16150 3950
rect 16200 3935 16300 3950
rect 16350 3935 16450 3950
rect 16500 3935 16600 3950
rect 16650 3935 16750 3950
rect 16800 3935 16900 3950
rect 16950 3935 17050 3950
rect 17100 3935 17200 3950
rect 17250 3935 17350 3950
rect 17400 3935 17500 3950
rect 17550 3935 17650 3950
rect 17700 3935 17800 3950
rect 17850 3935 17950 3950
rect 18000 3935 18100 3950
rect 18150 3935 18250 3950
rect 18300 3935 18400 3950
rect 18450 3935 18550 3950
rect 18600 3935 18700 3950
rect 18750 3935 18850 3950
rect 18900 3935 19000 3950
rect 19050 3935 19150 3950
rect 19200 3935 19300 3950
rect 19350 3935 19450 3950
rect 19500 3935 19600 3950
rect 19650 3935 19750 3950
rect 19800 3935 19900 3950
rect 19950 3935 20050 3950
rect 20100 3935 20200 3950
rect 20250 3935 20350 3950
rect -600 3800 -500 3815
rect -450 3800 -350 3815
rect -300 3800 -200 3815
rect -150 3800 -50 3815
rect 0 3800 100 3815
rect 150 3800 250 3815
rect 300 3800 400 3815
rect 450 3800 550 3815
rect 600 3800 700 3815
rect 750 3800 850 3815
rect 900 3800 1000 3815
rect 1050 3800 1150 3815
rect 1200 3800 1300 3815
rect 1350 3800 1450 3815
rect 1500 3800 1600 3815
rect 1650 3800 1750 3815
rect 1800 3800 1900 3815
rect 1950 3800 2050 3815
rect 2100 3800 2200 3815
rect 2250 3800 2350 3815
rect 2400 3800 2500 3815
rect 2550 3800 2650 3815
rect 2700 3800 2800 3815
rect 2850 3800 2950 3815
rect 3000 3800 3100 3815
rect 3150 3800 3250 3815
rect 3300 3800 3400 3815
rect 3450 3800 3550 3815
rect 3600 3800 3700 3815
rect 3750 3800 3850 3815
rect 3900 3800 4000 3815
rect 4050 3800 4150 3815
rect 4200 3800 4300 3815
rect 4350 3800 4450 3815
rect 4500 3800 4600 3815
rect 4650 3800 4750 3815
rect 4800 3800 4900 3815
rect 4950 3800 5050 3815
rect 5100 3800 5200 3815
rect 5250 3800 5350 3815
rect 5400 3800 5500 3815
rect 5550 3800 5650 3815
rect 5700 3800 5800 3815
rect 5850 3800 5950 3815
rect 6000 3800 6100 3815
rect 6150 3800 6250 3815
rect 6300 3800 6400 3815
rect 6450 3800 6550 3815
rect 6600 3800 6700 3815
rect 6750 3800 6850 3815
rect 6900 3800 7000 3815
rect 7050 3800 7150 3815
rect 7200 3800 7300 3815
rect 7350 3800 7450 3815
rect 7500 3800 7600 3815
rect 7650 3800 7750 3815
rect 7800 3800 7900 3815
rect 7950 3800 8050 3815
rect 8100 3800 8200 3815
rect 8250 3800 8350 3815
rect 8400 3800 8500 3815
rect 8550 3800 8650 3815
rect 8700 3800 8800 3815
rect 8850 3800 8950 3815
rect 9000 3800 9100 3815
rect 9150 3800 9250 3815
rect 9300 3800 9400 3815
rect 9450 3800 9550 3815
rect 9600 3800 9700 3815
rect 9750 3800 9850 3815
rect 9900 3800 10000 3815
rect 10050 3800 10150 3815
rect 10200 3800 10300 3815
rect 10350 3800 10450 3815
rect 10500 3800 10600 3815
rect 10650 3800 10750 3815
rect 10800 3800 10900 3815
rect 10950 3800 11050 3815
rect 11100 3800 11200 3815
rect 11250 3800 11350 3815
rect 11400 3800 11500 3815
rect 11550 3800 11650 3815
rect 11700 3800 11800 3815
rect 11850 3800 11950 3815
rect 12000 3800 12100 3815
rect 12150 3800 12250 3815
rect 12300 3800 12400 3815
rect 12450 3800 12550 3815
rect 12600 3800 12700 3815
rect 12750 3800 12850 3815
rect 12900 3800 13000 3815
rect 13050 3800 13150 3815
rect 13200 3800 13300 3815
rect 13350 3800 13450 3815
rect 13500 3800 13600 3815
rect 13650 3800 13750 3815
rect 13800 3800 13900 3815
rect 13950 3800 14050 3815
rect 14100 3800 14200 3815
rect 14250 3800 14350 3815
rect 14400 3800 14500 3815
rect 14550 3800 14650 3815
rect 14700 3800 14800 3815
rect 14850 3800 14950 3815
rect 15000 3800 15100 3815
rect 15150 3800 15250 3815
rect 15300 3800 15400 3815
rect 15450 3800 15550 3815
rect 15600 3800 15700 3815
rect 15750 3800 15850 3815
rect 15900 3800 16000 3815
rect 16050 3800 16150 3815
rect 16200 3800 16300 3815
rect 16350 3800 16450 3815
rect 16500 3800 16600 3815
rect 16650 3800 16750 3815
rect 16800 3800 16900 3815
rect 16950 3800 17050 3815
rect 17100 3800 17200 3815
rect 17250 3800 17350 3815
rect 17400 3800 17500 3815
rect 17550 3800 17650 3815
rect 17700 3800 17800 3815
rect 17850 3800 17950 3815
rect 18000 3800 18100 3815
rect 18150 3800 18250 3815
rect 18300 3800 18400 3815
rect 18450 3800 18550 3815
rect 18600 3800 18700 3815
rect 18750 3800 18850 3815
rect 18900 3800 19000 3815
rect 19050 3800 19150 3815
rect 19200 3800 19300 3815
rect 19350 3800 19450 3815
rect 19500 3800 19600 3815
rect 19650 3800 19750 3815
rect 19800 3800 19900 3815
rect 19950 3800 20050 3815
rect 20100 3800 20200 3815
rect 20250 3800 20350 3815
rect -600 3250 -500 3300
rect -450 3250 -350 3300
rect -600 3235 -350 3250
rect -600 3215 -585 3235
rect -565 3215 -535 3235
rect -515 3215 -485 3235
rect -465 3215 -435 3235
rect -415 3215 -385 3235
rect -365 3215 -350 3235
rect -600 3200 -350 3215
rect -600 3150 -500 3200
rect -450 3150 -350 3200
rect -300 3250 -200 3300
rect -150 3250 -50 3300
rect -300 3235 -50 3250
rect -300 3215 -285 3235
rect -265 3215 -235 3235
rect -215 3215 -185 3235
rect -165 3215 -135 3235
rect -115 3215 -85 3235
rect -65 3215 -50 3235
rect -300 3200 -50 3215
rect -300 3150 -200 3200
rect -150 3150 -50 3200
rect 0 3250 100 3300
rect 150 3250 250 3300
rect 0 3235 250 3250
rect 0 3215 15 3235
rect 35 3215 65 3235
rect 85 3215 115 3235
rect 135 3215 165 3235
rect 185 3215 215 3235
rect 235 3215 250 3235
rect 0 3200 250 3215
rect 0 3150 100 3200
rect 150 3150 250 3200
rect 300 3250 400 3300
rect 450 3250 550 3300
rect 300 3235 550 3250
rect 300 3215 315 3235
rect 335 3215 365 3235
rect 385 3215 415 3235
rect 435 3215 465 3235
rect 485 3215 515 3235
rect 535 3215 550 3235
rect 300 3200 550 3215
rect 300 3150 400 3200
rect 450 3150 550 3200
rect 600 3250 700 3300
rect 750 3250 850 3300
rect 600 3235 850 3250
rect 600 3215 615 3235
rect 635 3215 665 3235
rect 685 3215 715 3235
rect 735 3215 765 3235
rect 785 3215 815 3235
rect 835 3215 850 3235
rect 600 3200 850 3215
rect 600 3150 700 3200
rect 750 3150 850 3200
rect 900 3250 1000 3300
rect 1050 3250 1150 3300
rect 900 3235 1150 3250
rect 900 3215 915 3235
rect 935 3215 965 3235
rect 985 3215 1015 3235
rect 1035 3215 1065 3235
rect 1085 3215 1115 3235
rect 1135 3215 1150 3235
rect 900 3200 1150 3215
rect 900 3150 1000 3200
rect 1050 3150 1150 3200
rect 1200 3250 1300 3300
rect 1350 3250 1450 3300
rect 1200 3235 1450 3250
rect 1200 3215 1215 3235
rect 1235 3215 1265 3235
rect 1285 3215 1315 3235
rect 1335 3215 1365 3235
rect 1385 3215 1415 3235
rect 1435 3215 1450 3235
rect 1200 3200 1450 3215
rect 1200 3150 1300 3200
rect 1350 3150 1450 3200
rect 1500 3250 1600 3300
rect 1650 3250 1750 3300
rect 1500 3235 1750 3250
rect 1500 3215 1515 3235
rect 1535 3215 1565 3235
rect 1585 3215 1615 3235
rect 1635 3215 1665 3235
rect 1685 3215 1715 3235
rect 1735 3215 1750 3235
rect 1500 3200 1750 3215
rect 1500 3150 1600 3200
rect 1650 3150 1750 3200
rect 1800 3250 1900 3300
rect 1950 3250 2050 3300
rect 1800 3235 2050 3250
rect 1800 3215 1815 3235
rect 1835 3215 1865 3235
rect 1885 3215 1915 3235
rect 1935 3215 1965 3235
rect 1985 3215 2015 3235
rect 2035 3215 2050 3235
rect 1800 3200 2050 3215
rect 1800 3150 1900 3200
rect 1950 3150 2050 3200
rect 2100 3250 2200 3300
rect 2250 3250 2350 3300
rect 2100 3235 2350 3250
rect 2100 3215 2115 3235
rect 2135 3215 2165 3235
rect 2185 3215 2215 3235
rect 2235 3215 2265 3235
rect 2285 3215 2315 3235
rect 2335 3215 2350 3235
rect 2100 3200 2350 3215
rect 2100 3150 2200 3200
rect 2250 3150 2350 3200
rect 2400 3250 2500 3300
rect 2550 3250 2650 3300
rect 2400 3235 2650 3250
rect 2400 3215 2415 3235
rect 2435 3215 2465 3235
rect 2485 3215 2515 3235
rect 2535 3215 2565 3235
rect 2585 3215 2615 3235
rect 2635 3215 2650 3235
rect 2400 3200 2650 3215
rect 2400 3150 2500 3200
rect 2550 3150 2650 3200
rect 2700 3250 2800 3300
rect 2850 3250 2950 3300
rect 2700 3235 2950 3250
rect 2700 3215 2715 3235
rect 2735 3215 2765 3235
rect 2785 3215 2815 3235
rect 2835 3215 2865 3235
rect 2885 3215 2915 3235
rect 2935 3215 2950 3235
rect 2700 3200 2950 3215
rect 2700 3150 2800 3200
rect 2850 3150 2950 3200
rect 3000 3250 3100 3300
rect 3150 3250 3250 3300
rect 3000 3235 3250 3250
rect 3000 3215 3015 3235
rect 3035 3215 3065 3235
rect 3085 3215 3115 3235
rect 3135 3215 3165 3235
rect 3185 3215 3215 3235
rect 3235 3215 3250 3235
rect 3000 3200 3250 3215
rect 3000 3150 3100 3200
rect 3150 3150 3250 3200
rect 3300 3250 3400 3300
rect 3450 3250 3550 3300
rect 3300 3235 3550 3250
rect 3300 3215 3315 3235
rect 3335 3215 3365 3235
rect 3385 3215 3415 3235
rect 3435 3215 3465 3235
rect 3485 3215 3515 3235
rect 3535 3215 3550 3235
rect 3300 3200 3550 3215
rect 3300 3150 3400 3200
rect 3450 3150 3550 3200
rect 3600 3250 3700 3300
rect 3750 3250 3850 3300
rect 3600 3235 3850 3250
rect 3600 3215 3615 3235
rect 3635 3215 3665 3235
rect 3685 3215 3715 3235
rect 3735 3215 3765 3235
rect 3785 3215 3815 3235
rect 3835 3215 3850 3235
rect 3600 3200 3850 3215
rect 3600 3150 3700 3200
rect 3750 3150 3850 3200
rect 3900 3250 4000 3300
rect 4050 3250 4150 3300
rect 3900 3235 4150 3250
rect 3900 3215 3915 3235
rect 3935 3215 3965 3235
rect 3985 3215 4015 3235
rect 4035 3215 4065 3235
rect 4085 3215 4115 3235
rect 4135 3215 4150 3235
rect 3900 3200 4150 3215
rect 3900 3150 4000 3200
rect 4050 3150 4150 3200
rect 4200 3250 4300 3300
rect 4350 3250 4450 3300
rect 4200 3235 4450 3250
rect 4200 3215 4215 3235
rect 4235 3215 4265 3235
rect 4285 3215 4315 3235
rect 4335 3215 4365 3235
rect 4385 3215 4415 3235
rect 4435 3215 4450 3235
rect 4200 3200 4450 3215
rect 4200 3150 4300 3200
rect 4350 3150 4450 3200
rect 4500 3250 4600 3300
rect 4650 3250 4750 3300
rect 4500 3235 4750 3250
rect 4500 3215 4515 3235
rect 4535 3215 4565 3235
rect 4585 3215 4615 3235
rect 4635 3215 4665 3235
rect 4685 3215 4715 3235
rect 4735 3215 4750 3235
rect 4500 3200 4750 3215
rect 4500 3150 4600 3200
rect 4650 3150 4750 3200
rect 4800 3250 4900 3300
rect 4950 3250 5050 3300
rect 4800 3235 5050 3250
rect 4800 3215 4815 3235
rect 4835 3215 4865 3235
rect 4885 3215 4915 3235
rect 4935 3215 4965 3235
rect 4985 3215 5015 3235
rect 5035 3215 5050 3235
rect 4800 3200 5050 3215
rect 4800 3150 4900 3200
rect 4950 3150 5050 3200
rect 5100 3250 5200 3300
rect 5250 3250 5350 3300
rect 5100 3235 5350 3250
rect 5100 3215 5115 3235
rect 5135 3215 5165 3235
rect 5185 3215 5215 3235
rect 5235 3215 5265 3235
rect 5285 3215 5315 3235
rect 5335 3215 5350 3235
rect 5100 3200 5350 3215
rect 5100 3150 5200 3200
rect 5250 3150 5350 3200
rect 5400 3250 5500 3300
rect 5550 3250 5650 3300
rect 5400 3235 5650 3250
rect 5400 3215 5415 3235
rect 5435 3215 5465 3235
rect 5485 3215 5515 3235
rect 5535 3215 5565 3235
rect 5585 3215 5615 3235
rect 5635 3215 5650 3235
rect 5400 3200 5650 3215
rect 5400 3150 5500 3200
rect 5550 3150 5650 3200
rect 5700 3250 5800 3300
rect 5850 3250 5950 3300
rect 5700 3235 5950 3250
rect 5700 3215 5715 3235
rect 5735 3215 5765 3235
rect 5785 3215 5815 3235
rect 5835 3215 5865 3235
rect 5885 3215 5915 3235
rect 5935 3215 5950 3235
rect 5700 3200 5950 3215
rect 5700 3150 5800 3200
rect 5850 3150 5950 3200
rect 6000 3250 6100 3300
rect 6150 3250 6250 3300
rect 6000 3235 6250 3250
rect 6000 3215 6015 3235
rect 6035 3215 6065 3235
rect 6085 3215 6115 3235
rect 6135 3215 6165 3235
rect 6185 3215 6215 3235
rect 6235 3215 6250 3235
rect 6000 3200 6250 3215
rect 6000 3150 6100 3200
rect 6150 3150 6250 3200
rect 6300 3250 6400 3300
rect 6450 3250 6550 3300
rect 6300 3235 6550 3250
rect 6300 3215 6315 3235
rect 6335 3215 6365 3235
rect 6385 3215 6415 3235
rect 6435 3215 6465 3235
rect 6485 3215 6515 3235
rect 6535 3215 6550 3235
rect 6300 3200 6550 3215
rect 6300 3150 6400 3200
rect 6450 3150 6550 3200
rect 6600 3250 6700 3300
rect 6750 3250 6850 3300
rect 6600 3235 6850 3250
rect 6600 3215 6615 3235
rect 6635 3215 6665 3235
rect 6685 3215 6715 3235
rect 6735 3215 6765 3235
rect 6785 3215 6815 3235
rect 6835 3215 6850 3235
rect 6600 3200 6850 3215
rect 6600 3150 6700 3200
rect 6750 3150 6850 3200
rect 6900 3250 7000 3300
rect 7050 3250 7150 3300
rect 6900 3235 7150 3250
rect 6900 3215 6915 3235
rect 6935 3215 6965 3235
rect 6985 3215 7015 3235
rect 7035 3215 7065 3235
rect 7085 3215 7115 3235
rect 7135 3215 7150 3235
rect 6900 3200 7150 3215
rect 6900 3150 7000 3200
rect 7050 3150 7150 3200
rect 7200 3250 7300 3300
rect 7350 3250 7450 3300
rect 7200 3235 7450 3250
rect 7200 3215 7215 3235
rect 7235 3215 7265 3235
rect 7285 3215 7315 3235
rect 7335 3215 7365 3235
rect 7385 3215 7415 3235
rect 7435 3215 7450 3235
rect 7200 3200 7450 3215
rect 7200 3150 7300 3200
rect 7350 3150 7450 3200
rect 7500 3250 7600 3300
rect 7650 3250 7750 3300
rect 7500 3235 7750 3250
rect 7500 3215 7515 3235
rect 7535 3215 7565 3235
rect 7585 3215 7615 3235
rect 7635 3215 7665 3235
rect 7685 3215 7715 3235
rect 7735 3215 7750 3235
rect 7500 3200 7750 3215
rect 7500 3150 7600 3200
rect 7650 3150 7750 3200
rect 7800 3250 7900 3300
rect 7950 3250 8050 3300
rect 7800 3235 8050 3250
rect 7800 3215 7815 3235
rect 7835 3215 7865 3235
rect 7885 3215 7915 3235
rect 7935 3215 7965 3235
rect 7985 3215 8015 3235
rect 8035 3215 8050 3235
rect 7800 3200 8050 3215
rect 7800 3150 7900 3200
rect 7950 3150 8050 3200
rect 8100 3250 8200 3300
rect 8250 3250 8350 3300
rect 8100 3235 8350 3250
rect 8100 3215 8115 3235
rect 8135 3215 8165 3235
rect 8185 3215 8215 3235
rect 8235 3215 8265 3235
rect 8285 3215 8315 3235
rect 8335 3215 8350 3235
rect 8100 3200 8350 3215
rect 8100 3150 8200 3200
rect 8250 3150 8350 3200
rect 8400 3250 8500 3300
rect 8550 3250 8650 3300
rect 8400 3235 8650 3250
rect 8400 3215 8415 3235
rect 8435 3215 8465 3235
rect 8485 3215 8515 3235
rect 8535 3215 8565 3235
rect 8585 3215 8615 3235
rect 8635 3215 8650 3235
rect 8400 3200 8650 3215
rect 8400 3150 8500 3200
rect 8550 3150 8650 3200
rect 8700 3250 8800 3300
rect 8850 3250 8950 3300
rect 8700 3235 8950 3250
rect 8700 3215 8715 3235
rect 8735 3215 8765 3235
rect 8785 3215 8815 3235
rect 8835 3215 8865 3235
rect 8885 3215 8915 3235
rect 8935 3215 8950 3235
rect 8700 3200 8950 3215
rect 8700 3150 8800 3200
rect 8850 3150 8950 3200
rect 9000 3250 9100 3300
rect 9150 3250 9250 3300
rect 9000 3235 9250 3250
rect 9000 3215 9015 3235
rect 9035 3215 9065 3235
rect 9085 3215 9115 3235
rect 9135 3215 9165 3235
rect 9185 3215 9215 3235
rect 9235 3215 9250 3235
rect 9000 3200 9250 3215
rect 9000 3150 9100 3200
rect 9150 3150 9250 3200
rect 9300 3250 9400 3300
rect 9450 3250 9550 3300
rect 9300 3235 9550 3250
rect 9300 3215 9315 3235
rect 9335 3215 9365 3235
rect 9385 3215 9415 3235
rect 9435 3215 9465 3235
rect 9485 3215 9515 3235
rect 9535 3215 9550 3235
rect 9300 3200 9550 3215
rect 9300 3150 9400 3200
rect 9450 3150 9550 3200
rect 9600 3250 9700 3300
rect 9750 3250 9850 3300
rect 9600 3235 9850 3250
rect 9600 3215 9615 3235
rect 9635 3215 9665 3235
rect 9685 3215 9715 3235
rect 9735 3215 9765 3235
rect 9785 3215 9815 3235
rect 9835 3215 9850 3235
rect 9600 3200 9850 3215
rect 9600 3150 9700 3200
rect 9750 3150 9850 3200
rect 9900 3250 10000 3300
rect 10050 3250 10150 3300
rect 9900 3235 10150 3250
rect 9900 3215 9915 3235
rect 9935 3215 9965 3235
rect 9985 3215 10015 3235
rect 10035 3215 10065 3235
rect 10085 3215 10115 3235
rect 10135 3215 10150 3235
rect 9900 3200 10150 3215
rect 9900 3150 10000 3200
rect 10050 3150 10150 3200
rect 10200 3250 10300 3300
rect 10350 3250 10450 3300
rect 10200 3235 10450 3250
rect 10200 3215 10215 3235
rect 10235 3215 10265 3235
rect 10285 3215 10315 3235
rect 10335 3215 10365 3235
rect 10385 3215 10415 3235
rect 10435 3215 10450 3235
rect 10200 3200 10450 3215
rect 10200 3150 10300 3200
rect 10350 3150 10450 3200
rect 10500 3250 10600 3300
rect 10650 3250 10750 3300
rect 10500 3235 10750 3250
rect 10500 3215 10515 3235
rect 10535 3215 10565 3235
rect 10585 3215 10615 3235
rect 10635 3215 10665 3235
rect 10685 3215 10715 3235
rect 10735 3215 10750 3235
rect 10500 3200 10750 3215
rect 10500 3150 10600 3200
rect 10650 3150 10750 3200
rect 10800 3250 10900 3300
rect 10950 3250 11050 3300
rect 10800 3235 11050 3250
rect 10800 3215 10815 3235
rect 10835 3215 10865 3235
rect 10885 3215 10915 3235
rect 10935 3215 10965 3235
rect 10985 3215 11015 3235
rect 11035 3215 11050 3235
rect 10800 3200 11050 3215
rect 10800 3150 10900 3200
rect 10950 3150 11050 3200
rect 11100 3250 11200 3300
rect 11250 3250 11350 3300
rect 11100 3235 11350 3250
rect 11100 3215 11115 3235
rect 11135 3215 11165 3235
rect 11185 3215 11215 3235
rect 11235 3215 11265 3235
rect 11285 3215 11315 3235
rect 11335 3215 11350 3235
rect 11100 3200 11350 3215
rect 11100 3150 11200 3200
rect 11250 3150 11350 3200
rect 11400 3250 11500 3300
rect 11550 3250 11650 3300
rect 11400 3235 11650 3250
rect 11400 3215 11415 3235
rect 11435 3215 11465 3235
rect 11485 3215 11515 3235
rect 11535 3215 11565 3235
rect 11585 3215 11615 3235
rect 11635 3215 11650 3235
rect 11400 3200 11650 3215
rect 11400 3150 11500 3200
rect 11550 3150 11650 3200
rect 11700 3250 11800 3300
rect 11850 3250 11950 3300
rect 11700 3235 11950 3250
rect 11700 3215 11715 3235
rect 11735 3215 11765 3235
rect 11785 3215 11815 3235
rect 11835 3215 11865 3235
rect 11885 3215 11915 3235
rect 11935 3215 11950 3235
rect 11700 3200 11950 3215
rect 11700 3150 11800 3200
rect 11850 3150 11950 3200
rect 12000 3250 12100 3300
rect 12150 3250 12250 3300
rect 12000 3235 12250 3250
rect 12000 3215 12015 3235
rect 12035 3215 12065 3235
rect 12085 3215 12115 3235
rect 12135 3215 12165 3235
rect 12185 3215 12215 3235
rect 12235 3215 12250 3235
rect 12000 3200 12250 3215
rect 12000 3150 12100 3200
rect 12150 3150 12250 3200
rect 12300 3250 12400 3300
rect 12450 3250 12550 3300
rect 12300 3235 12550 3250
rect 12300 3215 12315 3235
rect 12335 3215 12365 3235
rect 12385 3215 12415 3235
rect 12435 3215 12465 3235
rect 12485 3215 12515 3235
rect 12535 3215 12550 3235
rect 12300 3200 12550 3215
rect 12300 3150 12400 3200
rect 12450 3150 12550 3200
rect 12600 3250 12700 3300
rect 12750 3250 12850 3300
rect 12600 3235 12850 3250
rect 12600 3215 12615 3235
rect 12635 3215 12665 3235
rect 12685 3215 12715 3235
rect 12735 3215 12765 3235
rect 12785 3215 12815 3235
rect 12835 3215 12850 3235
rect 12600 3200 12850 3215
rect 12600 3150 12700 3200
rect 12750 3150 12850 3200
rect 12900 3250 13000 3300
rect 13050 3250 13150 3300
rect 12900 3235 13150 3250
rect 12900 3215 12915 3235
rect 12935 3215 12965 3235
rect 12985 3215 13015 3235
rect 13035 3215 13065 3235
rect 13085 3215 13115 3235
rect 13135 3215 13150 3235
rect 12900 3200 13150 3215
rect 12900 3150 13000 3200
rect 13050 3150 13150 3200
rect 13200 3250 13300 3300
rect 13350 3250 13450 3300
rect 13200 3235 13450 3250
rect 13200 3215 13215 3235
rect 13235 3215 13265 3235
rect 13285 3215 13315 3235
rect 13335 3215 13365 3235
rect 13385 3215 13415 3235
rect 13435 3215 13450 3235
rect 13200 3200 13450 3215
rect 13200 3150 13300 3200
rect 13350 3150 13450 3200
rect 13500 3250 13600 3300
rect 13650 3250 13750 3300
rect 13500 3235 13750 3250
rect 13500 3215 13515 3235
rect 13535 3215 13565 3235
rect 13585 3215 13615 3235
rect 13635 3215 13665 3235
rect 13685 3215 13715 3235
rect 13735 3215 13750 3235
rect 13500 3200 13750 3215
rect 13500 3150 13600 3200
rect 13650 3150 13750 3200
rect 13800 3250 13900 3300
rect 13950 3250 14050 3300
rect 13800 3235 14050 3250
rect 13800 3215 13815 3235
rect 13835 3215 13865 3235
rect 13885 3215 13915 3235
rect 13935 3215 13965 3235
rect 13985 3215 14015 3235
rect 14035 3215 14050 3235
rect 13800 3200 14050 3215
rect 13800 3150 13900 3200
rect 13950 3150 14050 3200
rect 14100 3250 14200 3300
rect 14250 3250 14350 3300
rect 14100 3235 14350 3250
rect 14100 3215 14115 3235
rect 14135 3215 14165 3235
rect 14185 3215 14215 3235
rect 14235 3215 14265 3235
rect 14285 3215 14315 3235
rect 14335 3215 14350 3235
rect 14100 3200 14350 3215
rect 14100 3150 14200 3200
rect 14250 3150 14350 3200
rect 14400 3250 14500 3300
rect 14550 3250 14650 3300
rect 14400 3235 14650 3250
rect 14400 3215 14415 3235
rect 14435 3215 14465 3235
rect 14485 3215 14515 3235
rect 14535 3215 14565 3235
rect 14585 3215 14615 3235
rect 14635 3215 14650 3235
rect 14400 3200 14650 3215
rect 14400 3150 14500 3200
rect 14550 3150 14650 3200
rect 14700 3250 14800 3300
rect 14850 3250 14950 3300
rect 14700 3235 14950 3250
rect 14700 3215 14715 3235
rect 14735 3215 14765 3235
rect 14785 3215 14815 3235
rect 14835 3215 14865 3235
rect 14885 3215 14915 3235
rect 14935 3215 14950 3235
rect 14700 3200 14950 3215
rect 14700 3150 14800 3200
rect 14850 3150 14950 3200
rect 15000 3250 15100 3300
rect 15150 3250 15250 3300
rect 15000 3235 15250 3250
rect 15000 3215 15015 3235
rect 15035 3215 15065 3235
rect 15085 3215 15115 3235
rect 15135 3215 15165 3235
rect 15185 3215 15215 3235
rect 15235 3215 15250 3235
rect 15000 3200 15250 3215
rect 15000 3150 15100 3200
rect 15150 3150 15250 3200
rect 15300 3250 15400 3300
rect 15450 3250 15550 3300
rect 15300 3235 15550 3250
rect 15300 3215 15315 3235
rect 15335 3215 15365 3235
rect 15385 3215 15415 3235
rect 15435 3215 15465 3235
rect 15485 3215 15515 3235
rect 15535 3215 15550 3235
rect 15300 3200 15550 3215
rect 15300 3150 15400 3200
rect 15450 3150 15550 3200
rect 15600 3250 15700 3300
rect 15750 3250 15850 3300
rect 15600 3235 15850 3250
rect 15600 3215 15615 3235
rect 15635 3215 15665 3235
rect 15685 3215 15715 3235
rect 15735 3215 15765 3235
rect 15785 3215 15815 3235
rect 15835 3215 15850 3235
rect 15600 3200 15850 3215
rect 15600 3150 15700 3200
rect 15750 3150 15850 3200
rect 15900 3250 16000 3300
rect 16050 3250 16150 3300
rect 15900 3235 16150 3250
rect 15900 3215 15915 3235
rect 15935 3215 15965 3235
rect 15985 3215 16015 3235
rect 16035 3215 16065 3235
rect 16085 3215 16115 3235
rect 16135 3215 16150 3235
rect 15900 3200 16150 3215
rect 15900 3150 16000 3200
rect 16050 3150 16150 3200
rect 16200 3250 16300 3300
rect 16350 3250 16450 3300
rect 16200 3235 16450 3250
rect 16200 3215 16215 3235
rect 16235 3215 16265 3235
rect 16285 3215 16315 3235
rect 16335 3215 16365 3235
rect 16385 3215 16415 3235
rect 16435 3215 16450 3235
rect 16200 3200 16450 3215
rect 16200 3150 16300 3200
rect 16350 3150 16450 3200
rect 16500 3250 16600 3300
rect 16650 3250 16750 3300
rect 16500 3235 16750 3250
rect 16500 3215 16515 3235
rect 16535 3215 16565 3235
rect 16585 3215 16615 3235
rect 16635 3215 16665 3235
rect 16685 3215 16715 3235
rect 16735 3215 16750 3235
rect 16500 3200 16750 3215
rect 16500 3150 16600 3200
rect 16650 3150 16750 3200
rect 16800 3250 16900 3300
rect 16950 3250 17050 3300
rect 16800 3235 17050 3250
rect 16800 3215 16815 3235
rect 16835 3215 16865 3235
rect 16885 3215 16915 3235
rect 16935 3215 16965 3235
rect 16985 3215 17015 3235
rect 17035 3215 17050 3235
rect 16800 3200 17050 3215
rect 16800 3150 16900 3200
rect 16950 3150 17050 3200
rect 17100 3250 17200 3300
rect 17250 3250 17350 3300
rect 17100 3235 17350 3250
rect 17100 3215 17115 3235
rect 17135 3215 17165 3235
rect 17185 3215 17215 3235
rect 17235 3215 17265 3235
rect 17285 3215 17315 3235
rect 17335 3215 17350 3235
rect 17100 3200 17350 3215
rect 17100 3150 17200 3200
rect 17250 3150 17350 3200
rect 17400 3250 17500 3300
rect 17550 3250 17650 3300
rect 17400 3235 17650 3250
rect 17400 3215 17415 3235
rect 17435 3215 17465 3235
rect 17485 3215 17515 3235
rect 17535 3215 17565 3235
rect 17585 3215 17615 3235
rect 17635 3215 17650 3235
rect 17400 3200 17650 3215
rect 17400 3150 17500 3200
rect 17550 3150 17650 3200
rect 17700 3250 17800 3300
rect 17850 3250 17950 3300
rect 17700 3235 17950 3250
rect 17700 3215 17715 3235
rect 17735 3215 17765 3235
rect 17785 3215 17815 3235
rect 17835 3215 17865 3235
rect 17885 3215 17915 3235
rect 17935 3215 17950 3235
rect 17700 3200 17950 3215
rect 17700 3150 17800 3200
rect 17850 3150 17950 3200
rect 18000 3250 18100 3300
rect 18150 3250 18250 3300
rect 18000 3235 18250 3250
rect 18000 3215 18015 3235
rect 18035 3215 18065 3235
rect 18085 3215 18115 3235
rect 18135 3215 18165 3235
rect 18185 3215 18215 3235
rect 18235 3215 18250 3235
rect 18000 3200 18250 3215
rect 18000 3150 18100 3200
rect 18150 3150 18250 3200
rect 18300 3250 18400 3300
rect 18450 3250 18550 3300
rect 18300 3235 18550 3250
rect 18300 3215 18315 3235
rect 18335 3215 18365 3235
rect 18385 3215 18415 3235
rect 18435 3215 18465 3235
rect 18485 3215 18515 3235
rect 18535 3215 18550 3235
rect 18300 3200 18550 3215
rect 18300 3150 18400 3200
rect 18450 3150 18550 3200
rect 18600 3250 18700 3300
rect 18750 3250 18850 3300
rect 18600 3235 18850 3250
rect 18600 3215 18615 3235
rect 18635 3215 18665 3235
rect 18685 3215 18715 3235
rect 18735 3215 18765 3235
rect 18785 3215 18815 3235
rect 18835 3215 18850 3235
rect 18600 3200 18850 3215
rect 18600 3150 18700 3200
rect 18750 3150 18850 3200
rect 18900 3250 19000 3300
rect 19050 3250 19150 3300
rect 18900 3235 19150 3250
rect 18900 3215 18915 3235
rect 18935 3215 18965 3235
rect 18985 3215 19015 3235
rect 19035 3215 19065 3235
rect 19085 3215 19115 3235
rect 19135 3215 19150 3235
rect 18900 3200 19150 3215
rect 18900 3150 19000 3200
rect 19050 3150 19150 3200
rect 19200 3250 19300 3300
rect 19350 3250 19450 3300
rect 19200 3235 19450 3250
rect 19200 3215 19215 3235
rect 19235 3215 19265 3235
rect 19285 3215 19315 3235
rect 19335 3215 19365 3235
rect 19385 3215 19415 3235
rect 19435 3215 19450 3235
rect 19200 3200 19450 3215
rect 19200 3150 19300 3200
rect 19350 3150 19450 3200
rect 19500 3250 19600 3300
rect 19650 3250 19750 3300
rect 19500 3235 19750 3250
rect 19500 3215 19515 3235
rect 19535 3215 19565 3235
rect 19585 3215 19615 3235
rect 19635 3215 19665 3235
rect 19685 3215 19715 3235
rect 19735 3215 19750 3235
rect 19500 3200 19750 3215
rect 19500 3150 19600 3200
rect 19650 3150 19750 3200
rect 19800 3250 19900 3300
rect 19950 3250 20050 3300
rect 19800 3235 20050 3250
rect 19800 3215 19815 3235
rect 19835 3215 19865 3235
rect 19885 3215 19915 3235
rect 19935 3215 19965 3235
rect 19985 3215 20015 3235
rect 20035 3215 20050 3235
rect 19800 3200 20050 3215
rect 19800 3150 19900 3200
rect 19950 3150 20050 3200
rect 20100 3250 20200 3300
rect 20250 3250 20350 3300
rect 20100 3235 20350 3250
rect 20100 3215 20115 3235
rect 20135 3215 20165 3235
rect 20185 3215 20215 3235
rect 20235 3215 20265 3235
rect 20285 3215 20315 3235
rect 20335 3215 20350 3235
rect 20100 3200 20350 3215
rect 20100 3150 20200 3200
rect 20250 3150 20350 3200
rect -600 2635 -500 2650
rect -450 2635 -350 2650
rect -300 2635 -200 2650
rect -150 2635 -50 2650
rect 0 2635 100 2650
rect 150 2635 250 2650
rect 300 2635 400 2650
rect 450 2635 550 2650
rect 600 2635 700 2650
rect 750 2635 850 2650
rect 900 2635 1000 2650
rect 1050 2635 1150 2650
rect 1200 2635 1300 2650
rect 1350 2635 1450 2650
rect 1500 2635 1600 2650
rect 1650 2635 1750 2650
rect 1800 2635 1900 2650
rect 1950 2635 2050 2650
rect 2100 2635 2200 2650
rect 2250 2635 2350 2650
rect 2400 2635 2500 2650
rect 2550 2635 2650 2650
rect 2700 2635 2800 2650
rect 2850 2635 2950 2650
rect 3000 2635 3100 2650
rect 3150 2635 3250 2650
rect 3300 2635 3400 2650
rect 3450 2635 3550 2650
rect 3600 2635 3700 2650
rect 3750 2635 3850 2650
rect 3900 2635 4000 2650
rect 4050 2635 4150 2650
rect 4200 2635 4300 2650
rect 4350 2635 4450 2650
rect 4500 2635 4600 2650
rect 4650 2635 4750 2650
rect 4800 2635 4900 2650
rect 4950 2635 5050 2650
rect 5100 2635 5200 2650
rect 5250 2635 5350 2650
rect 5400 2635 5500 2650
rect 5550 2635 5650 2650
rect 5700 2635 5800 2650
rect 5850 2635 5950 2650
rect 6000 2635 6100 2650
rect 6150 2635 6250 2650
rect 6300 2635 6400 2650
rect 6450 2635 6550 2650
rect 6600 2635 6700 2650
rect 6750 2635 6850 2650
rect 6900 2635 7000 2650
rect 7050 2635 7150 2650
rect 7200 2635 7300 2650
rect 7350 2635 7450 2650
rect 7500 2635 7600 2650
rect 7650 2635 7750 2650
rect 7800 2635 7900 2650
rect 7950 2635 8050 2650
rect 8100 2635 8200 2650
rect 8250 2635 8350 2650
rect 8400 2635 8500 2650
rect 8550 2635 8650 2650
rect 8700 2635 8800 2650
rect 8850 2635 8950 2650
rect 9000 2635 9100 2650
rect 9150 2635 9250 2650
rect 9300 2635 9400 2650
rect 9450 2635 9550 2650
rect 9600 2635 9700 2650
rect 9750 2635 9850 2650
rect 9900 2635 10000 2650
rect 10050 2635 10150 2650
rect 10200 2635 10300 2650
rect 10350 2635 10450 2650
rect 10500 2635 10600 2650
rect 10650 2635 10750 2650
rect 10800 2635 10900 2650
rect 10950 2635 11050 2650
rect 11100 2635 11200 2650
rect 11250 2635 11350 2650
rect 11400 2635 11500 2650
rect 11550 2635 11650 2650
rect 11700 2635 11800 2650
rect 11850 2635 11950 2650
rect 12000 2635 12100 2650
rect 12150 2635 12250 2650
rect 12300 2635 12400 2650
rect 12450 2635 12550 2650
rect 12600 2635 12700 2650
rect 12750 2635 12850 2650
rect 12900 2635 13000 2650
rect 13050 2635 13150 2650
rect 13200 2635 13300 2650
rect 13350 2635 13450 2650
rect 13500 2635 13600 2650
rect 13650 2635 13750 2650
rect 13800 2635 13900 2650
rect 13950 2635 14050 2650
rect 14100 2635 14200 2650
rect 14250 2635 14350 2650
rect 14400 2635 14500 2650
rect 14550 2635 14650 2650
rect 14700 2635 14800 2650
rect 14850 2635 14950 2650
rect 15000 2635 15100 2650
rect 15150 2635 15250 2650
rect 15300 2635 15400 2650
rect 15450 2635 15550 2650
rect 15600 2635 15700 2650
rect 15750 2635 15850 2650
rect 15900 2635 16000 2650
rect 16050 2635 16150 2650
rect 16200 2635 16300 2650
rect 16350 2635 16450 2650
rect 16500 2635 16600 2650
rect 16650 2635 16750 2650
rect 16800 2635 16900 2650
rect 16950 2635 17050 2650
rect 17100 2635 17200 2650
rect 17250 2635 17350 2650
rect 17400 2635 17500 2650
rect 17550 2635 17650 2650
rect 17700 2635 17800 2650
rect 17850 2635 17950 2650
rect 18000 2635 18100 2650
rect 18150 2635 18250 2650
rect 18300 2635 18400 2650
rect 18450 2635 18550 2650
rect 18600 2635 18700 2650
rect 18750 2635 18850 2650
rect 18900 2635 19000 2650
rect 19050 2635 19150 2650
rect 19200 2635 19300 2650
rect 19350 2635 19450 2650
rect 19500 2635 19600 2650
rect 19650 2635 19750 2650
rect 19800 2635 19900 2650
rect 19950 2635 20050 2650
rect 20100 2635 20200 2650
rect 20250 2635 20350 2650
rect -600 1600 -500 1615
rect -450 1600 -350 1615
rect -300 1600 -200 1615
rect -150 1600 -50 1615
rect 0 1600 100 1615
rect 150 1600 250 1615
rect 300 1600 400 1615
rect 450 1600 550 1615
rect 600 1600 700 1615
rect 750 1600 850 1615
rect 900 1600 1000 1615
rect 1050 1600 1150 1615
rect 1200 1600 1300 1615
rect 1350 1600 1450 1615
rect 1500 1600 1600 1615
rect 1650 1600 1750 1615
rect 1800 1600 1900 1615
rect 1950 1600 2050 1615
rect 2100 1600 2200 1615
rect 2250 1600 2350 1615
rect 2400 1600 2500 1615
rect 2550 1600 2650 1615
rect 2700 1600 2800 1615
rect 2850 1600 2950 1615
rect 3000 1600 3100 1615
rect 3150 1600 3250 1615
rect 3300 1600 3400 1615
rect 3450 1600 3550 1615
rect 3600 1600 3700 1615
rect 3750 1600 3850 1615
rect 3900 1600 4000 1615
rect 4050 1600 4150 1615
rect 4200 1600 4300 1615
rect 4350 1600 4450 1615
rect 4500 1600 4600 1615
rect 4650 1600 4750 1615
rect 4800 1600 4900 1615
rect 4950 1600 5050 1615
rect 5100 1600 5200 1615
rect 5250 1600 5350 1615
rect 5400 1600 5500 1615
rect 5550 1600 5650 1615
rect 5700 1600 5800 1615
rect 5850 1600 5950 1615
rect 6000 1600 6100 1615
rect 6150 1600 6250 1615
rect 6300 1600 6400 1615
rect 6450 1600 6550 1615
rect 6600 1600 6700 1615
rect 6750 1600 6850 1615
rect 6900 1600 7000 1615
rect 7050 1600 7150 1615
rect 7200 1600 7300 1615
rect 7350 1600 7450 1615
rect 7500 1600 7600 1615
rect 7650 1600 7750 1615
rect 7800 1600 7900 1615
rect 7950 1600 8050 1615
rect 8100 1600 8200 1615
rect 8250 1600 8350 1615
rect 8400 1600 8500 1615
rect 8550 1600 8650 1615
rect 8700 1600 8800 1615
rect 8850 1600 8950 1615
rect 9000 1600 9100 1615
rect 9150 1600 9250 1615
rect 9300 1600 9400 1615
rect 9450 1600 9550 1615
rect 9600 1600 9700 1615
rect 9750 1600 9850 1615
rect 9900 1600 10000 1615
rect 10050 1600 10150 1615
rect 10200 1600 10300 1615
rect 10350 1600 10450 1615
rect 10500 1600 10600 1615
rect 10650 1600 10750 1615
rect 10800 1600 10900 1615
rect 10950 1600 11050 1615
rect 11100 1600 11200 1615
rect 11250 1600 11350 1615
rect 11400 1600 11500 1615
rect 11550 1600 11650 1615
rect 11700 1600 11800 1615
rect 11850 1600 11950 1615
rect 12000 1600 12100 1615
rect 12150 1600 12250 1615
rect 12300 1600 12400 1615
rect 12450 1600 12550 1615
rect 12600 1600 12700 1615
rect 12750 1600 12850 1615
rect 12900 1600 13000 1615
rect 13050 1600 13150 1615
rect 13200 1600 13300 1615
rect 13350 1600 13450 1615
rect 13500 1600 13600 1615
rect 13650 1600 13750 1615
rect 13800 1600 13900 1615
rect 13950 1600 14050 1615
rect 14100 1600 14200 1615
rect 14250 1600 14350 1615
rect 14400 1600 14500 1615
rect 14550 1600 14650 1615
rect 14700 1600 14800 1615
rect 14850 1600 14950 1615
rect 15000 1600 15100 1615
rect 15150 1600 15250 1615
rect 15300 1600 15400 1615
rect 15450 1600 15550 1615
rect 15600 1600 15700 1615
rect 15750 1600 15850 1615
rect 15900 1600 16000 1615
rect 16050 1600 16150 1615
rect 16200 1600 16300 1615
rect 16350 1600 16450 1615
rect 16500 1600 16600 1615
rect 16650 1600 16750 1615
rect 16800 1600 16900 1615
rect 16950 1600 17050 1615
rect 17100 1600 17200 1615
rect 17250 1600 17350 1615
rect 17400 1600 17500 1615
rect 17550 1600 17650 1615
rect 17700 1600 17800 1615
rect 17850 1600 17950 1615
rect 18000 1600 18100 1615
rect 18150 1600 18250 1615
rect 18300 1600 18400 1615
rect 18450 1600 18550 1615
rect 18600 1600 18700 1615
rect 18750 1600 18850 1615
rect 18900 1600 19000 1615
rect 19050 1600 19150 1615
rect 19200 1600 19300 1615
rect 19350 1600 19450 1615
rect 19500 1600 19600 1615
rect 19650 1600 19750 1615
rect 19800 1600 19900 1615
rect 19950 1600 20050 1615
rect 20100 1600 20200 1615
rect 20250 1600 20350 1615
rect -600 850 -500 900
rect -450 850 -350 900
rect -600 835 -350 850
rect -600 815 -585 835
rect -565 815 -535 835
rect -515 815 -485 835
rect -465 815 -435 835
rect -415 815 -385 835
rect -365 815 -350 835
rect -600 800 -350 815
rect -600 750 -500 800
rect -450 750 -350 800
rect -300 850 -200 900
rect -150 850 -50 900
rect -300 835 -50 850
rect -300 815 -285 835
rect -265 815 -235 835
rect -215 815 -185 835
rect -165 815 -135 835
rect -115 815 -85 835
rect -65 815 -50 835
rect -300 800 -50 815
rect -300 750 -200 800
rect -150 750 -50 800
rect 0 850 100 900
rect 150 850 250 900
rect 0 835 250 850
rect 0 815 15 835
rect 35 815 65 835
rect 85 815 115 835
rect 135 815 165 835
rect 185 815 215 835
rect 235 815 250 835
rect 0 800 250 815
rect 0 750 100 800
rect 150 750 250 800
rect 300 850 400 900
rect 450 850 550 900
rect 300 835 550 850
rect 300 815 315 835
rect 335 815 365 835
rect 385 815 415 835
rect 435 815 465 835
rect 485 815 515 835
rect 535 815 550 835
rect 300 800 550 815
rect 300 750 400 800
rect 450 750 550 800
rect 600 850 700 900
rect 750 850 850 900
rect 600 835 850 850
rect 600 815 615 835
rect 635 815 665 835
rect 685 815 715 835
rect 735 815 765 835
rect 785 815 815 835
rect 835 815 850 835
rect 600 800 850 815
rect 600 750 700 800
rect 750 750 850 800
rect 900 850 1000 900
rect 1050 850 1150 900
rect 900 835 1150 850
rect 900 815 915 835
rect 935 815 965 835
rect 985 815 1015 835
rect 1035 815 1065 835
rect 1085 815 1115 835
rect 1135 815 1150 835
rect 900 800 1150 815
rect 900 750 1000 800
rect 1050 750 1150 800
rect 1200 850 1300 900
rect 1350 850 1450 900
rect 1200 835 1450 850
rect 1200 815 1215 835
rect 1235 815 1265 835
rect 1285 815 1315 835
rect 1335 815 1365 835
rect 1385 815 1415 835
rect 1435 815 1450 835
rect 1200 800 1450 815
rect 1200 750 1300 800
rect 1350 750 1450 800
rect 1500 850 1600 900
rect 1650 850 1750 900
rect 1500 835 1750 850
rect 1500 815 1515 835
rect 1535 815 1565 835
rect 1585 815 1615 835
rect 1635 815 1665 835
rect 1685 815 1715 835
rect 1735 815 1750 835
rect 1500 800 1750 815
rect 1500 750 1600 800
rect 1650 750 1750 800
rect 1800 850 1900 900
rect 1950 850 2050 900
rect 1800 835 2050 850
rect 1800 815 1815 835
rect 1835 815 1865 835
rect 1885 815 1915 835
rect 1935 815 1965 835
rect 1985 815 2015 835
rect 2035 815 2050 835
rect 1800 800 2050 815
rect 1800 750 1900 800
rect 1950 750 2050 800
rect 2100 850 2200 900
rect 2250 850 2350 900
rect 2100 835 2350 850
rect 2100 815 2115 835
rect 2135 815 2165 835
rect 2185 815 2215 835
rect 2235 815 2265 835
rect 2285 815 2315 835
rect 2335 815 2350 835
rect 2100 800 2350 815
rect 2100 750 2200 800
rect 2250 750 2350 800
rect 2400 850 2500 900
rect 2550 850 2650 900
rect 2400 835 2650 850
rect 2400 815 2415 835
rect 2435 815 2465 835
rect 2485 815 2515 835
rect 2535 815 2565 835
rect 2585 815 2615 835
rect 2635 815 2650 835
rect 2400 800 2650 815
rect 2400 750 2500 800
rect 2550 750 2650 800
rect 2700 850 2800 900
rect 2850 850 2950 900
rect 2700 835 2950 850
rect 2700 815 2715 835
rect 2735 815 2765 835
rect 2785 815 2815 835
rect 2835 815 2865 835
rect 2885 815 2915 835
rect 2935 815 2950 835
rect 2700 800 2950 815
rect 2700 750 2800 800
rect 2850 750 2950 800
rect 3000 850 3100 900
rect 3150 850 3250 900
rect 3000 835 3250 850
rect 3000 815 3015 835
rect 3035 815 3065 835
rect 3085 815 3115 835
rect 3135 815 3165 835
rect 3185 815 3215 835
rect 3235 815 3250 835
rect 3000 800 3250 815
rect 3000 750 3100 800
rect 3150 750 3250 800
rect 3300 850 3400 900
rect 3450 850 3550 900
rect 3300 835 3550 850
rect 3300 815 3315 835
rect 3335 815 3365 835
rect 3385 815 3415 835
rect 3435 815 3465 835
rect 3485 815 3515 835
rect 3535 815 3550 835
rect 3300 800 3550 815
rect 3300 750 3400 800
rect 3450 750 3550 800
rect 3600 850 3700 900
rect 3750 850 3850 900
rect 3600 835 3850 850
rect 3600 815 3615 835
rect 3635 815 3665 835
rect 3685 815 3715 835
rect 3735 815 3765 835
rect 3785 815 3815 835
rect 3835 815 3850 835
rect 3600 800 3850 815
rect 3600 750 3700 800
rect 3750 750 3850 800
rect 3900 850 4000 900
rect 4050 850 4150 900
rect 3900 835 4150 850
rect 3900 815 3915 835
rect 3935 815 3965 835
rect 3985 815 4015 835
rect 4035 815 4065 835
rect 4085 815 4115 835
rect 4135 815 4150 835
rect 3900 800 4150 815
rect 3900 750 4000 800
rect 4050 750 4150 800
rect 4200 850 4300 900
rect 4350 850 4450 900
rect 4200 835 4450 850
rect 4200 815 4215 835
rect 4235 815 4265 835
rect 4285 815 4315 835
rect 4335 815 4365 835
rect 4385 815 4415 835
rect 4435 815 4450 835
rect 4200 800 4450 815
rect 4200 750 4300 800
rect 4350 750 4450 800
rect 4500 850 4600 900
rect 4650 850 4750 900
rect 4500 835 4750 850
rect 4500 815 4515 835
rect 4535 815 4565 835
rect 4585 815 4615 835
rect 4635 815 4665 835
rect 4685 815 4715 835
rect 4735 815 4750 835
rect 4500 800 4750 815
rect 4500 750 4600 800
rect 4650 750 4750 800
rect 4800 850 4900 900
rect 4950 850 5050 900
rect 4800 835 5050 850
rect 4800 815 4815 835
rect 4835 815 4865 835
rect 4885 815 4915 835
rect 4935 815 4965 835
rect 4985 815 5015 835
rect 5035 815 5050 835
rect 4800 800 5050 815
rect 4800 750 4900 800
rect 4950 750 5050 800
rect 5100 850 5200 900
rect 5250 850 5350 900
rect 5100 835 5350 850
rect 5100 815 5115 835
rect 5135 815 5165 835
rect 5185 815 5215 835
rect 5235 815 5265 835
rect 5285 815 5315 835
rect 5335 815 5350 835
rect 5100 800 5350 815
rect 5100 750 5200 800
rect 5250 750 5350 800
rect 5400 850 5500 900
rect 5550 850 5650 900
rect 5400 835 5650 850
rect 5400 815 5415 835
rect 5435 815 5465 835
rect 5485 815 5515 835
rect 5535 815 5565 835
rect 5585 815 5615 835
rect 5635 815 5650 835
rect 5400 800 5650 815
rect 5400 750 5500 800
rect 5550 750 5650 800
rect 5700 850 5800 900
rect 5850 850 5950 900
rect 5700 835 5950 850
rect 5700 815 5715 835
rect 5735 815 5765 835
rect 5785 815 5815 835
rect 5835 815 5865 835
rect 5885 815 5915 835
rect 5935 815 5950 835
rect 5700 800 5950 815
rect 5700 750 5800 800
rect 5850 750 5950 800
rect 6000 850 6100 900
rect 6150 850 6250 900
rect 6000 835 6250 850
rect 6000 815 6015 835
rect 6035 815 6065 835
rect 6085 815 6115 835
rect 6135 815 6165 835
rect 6185 815 6215 835
rect 6235 815 6250 835
rect 6000 800 6250 815
rect 6000 750 6100 800
rect 6150 750 6250 800
rect 6300 850 6400 900
rect 6450 850 6550 900
rect 6300 835 6550 850
rect 6300 815 6315 835
rect 6335 815 6365 835
rect 6385 815 6415 835
rect 6435 815 6465 835
rect 6485 815 6515 835
rect 6535 815 6550 835
rect 6300 800 6550 815
rect 6300 750 6400 800
rect 6450 750 6550 800
rect 6600 850 6700 900
rect 6750 850 6850 900
rect 6600 835 6850 850
rect 6600 815 6615 835
rect 6635 815 6665 835
rect 6685 815 6715 835
rect 6735 815 6765 835
rect 6785 815 6815 835
rect 6835 815 6850 835
rect 6600 800 6850 815
rect 6600 750 6700 800
rect 6750 750 6850 800
rect 6900 850 7000 900
rect 7050 850 7150 900
rect 6900 835 7150 850
rect 6900 815 6915 835
rect 6935 815 6965 835
rect 6985 815 7015 835
rect 7035 815 7065 835
rect 7085 815 7115 835
rect 7135 815 7150 835
rect 6900 800 7150 815
rect 6900 750 7000 800
rect 7050 750 7150 800
rect 7200 850 7300 900
rect 7350 850 7450 900
rect 7200 835 7450 850
rect 7200 815 7215 835
rect 7235 815 7265 835
rect 7285 815 7315 835
rect 7335 815 7365 835
rect 7385 815 7415 835
rect 7435 815 7450 835
rect 7200 800 7450 815
rect 7200 750 7300 800
rect 7350 750 7450 800
rect 7500 850 7600 900
rect 7650 850 7750 900
rect 7500 835 7750 850
rect 7500 815 7515 835
rect 7535 815 7565 835
rect 7585 815 7615 835
rect 7635 815 7665 835
rect 7685 815 7715 835
rect 7735 815 7750 835
rect 7500 800 7750 815
rect 7500 750 7600 800
rect 7650 750 7750 800
rect 7800 850 7900 900
rect 7950 850 8050 900
rect 7800 835 8050 850
rect 7800 815 7815 835
rect 7835 815 7865 835
rect 7885 815 7915 835
rect 7935 815 7965 835
rect 7985 815 8015 835
rect 8035 815 8050 835
rect 7800 800 8050 815
rect 7800 750 7900 800
rect 7950 750 8050 800
rect 8100 850 8200 900
rect 8250 850 8350 900
rect 8100 835 8350 850
rect 8100 815 8115 835
rect 8135 815 8165 835
rect 8185 815 8215 835
rect 8235 815 8265 835
rect 8285 815 8315 835
rect 8335 815 8350 835
rect 8100 800 8350 815
rect 8100 750 8200 800
rect 8250 750 8350 800
rect 8400 850 8500 900
rect 8550 850 8650 900
rect 8400 835 8650 850
rect 8400 815 8415 835
rect 8435 815 8465 835
rect 8485 815 8515 835
rect 8535 815 8565 835
rect 8585 815 8615 835
rect 8635 815 8650 835
rect 8400 800 8650 815
rect 8400 750 8500 800
rect 8550 750 8650 800
rect 8700 850 8800 900
rect 8850 850 8950 900
rect 8700 835 8950 850
rect 8700 815 8715 835
rect 8735 815 8765 835
rect 8785 815 8815 835
rect 8835 815 8865 835
rect 8885 815 8915 835
rect 8935 815 8950 835
rect 8700 800 8950 815
rect 8700 750 8800 800
rect 8850 750 8950 800
rect 9000 850 9100 900
rect 9150 850 9250 900
rect 9000 835 9250 850
rect 9000 815 9015 835
rect 9035 815 9065 835
rect 9085 815 9115 835
rect 9135 815 9165 835
rect 9185 815 9215 835
rect 9235 815 9250 835
rect 9000 800 9250 815
rect 9000 750 9100 800
rect 9150 750 9250 800
rect 9300 850 9400 900
rect 9450 850 9550 900
rect 9300 835 9550 850
rect 9300 815 9315 835
rect 9335 815 9365 835
rect 9385 815 9415 835
rect 9435 815 9465 835
rect 9485 815 9515 835
rect 9535 815 9550 835
rect 9300 800 9550 815
rect 9300 750 9400 800
rect 9450 750 9550 800
rect 9600 850 9700 900
rect 9750 850 9850 900
rect 9600 835 9850 850
rect 9600 815 9615 835
rect 9635 815 9665 835
rect 9685 815 9715 835
rect 9735 815 9765 835
rect 9785 815 9815 835
rect 9835 815 9850 835
rect 9600 800 9850 815
rect 9600 750 9700 800
rect 9750 750 9850 800
rect 9900 850 10000 900
rect 10050 850 10150 900
rect 9900 835 10150 850
rect 9900 815 9915 835
rect 9935 815 9965 835
rect 9985 815 10015 835
rect 10035 815 10065 835
rect 10085 815 10115 835
rect 10135 815 10150 835
rect 9900 800 10150 815
rect 9900 750 10000 800
rect 10050 750 10150 800
rect 10200 850 10300 900
rect 10350 850 10450 900
rect 10200 835 10450 850
rect 10200 815 10215 835
rect 10235 815 10265 835
rect 10285 815 10315 835
rect 10335 815 10365 835
rect 10385 815 10415 835
rect 10435 815 10450 835
rect 10200 800 10450 815
rect 10200 750 10300 800
rect 10350 750 10450 800
rect 10500 850 10600 900
rect 10650 850 10750 900
rect 10500 835 10750 850
rect 10500 815 10515 835
rect 10535 815 10565 835
rect 10585 815 10615 835
rect 10635 815 10665 835
rect 10685 815 10715 835
rect 10735 815 10750 835
rect 10500 800 10750 815
rect 10500 750 10600 800
rect 10650 750 10750 800
rect 10800 850 10900 900
rect 10950 850 11050 900
rect 10800 835 11050 850
rect 10800 815 10815 835
rect 10835 815 10865 835
rect 10885 815 10915 835
rect 10935 815 10965 835
rect 10985 815 11015 835
rect 11035 815 11050 835
rect 10800 800 11050 815
rect 10800 750 10900 800
rect 10950 750 11050 800
rect 11100 850 11200 900
rect 11250 850 11350 900
rect 11100 835 11350 850
rect 11100 815 11115 835
rect 11135 815 11165 835
rect 11185 815 11215 835
rect 11235 815 11265 835
rect 11285 815 11315 835
rect 11335 815 11350 835
rect 11100 800 11350 815
rect 11100 750 11200 800
rect 11250 750 11350 800
rect 11400 850 11500 900
rect 11550 850 11650 900
rect 11400 835 11650 850
rect 11400 815 11415 835
rect 11435 815 11465 835
rect 11485 815 11515 835
rect 11535 815 11565 835
rect 11585 815 11615 835
rect 11635 815 11650 835
rect 11400 800 11650 815
rect 11400 750 11500 800
rect 11550 750 11650 800
rect 11700 850 11800 900
rect 11850 850 11950 900
rect 11700 835 11950 850
rect 11700 815 11715 835
rect 11735 815 11765 835
rect 11785 815 11815 835
rect 11835 815 11865 835
rect 11885 815 11915 835
rect 11935 815 11950 835
rect 11700 800 11950 815
rect 11700 750 11800 800
rect 11850 750 11950 800
rect 12000 850 12100 900
rect 12150 850 12250 900
rect 12000 835 12250 850
rect 12000 815 12015 835
rect 12035 815 12065 835
rect 12085 815 12115 835
rect 12135 815 12165 835
rect 12185 815 12215 835
rect 12235 815 12250 835
rect 12000 800 12250 815
rect 12000 750 12100 800
rect 12150 750 12250 800
rect 12300 850 12400 900
rect 12450 850 12550 900
rect 12300 835 12550 850
rect 12300 815 12315 835
rect 12335 815 12365 835
rect 12385 815 12415 835
rect 12435 815 12465 835
rect 12485 815 12515 835
rect 12535 815 12550 835
rect 12300 800 12550 815
rect 12300 750 12400 800
rect 12450 750 12550 800
rect 12600 850 12700 900
rect 12750 850 12850 900
rect 12600 835 12850 850
rect 12600 815 12615 835
rect 12635 815 12665 835
rect 12685 815 12715 835
rect 12735 815 12765 835
rect 12785 815 12815 835
rect 12835 815 12850 835
rect 12600 800 12850 815
rect 12600 750 12700 800
rect 12750 750 12850 800
rect 12900 850 13000 900
rect 13050 850 13150 900
rect 12900 835 13150 850
rect 12900 815 12915 835
rect 12935 815 12965 835
rect 12985 815 13015 835
rect 13035 815 13065 835
rect 13085 815 13115 835
rect 13135 815 13150 835
rect 12900 800 13150 815
rect 12900 750 13000 800
rect 13050 750 13150 800
rect 13200 850 13300 900
rect 13350 850 13450 900
rect 13200 835 13450 850
rect 13200 815 13215 835
rect 13235 815 13265 835
rect 13285 815 13315 835
rect 13335 815 13365 835
rect 13385 815 13415 835
rect 13435 815 13450 835
rect 13200 800 13450 815
rect 13200 750 13300 800
rect 13350 750 13450 800
rect 13500 850 13600 900
rect 13650 850 13750 900
rect 13500 835 13750 850
rect 13500 815 13515 835
rect 13535 815 13565 835
rect 13585 815 13615 835
rect 13635 815 13665 835
rect 13685 815 13715 835
rect 13735 815 13750 835
rect 13500 800 13750 815
rect 13500 750 13600 800
rect 13650 750 13750 800
rect 13800 850 13900 900
rect 13950 850 14050 900
rect 13800 835 14050 850
rect 13800 815 13815 835
rect 13835 815 13865 835
rect 13885 815 13915 835
rect 13935 815 13965 835
rect 13985 815 14015 835
rect 14035 815 14050 835
rect 13800 800 14050 815
rect 13800 750 13900 800
rect 13950 750 14050 800
rect 14100 850 14200 900
rect 14250 850 14350 900
rect 14100 835 14350 850
rect 14100 815 14115 835
rect 14135 815 14165 835
rect 14185 815 14215 835
rect 14235 815 14265 835
rect 14285 815 14315 835
rect 14335 815 14350 835
rect 14100 800 14350 815
rect 14100 750 14200 800
rect 14250 750 14350 800
rect 14400 850 14500 900
rect 14550 850 14650 900
rect 14400 835 14650 850
rect 14400 815 14415 835
rect 14435 815 14465 835
rect 14485 815 14515 835
rect 14535 815 14565 835
rect 14585 815 14615 835
rect 14635 815 14650 835
rect 14400 800 14650 815
rect 14400 750 14500 800
rect 14550 750 14650 800
rect 14700 850 14800 900
rect 14850 850 14950 900
rect 14700 835 14950 850
rect 14700 815 14715 835
rect 14735 815 14765 835
rect 14785 815 14815 835
rect 14835 815 14865 835
rect 14885 815 14915 835
rect 14935 815 14950 835
rect 14700 800 14950 815
rect 14700 750 14800 800
rect 14850 750 14950 800
rect 15000 850 15100 900
rect 15150 850 15250 900
rect 15000 835 15250 850
rect 15000 815 15015 835
rect 15035 815 15065 835
rect 15085 815 15115 835
rect 15135 815 15165 835
rect 15185 815 15215 835
rect 15235 815 15250 835
rect 15000 800 15250 815
rect 15000 750 15100 800
rect 15150 750 15250 800
rect 15300 850 15400 900
rect 15450 850 15550 900
rect 15300 835 15550 850
rect 15300 815 15315 835
rect 15335 815 15365 835
rect 15385 815 15415 835
rect 15435 815 15465 835
rect 15485 815 15515 835
rect 15535 815 15550 835
rect 15300 800 15550 815
rect 15300 750 15400 800
rect 15450 750 15550 800
rect 15600 850 15700 900
rect 15750 850 15850 900
rect 15600 835 15850 850
rect 15600 815 15615 835
rect 15635 815 15665 835
rect 15685 815 15715 835
rect 15735 815 15765 835
rect 15785 815 15815 835
rect 15835 815 15850 835
rect 15600 800 15850 815
rect 15600 750 15700 800
rect 15750 750 15850 800
rect 15900 850 16000 900
rect 16050 850 16150 900
rect 15900 835 16150 850
rect 15900 815 15915 835
rect 15935 815 15965 835
rect 15985 815 16015 835
rect 16035 815 16065 835
rect 16085 815 16115 835
rect 16135 815 16150 835
rect 15900 800 16150 815
rect 15900 750 16000 800
rect 16050 750 16150 800
rect 16200 850 16300 900
rect 16350 850 16450 900
rect 16200 835 16450 850
rect 16200 815 16215 835
rect 16235 815 16265 835
rect 16285 815 16315 835
rect 16335 815 16365 835
rect 16385 815 16415 835
rect 16435 815 16450 835
rect 16200 800 16450 815
rect 16200 750 16300 800
rect 16350 750 16450 800
rect 16500 850 16600 900
rect 16650 850 16750 900
rect 16500 835 16750 850
rect 16500 815 16515 835
rect 16535 815 16565 835
rect 16585 815 16615 835
rect 16635 815 16665 835
rect 16685 815 16715 835
rect 16735 815 16750 835
rect 16500 800 16750 815
rect 16500 750 16600 800
rect 16650 750 16750 800
rect 16800 850 16900 900
rect 16950 850 17050 900
rect 16800 835 17050 850
rect 16800 815 16815 835
rect 16835 815 16865 835
rect 16885 815 16915 835
rect 16935 815 16965 835
rect 16985 815 17015 835
rect 17035 815 17050 835
rect 16800 800 17050 815
rect 16800 750 16900 800
rect 16950 750 17050 800
rect 17100 850 17200 900
rect 17250 850 17350 900
rect 17100 835 17350 850
rect 17100 815 17115 835
rect 17135 815 17165 835
rect 17185 815 17215 835
rect 17235 815 17265 835
rect 17285 815 17315 835
rect 17335 815 17350 835
rect 17100 800 17350 815
rect 17100 750 17200 800
rect 17250 750 17350 800
rect 17400 850 17500 900
rect 17550 850 17650 900
rect 17400 835 17650 850
rect 17400 815 17415 835
rect 17435 815 17465 835
rect 17485 815 17515 835
rect 17535 815 17565 835
rect 17585 815 17615 835
rect 17635 815 17650 835
rect 17400 800 17650 815
rect 17400 750 17500 800
rect 17550 750 17650 800
rect 17700 850 17800 900
rect 17850 850 17950 900
rect 17700 835 17950 850
rect 17700 815 17715 835
rect 17735 815 17765 835
rect 17785 815 17815 835
rect 17835 815 17865 835
rect 17885 815 17915 835
rect 17935 815 17950 835
rect 17700 800 17950 815
rect 17700 750 17800 800
rect 17850 750 17950 800
rect 18000 850 18100 900
rect 18150 850 18250 900
rect 18000 835 18250 850
rect 18000 815 18015 835
rect 18035 815 18065 835
rect 18085 815 18115 835
rect 18135 815 18165 835
rect 18185 815 18215 835
rect 18235 815 18250 835
rect 18000 800 18250 815
rect 18000 750 18100 800
rect 18150 750 18250 800
rect 18300 850 18400 900
rect 18450 850 18550 900
rect 18300 835 18550 850
rect 18300 815 18315 835
rect 18335 815 18365 835
rect 18385 815 18415 835
rect 18435 815 18465 835
rect 18485 815 18515 835
rect 18535 815 18550 835
rect 18300 800 18550 815
rect 18300 750 18400 800
rect 18450 750 18550 800
rect 18600 850 18700 900
rect 18750 850 18850 900
rect 18600 835 18850 850
rect 18600 815 18615 835
rect 18635 815 18665 835
rect 18685 815 18715 835
rect 18735 815 18765 835
rect 18785 815 18815 835
rect 18835 815 18850 835
rect 18600 800 18850 815
rect 18600 750 18700 800
rect 18750 750 18850 800
rect 18900 850 19000 900
rect 19050 850 19150 900
rect 18900 835 19150 850
rect 18900 815 18915 835
rect 18935 815 18965 835
rect 18985 815 19015 835
rect 19035 815 19065 835
rect 19085 815 19115 835
rect 19135 815 19150 835
rect 18900 800 19150 815
rect 18900 750 19000 800
rect 19050 750 19150 800
rect 19200 850 19300 900
rect 19350 850 19450 900
rect 19200 835 19450 850
rect 19200 815 19215 835
rect 19235 815 19265 835
rect 19285 815 19315 835
rect 19335 815 19365 835
rect 19385 815 19415 835
rect 19435 815 19450 835
rect 19200 800 19450 815
rect 19200 750 19300 800
rect 19350 750 19450 800
rect 19500 850 19600 900
rect 19650 850 19750 900
rect 19500 835 19750 850
rect 19500 815 19515 835
rect 19535 815 19565 835
rect 19585 815 19615 835
rect 19635 815 19665 835
rect 19685 815 19715 835
rect 19735 815 19750 835
rect 19500 800 19750 815
rect 19500 750 19600 800
rect 19650 750 19750 800
rect 19800 850 19900 900
rect 19950 850 20050 900
rect 19800 835 20050 850
rect 19800 815 19815 835
rect 19835 815 19865 835
rect 19885 815 19915 835
rect 19935 815 19965 835
rect 19985 815 20015 835
rect 20035 815 20050 835
rect 19800 800 20050 815
rect 19800 750 19900 800
rect 19950 750 20050 800
rect 20100 850 20200 900
rect 20250 850 20350 900
rect 20100 835 20350 850
rect 20100 815 20115 835
rect 20135 815 20165 835
rect 20185 815 20215 835
rect 20235 815 20265 835
rect 20285 815 20315 835
rect 20335 815 20350 835
rect 20100 800 20350 815
rect 20100 750 20200 800
rect 20250 750 20350 800
rect -600 35 -500 50
rect -450 35 -350 50
rect -300 35 -200 50
rect -150 35 -50 50
rect 0 35 100 50
rect 150 35 250 50
rect 300 35 400 50
rect 450 35 550 50
rect 600 35 700 50
rect 750 35 850 50
rect 900 35 1000 50
rect 1050 35 1150 50
rect 1200 35 1300 50
rect 1350 35 1450 50
rect 1500 35 1600 50
rect 1650 35 1750 50
rect 1800 35 1900 50
rect 1950 35 2050 50
rect 2100 35 2200 50
rect 2250 35 2350 50
rect 2400 35 2500 50
rect 2550 35 2650 50
rect 2700 35 2800 50
rect 2850 35 2950 50
rect 3000 35 3100 50
rect 3150 35 3250 50
rect 3300 35 3400 50
rect 3450 35 3550 50
rect 3600 35 3700 50
rect 3750 35 3850 50
rect 3900 35 4000 50
rect 4050 35 4150 50
rect 4200 35 4300 50
rect 4350 35 4450 50
rect 4500 35 4600 50
rect 4650 35 4750 50
rect 4800 35 4900 50
rect 4950 35 5050 50
rect 5100 35 5200 50
rect 5250 35 5350 50
rect 5400 35 5500 50
rect 5550 35 5650 50
rect 5700 35 5800 50
rect 5850 35 5950 50
rect 6000 35 6100 50
rect 6150 35 6250 50
rect 6300 35 6400 50
rect 6450 35 6550 50
rect 6600 35 6700 50
rect 6750 35 6850 50
rect 6900 35 7000 50
rect 7050 35 7150 50
rect 7200 35 7300 50
rect 7350 35 7450 50
rect 7500 35 7600 50
rect 7650 35 7750 50
rect 7800 35 7900 50
rect 7950 35 8050 50
rect 8100 35 8200 50
rect 8250 35 8350 50
rect 8400 35 8500 50
rect 8550 35 8650 50
rect 8700 35 8800 50
rect 8850 35 8950 50
rect 9000 35 9100 50
rect 9150 35 9250 50
rect 9300 35 9400 50
rect 9450 35 9550 50
rect 9600 35 9700 50
rect 9750 35 9850 50
rect 9900 35 10000 50
rect 10050 35 10150 50
rect 10200 35 10300 50
rect 10350 35 10450 50
rect 10500 35 10600 50
rect 10650 35 10750 50
rect 10800 35 10900 50
rect 10950 35 11050 50
rect 11100 35 11200 50
rect 11250 35 11350 50
rect 11400 35 11500 50
rect 11550 35 11650 50
rect 11700 35 11800 50
rect 11850 35 11950 50
rect 12000 35 12100 50
rect 12150 35 12250 50
rect 12300 35 12400 50
rect 12450 35 12550 50
rect 12600 35 12700 50
rect 12750 35 12850 50
rect 12900 35 13000 50
rect 13050 35 13150 50
rect 13200 35 13300 50
rect 13350 35 13450 50
rect 13500 35 13600 50
rect 13650 35 13750 50
rect 13800 35 13900 50
rect 13950 35 14050 50
rect 14100 35 14200 50
rect 14250 35 14350 50
rect 14400 35 14500 50
rect 14550 35 14650 50
rect 14700 35 14800 50
rect 14850 35 14950 50
rect 15000 35 15100 50
rect 15150 35 15250 50
rect 15300 35 15400 50
rect 15450 35 15550 50
rect 15600 35 15700 50
rect 15750 35 15850 50
rect 15900 35 16000 50
rect 16050 35 16150 50
rect 16200 35 16300 50
rect 16350 35 16450 50
rect 16500 35 16600 50
rect 16650 35 16750 50
rect 16800 35 16900 50
rect 16950 35 17050 50
rect 17100 35 17200 50
rect 17250 35 17350 50
rect 17400 35 17500 50
rect 17550 35 17650 50
rect 17700 35 17800 50
rect 17850 35 17950 50
rect 18000 35 18100 50
rect 18150 35 18250 50
rect 18300 35 18400 50
rect 18450 35 18550 50
rect 18600 35 18700 50
rect 18750 35 18850 50
rect 18900 35 19000 50
rect 19050 35 19150 50
rect 19200 35 19300 50
rect 19350 35 19450 50
rect 19500 35 19600 50
rect 19650 35 19750 50
rect 19800 35 19900 50
rect 19950 35 20050 50
rect 20100 35 20200 50
rect 20250 35 20350 50
rect -600 -100 -500 -85
rect -450 -100 -350 -85
rect -300 -100 -200 -85
rect -150 -100 -50 -85
rect 0 -100 100 -85
rect 150 -100 250 -85
rect 300 -100 400 -85
rect 450 -100 550 -85
rect 600 -100 700 -85
rect 750 -100 850 -85
rect 900 -100 1000 -85
rect 1050 -100 1150 -85
rect 1200 -100 1300 -85
rect 1350 -100 1450 -85
rect 1500 -100 1600 -85
rect 1650 -100 1750 -85
rect 1800 -100 1900 -85
rect 1950 -100 2050 -85
rect 2100 -100 2200 -85
rect 2250 -100 2350 -85
rect 2400 -100 2500 -85
rect 2550 -100 2650 -85
rect 2700 -100 2800 -85
rect 2850 -100 2950 -85
rect 3000 -100 3100 -85
rect 3150 -100 3250 -85
rect 3300 -100 3400 -85
rect 3450 -100 3550 -85
rect 3600 -100 3700 -85
rect 3750 -100 3850 -85
rect 3900 -100 4000 -85
rect 4050 -100 4150 -85
rect 4200 -100 4300 -85
rect 4350 -100 4450 -85
rect 4500 -100 4600 -85
rect 4650 -100 4750 -85
rect 4800 -100 4900 -85
rect 4950 -100 5050 -85
rect 5100 -100 5200 -85
rect 5250 -100 5350 -85
rect 5400 -100 5500 -85
rect 5550 -100 5650 -85
rect 5700 -100 5800 -85
rect 5850 -100 5950 -85
rect 6000 -100 6100 -85
rect 6150 -100 6250 -85
rect 6300 -100 6400 -85
rect 6450 -100 6550 -85
rect 6600 -100 6700 -85
rect 6750 -100 6850 -85
rect 6900 -100 7000 -85
rect 7050 -100 7150 -85
rect 7200 -100 7300 -85
rect 7350 -100 7450 -85
rect 7500 -100 7600 -85
rect 7650 -100 7750 -85
rect 7800 -100 7900 -85
rect 7950 -100 8050 -85
rect 8100 -100 8200 -85
rect 8250 -100 8350 -85
rect 8400 -100 8500 -85
rect 8550 -100 8650 -85
rect 8700 -100 8800 -85
rect 8850 -100 8950 -85
rect 9000 -100 9100 -85
rect 9150 -100 9250 -85
rect 9300 -100 9400 -85
rect 9450 -100 9550 -85
rect 9600 -100 9700 -85
rect 9750 -100 9850 -85
rect 9900 -100 10000 -85
rect 10050 -100 10150 -85
rect 10200 -100 10300 -85
rect 10350 -100 10450 -85
rect 10500 -100 10600 -85
rect 10650 -100 10750 -85
rect 10800 -100 10900 -85
rect 10950 -100 11050 -85
rect 11100 -100 11200 -85
rect 11250 -100 11350 -85
rect 11400 -100 11500 -85
rect 11550 -100 11650 -85
rect 11700 -100 11800 -85
rect 11850 -100 11950 -85
rect 12000 -100 12100 -85
rect 12150 -100 12250 -85
rect 12300 -100 12400 -85
rect 12450 -100 12550 -85
rect 12600 -100 12700 -85
rect 12750 -100 12850 -85
rect 12900 -100 13000 -85
rect 13050 -100 13150 -85
rect 13200 -100 13300 -85
rect 13350 -100 13450 -85
rect 13500 -100 13600 -85
rect 13650 -100 13750 -85
rect 13800 -100 13900 -85
rect 13950 -100 14050 -85
rect 14100 -100 14200 -85
rect 14250 -100 14350 -85
rect 14400 -100 14500 -85
rect 14550 -100 14650 -85
rect 14700 -100 14800 -85
rect 14850 -100 14950 -85
rect 15000 -100 15100 -85
rect 15150 -100 15250 -85
rect 15300 -100 15400 -85
rect 15450 -100 15550 -85
rect 15600 -100 15700 -85
rect 15750 -100 15850 -85
rect 15900 -100 16000 -85
rect 16050 -100 16150 -85
rect 16200 -100 16300 -85
rect 16350 -100 16450 -85
rect 16500 -100 16600 -85
rect 16650 -100 16750 -85
rect 16800 -100 16900 -85
rect 16950 -100 17050 -85
rect 17100 -100 17200 -85
rect 17250 -100 17350 -85
rect 17400 -100 17500 -85
rect 17550 -100 17650 -85
rect 17700 -100 17800 -85
rect 17850 -100 17950 -85
rect 18000 -100 18100 -85
rect 18150 -100 18250 -85
rect 18300 -100 18400 -85
rect 18450 -100 18550 -85
rect 18600 -100 18700 -85
rect 18750 -100 18850 -85
rect 18900 -100 19000 -85
rect 19050 -100 19150 -85
rect 19200 -100 19300 -85
rect 19350 -100 19450 -85
rect 19500 -100 19600 -85
rect 19650 -100 19750 -85
rect 19800 -100 19900 -85
rect 19950 -100 20050 -85
rect 20100 -100 20200 -85
rect 20250 -100 20350 -85
rect -600 -850 -500 -800
rect -450 -850 -350 -800
rect -600 -865 -350 -850
rect -600 -885 -585 -865
rect -565 -885 -535 -865
rect -515 -885 -485 -865
rect -465 -885 -435 -865
rect -415 -885 -385 -865
rect -365 -885 -350 -865
rect -600 -900 -350 -885
rect -600 -950 -500 -900
rect -450 -950 -350 -900
rect -300 -850 -200 -800
rect -150 -850 -50 -800
rect -300 -865 -50 -850
rect -300 -885 -285 -865
rect -265 -885 -235 -865
rect -215 -885 -185 -865
rect -165 -885 -135 -865
rect -115 -885 -85 -865
rect -65 -885 -50 -865
rect -300 -900 -50 -885
rect -300 -950 -200 -900
rect -150 -950 -50 -900
rect 0 -850 100 -800
rect 150 -850 250 -800
rect 0 -865 250 -850
rect 0 -885 15 -865
rect 35 -885 65 -865
rect 85 -885 115 -865
rect 135 -885 165 -865
rect 185 -885 215 -865
rect 235 -885 250 -865
rect 0 -900 250 -885
rect 0 -950 100 -900
rect 150 -950 250 -900
rect 300 -850 400 -800
rect 450 -850 550 -800
rect 300 -865 550 -850
rect 300 -885 315 -865
rect 335 -885 365 -865
rect 385 -885 415 -865
rect 435 -885 465 -865
rect 485 -885 515 -865
rect 535 -885 550 -865
rect 300 -900 550 -885
rect 300 -950 400 -900
rect 450 -950 550 -900
rect 600 -850 700 -800
rect 750 -850 850 -800
rect 600 -865 850 -850
rect 600 -885 615 -865
rect 635 -885 665 -865
rect 685 -885 715 -865
rect 735 -885 765 -865
rect 785 -885 815 -865
rect 835 -885 850 -865
rect 600 -900 850 -885
rect 600 -950 700 -900
rect 750 -950 850 -900
rect 900 -850 1000 -800
rect 1050 -850 1150 -800
rect 900 -865 1150 -850
rect 900 -885 915 -865
rect 935 -885 965 -865
rect 985 -885 1015 -865
rect 1035 -885 1065 -865
rect 1085 -885 1115 -865
rect 1135 -885 1150 -865
rect 900 -900 1150 -885
rect 900 -950 1000 -900
rect 1050 -950 1150 -900
rect 1200 -850 1300 -800
rect 1350 -850 1450 -800
rect 1200 -865 1450 -850
rect 1200 -885 1215 -865
rect 1235 -885 1265 -865
rect 1285 -885 1315 -865
rect 1335 -885 1365 -865
rect 1385 -885 1415 -865
rect 1435 -885 1450 -865
rect 1200 -900 1450 -885
rect 1200 -950 1300 -900
rect 1350 -950 1450 -900
rect 1500 -850 1600 -800
rect 1650 -850 1750 -800
rect 1500 -865 1750 -850
rect 1500 -885 1515 -865
rect 1535 -885 1565 -865
rect 1585 -885 1615 -865
rect 1635 -885 1665 -865
rect 1685 -885 1715 -865
rect 1735 -885 1750 -865
rect 1500 -900 1750 -885
rect 1500 -950 1600 -900
rect 1650 -950 1750 -900
rect 1800 -850 1900 -800
rect 1950 -850 2050 -800
rect 1800 -865 2050 -850
rect 1800 -885 1815 -865
rect 1835 -885 1865 -865
rect 1885 -885 1915 -865
rect 1935 -885 1965 -865
rect 1985 -885 2015 -865
rect 2035 -885 2050 -865
rect 1800 -900 2050 -885
rect 1800 -950 1900 -900
rect 1950 -950 2050 -900
rect 2100 -850 2200 -800
rect 2250 -850 2350 -800
rect 2100 -865 2350 -850
rect 2100 -885 2115 -865
rect 2135 -885 2165 -865
rect 2185 -885 2215 -865
rect 2235 -885 2265 -865
rect 2285 -885 2315 -865
rect 2335 -885 2350 -865
rect 2100 -900 2350 -885
rect 2100 -950 2200 -900
rect 2250 -950 2350 -900
rect 2400 -850 2500 -800
rect 2550 -850 2650 -800
rect 2400 -865 2650 -850
rect 2400 -885 2415 -865
rect 2435 -885 2465 -865
rect 2485 -885 2515 -865
rect 2535 -885 2565 -865
rect 2585 -885 2615 -865
rect 2635 -885 2650 -865
rect 2400 -900 2650 -885
rect 2400 -950 2500 -900
rect 2550 -950 2650 -900
rect 2700 -850 2800 -800
rect 2850 -850 2950 -800
rect 2700 -865 2950 -850
rect 2700 -885 2715 -865
rect 2735 -885 2765 -865
rect 2785 -885 2815 -865
rect 2835 -885 2865 -865
rect 2885 -885 2915 -865
rect 2935 -885 2950 -865
rect 2700 -900 2950 -885
rect 2700 -950 2800 -900
rect 2850 -950 2950 -900
rect 3000 -850 3100 -800
rect 3150 -850 3250 -800
rect 3000 -865 3250 -850
rect 3000 -885 3015 -865
rect 3035 -885 3065 -865
rect 3085 -885 3115 -865
rect 3135 -885 3165 -865
rect 3185 -885 3215 -865
rect 3235 -885 3250 -865
rect 3000 -900 3250 -885
rect 3000 -950 3100 -900
rect 3150 -950 3250 -900
rect 3300 -850 3400 -800
rect 3450 -850 3550 -800
rect 3300 -865 3550 -850
rect 3300 -885 3315 -865
rect 3335 -885 3365 -865
rect 3385 -885 3415 -865
rect 3435 -885 3465 -865
rect 3485 -885 3515 -865
rect 3535 -885 3550 -865
rect 3300 -900 3550 -885
rect 3300 -950 3400 -900
rect 3450 -950 3550 -900
rect 3600 -850 3700 -800
rect 3750 -850 3850 -800
rect 3600 -865 3850 -850
rect 3600 -885 3615 -865
rect 3635 -885 3665 -865
rect 3685 -885 3715 -865
rect 3735 -885 3765 -865
rect 3785 -885 3815 -865
rect 3835 -885 3850 -865
rect 3600 -900 3850 -885
rect 3600 -950 3700 -900
rect 3750 -950 3850 -900
rect 3900 -850 4000 -800
rect 4050 -850 4150 -800
rect 3900 -865 4150 -850
rect 3900 -885 3915 -865
rect 3935 -885 3965 -865
rect 3985 -885 4015 -865
rect 4035 -885 4065 -865
rect 4085 -885 4115 -865
rect 4135 -885 4150 -865
rect 3900 -900 4150 -885
rect 3900 -950 4000 -900
rect 4050 -950 4150 -900
rect 4200 -850 4300 -800
rect 4350 -850 4450 -800
rect 4200 -865 4450 -850
rect 4200 -885 4215 -865
rect 4235 -885 4265 -865
rect 4285 -885 4315 -865
rect 4335 -885 4365 -865
rect 4385 -885 4415 -865
rect 4435 -885 4450 -865
rect 4200 -900 4450 -885
rect 4200 -950 4300 -900
rect 4350 -950 4450 -900
rect 4500 -850 4600 -800
rect 4650 -850 4750 -800
rect 4500 -865 4750 -850
rect 4500 -885 4515 -865
rect 4535 -885 4565 -865
rect 4585 -885 4615 -865
rect 4635 -885 4665 -865
rect 4685 -885 4715 -865
rect 4735 -885 4750 -865
rect 4500 -900 4750 -885
rect 4500 -950 4600 -900
rect 4650 -950 4750 -900
rect 4800 -850 4900 -800
rect 4950 -850 5050 -800
rect 4800 -865 5050 -850
rect 4800 -885 4815 -865
rect 4835 -885 4865 -865
rect 4885 -885 4915 -865
rect 4935 -885 4965 -865
rect 4985 -885 5015 -865
rect 5035 -885 5050 -865
rect 4800 -900 5050 -885
rect 4800 -950 4900 -900
rect 4950 -950 5050 -900
rect 5100 -850 5200 -800
rect 5250 -850 5350 -800
rect 5100 -865 5350 -850
rect 5100 -885 5115 -865
rect 5135 -885 5165 -865
rect 5185 -885 5215 -865
rect 5235 -885 5265 -865
rect 5285 -885 5315 -865
rect 5335 -885 5350 -865
rect 5100 -900 5350 -885
rect 5100 -950 5200 -900
rect 5250 -950 5350 -900
rect 5400 -850 5500 -800
rect 5550 -850 5650 -800
rect 5400 -865 5650 -850
rect 5400 -885 5415 -865
rect 5435 -885 5465 -865
rect 5485 -885 5515 -865
rect 5535 -885 5565 -865
rect 5585 -885 5615 -865
rect 5635 -885 5650 -865
rect 5400 -900 5650 -885
rect 5400 -950 5500 -900
rect 5550 -950 5650 -900
rect 5700 -850 5800 -800
rect 5850 -850 5950 -800
rect 5700 -865 5950 -850
rect 5700 -885 5715 -865
rect 5735 -885 5765 -865
rect 5785 -885 5815 -865
rect 5835 -885 5865 -865
rect 5885 -885 5915 -865
rect 5935 -885 5950 -865
rect 5700 -900 5950 -885
rect 5700 -950 5800 -900
rect 5850 -950 5950 -900
rect 6000 -850 6100 -800
rect 6150 -850 6250 -800
rect 6000 -865 6250 -850
rect 6000 -885 6015 -865
rect 6035 -885 6065 -865
rect 6085 -885 6115 -865
rect 6135 -885 6165 -865
rect 6185 -885 6215 -865
rect 6235 -885 6250 -865
rect 6000 -900 6250 -885
rect 6000 -950 6100 -900
rect 6150 -950 6250 -900
rect 6300 -850 6400 -800
rect 6450 -850 6550 -800
rect 6300 -865 6550 -850
rect 6300 -885 6315 -865
rect 6335 -885 6365 -865
rect 6385 -885 6415 -865
rect 6435 -885 6465 -865
rect 6485 -885 6515 -865
rect 6535 -885 6550 -865
rect 6300 -900 6550 -885
rect 6300 -950 6400 -900
rect 6450 -950 6550 -900
rect 6600 -850 6700 -800
rect 6750 -850 6850 -800
rect 6600 -865 6850 -850
rect 6600 -885 6615 -865
rect 6635 -885 6665 -865
rect 6685 -885 6715 -865
rect 6735 -885 6765 -865
rect 6785 -885 6815 -865
rect 6835 -885 6850 -865
rect 6600 -900 6850 -885
rect 6600 -950 6700 -900
rect 6750 -950 6850 -900
rect 6900 -850 7000 -800
rect 7050 -850 7150 -800
rect 6900 -865 7150 -850
rect 6900 -885 6915 -865
rect 6935 -885 6965 -865
rect 6985 -885 7015 -865
rect 7035 -885 7065 -865
rect 7085 -885 7115 -865
rect 7135 -885 7150 -865
rect 6900 -900 7150 -885
rect 6900 -950 7000 -900
rect 7050 -950 7150 -900
rect 7200 -850 7300 -800
rect 7350 -850 7450 -800
rect 7200 -865 7450 -850
rect 7200 -885 7215 -865
rect 7235 -885 7265 -865
rect 7285 -885 7315 -865
rect 7335 -885 7365 -865
rect 7385 -885 7415 -865
rect 7435 -885 7450 -865
rect 7200 -900 7450 -885
rect 7200 -950 7300 -900
rect 7350 -950 7450 -900
rect 7500 -850 7600 -800
rect 7650 -850 7750 -800
rect 7500 -865 7750 -850
rect 7500 -885 7515 -865
rect 7535 -885 7565 -865
rect 7585 -885 7615 -865
rect 7635 -885 7665 -865
rect 7685 -885 7715 -865
rect 7735 -885 7750 -865
rect 7500 -900 7750 -885
rect 7500 -950 7600 -900
rect 7650 -950 7750 -900
rect 7800 -850 7900 -800
rect 7950 -850 8050 -800
rect 7800 -865 8050 -850
rect 7800 -885 7815 -865
rect 7835 -885 7865 -865
rect 7885 -885 7915 -865
rect 7935 -885 7965 -865
rect 7985 -885 8015 -865
rect 8035 -885 8050 -865
rect 7800 -900 8050 -885
rect 7800 -950 7900 -900
rect 7950 -950 8050 -900
rect 8100 -850 8200 -800
rect 8250 -850 8350 -800
rect 8100 -865 8350 -850
rect 8100 -885 8115 -865
rect 8135 -885 8165 -865
rect 8185 -885 8215 -865
rect 8235 -885 8265 -865
rect 8285 -885 8315 -865
rect 8335 -885 8350 -865
rect 8100 -900 8350 -885
rect 8100 -950 8200 -900
rect 8250 -950 8350 -900
rect 8400 -850 8500 -800
rect 8550 -850 8650 -800
rect 8400 -865 8650 -850
rect 8400 -885 8415 -865
rect 8435 -885 8465 -865
rect 8485 -885 8515 -865
rect 8535 -885 8565 -865
rect 8585 -885 8615 -865
rect 8635 -885 8650 -865
rect 8400 -900 8650 -885
rect 8400 -950 8500 -900
rect 8550 -950 8650 -900
rect 8700 -850 8800 -800
rect 8850 -850 8950 -800
rect 8700 -865 8950 -850
rect 8700 -885 8715 -865
rect 8735 -885 8765 -865
rect 8785 -885 8815 -865
rect 8835 -885 8865 -865
rect 8885 -885 8915 -865
rect 8935 -885 8950 -865
rect 8700 -900 8950 -885
rect 8700 -950 8800 -900
rect 8850 -950 8950 -900
rect 9000 -850 9100 -800
rect 9150 -850 9250 -800
rect 9000 -865 9250 -850
rect 9000 -885 9015 -865
rect 9035 -885 9065 -865
rect 9085 -885 9115 -865
rect 9135 -885 9165 -865
rect 9185 -885 9215 -865
rect 9235 -885 9250 -865
rect 9000 -900 9250 -885
rect 9000 -950 9100 -900
rect 9150 -950 9250 -900
rect 9300 -850 9400 -800
rect 9450 -850 9550 -800
rect 9300 -865 9550 -850
rect 9300 -885 9315 -865
rect 9335 -885 9365 -865
rect 9385 -885 9415 -865
rect 9435 -885 9465 -865
rect 9485 -885 9515 -865
rect 9535 -885 9550 -865
rect 9300 -900 9550 -885
rect 9300 -950 9400 -900
rect 9450 -950 9550 -900
rect 9600 -850 9700 -800
rect 9750 -850 9850 -800
rect 9600 -865 9850 -850
rect 9600 -885 9615 -865
rect 9635 -885 9665 -865
rect 9685 -885 9715 -865
rect 9735 -885 9765 -865
rect 9785 -885 9815 -865
rect 9835 -885 9850 -865
rect 9600 -900 9850 -885
rect 9600 -950 9700 -900
rect 9750 -950 9850 -900
rect 9900 -850 10000 -800
rect 10050 -850 10150 -800
rect 9900 -865 10150 -850
rect 9900 -885 9915 -865
rect 9935 -885 9965 -865
rect 9985 -885 10015 -865
rect 10035 -885 10065 -865
rect 10085 -885 10115 -865
rect 10135 -885 10150 -865
rect 9900 -900 10150 -885
rect 9900 -950 10000 -900
rect 10050 -950 10150 -900
rect 10200 -850 10300 -800
rect 10350 -850 10450 -800
rect 10200 -865 10450 -850
rect 10200 -885 10215 -865
rect 10235 -885 10265 -865
rect 10285 -885 10315 -865
rect 10335 -885 10365 -865
rect 10385 -885 10415 -865
rect 10435 -885 10450 -865
rect 10200 -900 10450 -885
rect 10200 -950 10300 -900
rect 10350 -950 10450 -900
rect 10500 -850 10600 -800
rect 10650 -850 10750 -800
rect 10500 -865 10750 -850
rect 10500 -885 10515 -865
rect 10535 -885 10565 -865
rect 10585 -885 10615 -865
rect 10635 -885 10665 -865
rect 10685 -885 10715 -865
rect 10735 -885 10750 -865
rect 10500 -900 10750 -885
rect 10500 -950 10600 -900
rect 10650 -950 10750 -900
rect 10800 -850 10900 -800
rect 10950 -850 11050 -800
rect 10800 -865 11050 -850
rect 10800 -885 10815 -865
rect 10835 -885 10865 -865
rect 10885 -885 10915 -865
rect 10935 -885 10965 -865
rect 10985 -885 11015 -865
rect 11035 -885 11050 -865
rect 10800 -900 11050 -885
rect 10800 -950 10900 -900
rect 10950 -950 11050 -900
rect 11100 -850 11200 -800
rect 11250 -850 11350 -800
rect 11100 -865 11350 -850
rect 11100 -885 11115 -865
rect 11135 -885 11165 -865
rect 11185 -885 11215 -865
rect 11235 -885 11265 -865
rect 11285 -885 11315 -865
rect 11335 -885 11350 -865
rect 11100 -900 11350 -885
rect 11100 -950 11200 -900
rect 11250 -950 11350 -900
rect 11400 -850 11500 -800
rect 11550 -850 11650 -800
rect 11400 -865 11650 -850
rect 11400 -885 11415 -865
rect 11435 -885 11465 -865
rect 11485 -885 11515 -865
rect 11535 -885 11565 -865
rect 11585 -885 11615 -865
rect 11635 -885 11650 -865
rect 11400 -900 11650 -885
rect 11400 -950 11500 -900
rect 11550 -950 11650 -900
rect 11700 -850 11800 -800
rect 11850 -850 11950 -800
rect 11700 -865 11950 -850
rect 11700 -885 11715 -865
rect 11735 -885 11765 -865
rect 11785 -885 11815 -865
rect 11835 -885 11865 -865
rect 11885 -885 11915 -865
rect 11935 -885 11950 -865
rect 11700 -900 11950 -885
rect 11700 -950 11800 -900
rect 11850 -950 11950 -900
rect 12000 -850 12100 -800
rect 12150 -850 12250 -800
rect 12000 -865 12250 -850
rect 12000 -885 12015 -865
rect 12035 -885 12065 -865
rect 12085 -885 12115 -865
rect 12135 -885 12165 -865
rect 12185 -885 12215 -865
rect 12235 -885 12250 -865
rect 12000 -900 12250 -885
rect 12000 -950 12100 -900
rect 12150 -950 12250 -900
rect 12300 -850 12400 -800
rect 12450 -850 12550 -800
rect 12300 -865 12550 -850
rect 12300 -885 12315 -865
rect 12335 -885 12365 -865
rect 12385 -885 12415 -865
rect 12435 -885 12465 -865
rect 12485 -885 12515 -865
rect 12535 -885 12550 -865
rect 12300 -900 12550 -885
rect 12300 -950 12400 -900
rect 12450 -950 12550 -900
rect 12600 -850 12700 -800
rect 12750 -850 12850 -800
rect 12600 -865 12850 -850
rect 12600 -885 12615 -865
rect 12635 -885 12665 -865
rect 12685 -885 12715 -865
rect 12735 -885 12765 -865
rect 12785 -885 12815 -865
rect 12835 -885 12850 -865
rect 12600 -900 12850 -885
rect 12600 -950 12700 -900
rect 12750 -950 12850 -900
rect 12900 -850 13000 -800
rect 13050 -850 13150 -800
rect 12900 -865 13150 -850
rect 12900 -885 12915 -865
rect 12935 -885 12965 -865
rect 12985 -885 13015 -865
rect 13035 -885 13065 -865
rect 13085 -885 13115 -865
rect 13135 -885 13150 -865
rect 12900 -900 13150 -885
rect 12900 -950 13000 -900
rect 13050 -950 13150 -900
rect 13200 -850 13300 -800
rect 13350 -850 13450 -800
rect 13200 -865 13450 -850
rect 13200 -885 13215 -865
rect 13235 -885 13265 -865
rect 13285 -885 13315 -865
rect 13335 -885 13365 -865
rect 13385 -885 13415 -865
rect 13435 -885 13450 -865
rect 13200 -900 13450 -885
rect 13200 -950 13300 -900
rect 13350 -950 13450 -900
rect 13500 -850 13600 -800
rect 13650 -850 13750 -800
rect 13500 -865 13750 -850
rect 13500 -885 13515 -865
rect 13535 -885 13565 -865
rect 13585 -885 13615 -865
rect 13635 -885 13665 -865
rect 13685 -885 13715 -865
rect 13735 -885 13750 -865
rect 13500 -900 13750 -885
rect 13500 -950 13600 -900
rect 13650 -950 13750 -900
rect 13800 -850 13900 -800
rect 13950 -850 14050 -800
rect 13800 -865 14050 -850
rect 13800 -885 13815 -865
rect 13835 -885 13865 -865
rect 13885 -885 13915 -865
rect 13935 -885 13965 -865
rect 13985 -885 14015 -865
rect 14035 -885 14050 -865
rect 13800 -900 14050 -885
rect 13800 -950 13900 -900
rect 13950 -950 14050 -900
rect 14100 -850 14200 -800
rect 14250 -850 14350 -800
rect 14100 -865 14350 -850
rect 14100 -885 14115 -865
rect 14135 -885 14165 -865
rect 14185 -885 14215 -865
rect 14235 -885 14265 -865
rect 14285 -885 14315 -865
rect 14335 -885 14350 -865
rect 14100 -900 14350 -885
rect 14100 -950 14200 -900
rect 14250 -950 14350 -900
rect 14400 -850 14500 -800
rect 14550 -850 14650 -800
rect 14400 -865 14650 -850
rect 14400 -885 14415 -865
rect 14435 -885 14465 -865
rect 14485 -885 14515 -865
rect 14535 -885 14565 -865
rect 14585 -885 14615 -865
rect 14635 -885 14650 -865
rect 14400 -900 14650 -885
rect 14400 -950 14500 -900
rect 14550 -950 14650 -900
rect 14700 -850 14800 -800
rect 14850 -850 14950 -800
rect 14700 -865 14950 -850
rect 14700 -885 14715 -865
rect 14735 -885 14765 -865
rect 14785 -885 14815 -865
rect 14835 -885 14865 -865
rect 14885 -885 14915 -865
rect 14935 -885 14950 -865
rect 14700 -900 14950 -885
rect 14700 -950 14800 -900
rect 14850 -950 14950 -900
rect 15000 -850 15100 -800
rect 15150 -850 15250 -800
rect 15000 -865 15250 -850
rect 15000 -885 15015 -865
rect 15035 -885 15065 -865
rect 15085 -885 15115 -865
rect 15135 -885 15165 -865
rect 15185 -885 15215 -865
rect 15235 -885 15250 -865
rect 15000 -900 15250 -885
rect 15000 -950 15100 -900
rect 15150 -950 15250 -900
rect 15300 -850 15400 -800
rect 15450 -850 15550 -800
rect 15300 -865 15550 -850
rect 15300 -885 15315 -865
rect 15335 -885 15365 -865
rect 15385 -885 15415 -865
rect 15435 -885 15465 -865
rect 15485 -885 15515 -865
rect 15535 -885 15550 -865
rect 15300 -900 15550 -885
rect 15300 -950 15400 -900
rect 15450 -950 15550 -900
rect 15600 -850 15700 -800
rect 15750 -850 15850 -800
rect 15600 -865 15850 -850
rect 15600 -885 15615 -865
rect 15635 -885 15665 -865
rect 15685 -885 15715 -865
rect 15735 -885 15765 -865
rect 15785 -885 15815 -865
rect 15835 -885 15850 -865
rect 15600 -900 15850 -885
rect 15600 -950 15700 -900
rect 15750 -950 15850 -900
rect 15900 -850 16000 -800
rect 16050 -850 16150 -800
rect 15900 -865 16150 -850
rect 15900 -885 15915 -865
rect 15935 -885 15965 -865
rect 15985 -885 16015 -865
rect 16035 -885 16065 -865
rect 16085 -885 16115 -865
rect 16135 -885 16150 -865
rect 15900 -900 16150 -885
rect 15900 -950 16000 -900
rect 16050 -950 16150 -900
rect 16200 -850 16300 -800
rect 16350 -850 16450 -800
rect 16200 -865 16450 -850
rect 16200 -885 16215 -865
rect 16235 -885 16265 -865
rect 16285 -885 16315 -865
rect 16335 -885 16365 -865
rect 16385 -885 16415 -865
rect 16435 -885 16450 -865
rect 16200 -900 16450 -885
rect 16200 -950 16300 -900
rect 16350 -950 16450 -900
rect 16500 -850 16600 -800
rect 16650 -850 16750 -800
rect 16500 -865 16750 -850
rect 16500 -885 16515 -865
rect 16535 -885 16565 -865
rect 16585 -885 16615 -865
rect 16635 -885 16665 -865
rect 16685 -885 16715 -865
rect 16735 -885 16750 -865
rect 16500 -900 16750 -885
rect 16500 -950 16600 -900
rect 16650 -950 16750 -900
rect 16800 -850 16900 -800
rect 16950 -850 17050 -800
rect 16800 -865 17050 -850
rect 16800 -885 16815 -865
rect 16835 -885 16865 -865
rect 16885 -885 16915 -865
rect 16935 -885 16965 -865
rect 16985 -885 17015 -865
rect 17035 -885 17050 -865
rect 16800 -900 17050 -885
rect 16800 -950 16900 -900
rect 16950 -950 17050 -900
rect 17100 -850 17200 -800
rect 17250 -850 17350 -800
rect 17100 -865 17350 -850
rect 17100 -885 17115 -865
rect 17135 -885 17165 -865
rect 17185 -885 17215 -865
rect 17235 -885 17265 -865
rect 17285 -885 17315 -865
rect 17335 -885 17350 -865
rect 17100 -900 17350 -885
rect 17100 -950 17200 -900
rect 17250 -950 17350 -900
rect 17400 -850 17500 -800
rect 17550 -850 17650 -800
rect 17400 -865 17650 -850
rect 17400 -885 17415 -865
rect 17435 -885 17465 -865
rect 17485 -885 17515 -865
rect 17535 -885 17565 -865
rect 17585 -885 17615 -865
rect 17635 -885 17650 -865
rect 17400 -900 17650 -885
rect 17400 -950 17500 -900
rect 17550 -950 17650 -900
rect 17700 -850 17800 -800
rect 17850 -850 17950 -800
rect 17700 -865 17950 -850
rect 17700 -885 17715 -865
rect 17735 -885 17765 -865
rect 17785 -885 17815 -865
rect 17835 -885 17865 -865
rect 17885 -885 17915 -865
rect 17935 -885 17950 -865
rect 17700 -900 17950 -885
rect 17700 -950 17800 -900
rect 17850 -950 17950 -900
rect 18000 -850 18100 -800
rect 18150 -850 18250 -800
rect 18000 -865 18250 -850
rect 18000 -885 18015 -865
rect 18035 -885 18065 -865
rect 18085 -885 18115 -865
rect 18135 -885 18165 -865
rect 18185 -885 18215 -865
rect 18235 -885 18250 -865
rect 18000 -900 18250 -885
rect 18000 -950 18100 -900
rect 18150 -950 18250 -900
rect 18300 -850 18400 -800
rect 18450 -850 18550 -800
rect 18300 -865 18550 -850
rect 18300 -885 18315 -865
rect 18335 -885 18365 -865
rect 18385 -885 18415 -865
rect 18435 -885 18465 -865
rect 18485 -885 18515 -865
rect 18535 -885 18550 -865
rect 18300 -900 18550 -885
rect 18300 -950 18400 -900
rect 18450 -950 18550 -900
rect 18600 -850 18700 -800
rect 18750 -850 18850 -800
rect 18600 -865 18850 -850
rect 18600 -885 18615 -865
rect 18635 -885 18665 -865
rect 18685 -885 18715 -865
rect 18735 -885 18765 -865
rect 18785 -885 18815 -865
rect 18835 -885 18850 -865
rect 18600 -900 18850 -885
rect 18600 -950 18700 -900
rect 18750 -950 18850 -900
rect 18900 -850 19000 -800
rect 19050 -850 19150 -800
rect 18900 -865 19150 -850
rect 18900 -885 18915 -865
rect 18935 -885 18965 -865
rect 18985 -885 19015 -865
rect 19035 -885 19065 -865
rect 19085 -885 19115 -865
rect 19135 -885 19150 -865
rect 18900 -900 19150 -885
rect 18900 -950 19000 -900
rect 19050 -950 19150 -900
rect 19200 -850 19300 -800
rect 19350 -850 19450 -800
rect 19200 -865 19450 -850
rect 19200 -885 19215 -865
rect 19235 -885 19265 -865
rect 19285 -885 19315 -865
rect 19335 -885 19365 -865
rect 19385 -885 19415 -865
rect 19435 -885 19450 -865
rect 19200 -900 19450 -885
rect 19200 -950 19300 -900
rect 19350 -950 19450 -900
rect 19500 -850 19600 -800
rect 19650 -850 19750 -800
rect 19500 -865 19750 -850
rect 19500 -885 19515 -865
rect 19535 -885 19565 -865
rect 19585 -885 19615 -865
rect 19635 -885 19665 -865
rect 19685 -885 19715 -865
rect 19735 -885 19750 -865
rect 19500 -900 19750 -885
rect 19500 -950 19600 -900
rect 19650 -950 19750 -900
rect 19800 -850 19900 -800
rect 19950 -850 20050 -800
rect 19800 -865 20050 -850
rect 19800 -885 19815 -865
rect 19835 -885 19865 -865
rect 19885 -885 19915 -865
rect 19935 -885 19965 -865
rect 19985 -885 20015 -865
rect 20035 -885 20050 -865
rect 19800 -900 20050 -885
rect 19800 -950 19900 -900
rect 19950 -950 20050 -900
rect 20100 -850 20200 -800
rect 20250 -850 20350 -800
rect 20100 -865 20350 -850
rect 20100 -885 20115 -865
rect 20135 -885 20165 -865
rect 20185 -885 20215 -865
rect 20235 -885 20265 -865
rect 20285 -885 20315 -865
rect 20335 -885 20350 -865
rect 20100 -900 20350 -885
rect 20100 -950 20200 -900
rect 20250 -950 20350 -900
rect -600 -1665 -500 -1650
rect -450 -1665 -350 -1650
rect -300 -1665 -200 -1650
rect -150 -1665 -50 -1650
rect 0 -1665 100 -1650
rect 150 -1665 250 -1650
rect 300 -1665 400 -1650
rect 450 -1665 550 -1650
rect 600 -1665 700 -1650
rect 750 -1665 850 -1650
rect 900 -1665 1000 -1650
rect 1050 -1665 1150 -1650
rect 1200 -1665 1300 -1650
rect 1350 -1665 1450 -1650
rect 1500 -1665 1600 -1650
rect 1650 -1665 1750 -1650
rect 1800 -1665 1900 -1650
rect 1950 -1665 2050 -1650
rect 2100 -1665 2200 -1650
rect 2250 -1665 2350 -1650
rect 2400 -1665 2500 -1650
rect 2550 -1665 2650 -1650
rect 2700 -1665 2800 -1650
rect 2850 -1665 2950 -1650
rect 3000 -1665 3100 -1650
rect 3150 -1665 3250 -1650
rect 3300 -1665 3400 -1650
rect 3450 -1665 3550 -1650
rect 3600 -1665 3700 -1650
rect 3750 -1665 3850 -1650
rect 3900 -1665 4000 -1650
rect 4050 -1665 4150 -1650
rect 4200 -1665 4300 -1650
rect 4350 -1665 4450 -1650
rect 4500 -1665 4600 -1650
rect 4650 -1665 4750 -1650
rect 4800 -1665 4900 -1650
rect 4950 -1665 5050 -1650
rect 5100 -1665 5200 -1650
rect 5250 -1665 5350 -1650
rect 5400 -1665 5500 -1650
rect 5550 -1665 5650 -1650
rect 5700 -1665 5800 -1650
rect 5850 -1665 5950 -1650
rect 6000 -1665 6100 -1650
rect 6150 -1665 6250 -1650
rect 6300 -1665 6400 -1650
rect 6450 -1665 6550 -1650
rect 6600 -1665 6700 -1650
rect 6750 -1665 6850 -1650
rect 6900 -1665 7000 -1650
rect 7050 -1665 7150 -1650
rect 7200 -1665 7300 -1650
rect 7350 -1665 7450 -1650
rect 7500 -1665 7600 -1650
rect 7650 -1665 7750 -1650
rect 7800 -1665 7900 -1650
rect 7950 -1665 8050 -1650
rect 8100 -1665 8200 -1650
rect 8250 -1665 8350 -1650
rect 8400 -1665 8500 -1650
rect 8550 -1665 8650 -1650
rect 8700 -1665 8800 -1650
rect 8850 -1665 8950 -1650
rect 9000 -1665 9100 -1650
rect 9150 -1665 9250 -1650
rect 9300 -1665 9400 -1650
rect 9450 -1665 9550 -1650
rect 9600 -1665 9700 -1650
rect 9750 -1665 9850 -1650
rect 9900 -1665 10000 -1650
rect 10050 -1665 10150 -1650
rect 10200 -1665 10300 -1650
rect 10350 -1665 10450 -1650
rect 10500 -1665 10600 -1650
rect 10650 -1665 10750 -1650
rect 10800 -1665 10900 -1650
rect 10950 -1665 11050 -1650
rect 11100 -1665 11200 -1650
rect 11250 -1665 11350 -1650
rect 11400 -1665 11500 -1650
rect 11550 -1665 11650 -1650
rect 11700 -1665 11800 -1650
rect 11850 -1665 11950 -1650
rect 12000 -1665 12100 -1650
rect 12150 -1665 12250 -1650
rect 12300 -1665 12400 -1650
rect 12450 -1665 12550 -1650
rect 12600 -1665 12700 -1650
rect 12750 -1665 12850 -1650
rect 12900 -1665 13000 -1650
rect 13050 -1665 13150 -1650
rect 13200 -1665 13300 -1650
rect 13350 -1665 13450 -1650
rect 13500 -1665 13600 -1650
rect 13650 -1665 13750 -1650
rect 13800 -1665 13900 -1650
rect 13950 -1665 14050 -1650
rect 14100 -1665 14200 -1650
rect 14250 -1665 14350 -1650
rect 14400 -1665 14500 -1650
rect 14550 -1665 14650 -1650
rect 14700 -1665 14800 -1650
rect 14850 -1665 14950 -1650
rect 15000 -1665 15100 -1650
rect 15150 -1665 15250 -1650
rect 15300 -1665 15400 -1650
rect 15450 -1665 15550 -1650
rect 15600 -1665 15700 -1650
rect 15750 -1665 15850 -1650
rect 15900 -1665 16000 -1650
rect 16050 -1665 16150 -1650
rect 16200 -1665 16300 -1650
rect 16350 -1665 16450 -1650
rect 16500 -1665 16600 -1650
rect 16650 -1665 16750 -1650
rect 16800 -1665 16900 -1650
rect 16950 -1665 17050 -1650
rect 17100 -1665 17200 -1650
rect 17250 -1665 17350 -1650
rect 17400 -1665 17500 -1650
rect 17550 -1665 17650 -1650
rect 17700 -1665 17800 -1650
rect 17850 -1665 17950 -1650
rect 18000 -1665 18100 -1650
rect 18150 -1665 18250 -1650
rect 18300 -1665 18400 -1650
rect 18450 -1665 18550 -1650
rect 18600 -1665 18700 -1650
rect 18750 -1665 18850 -1650
rect 18900 -1665 19000 -1650
rect 19050 -1665 19150 -1650
rect 19200 -1665 19300 -1650
rect 19350 -1665 19450 -1650
rect 19500 -1665 19600 -1650
rect 19650 -1665 19750 -1650
rect 19800 -1665 19900 -1650
rect 19950 -1665 20050 -1650
rect 20100 -1665 20200 -1650
rect 20250 -1665 20350 -1650
<< polycont >>
rect -585 4515 -565 4535
rect -535 4515 -515 4535
rect -485 4515 -465 4535
rect -435 4515 -415 4535
rect -385 4515 -365 4535
rect -285 4515 -265 4535
rect -235 4515 -215 4535
rect -185 4515 -165 4535
rect -135 4515 -115 4535
rect -85 4515 -65 4535
rect 15 4515 35 4535
rect 65 4515 85 4535
rect 115 4515 135 4535
rect 165 4515 185 4535
rect 215 4515 235 4535
rect 315 4515 335 4535
rect 365 4515 385 4535
rect 415 4515 435 4535
rect 465 4515 485 4535
rect 515 4515 535 4535
rect 615 4515 635 4535
rect 665 4515 685 4535
rect 715 4515 735 4535
rect 765 4515 785 4535
rect 815 4515 835 4535
rect 915 4515 935 4535
rect 965 4515 985 4535
rect 1015 4515 1035 4535
rect 1065 4515 1085 4535
rect 1115 4515 1135 4535
rect 1215 4515 1235 4535
rect 1265 4515 1285 4535
rect 1315 4515 1335 4535
rect 1365 4515 1385 4535
rect 1415 4515 1435 4535
rect 1515 4515 1535 4535
rect 1565 4515 1585 4535
rect 1615 4515 1635 4535
rect 1665 4515 1685 4535
rect 1715 4515 1735 4535
rect 1815 4515 1835 4535
rect 1865 4515 1885 4535
rect 1915 4515 1935 4535
rect 1965 4515 1985 4535
rect 2015 4515 2035 4535
rect 2115 4515 2135 4535
rect 2165 4515 2185 4535
rect 2215 4515 2235 4535
rect 2265 4515 2285 4535
rect 2315 4515 2335 4535
rect 2415 4515 2435 4535
rect 2465 4515 2485 4535
rect 2515 4515 2535 4535
rect 2565 4515 2585 4535
rect 2615 4515 2635 4535
rect 2715 4515 2735 4535
rect 2765 4515 2785 4535
rect 2815 4515 2835 4535
rect 2865 4515 2885 4535
rect 2915 4515 2935 4535
rect 3015 4515 3035 4535
rect 3065 4515 3085 4535
rect 3115 4515 3135 4535
rect 3165 4515 3185 4535
rect 3215 4515 3235 4535
rect 3315 4515 3335 4535
rect 3365 4515 3385 4535
rect 3415 4515 3435 4535
rect 3465 4515 3485 4535
rect 3515 4515 3535 4535
rect 3615 4515 3635 4535
rect 3665 4515 3685 4535
rect 3715 4515 3735 4535
rect 3765 4515 3785 4535
rect 3815 4515 3835 4535
rect 3915 4515 3935 4535
rect 3965 4515 3985 4535
rect 4015 4515 4035 4535
rect 4065 4515 4085 4535
rect 4115 4515 4135 4535
rect 4215 4515 4235 4535
rect 4265 4515 4285 4535
rect 4315 4515 4335 4535
rect 4365 4515 4385 4535
rect 4415 4515 4435 4535
rect 4515 4515 4535 4535
rect 4565 4515 4585 4535
rect 4615 4515 4635 4535
rect 4665 4515 4685 4535
rect 4715 4515 4735 4535
rect 4815 4515 4835 4535
rect 4865 4515 4885 4535
rect 4915 4515 4935 4535
rect 4965 4515 4985 4535
rect 5015 4515 5035 4535
rect 5115 4515 5135 4535
rect 5165 4515 5185 4535
rect 5215 4515 5235 4535
rect 5265 4515 5285 4535
rect 5315 4515 5335 4535
rect 5415 4515 5435 4535
rect 5465 4515 5485 4535
rect 5515 4515 5535 4535
rect 5565 4515 5585 4535
rect 5615 4515 5635 4535
rect 5715 4515 5735 4535
rect 5765 4515 5785 4535
rect 5815 4515 5835 4535
rect 5865 4515 5885 4535
rect 5915 4515 5935 4535
rect 6015 4515 6035 4535
rect 6065 4515 6085 4535
rect 6115 4515 6135 4535
rect 6165 4515 6185 4535
rect 6215 4515 6235 4535
rect 6315 4515 6335 4535
rect 6365 4515 6385 4535
rect 6415 4515 6435 4535
rect 6465 4515 6485 4535
rect 6515 4515 6535 4535
rect 6615 4515 6635 4535
rect 6665 4515 6685 4535
rect 6715 4515 6735 4535
rect 6765 4515 6785 4535
rect 6815 4515 6835 4535
rect 6915 4515 6935 4535
rect 6965 4515 6985 4535
rect 7015 4515 7035 4535
rect 7065 4515 7085 4535
rect 7115 4515 7135 4535
rect 7215 4515 7235 4535
rect 7265 4515 7285 4535
rect 7315 4515 7335 4535
rect 7365 4515 7385 4535
rect 7415 4515 7435 4535
rect 7515 4515 7535 4535
rect 7565 4515 7585 4535
rect 7615 4515 7635 4535
rect 7665 4515 7685 4535
rect 7715 4515 7735 4535
rect 7815 4515 7835 4535
rect 7865 4515 7885 4535
rect 7915 4515 7935 4535
rect 7965 4515 7985 4535
rect 8015 4515 8035 4535
rect 8115 4515 8135 4535
rect 8165 4515 8185 4535
rect 8215 4515 8235 4535
rect 8265 4515 8285 4535
rect 8315 4515 8335 4535
rect 8415 4515 8435 4535
rect 8465 4515 8485 4535
rect 8515 4515 8535 4535
rect 8565 4515 8585 4535
rect 8615 4515 8635 4535
rect 8715 4515 8735 4535
rect 8765 4515 8785 4535
rect 8815 4515 8835 4535
rect 8865 4515 8885 4535
rect 8915 4515 8935 4535
rect 9015 4515 9035 4535
rect 9065 4515 9085 4535
rect 9115 4515 9135 4535
rect 9165 4515 9185 4535
rect 9215 4515 9235 4535
rect 9315 4515 9335 4535
rect 9365 4515 9385 4535
rect 9415 4515 9435 4535
rect 9465 4515 9485 4535
rect 9515 4515 9535 4535
rect 9615 4515 9635 4535
rect 9665 4515 9685 4535
rect 9715 4515 9735 4535
rect 9765 4515 9785 4535
rect 9815 4515 9835 4535
rect 9915 4515 9935 4535
rect 9965 4515 9985 4535
rect 10015 4515 10035 4535
rect 10065 4515 10085 4535
rect 10115 4515 10135 4535
rect 10215 4515 10235 4535
rect 10265 4515 10285 4535
rect 10315 4515 10335 4535
rect 10365 4515 10385 4535
rect 10415 4515 10435 4535
rect 10515 4515 10535 4535
rect 10565 4515 10585 4535
rect 10615 4515 10635 4535
rect 10665 4515 10685 4535
rect 10715 4515 10735 4535
rect 10815 4515 10835 4535
rect 10865 4515 10885 4535
rect 10915 4515 10935 4535
rect 10965 4515 10985 4535
rect 11015 4515 11035 4535
rect 11115 4515 11135 4535
rect 11165 4515 11185 4535
rect 11215 4515 11235 4535
rect 11265 4515 11285 4535
rect 11315 4515 11335 4535
rect 11415 4515 11435 4535
rect 11465 4515 11485 4535
rect 11515 4515 11535 4535
rect 11565 4515 11585 4535
rect 11615 4515 11635 4535
rect 11715 4515 11735 4535
rect 11765 4515 11785 4535
rect 11815 4515 11835 4535
rect 11865 4515 11885 4535
rect 11915 4515 11935 4535
rect 12015 4515 12035 4535
rect 12065 4515 12085 4535
rect 12115 4515 12135 4535
rect 12165 4515 12185 4535
rect 12215 4515 12235 4535
rect 12315 4515 12335 4535
rect 12365 4515 12385 4535
rect 12415 4515 12435 4535
rect 12465 4515 12485 4535
rect 12515 4515 12535 4535
rect 12615 4515 12635 4535
rect 12665 4515 12685 4535
rect 12715 4515 12735 4535
rect 12765 4515 12785 4535
rect 12815 4515 12835 4535
rect 12915 4515 12935 4535
rect 12965 4515 12985 4535
rect 13015 4515 13035 4535
rect 13065 4515 13085 4535
rect 13115 4515 13135 4535
rect 13215 4515 13235 4535
rect 13265 4515 13285 4535
rect 13315 4515 13335 4535
rect 13365 4515 13385 4535
rect 13415 4515 13435 4535
rect 13515 4515 13535 4535
rect 13565 4515 13585 4535
rect 13615 4515 13635 4535
rect 13665 4515 13685 4535
rect 13715 4515 13735 4535
rect 13815 4515 13835 4535
rect 13865 4515 13885 4535
rect 13915 4515 13935 4535
rect 13965 4515 13985 4535
rect 14015 4515 14035 4535
rect 14115 4515 14135 4535
rect 14165 4515 14185 4535
rect 14215 4515 14235 4535
rect 14265 4515 14285 4535
rect 14315 4515 14335 4535
rect 14415 4515 14435 4535
rect 14465 4515 14485 4535
rect 14515 4515 14535 4535
rect 14565 4515 14585 4535
rect 14615 4515 14635 4535
rect 14715 4515 14735 4535
rect 14765 4515 14785 4535
rect 14815 4515 14835 4535
rect 14865 4515 14885 4535
rect 14915 4515 14935 4535
rect 15015 4515 15035 4535
rect 15065 4515 15085 4535
rect 15115 4515 15135 4535
rect 15165 4515 15185 4535
rect 15215 4515 15235 4535
rect 15315 4515 15335 4535
rect 15365 4515 15385 4535
rect 15415 4515 15435 4535
rect 15465 4515 15485 4535
rect 15515 4515 15535 4535
rect 15615 4515 15635 4535
rect 15665 4515 15685 4535
rect 15715 4515 15735 4535
rect 15765 4515 15785 4535
rect 15815 4515 15835 4535
rect 15915 4515 15935 4535
rect 15965 4515 15985 4535
rect 16015 4515 16035 4535
rect 16065 4515 16085 4535
rect 16115 4515 16135 4535
rect 16215 4515 16235 4535
rect 16265 4515 16285 4535
rect 16315 4515 16335 4535
rect 16365 4515 16385 4535
rect 16415 4515 16435 4535
rect 16515 4515 16535 4535
rect 16565 4515 16585 4535
rect 16615 4515 16635 4535
rect 16665 4515 16685 4535
rect 16715 4515 16735 4535
rect 16815 4515 16835 4535
rect 16865 4515 16885 4535
rect 16915 4515 16935 4535
rect 16965 4515 16985 4535
rect 17015 4515 17035 4535
rect 17115 4515 17135 4535
rect 17165 4515 17185 4535
rect 17215 4515 17235 4535
rect 17265 4515 17285 4535
rect 17315 4515 17335 4535
rect 17415 4515 17435 4535
rect 17465 4515 17485 4535
rect 17515 4515 17535 4535
rect 17565 4515 17585 4535
rect 17615 4515 17635 4535
rect 17715 4515 17735 4535
rect 17765 4515 17785 4535
rect 17815 4515 17835 4535
rect 17865 4515 17885 4535
rect 17915 4515 17935 4535
rect 18015 4515 18035 4535
rect 18065 4515 18085 4535
rect 18115 4515 18135 4535
rect 18165 4515 18185 4535
rect 18215 4515 18235 4535
rect 18315 4515 18335 4535
rect 18365 4515 18385 4535
rect 18415 4515 18435 4535
rect 18465 4515 18485 4535
rect 18515 4515 18535 4535
rect 18615 4515 18635 4535
rect 18665 4515 18685 4535
rect 18715 4515 18735 4535
rect 18765 4515 18785 4535
rect 18815 4515 18835 4535
rect 18915 4515 18935 4535
rect 18965 4515 18985 4535
rect 19015 4515 19035 4535
rect 19065 4515 19085 4535
rect 19115 4515 19135 4535
rect 19215 4515 19235 4535
rect 19265 4515 19285 4535
rect 19315 4515 19335 4535
rect 19365 4515 19385 4535
rect 19415 4515 19435 4535
rect 19515 4515 19535 4535
rect 19565 4515 19585 4535
rect 19615 4515 19635 4535
rect 19665 4515 19685 4535
rect 19715 4515 19735 4535
rect 19815 4515 19835 4535
rect 19865 4515 19885 4535
rect 19915 4515 19935 4535
rect 19965 4515 19985 4535
rect 20015 4515 20035 4535
rect 20115 4515 20135 4535
rect 20165 4515 20185 4535
rect 20215 4515 20235 4535
rect 20265 4515 20285 4535
rect 20315 4515 20335 4535
rect -585 3215 -565 3235
rect -535 3215 -515 3235
rect -485 3215 -465 3235
rect -435 3215 -415 3235
rect -385 3215 -365 3235
rect -285 3215 -265 3235
rect -235 3215 -215 3235
rect -185 3215 -165 3235
rect -135 3215 -115 3235
rect -85 3215 -65 3235
rect 15 3215 35 3235
rect 65 3215 85 3235
rect 115 3215 135 3235
rect 165 3215 185 3235
rect 215 3215 235 3235
rect 315 3215 335 3235
rect 365 3215 385 3235
rect 415 3215 435 3235
rect 465 3215 485 3235
rect 515 3215 535 3235
rect 615 3215 635 3235
rect 665 3215 685 3235
rect 715 3215 735 3235
rect 765 3215 785 3235
rect 815 3215 835 3235
rect 915 3215 935 3235
rect 965 3215 985 3235
rect 1015 3215 1035 3235
rect 1065 3215 1085 3235
rect 1115 3215 1135 3235
rect 1215 3215 1235 3235
rect 1265 3215 1285 3235
rect 1315 3215 1335 3235
rect 1365 3215 1385 3235
rect 1415 3215 1435 3235
rect 1515 3215 1535 3235
rect 1565 3215 1585 3235
rect 1615 3215 1635 3235
rect 1665 3215 1685 3235
rect 1715 3215 1735 3235
rect 1815 3215 1835 3235
rect 1865 3215 1885 3235
rect 1915 3215 1935 3235
rect 1965 3215 1985 3235
rect 2015 3215 2035 3235
rect 2115 3215 2135 3235
rect 2165 3215 2185 3235
rect 2215 3215 2235 3235
rect 2265 3215 2285 3235
rect 2315 3215 2335 3235
rect 2415 3215 2435 3235
rect 2465 3215 2485 3235
rect 2515 3215 2535 3235
rect 2565 3215 2585 3235
rect 2615 3215 2635 3235
rect 2715 3215 2735 3235
rect 2765 3215 2785 3235
rect 2815 3215 2835 3235
rect 2865 3215 2885 3235
rect 2915 3215 2935 3235
rect 3015 3215 3035 3235
rect 3065 3215 3085 3235
rect 3115 3215 3135 3235
rect 3165 3215 3185 3235
rect 3215 3215 3235 3235
rect 3315 3215 3335 3235
rect 3365 3215 3385 3235
rect 3415 3215 3435 3235
rect 3465 3215 3485 3235
rect 3515 3215 3535 3235
rect 3615 3215 3635 3235
rect 3665 3215 3685 3235
rect 3715 3215 3735 3235
rect 3765 3215 3785 3235
rect 3815 3215 3835 3235
rect 3915 3215 3935 3235
rect 3965 3215 3985 3235
rect 4015 3215 4035 3235
rect 4065 3215 4085 3235
rect 4115 3215 4135 3235
rect 4215 3215 4235 3235
rect 4265 3215 4285 3235
rect 4315 3215 4335 3235
rect 4365 3215 4385 3235
rect 4415 3215 4435 3235
rect 4515 3215 4535 3235
rect 4565 3215 4585 3235
rect 4615 3215 4635 3235
rect 4665 3215 4685 3235
rect 4715 3215 4735 3235
rect 4815 3215 4835 3235
rect 4865 3215 4885 3235
rect 4915 3215 4935 3235
rect 4965 3215 4985 3235
rect 5015 3215 5035 3235
rect 5115 3215 5135 3235
rect 5165 3215 5185 3235
rect 5215 3215 5235 3235
rect 5265 3215 5285 3235
rect 5315 3215 5335 3235
rect 5415 3215 5435 3235
rect 5465 3215 5485 3235
rect 5515 3215 5535 3235
rect 5565 3215 5585 3235
rect 5615 3215 5635 3235
rect 5715 3215 5735 3235
rect 5765 3215 5785 3235
rect 5815 3215 5835 3235
rect 5865 3215 5885 3235
rect 5915 3215 5935 3235
rect 6015 3215 6035 3235
rect 6065 3215 6085 3235
rect 6115 3215 6135 3235
rect 6165 3215 6185 3235
rect 6215 3215 6235 3235
rect 6315 3215 6335 3235
rect 6365 3215 6385 3235
rect 6415 3215 6435 3235
rect 6465 3215 6485 3235
rect 6515 3215 6535 3235
rect 6615 3215 6635 3235
rect 6665 3215 6685 3235
rect 6715 3215 6735 3235
rect 6765 3215 6785 3235
rect 6815 3215 6835 3235
rect 6915 3215 6935 3235
rect 6965 3215 6985 3235
rect 7015 3215 7035 3235
rect 7065 3215 7085 3235
rect 7115 3215 7135 3235
rect 7215 3215 7235 3235
rect 7265 3215 7285 3235
rect 7315 3215 7335 3235
rect 7365 3215 7385 3235
rect 7415 3215 7435 3235
rect 7515 3215 7535 3235
rect 7565 3215 7585 3235
rect 7615 3215 7635 3235
rect 7665 3215 7685 3235
rect 7715 3215 7735 3235
rect 7815 3215 7835 3235
rect 7865 3215 7885 3235
rect 7915 3215 7935 3235
rect 7965 3215 7985 3235
rect 8015 3215 8035 3235
rect 8115 3215 8135 3235
rect 8165 3215 8185 3235
rect 8215 3215 8235 3235
rect 8265 3215 8285 3235
rect 8315 3215 8335 3235
rect 8415 3215 8435 3235
rect 8465 3215 8485 3235
rect 8515 3215 8535 3235
rect 8565 3215 8585 3235
rect 8615 3215 8635 3235
rect 8715 3215 8735 3235
rect 8765 3215 8785 3235
rect 8815 3215 8835 3235
rect 8865 3215 8885 3235
rect 8915 3215 8935 3235
rect 9015 3215 9035 3235
rect 9065 3215 9085 3235
rect 9115 3215 9135 3235
rect 9165 3215 9185 3235
rect 9215 3215 9235 3235
rect 9315 3215 9335 3235
rect 9365 3215 9385 3235
rect 9415 3215 9435 3235
rect 9465 3215 9485 3235
rect 9515 3215 9535 3235
rect 9615 3215 9635 3235
rect 9665 3215 9685 3235
rect 9715 3215 9735 3235
rect 9765 3215 9785 3235
rect 9815 3215 9835 3235
rect 9915 3215 9935 3235
rect 9965 3215 9985 3235
rect 10015 3215 10035 3235
rect 10065 3215 10085 3235
rect 10115 3215 10135 3235
rect 10215 3215 10235 3235
rect 10265 3215 10285 3235
rect 10315 3215 10335 3235
rect 10365 3215 10385 3235
rect 10415 3215 10435 3235
rect 10515 3215 10535 3235
rect 10565 3215 10585 3235
rect 10615 3215 10635 3235
rect 10665 3215 10685 3235
rect 10715 3215 10735 3235
rect 10815 3215 10835 3235
rect 10865 3215 10885 3235
rect 10915 3215 10935 3235
rect 10965 3215 10985 3235
rect 11015 3215 11035 3235
rect 11115 3215 11135 3235
rect 11165 3215 11185 3235
rect 11215 3215 11235 3235
rect 11265 3215 11285 3235
rect 11315 3215 11335 3235
rect 11415 3215 11435 3235
rect 11465 3215 11485 3235
rect 11515 3215 11535 3235
rect 11565 3215 11585 3235
rect 11615 3215 11635 3235
rect 11715 3215 11735 3235
rect 11765 3215 11785 3235
rect 11815 3215 11835 3235
rect 11865 3215 11885 3235
rect 11915 3215 11935 3235
rect 12015 3215 12035 3235
rect 12065 3215 12085 3235
rect 12115 3215 12135 3235
rect 12165 3215 12185 3235
rect 12215 3215 12235 3235
rect 12315 3215 12335 3235
rect 12365 3215 12385 3235
rect 12415 3215 12435 3235
rect 12465 3215 12485 3235
rect 12515 3215 12535 3235
rect 12615 3215 12635 3235
rect 12665 3215 12685 3235
rect 12715 3215 12735 3235
rect 12765 3215 12785 3235
rect 12815 3215 12835 3235
rect 12915 3215 12935 3235
rect 12965 3215 12985 3235
rect 13015 3215 13035 3235
rect 13065 3215 13085 3235
rect 13115 3215 13135 3235
rect 13215 3215 13235 3235
rect 13265 3215 13285 3235
rect 13315 3215 13335 3235
rect 13365 3215 13385 3235
rect 13415 3215 13435 3235
rect 13515 3215 13535 3235
rect 13565 3215 13585 3235
rect 13615 3215 13635 3235
rect 13665 3215 13685 3235
rect 13715 3215 13735 3235
rect 13815 3215 13835 3235
rect 13865 3215 13885 3235
rect 13915 3215 13935 3235
rect 13965 3215 13985 3235
rect 14015 3215 14035 3235
rect 14115 3215 14135 3235
rect 14165 3215 14185 3235
rect 14215 3215 14235 3235
rect 14265 3215 14285 3235
rect 14315 3215 14335 3235
rect 14415 3215 14435 3235
rect 14465 3215 14485 3235
rect 14515 3215 14535 3235
rect 14565 3215 14585 3235
rect 14615 3215 14635 3235
rect 14715 3215 14735 3235
rect 14765 3215 14785 3235
rect 14815 3215 14835 3235
rect 14865 3215 14885 3235
rect 14915 3215 14935 3235
rect 15015 3215 15035 3235
rect 15065 3215 15085 3235
rect 15115 3215 15135 3235
rect 15165 3215 15185 3235
rect 15215 3215 15235 3235
rect 15315 3215 15335 3235
rect 15365 3215 15385 3235
rect 15415 3215 15435 3235
rect 15465 3215 15485 3235
rect 15515 3215 15535 3235
rect 15615 3215 15635 3235
rect 15665 3215 15685 3235
rect 15715 3215 15735 3235
rect 15765 3215 15785 3235
rect 15815 3215 15835 3235
rect 15915 3215 15935 3235
rect 15965 3215 15985 3235
rect 16015 3215 16035 3235
rect 16065 3215 16085 3235
rect 16115 3215 16135 3235
rect 16215 3215 16235 3235
rect 16265 3215 16285 3235
rect 16315 3215 16335 3235
rect 16365 3215 16385 3235
rect 16415 3215 16435 3235
rect 16515 3215 16535 3235
rect 16565 3215 16585 3235
rect 16615 3215 16635 3235
rect 16665 3215 16685 3235
rect 16715 3215 16735 3235
rect 16815 3215 16835 3235
rect 16865 3215 16885 3235
rect 16915 3215 16935 3235
rect 16965 3215 16985 3235
rect 17015 3215 17035 3235
rect 17115 3215 17135 3235
rect 17165 3215 17185 3235
rect 17215 3215 17235 3235
rect 17265 3215 17285 3235
rect 17315 3215 17335 3235
rect 17415 3215 17435 3235
rect 17465 3215 17485 3235
rect 17515 3215 17535 3235
rect 17565 3215 17585 3235
rect 17615 3215 17635 3235
rect 17715 3215 17735 3235
rect 17765 3215 17785 3235
rect 17815 3215 17835 3235
rect 17865 3215 17885 3235
rect 17915 3215 17935 3235
rect 18015 3215 18035 3235
rect 18065 3215 18085 3235
rect 18115 3215 18135 3235
rect 18165 3215 18185 3235
rect 18215 3215 18235 3235
rect 18315 3215 18335 3235
rect 18365 3215 18385 3235
rect 18415 3215 18435 3235
rect 18465 3215 18485 3235
rect 18515 3215 18535 3235
rect 18615 3215 18635 3235
rect 18665 3215 18685 3235
rect 18715 3215 18735 3235
rect 18765 3215 18785 3235
rect 18815 3215 18835 3235
rect 18915 3215 18935 3235
rect 18965 3215 18985 3235
rect 19015 3215 19035 3235
rect 19065 3215 19085 3235
rect 19115 3215 19135 3235
rect 19215 3215 19235 3235
rect 19265 3215 19285 3235
rect 19315 3215 19335 3235
rect 19365 3215 19385 3235
rect 19415 3215 19435 3235
rect 19515 3215 19535 3235
rect 19565 3215 19585 3235
rect 19615 3215 19635 3235
rect 19665 3215 19685 3235
rect 19715 3215 19735 3235
rect 19815 3215 19835 3235
rect 19865 3215 19885 3235
rect 19915 3215 19935 3235
rect 19965 3215 19985 3235
rect 20015 3215 20035 3235
rect 20115 3215 20135 3235
rect 20165 3215 20185 3235
rect 20215 3215 20235 3235
rect 20265 3215 20285 3235
rect 20315 3215 20335 3235
rect -585 815 -565 835
rect -535 815 -515 835
rect -485 815 -465 835
rect -435 815 -415 835
rect -385 815 -365 835
rect -285 815 -265 835
rect -235 815 -215 835
rect -185 815 -165 835
rect -135 815 -115 835
rect -85 815 -65 835
rect 15 815 35 835
rect 65 815 85 835
rect 115 815 135 835
rect 165 815 185 835
rect 215 815 235 835
rect 315 815 335 835
rect 365 815 385 835
rect 415 815 435 835
rect 465 815 485 835
rect 515 815 535 835
rect 615 815 635 835
rect 665 815 685 835
rect 715 815 735 835
rect 765 815 785 835
rect 815 815 835 835
rect 915 815 935 835
rect 965 815 985 835
rect 1015 815 1035 835
rect 1065 815 1085 835
rect 1115 815 1135 835
rect 1215 815 1235 835
rect 1265 815 1285 835
rect 1315 815 1335 835
rect 1365 815 1385 835
rect 1415 815 1435 835
rect 1515 815 1535 835
rect 1565 815 1585 835
rect 1615 815 1635 835
rect 1665 815 1685 835
rect 1715 815 1735 835
rect 1815 815 1835 835
rect 1865 815 1885 835
rect 1915 815 1935 835
rect 1965 815 1985 835
rect 2015 815 2035 835
rect 2115 815 2135 835
rect 2165 815 2185 835
rect 2215 815 2235 835
rect 2265 815 2285 835
rect 2315 815 2335 835
rect 2415 815 2435 835
rect 2465 815 2485 835
rect 2515 815 2535 835
rect 2565 815 2585 835
rect 2615 815 2635 835
rect 2715 815 2735 835
rect 2765 815 2785 835
rect 2815 815 2835 835
rect 2865 815 2885 835
rect 2915 815 2935 835
rect 3015 815 3035 835
rect 3065 815 3085 835
rect 3115 815 3135 835
rect 3165 815 3185 835
rect 3215 815 3235 835
rect 3315 815 3335 835
rect 3365 815 3385 835
rect 3415 815 3435 835
rect 3465 815 3485 835
rect 3515 815 3535 835
rect 3615 815 3635 835
rect 3665 815 3685 835
rect 3715 815 3735 835
rect 3765 815 3785 835
rect 3815 815 3835 835
rect 3915 815 3935 835
rect 3965 815 3985 835
rect 4015 815 4035 835
rect 4065 815 4085 835
rect 4115 815 4135 835
rect 4215 815 4235 835
rect 4265 815 4285 835
rect 4315 815 4335 835
rect 4365 815 4385 835
rect 4415 815 4435 835
rect 4515 815 4535 835
rect 4565 815 4585 835
rect 4615 815 4635 835
rect 4665 815 4685 835
rect 4715 815 4735 835
rect 4815 815 4835 835
rect 4865 815 4885 835
rect 4915 815 4935 835
rect 4965 815 4985 835
rect 5015 815 5035 835
rect 5115 815 5135 835
rect 5165 815 5185 835
rect 5215 815 5235 835
rect 5265 815 5285 835
rect 5315 815 5335 835
rect 5415 815 5435 835
rect 5465 815 5485 835
rect 5515 815 5535 835
rect 5565 815 5585 835
rect 5615 815 5635 835
rect 5715 815 5735 835
rect 5765 815 5785 835
rect 5815 815 5835 835
rect 5865 815 5885 835
rect 5915 815 5935 835
rect 6015 815 6035 835
rect 6065 815 6085 835
rect 6115 815 6135 835
rect 6165 815 6185 835
rect 6215 815 6235 835
rect 6315 815 6335 835
rect 6365 815 6385 835
rect 6415 815 6435 835
rect 6465 815 6485 835
rect 6515 815 6535 835
rect 6615 815 6635 835
rect 6665 815 6685 835
rect 6715 815 6735 835
rect 6765 815 6785 835
rect 6815 815 6835 835
rect 6915 815 6935 835
rect 6965 815 6985 835
rect 7015 815 7035 835
rect 7065 815 7085 835
rect 7115 815 7135 835
rect 7215 815 7235 835
rect 7265 815 7285 835
rect 7315 815 7335 835
rect 7365 815 7385 835
rect 7415 815 7435 835
rect 7515 815 7535 835
rect 7565 815 7585 835
rect 7615 815 7635 835
rect 7665 815 7685 835
rect 7715 815 7735 835
rect 7815 815 7835 835
rect 7865 815 7885 835
rect 7915 815 7935 835
rect 7965 815 7985 835
rect 8015 815 8035 835
rect 8115 815 8135 835
rect 8165 815 8185 835
rect 8215 815 8235 835
rect 8265 815 8285 835
rect 8315 815 8335 835
rect 8415 815 8435 835
rect 8465 815 8485 835
rect 8515 815 8535 835
rect 8565 815 8585 835
rect 8615 815 8635 835
rect 8715 815 8735 835
rect 8765 815 8785 835
rect 8815 815 8835 835
rect 8865 815 8885 835
rect 8915 815 8935 835
rect 9015 815 9035 835
rect 9065 815 9085 835
rect 9115 815 9135 835
rect 9165 815 9185 835
rect 9215 815 9235 835
rect 9315 815 9335 835
rect 9365 815 9385 835
rect 9415 815 9435 835
rect 9465 815 9485 835
rect 9515 815 9535 835
rect 9615 815 9635 835
rect 9665 815 9685 835
rect 9715 815 9735 835
rect 9765 815 9785 835
rect 9815 815 9835 835
rect 9915 815 9935 835
rect 9965 815 9985 835
rect 10015 815 10035 835
rect 10065 815 10085 835
rect 10115 815 10135 835
rect 10215 815 10235 835
rect 10265 815 10285 835
rect 10315 815 10335 835
rect 10365 815 10385 835
rect 10415 815 10435 835
rect 10515 815 10535 835
rect 10565 815 10585 835
rect 10615 815 10635 835
rect 10665 815 10685 835
rect 10715 815 10735 835
rect 10815 815 10835 835
rect 10865 815 10885 835
rect 10915 815 10935 835
rect 10965 815 10985 835
rect 11015 815 11035 835
rect 11115 815 11135 835
rect 11165 815 11185 835
rect 11215 815 11235 835
rect 11265 815 11285 835
rect 11315 815 11335 835
rect 11415 815 11435 835
rect 11465 815 11485 835
rect 11515 815 11535 835
rect 11565 815 11585 835
rect 11615 815 11635 835
rect 11715 815 11735 835
rect 11765 815 11785 835
rect 11815 815 11835 835
rect 11865 815 11885 835
rect 11915 815 11935 835
rect 12015 815 12035 835
rect 12065 815 12085 835
rect 12115 815 12135 835
rect 12165 815 12185 835
rect 12215 815 12235 835
rect 12315 815 12335 835
rect 12365 815 12385 835
rect 12415 815 12435 835
rect 12465 815 12485 835
rect 12515 815 12535 835
rect 12615 815 12635 835
rect 12665 815 12685 835
rect 12715 815 12735 835
rect 12765 815 12785 835
rect 12815 815 12835 835
rect 12915 815 12935 835
rect 12965 815 12985 835
rect 13015 815 13035 835
rect 13065 815 13085 835
rect 13115 815 13135 835
rect 13215 815 13235 835
rect 13265 815 13285 835
rect 13315 815 13335 835
rect 13365 815 13385 835
rect 13415 815 13435 835
rect 13515 815 13535 835
rect 13565 815 13585 835
rect 13615 815 13635 835
rect 13665 815 13685 835
rect 13715 815 13735 835
rect 13815 815 13835 835
rect 13865 815 13885 835
rect 13915 815 13935 835
rect 13965 815 13985 835
rect 14015 815 14035 835
rect 14115 815 14135 835
rect 14165 815 14185 835
rect 14215 815 14235 835
rect 14265 815 14285 835
rect 14315 815 14335 835
rect 14415 815 14435 835
rect 14465 815 14485 835
rect 14515 815 14535 835
rect 14565 815 14585 835
rect 14615 815 14635 835
rect 14715 815 14735 835
rect 14765 815 14785 835
rect 14815 815 14835 835
rect 14865 815 14885 835
rect 14915 815 14935 835
rect 15015 815 15035 835
rect 15065 815 15085 835
rect 15115 815 15135 835
rect 15165 815 15185 835
rect 15215 815 15235 835
rect 15315 815 15335 835
rect 15365 815 15385 835
rect 15415 815 15435 835
rect 15465 815 15485 835
rect 15515 815 15535 835
rect 15615 815 15635 835
rect 15665 815 15685 835
rect 15715 815 15735 835
rect 15765 815 15785 835
rect 15815 815 15835 835
rect 15915 815 15935 835
rect 15965 815 15985 835
rect 16015 815 16035 835
rect 16065 815 16085 835
rect 16115 815 16135 835
rect 16215 815 16235 835
rect 16265 815 16285 835
rect 16315 815 16335 835
rect 16365 815 16385 835
rect 16415 815 16435 835
rect 16515 815 16535 835
rect 16565 815 16585 835
rect 16615 815 16635 835
rect 16665 815 16685 835
rect 16715 815 16735 835
rect 16815 815 16835 835
rect 16865 815 16885 835
rect 16915 815 16935 835
rect 16965 815 16985 835
rect 17015 815 17035 835
rect 17115 815 17135 835
rect 17165 815 17185 835
rect 17215 815 17235 835
rect 17265 815 17285 835
rect 17315 815 17335 835
rect 17415 815 17435 835
rect 17465 815 17485 835
rect 17515 815 17535 835
rect 17565 815 17585 835
rect 17615 815 17635 835
rect 17715 815 17735 835
rect 17765 815 17785 835
rect 17815 815 17835 835
rect 17865 815 17885 835
rect 17915 815 17935 835
rect 18015 815 18035 835
rect 18065 815 18085 835
rect 18115 815 18135 835
rect 18165 815 18185 835
rect 18215 815 18235 835
rect 18315 815 18335 835
rect 18365 815 18385 835
rect 18415 815 18435 835
rect 18465 815 18485 835
rect 18515 815 18535 835
rect 18615 815 18635 835
rect 18665 815 18685 835
rect 18715 815 18735 835
rect 18765 815 18785 835
rect 18815 815 18835 835
rect 18915 815 18935 835
rect 18965 815 18985 835
rect 19015 815 19035 835
rect 19065 815 19085 835
rect 19115 815 19135 835
rect 19215 815 19235 835
rect 19265 815 19285 835
rect 19315 815 19335 835
rect 19365 815 19385 835
rect 19415 815 19435 835
rect 19515 815 19535 835
rect 19565 815 19585 835
rect 19615 815 19635 835
rect 19665 815 19685 835
rect 19715 815 19735 835
rect 19815 815 19835 835
rect 19865 815 19885 835
rect 19915 815 19935 835
rect 19965 815 19985 835
rect 20015 815 20035 835
rect 20115 815 20135 835
rect 20165 815 20185 835
rect 20215 815 20235 835
rect 20265 815 20285 835
rect 20315 815 20335 835
rect -585 -885 -565 -865
rect -535 -885 -515 -865
rect -485 -885 -465 -865
rect -435 -885 -415 -865
rect -385 -885 -365 -865
rect -285 -885 -265 -865
rect -235 -885 -215 -865
rect -185 -885 -165 -865
rect -135 -885 -115 -865
rect -85 -885 -65 -865
rect 15 -885 35 -865
rect 65 -885 85 -865
rect 115 -885 135 -865
rect 165 -885 185 -865
rect 215 -885 235 -865
rect 315 -885 335 -865
rect 365 -885 385 -865
rect 415 -885 435 -865
rect 465 -885 485 -865
rect 515 -885 535 -865
rect 615 -885 635 -865
rect 665 -885 685 -865
rect 715 -885 735 -865
rect 765 -885 785 -865
rect 815 -885 835 -865
rect 915 -885 935 -865
rect 965 -885 985 -865
rect 1015 -885 1035 -865
rect 1065 -885 1085 -865
rect 1115 -885 1135 -865
rect 1215 -885 1235 -865
rect 1265 -885 1285 -865
rect 1315 -885 1335 -865
rect 1365 -885 1385 -865
rect 1415 -885 1435 -865
rect 1515 -885 1535 -865
rect 1565 -885 1585 -865
rect 1615 -885 1635 -865
rect 1665 -885 1685 -865
rect 1715 -885 1735 -865
rect 1815 -885 1835 -865
rect 1865 -885 1885 -865
rect 1915 -885 1935 -865
rect 1965 -885 1985 -865
rect 2015 -885 2035 -865
rect 2115 -885 2135 -865
rect 2165 -885 2185 -865
rect 2215 -885 2235 -865
rect 2265 -885 2285 -865
rect 2315 -885 2335 -865
rect 2415 -885 2435 -865
rect 2465 -885 2485 -865
rect 2515 -885 2535 -865
rect 2565 -885 2585 -865
rect 2615 -885 2635 -865
rect 2715 -885 2735 -865
rect 2765 -885 2785 -865
rect 2815 -885 2835 -865
rect 2865 -885 2885 -865
rect 2915 -885 2935 -865
rect 3015 -885 3035 -865
rect 3065 -885 3085 -865
rect 3115 -885 3135 -865
rect 3165 -885 3185 -865
rect 3215 -885 3235 -865
rect 3315 -885 3335 -865
rect 3365 -885 3385 -865
rect 3415 -885 3435 -865
rect 3465 -885 3485 -865
rect 3515 -885 3535 -865
rect 3615 -885 3635 -865
rect 3665 -885 3685 -865
rect 3715 -885 3735 -865
rect 3765 -885 3785 -865
rect 3815 -885 3835 -865
rect 3915 -885 3935 -865
rect 3965 -885 3985 -865
rect 4015 -885 4035 -865
rect 4065 -885 4085 -865
rect 4115 -885 4135 -865
rect 4215 -885 4235 -865
rect 4265 -885 4285 -865
rect 4315 -885 4335 -865
rect 4365 -885 4385 -865
rect 4415 -885 4435 -865
rect 4515 -885 4535 -865
rect 4565 -885 4585 -865
rect 4615 -885 4635 -865
rect 4665 -885 4685 -865
rect 4715 -885 4735 -865
rect 4815 -885 4835 -865
rect 4865 -885 4885 -865
rect 4915 -885 4935 -865
rect 4965 -885 4985 -865
rect 5015 -885 5035 -865
rect 5115 -885 5135 -865
rect 5165 -885 5185 -865
rect 5215 -885 5235 -865
rect 5265 -885 5285 -865
rect 5315 -885 5335 -865
rect 5415 -885 5435 -865
rect 5465 -885 5485 -865
rect 5515 -885 5535 -865
rect 5565 -885 5585 -865
rect 5615 -885 5635 -865
rect 5715 -885 5735 -865
rect 5765 -885 5785 -865
rect 5815 -885 5835 -865
rect 5865 -885 5885 -865
rect 5915 -885 5935 -865
rect 6015 -885 6035 -865
rect 6065 -885 6085 -865
rect 6115 -885 6135 -865
rect 6165 -885 6185 -865
rect 6215 -885 6235 -865
rect 6315 -885 6335 -865
rect 6365 -885 6385 -865
rect 6415 -885 6435 -865
rect 6465 -885 6485 -865
rect 6515 -885 6535 -865
rect 6615 -885 6635 -865
rect 6665 -885 6685 -865
rect 6715 -885 6735 -865
rect 6765 -885 6785 -865
rect 6815 -885 6835 -865
rect 6915 -885 6935 -865
rect 6965 -885 6985 -865
rect 7015 -885 7035 -865
rect 7065 -885 7085 -865
rect 7115 -885 7135 -865
rect 7215 -885 7235 -865
rect 7265 -885 7285 -865
rect 7315 -885 7335 -865
rect 7365 -885 7385 -865
rect 7415 -885 7435 -865
rect 7515 -885 7535 -865
rect 7565 -885 7585 -865
rect 7615 -885 7635 -865
rect 7665 -885 7685 -865
rect 7715 -885 7735 -865
rect 7815 -885 7835 -865
rect 7865 -885 7885 -865
rect 7915 -885 7935 -865
rect 7965 -885 7985 -865
rect 8015 -885 8035 -865
rect 8115 -885 8135 -865
rect 8165 -885 8185 -865
rect 8215 -885 8235 -865
rect 8265 -885 8285 -865
rect 8315 -885 8335 -865
rect 8415 -885 8435 -865
rect 8465 -885 8485 -865
rect 8515 -885 8535 -865
rect 8565 -885 8585 -865
rect 8615 -885 8635 -865
rect 8715 -885 8735 -865
rect 8765 -885 8785 -865
rect 8815 -885 8835 -865
rect 8865 -885 8885 -865
rect 8915 -885 8935 -865
rect 9015 -885 9035 -865
rect 9065 -885 9085 -865
rect 9115 -885 9135 -865
rect 9165 -885 9185 -865
rect 9215 -885 9235 -865
rect 9315 -885 9335 -865
rect 9365 -885 9385 -865
rect 9415 -885 9435 -865
rect 9465 -885 9485 -865
rect 9515 -885 9535 -865
rect 9615 -885 9635 -865
rect 9665 -885 9685 -865
rect 9715 -885 9735 -865
rect 9765 -885 9785 -865
rect 9815 -885 9835 -865
rect 9915 -885 9935 -865
rect 9965 -885 9985 -865
rect 10015 -885 10035 -865
rect 10065 -885 10085 -865
rect 10115 -885 10135 -865
rect 10215 -885 10235 -865
rect 10265 -885 10285 -865
rect 10315 -885 10335 -865
rect 10365 -885 10385 -865
rect 10415 -885 10435 -865
rect 10515 -885 10535 -865
rect 10565 -885 10585 -865
rect 10615 -885 10635 -865
rect 10665 -885 10685 -865
rect 10715 -885 10735 -865
rect 10815 -885 10835 -865
rect 10865 -885 10885 -865
rect 10915 -885 10935 -865
rect 10965 -885 10985 -865
rect 11015 -885 11035 -865
rect 11115 -885 11135 -865
rect 11165 -885 11185 -865
rect 11215 -885 11235 -865
rect 11265 -885 11285 -865
rect 11315 -885 11335 -865
rect 11415 -885 11435 -865
rect 11465 -885 11485 -865
rect 11515 -885 11535 -865
rect 11565 -885 11585 -865
rect 11615 -885 11635 -865
rect 11715 -885 11735 -865
rect 11765 -885 11785 -865
rect 11815 -885 11835 -865
rect 11865 -885 11885 -865
rect 11915 -885 11935 -865
rect 12015 -885 12035 -865
rect 12065 -885 12085 -865
rect 12115 -885 12135 -865
rect 12165 -885 12185 -865
rect 12215 -885 12235 -865
rect 12315 -885 12335 -865
rect 12365 -885 12385 -865
rect 12415 -885 12435 -865
rect 12465 -885 12485 -865
rect 12515 -885 12535 -865
rect 12615 -885 12635 -865
rect 12665 -885 12685 -865
rect 12715 -885 12735 -865
rect 12765 -885 12785 -865
rect 12815 -885 12835 -865
rect 12915 -885 12935 -865
rect 12965 -885 12985 -865
rect 13015 -885 13035 -865
rect 13065 -885 13085 -865
rect 13115 -885 13135 -865
rect 13215 -885 13235 -865
rect 13265 -885 13285 -865
rect 13315 -885 13335 -865
rect 13365 -885 13385 -865
rect 13415 -885 13435 -865
rect 13515 -885 13535 -865
rect 13565 -885 13585 -865
rect 13615 -885 13635 -865
rect 13665 -885 13685 -865
rect 13715 -885 13735 -865
rect 13815 -885 13835 -865
rect 13865 -885 13885 -865
rect 13915 -885 13935 -865
rect 13965 -885 13985 -865
rect 14015 -885 14035 -865
rect 14115 -885 14135 -865
rect 14165 -885 14185 -865
rect 14215 -885 14235 -865
rect 14265 -885 14285 -865
rect 14315 -885 14335 -865
rect 14415 -885 14435 -865
rect 14465 -885 14485 -865
rect 14515 -885 14535 -865
rect 14565 -885 14585 -865
rect 14615 -885 14635 -865
rect 14715 -885 14735 -865
rect 14765 -885 14785 -865
rect 14815 -885 14835 -865
rect 14865 -885 14885 -865
rect 14915 -885 14935 -865
rect 15015 -885 15035 -865
rect 15065 -885 15085 -865
rect 15115 -885 15135 -865
rect 15165 -885 15185 -865
rect 15215 -885 15235 -865
rect 15315 -885 15335 -865
rect 15365 -885 15385 -865
rect 15415 -885 15435 -865
rect 15465 -885 15485 -865
rect 15515 -885 15535 -865
rect 15615 -885 15635 -865
rect 15665 -885 15685 -865
rect 15715 -885 15735 -865
rect 15765 -885 15785 -865
rect 15815 -885 15835 -865
rect 15915 -885 15935 -865
rect 15965 -885 15985 -865
rect 16015 -885 16035 -865
rect 16065 -885 16085 -865
rect 16115 -885 16135 -865
rect 16215 -885 16235 -865
rect 16265 -885 16285 -865
rect 16315 -885 16335 -865
rect 16365 -885 16385 -865
rect 16415 -885 16435 -865
rect 16515 -885 16535 -865
rect 16565 -885 16585 -865
rect 16615 -885 16635 -865
rect 16665 -885 16685 -865
rect 16715 -885 16735 -865
rect 16815 -885 16835 -865
rect 16865 -885 16885 -865
rect 16915 -885 16935 -865
rect 16965 -885 16985 -865
rect 17015 -885 17035 -865
rect 17115 -885 17135 -865
rect 17165 -885 17185 -865
rect 17215 -885 17235 -865
rect 17265 -885 17285 -865
rect 17315 -885 17335 -865
rect 17415 -885 17435 -865
rect 17465 -885 17485 -865
rect 17515 -885 17535 -865
rect 17565 -885 17585 -865
rect 17615 -885 17635 -865
rect 17715 -885 17735 -865
rect 17765 -885 17785 -865
rect 17815 -885 17835 -865
rect 17865 -885 17885 -865
rect 17915 -885 17935 -865
rect 18015 -885 18035 -865
rect 18065 -885 18085 -865
rect 18115 -885 18135 -865
rect 18165 -885 18185 -865
rect 18215 -885 18235 -865
rect 18315 -885 18335 -865
rect 18365 -885 18385 -865
rect 18415 -885 18435 -865
rect 18465 -885 18485 -865
rect 18515 -885 18535 -865
rect 18615 -885 18635 -865
rect 18665 -885 18685 -865
rect 18715 -885 18735 -865
rect 18765 -885 18785 -865
rect 18815 -885 18835 -865
rect 18915 -885 18935 -865
rect 18965 -885 18985 -865
rect 19015 -885 19035 -865
rect 19065 -885 19085 -865
rect 19115 -885 19135 -865
rect 19215 -885 19235 -865
rect 19265 -885 19285 -865
rect 19315 -885 19335 -865
rect 19365 -885 19385 -865
rect 19415 -885 19435 -865
rect 19515 -885 19535 -865
rect 19565 -885 19585 -865
rect 19615 -885 19635 -865
rect 19665 -885 19685 -865
rect 19715 -885 19735 -865
rect 19815 -885 19835 -865
rect 19865 -885 19885 -865
rect 19915 -885 19935 -865
rect 19965 -885 19985 -865
rect 20015 -885 20035 -865
rect 20115 -885 20135 -865
rect 20165 -885 20185 -865
rect 20215 -885 20235 -865
rect 20265 -885 20285 -865
rect 20315 -885 20335 -865
<< locali >>
rect -650 5185 20400 5200
rect -650 5165 -635 5185
rect -615 5165 -585 5185
rect -565 5165 -535 5185
rect -515 5165 -485 5185
rect -465 5165 -435 5185
rect -415 5165 -385 5185
rect -365 5165 -335 5185
rect -315 5165 -285 5185
rect -265 5165 -235 5185
rect -215 5165 -185 5185
rect -165 5165 -135 5185
rect -115 5165 -85 5185
rect -65 5165 -35 5185
rect -15 5165 15 5185
rect 35 5165 65 5185
rect 85 5165 115 5185
rect 135 5165 165 5185
rect 185 5165 215 5185
rect 235 5165 265 5185
rect 285 5165 315 5185
rect 335 5165 365 5185
rect 385 5165 415 5185
rect 435 5165 465 5185
rect 485 5165 515 5185
rect 535 5165 565 5185
rect 585 5165 615 5185
rect 635 5165 665 5185
rect 685 5165 715 5185
rect 735 5165 765 5185
rect 785 5165 815 5185
rect 835 5165 865 5185
rect 885 5165 915 5185
rect 935 5165 965 5185
rect 985 5165 1015 5185
rect 1035 5165 1065 5185
rect 1085 5165 1115 5185
rect 1135 5165 1165 5185
rect 1185 5165 1215 5185
rect 1235 5165 1265 5185
rect 1285 5165 1315 5185
rect 1335 5165 1365 5185
rect 1385 5165 1415 5185
rect 1435 5165 1465 5185
rect 1485 5165 1515 5185
rect 1535 5165 1565 5185
rect 1585 5165 1615 5185
rect 1635 5165 1665 5185
rect 1685 5165 1715 5185
rect 1735 5165 1765 5185
rect 1785 5165 1815 5185
rect 1835 5165 1865 5185
rect 1885 5165 1915 5185
rect 1935 5165 1965 5185
rect 1985 5165 2015 5185
rect 2035 5165 2065 5185
rect 2085 5165 2115 5185
rect 2135 5165 2165 5185
rect 2185 5165 2215 5185
rect 2235 5165 2265 5185
rect 2285 5165 2315 5185
rect 2335 5165 2365 5185
rect 2385 5165 2415 5185
rect 2435 5165 2465 5185
rect 2485 5165 2515 5185
rect 2535 5165 2565 5185
rect 2585 5165 2615 5185
rect 2635 5165 2665 5185
rect 2685 5165 2715 5185
rect 2735 5165 2765 5185
rect 2785 5165 2815 5185
rect 2835 5165 2865 5185
rect 2885 5165 2915 5185
rect 2935 5165 2965 5185
rect 2985 5165 3015 5185
rect 3035 5165 3065 5185
rect 3085 5165 3115 5185
rect 3135 5165 3165 5185
rect 3185 5165 3215 5185
rect 3235 5165 3265 5185
rect 3285 5165 3315 5185
rect 3335 5165 3365 5185
rect 3385 5165 3415 5185
rect 3435 5165 3465 5185
rect 3485 5165 3515 5185
rect 3535 5165 3565 5185
rect 3585 5165 3615 5185
rect 3635 5165 3665 5185
rect 3685 5165 3715 5185
rect 3735 5165 3765 5185
rect 3785 5165 3815 5185
rect 3835 5165 3865 5185
rect 3885 5165 3915 5185
rect 3935 5165 3965 5185
rect 3985 5165 4015 5185
rect 4035 5165 4065 5185
rect 4085 5165 4115 5185
rect 4135 5165 4165 5185
rect 4185 5165 4215 5185
rect 4235 5165 4265 5185
rect 4285 5165 4315 5185
rect 4335 5165 4365 5185
rect 4385 5165 4415 5185
rect 4435 5165 4465 5185
rect 4485 5165 4515 5185
rect 4535 5165 4565 5185
rect 4585 5165 4615 5185
rect 4635 5165 4665 5185
rect 4685 5165 4715 5185
rect 4735 5165 4765 5185
rect 4785 5165 4815 5185
rect 4835 5165 4865 5185
rect 4885 5165 4915 5185
rect 4935 5165 4965 5185
rect 4985 5165 5015 5185
rect 5035 5165 5065 5185
rect 5085 5165 5115 5185
rect 5135 5165 5165 5185
rect 5185 5165 5215 5185
rect 5235 5165 5265 5185
rect 5285 5165 5315 5185
rect 5335 5165 5365 5185
rect 5385 5165 5415 5185
rect 5435 5165 5465 5185
rect 5485 5165 5515 5185
rect 5535 5165 5565 5185
rect 5585 5165 5615 5185
rect 5635 5165 5665 5185
rect 5685 5165 5715 5185
rect 5735 5165 5765 5185
rect 5785 5165 5815 5185
rect 5835 5165 5865 5185
rect 5885 5165 5915 5185
rect 5935 5165 5965 5185
rect 5985 5165 6015 5185
rect 6035 5165 6065 5185
rect 6085 5165 6115 5185
rect 6135 5165 6165 5185
rect 6185 5165 6215 5185
rect 6235 5165 6265 5185
rect 6285 5165 6315 5185
rect 6335 5165 6365 5185
rect 6385 5165 6415 5185
rect 6435 5165 6465 5185
rect 6485 5165 6515 5185
rect 6535 5165 6565 5185
rect 6585 5165 6615 5185
rect 6635 5165 6665 5185
rect 6685 5165 6715 5185
rect 6735 5165 6765 5185
rect 6785 5165 6815 5185
rect 6835 5165 6865 5185
rect 6885 5165 6915 5185
rect 6935 5165 6965 5185
rect 6985 5165 7015 5185
rect 7035 5165 7065 5185
rect 7085 5165 7115 5185
rect 7135 5165 7165 5185
rect 7185 5165 7215 5185
rect 7235 5165 7265 5185
rect 7285 5165 7315 5185
rect 7335 5165 7365 5185
rect 7385 5165 7415 5185
rect 7435 5165 7465 5185
rect 7485 5165 7515 5185
rect 7535 5165 7565 5185
rect 7585 5165 7615 5185
rect 7635 5165 7665 5185
rect 7685 5165 7715 5185
rect 7735 5165 7765 5185
rect 7785 5165 7815 5185
rect 7835 5165 7865 5185
rect 7885 5165 7915 5185
rect 7935 5165 7965 5185
rect 7985 5165 8015 5185
rect 8035 5165 8065 5185
rect 8085 5165 8115 5185
rect 8135 5165 8165 5185
rect 8185 5165 8215 5185
rect 8235 5165 8265 5185
rect 8285 5165 8315 5185
rect 8335 5165 8365 5185
rect 8385 5165 8415 5185
rect 8435 5165 8465 5185
rect 8485 5165 8515 5185
rect 8535 5165 8565 5185
rect 8585 5165 8615 5185
rect 8635 5165 8665 5185
rect 8685 5165 8715 5185
rect 8735 5165 8765 5185
rect 8785 5165 8815 5185
rect 8835 5165 8865 5185
rect 8885 5165 8915 5185
rect 8935 5165 8965 5185
rect 8985 5165 9015 5185
rect 9035 5165 9065 5185
rect 9085 5165 9115 5185
rect 9135 5165 9165 5185
rect 9185 5165 9215 5185
rect 9235 5165 9265 5185
rect 9285 5165 9315 5185
rect 9335 5165 9365 5185
rect 9385 5165 9415 5185
rect 9435 5165 9465 5185
rect 9485 5165 9515 5185
rect 9535 5165 9565 5185
rect 9585 5165 9615 5185
rect 9635 5165 9665 5185
rect 9685 5165 9715 5185
rect 9735 5165 9765 5185
rect 9785 5165 9815 5185
rect 9835 5165 9865 5185
rect 9885 5165 9915 5185
rect 9935 5165 9965 5185
rect 9985 5165 10015 5185
rect 10035 5165 10065 5185
rect 10085 5165 10115 5185
rect 10135 5165 10165 5185
rect 10185 5165 10215 5185
rect 10235 5165 10265 5185
rect 10285 5165 10315 5185
rect 10335 5165 10365 5185
rect 10385 5165 10415 5185
rect 10435 5165 10465 5185
rect 10485 5165 10515 5185
rect 10535 5165 10565 5185
rect 10585 5165 10615 5185
rect 10635 5165 10665 5185
rect 10685 5165 10715 5185
rect 10735 5165 10765 5185
rect 10785 5165 10815 5185
rect 10835 5165 10865 5185
rect 10885 5165 10915 5185
rect 10935 5165 10965 5185
rect 10985 5165 11015 5185
rect 11035 5165 11065 5185
rect 11085 5165 11115 5185
rect 11135 5165 11165 5185
rect 11185 5165 11215 5185
rect 11235 5165 11265 5185
rect 11285 5165 11315 5185
rect 11335 5165 11365 5185
rect 11385 5165 11415 5185
rect 11435 5165 11465 5185
rect 11485 5165 11515 5185
rect 11535 5165 11565 5185
rect 11585 5165 11615 5185
rect 11635 5165 11665 5185
rect 11685 5165 11715 5185
rect 11735 5165 11765 5185
rect 11785 5165 11815 5185
rect 11835 5165 11865 5185
rect 11885 5165 11915 5185
rect 11935 5165 11965 5185
rect 11985 5165 12015 5185
rect 12035 5165 12065 5185
rect 12085 5165 12115 5185
rect 12135 5165 12165 5185
rect 12185 5165 12215 5185
rect 12235 5165 12265 5185
rect 12285 5165 12315 5185
rect 12335 5165 12365 5185
rect 12385 5165 12415 5185
rect 12435 5165 12465 5185
rect 12485 5165 12515 5185
rect 12535 5165 12565 5185
rect 12585 5165 12615 5185
rect 12635 5165 12665 5185
rect 12685 5165 12715 5185
rect 12735 5165 12765 5185
rect 12785 5165 12815 5185
rect 12835 5165 12865 5185
rect 12885 5165 12915 5185
rect 12935 5165 12965 5185
rect 12985 5165 13015 5185
rect 13035 5165 13065 5185
rect 13085 5165 13115 5185
rect 13135 5165 13165 5185
rect 13185 5165 13215 5185
rect 13235 5165 13265 5185
rect 13285 5165 13315 5185
rect 13335 5165 13365 5185
rect 13385 5165 13415 5185
rect 13435 5165 13465 5185
rect 13485 5165 13515 5185
rect 13535 5165 13565 5185
rect 13585 5165 13615 5185
rect 13635 5165 13665 5185
rect 13685 5165 13715 5185
rect 13735 5165 13765 5185
rect 13785 5165 13815 5185
rect 13835 5165 13865 5185
rect 13885 5165 13915 5185
rect 13935 5165 13965 5185
rect 13985 5165 14015 5185
rect 14035 5165 14065 5185
rect 14085 5165 14115 5185
rect 14135 5165 14165 5185
rect 14185 5165 14215 5185
rect 14235 5165 14265 5185
rect 14285 5165 14315 5185
rect 14335 5165 14365 5185
rect 14385 5165 14415 5185
rect 14435 5165 14465 5185
rect 14485 5165 14515 5185
rect 14535 5165 14565 5185
rect 14585 5165 14615 5185
rect 14635 5165 14665 5185
rect 14685 5165 14715 5185
rect 14735 5165 14765 5185
rect 14785 5165 14815 5185
rect 14835 5165 14865 5185
rect 14885 5165 14915 5185
rect 14935 5165 14965 5185
rect 14985 5165 15015 5185
rect 15035 5165 15065 5185
rect 15085 5165 15115 5185
rect 15135 5165 15165 5185
rect 15185 5165 15215 5185
rect 15235 5165 15265 5185
rect 15285 5165 15315 5185
rect 15335 5165 15365 5185
rect 15385 5165 15415 5185
rect 15435 5165 15465 5185
rect 15485 5165 15515 5185
rect 15535 5165 15565 5185
rect 15585 5165 15615 5185
rect 15635 5165 15665 5185
rect 15685 5165 15715 5185
rect 15735 5165 15765 5185
rect 15785 5165 15815 5185
rect 15835 5165 15865 5185
rect 15885 5165 15915 5185
rect 15935 5165 15965 5185
rect 15985 5165 16015 5185
rect 16035 5165 16065 5185
rect 16085 5165 16115 5185
rect 16135 5165 16165 5185
rect 16185 5165 16215 5185
rect 16235 5165 16265 5185
rect 16285 5165 16315 5185
rect 16335 5165 16365 5185
rect 16385 5165 16415 5185
rect 16435 5165 16465 5185
rect 16485 5165 16515 5185
rect 16535 5165 16565 5185
rect 16585 5165 16615 5185
rect 16635 5165 16665 5185
rect 16685 5165 16715 5185
rect 16735 5165 16765 5185
rect 16785 5165 16815 5185
rect 16835 5165 16865 5185
rect 16885 5165 16915 5185
rect 16935 5165 16965 5185
rect 16985 5165 17015 5185
rect 17035 5165 17065 5185
rect 17085 5165 17115 5185
rect 17135 5165 17165 5185
rect 17185 5165 17215 5185
rect 17235 5165 17265 5185
rect 17285 5165 17315 5185
rect 17335 5165 17365 5185
rect 17385 5165 17415 5185
rect 17435 5165 17465 5185
rect 17485 5165 17515 5185
rect 17535 5165 17565 5185
rect 17585 5165 17615 5185
rect 17635 5165 17665 5185
rect 17685 5165 17715 5185
rect 17735 5165 17765 5185
rect 17785 5165 17815 5185
rect 17835 5165 17865 5185
rect 17885 5165 17915 5185
rect 17935 5165 17965 5185
rect 17985 5165 18015 5185
rect 18035 5165 18065 5185
rect 18085 5165 18115 5185
rect 18135 5165 18165 5185
rect 18185 5165 18215 5185
rect 18235 5165 18265 5185
rect 18285 5165 18315 5185
rect 18335 5165 18365 5185
rect 18385 5165 18415 5185
rect 18435 5165 18465 5185
rect 18485 5165 18515 5185
rect 18535 5165 18565 5185
rect 18585 5165 18615 5185
rect 18635 5165 18665 5185
rect 18685 5165 18715 5185
rect 18735 5165 18765 5185
rect 18785 5165 18815 5185
rect 18835 5165 18865 5185
rect 18885 5165 18915 5185
rect 18935 5165 18965 5185
rect 18985 5165 19015 5185
rect 19035 5165 19065 5185
rect 19085 5165 19115 5185
rect 19135 5165 19165 5185
rect 19185 5165 19215 5185
rect 19235 5165 19265 5185
rect 19285 5165 19315 5185
rect 19335 5165 19365 5185
rect 19385 5165 19415 5185
rect 19435 5165 19465 5185
rect 19485 5165 19515 5185
rect 19535 5165 19565 5185
rect 19585 5165 19615 5185
rect 19635 5165 19665 5185
rect 19685 5165 19715 5185
rect 19735 5165 19765 5185
rect 19785 5165 19815 5185
rect 19835 5165 19865 5185
rect 19885 5165 19915 5185
rect 19935 5165 19965 5185
rect 19985 5165 20015 5185
rect 20035 5165 20065 5185
rect 20085 5165 20115 5185
rect 20135 5165 20165 5185
rect 20185 5165 20215 5185
rect 20235 5165 20265 5185
rect 20285 5165 20315 5185
rect 20335 5165 20365 5185
rect 20385 5165 20400 5185
rect -650 5150 20400 5165
rect -650 5085 -600 5100
rect -650 5065 -635 5085
rect -615 5065 -600 5085
rect -650 5035 -600 5065
rect -650 5015 -635 5035
rect -615 5015 -600 5035
rect -650 4985 -600 5015
rect -650 4965 -635 4985
rect -615 4965 -600 4985
rect -650 4935 -600 4965
rect -650 4915 -635 4935
rect -615 4915 -600 4935
rect -650 4885 -600 4915
rect -650 4865 -635 4885
rect -615 4865 -600 4885
rect -650 4835 -600 4865
rect -650 4815 -635 4835
rect -615 4815 -600 4835
rect -650 4785 -600 4815
rect -650 4765 -635 4785
rect -615 4765 -600 4785
rect -650 4735 -600 4765
rect -650 4715 -635 4735
rect -615 4715 -600 4735
rect -650 4685 -600 4715
rect -650 4665 -635 4685
rect -615 4665 -600 4685
rect -650 4635 -600 4665
rect -650 4615 -635 4635
rect -615 4615 -600 4635
rect -650 4600 -600 4615
rect -500 5085 -450 5100
rect -500 5065 -485 5085
rect -465 5065 -450 5085
rect -500 5035 -450 5065
rect -500 5015 -485 5035
rect -465 5015 -450 5035
rect -500 4985 -450 5015
rect -500 4965 -485 4985
rect -465 4965 -450 4985
rect -500 4935 -450 4965
rect -500 4915 -485 4935
rect -465 4915 -450 4935
rect -500 4885 -450 4915
rect -500 4865 -485 4885
rect -465 4865 -450 4885
rect -500 4835 -450 4865
rect -500 4815 -485 4835
rect -465 4815 -450 4835
rect -500 4785 -450 4815
rect -500 4765 -485 4785
rect -465 4765 -450 4785
rect -500 4735 -450 4765
rect -500 4715 -485 4735
rect -465 4715 -450 4735
rect -500 4685 -450 4715
rect -500 4665 -485 4685
rect -465 4665 -450 4685
rect -500 4635 -450 4665
rect -500 4615 -485 4635
rect -465 4615 -450 4635
rect -500 4600 -450 4615
rect -350 5085 -300 5100
rect -350 5065 -335 5085
rect -315 5065 -300 5085
rect -350 5035 -300 5065
rect -350 5015 -335 5035
rect -315 5015 -300 5035
rect -350 4985 -300 5015
rect -350 4965 -335 4985
rect -315 4965 -300 4985
rect -350 4935 -300 4965
rect -350 4915 -335 4935
rect -315 4915 -300 4935
rect -350 4885 -300 4915
rect -350 4865 -335 4885
rect -315 4865 -300 4885
rect -350 4835 -300 4865
rect -350 4815 -335 4835
rect -315 4815 -300 4835
rect -350 4785 -300 4815
rect -350 4765 -335 4785
rect -315 4765 -300 4785
rect -350 4735 -300 4765
rect -350 4715 -335 4735
rect -315 4715 -300 4735
rect -350 4685 -300 4715
rect -350 4665 -335 4685
rect -315 4665 -300 4685
rect -350 4635 -300 4665
rect -350 4615 -335 4635
rect -315 4615 -300 4635
rect -350 4600 -300 4615
rect -200 5085 -150 5100
rect -200 5065 -185 5085
rect -165 5065 -150 5085
rect -200 5035 -150 5065
rect -200 5015 -185 5035
rect -165 5015 -150 5035
rect -200 4985 -150 5015
rect -200 4965 -185 4985
rect -165 4965 -150 4985
rect -200 4935 -150 4965
rect -200 4915 -185 4935
rect -165 4915 -150 4935
rect -200 4885 -150 4915
rect -200 4865 -185 4885
rect -165 4865 -150 4885
rect -200 4835 -150 4865
rect -200 4815 -185 4835
rect -165 4815 -150 4835
rect -200 4785 -150 4815
rect -200 4765 -185 4785
rect -165 4765 -150 4785
rect -200 4735 -150 4765
rect -200 4715 -185 4735
rect -165 4715 -150 4735
rect -200 4685 -150 4715
rect -200 4665 -185 4685
rect -165 4665 -150 4685
rect -200 4635 -150 4665
rect -200 4615 -185 4635
rect -165 4615 -150 4635
rect -200 4600 -150 4615
rect -50 5085 0 5100
rect -50 5065 -35 5085
rect -15 5065 0 5085
rect -50 5035 0 5065
rect -50 5015 -35 5035
rect -15 5015 0 5035
rect -50 4985 0 5015
rect -50 4965 -35 4985
rect -15 4965 0 4985
rect -50 4935 0 4965
rect -50 4915 -35 4935
rect -15 4915 0 4935
rect -50 4885 0 4915
rect -50 4865 -35 4885
rect -15 4865 0 4885
rect -50 4835 0 4865
rect -50 4815 -35 4835
rect -15 4815 0 4835
rect -50 4785 0 4815
rect -50 4765 -35 4785
rect -15 4765 0 4785
rect -50 4735 0 4765
rect -50 4715 -35 4735
rect -15 4715 0 4735
rect -50 4685 0 4715
rect -50 4665 -35 4685
rect -15 4665 0 4685
rect -50 4635 0 4665
rect -50 4615 -35 4635
rect -15 4615 0 4635
rect -50 4600 0 4615
rect 550 5085 600 5100
rect 550 5065 565 5085
rect 585 5065 600 5085
rect 550 5035 600 5065
rect 550 5015 565 5035
rect 585 5015 600 5035
rect 550 4985 600 5015
rect 550 4965 565 4985
rect 585 4965 600 4985
rect 550 4935 600 4965
rect 550 4915 565 4935
rect 585 4915 600 4935
rect 550 4885 600 4915
rect 550 4865 565 4885
rect 585 4865 600 4885
rect 550 4835 600 4865
rect 550 4815 565 4835
rect 585 4815 600 4835
rect 550 4785 600 4815
rect 550 4765 565 4785
rect 585 4765 600 4785
rect 550 4735 600 4765
rect 550 4715 565 4735
rect 585 4715 600 4735
rect 550 4685 600 4715
rect 550 4665 565 4685
rect 585 4665 600 4685
rect 550 4635 600 4665
rect 550 4615 565 4635
rect 585 4615 600 4635
rect 550 4600 600 4615
rect 700 5085 750 5100
rect 700 5065 715 5085
rect 735 5065 750 5085
rect 700 5035 750 5065
rect 700 5015 715 5035
rect 735 5015 750 5035
rect 700 4985 750 5015
rect 700 4965 715 4985
rect 735 4965 750 4985
rect 700 4935 750 4965
rect 700 4915 715 4935
rect 735 4915 750 4935
rect 700 4885 750 4915
rect 700 4865 715 4885
rect 735 4865 750 4885
rect 700 4835 750 4865
rect 700 4815 715 4835
rect 735 4815 750 4835
rect 700 4785 750 4815
rect 700 4765 715 4785
rect 735 4765 750 4785
rect 700 4735 750 4765
rect 700 4715 715 4735
rect 735 4715 750 4735
rect 700 4685 750 4715
rect 700 4665 715 4685
rect 735 4665 750 4685
rect 700 4635 750 4665
rect 700 4615 715 4635
rect 735 4615 750 4635
rect 700 4600 750 4615
rect 850 5085 900 5100
rect 850 5065 865 5085
rect 885 5065 900 5085
rect 850 5035 900 5065
rect 850 5015 865 5035
rect 885 5015 900 5035
rect 850 4985 900 5015
rect 850 4965 865 4985
rect 885 4965 900 4985
rect 850 4935 900 4965
rect 850 4915 865 4935
rect 885 4915 900 4935
rect 850 4885 900 4915
rect 850 4865 865 4885
rect 885 4865 900 4885
rect 850 4835 900 4865
rect 850 4815 865 4835
rect 885 4815 900 4835
rect 850 4785 900 4815
rect 850 4765 865 4785
rect 885 4765 900 4785
rect 850 4735 900 4765
rect 850 4715 865 4735
rect 885 4715 900 4735
rect 850 4685 900 4715
rect 850 4665 865 4685
rect 885 4665 900 4685
rect 850 4635 900 4665
rect 850 4615 865 4635
rect 885 4615 900 4635
rect 850 4600 900 4615
rect 1000 5085 1050 5100
rect 1000 5065 1015 5085
rect 1035 5065 1050 5085
rect 1000 5035 1050 5065
rect 1000 5015 1015 5035
rect 1035 5015 1050 5035
rect 1000 4985 1050 5015
rect 1000 4965 1015 4985
rect 1035 4965 1050 4985
rect 1000 4935 1050 4965
rect 1000 4915 1015 4935
rect 1035 4915 1050 4935
rect 1000 4885 1050 4915
rect 1000 4865 1015 4885
rect 1035 4865 1050 4885
rect 1000 4835 1050 4865
rect 1000 4815 1015 4835
rect 1035 4815 1050 4835
rect 1000 4785 1050 4815
rect 1000 4765 1015 4785
rect 1035 4765 1050 4785
rect 1000 4735 1050 4765
rect 1000 4715 1015 4735
rect 1035 4715 1050 4735
rect 1000 4685 1050 4715
rect 1000 4665 1015 4685
rect 1035 4665 1050 4685
rect 1000 4635 1050 4665
rect 1000 4615 1015 4635
rect 1035 4615 1050 4635
rect 1000 4600 1050 4615
rect 1150 5085 1200 5100
rect 1150 5065 1165 5085
rect 1185 5065 1200 5085
rect 1150 5035 1200 5065
rect 1150 5015 1165 5035
rect 1185 5015 1200 5035
rect 1150 4985 1200 5015
rect 1150 4965 1165 4985
rect 1185 4965 1200 4985
rect 1150 4935 1200 4965
rect 1150 4915 1165 4935
rect 1185 4915 1200 4935
rect 1150 4885 1200 4915
rect 1150 4865 1165 4885
rect 1185 4865 1200 4885
rect 1150 4835 1200 4865
rect 1150 4815 1165 4835
rect 1185 4815 1200 4835
rect 1150 4785 1200 4815
rect 1150 4765 1165 4785
rect 1185 4765 1200 4785
rect 1150 4735 1200 4765
rect 1150 4715 1165 4735
rect 1185 4715 1200 4735
rect 1150 4685 1200 4715
rect 1150 4665 1165 4685
rect 1185 4665 1200 4685
rect 1150 4635 1200 4665
rect 1150 4615 1165 4635
rect 1185 4615 1200 4635
rect 1150 4600 1200 4615
rect 1300 5085 1350 5100
rect 1300 5065 1315 5085
rect 1335 5065 1350 5085
rect 1300 5035 1350 5065
rect 1300 5015 1315 5035
rect 1335 5015 1350 5035
rect 1300 4985 1350 5015
rect 1300 4965 1315 4985
rect 1335 4965 1350 4985
rect 1300 4935 1350 4965
rect 1300 4915 1315 4935
rect 1335 4915 1350 4935
rect 1300 4885 1350 4915
rect 1300 4865 1315 4885
rect 1335 4865 1350 4885
rect 1300 4835 1350 4865
rect 1300 4815 1315 4835
rect 1335 4815 1350 4835
rect 1300 4785 1350 4815
rect 1300 4765 1315 4785
rect 1335 4765 1350 4785
rect 1300 4735 1350 4765
rect 1300 4715 1315 4735
rect 1335 4715 1350 4735
rect 1300 4685 1350 4715
rect 1300 4665 1315 4685
rect 1335 4665 1350 4685
rect 1300 4635 1350 4665
rect 1300 4615 1315 4635
rect 1335 4615 1350 4635
rect 1300 4600 1350 4615
rect 1450 5085 1500 5100
rect 1450 5065 1465 5085
rect 1485 5065 1500 5085
rect 1450 5035 1500 5065
rect 1450 5015 1465 5035
rect 1485 5015 1500 5035
rect 1450 4985 1500 5015
rect 1450 4965 1465 4985
rect 1485 4965 1500 4985
rect 1450 4935 1500 4965
rect 1450 4915 1465 4935
rect 1485 4915 1500 4935
rect 1450 4885 1500 4915
rect 1450 4865 1465 4885
rect 1485 4865 1500 4885
rect 1450 4835 1500 4865
rect 1450 4815 1465 4835
rect 1485 4815 1500 4835
rect 1450 4785 1500 4815
rect 1450 4765 1465 4785
rect 1485 4765 1500 4785
rect 1450 4735 1500 4765
rect 1450 4715 1465 4735
rect 1485 4715 1500 4735
rect 1450 4685 1500 4715
rect 1450 4665 1465 4685
rect 1485 4665 1500 4685
rect 1450 4635 1500 4665
rect 1450 4615 1465 4635
rect 1485 4615 1500 4635
rect 1450 4600 1500 4615
rect 1600 5085 1650 5100
rect 1600 5065 1615 5085
rect 1635 5065 1650 5085
rect 1600 5035 1650 5065
rect 1600 5015 1615 5035
rect 1635 5015 1650 5035
rect 1600 4985 1650 5015
rect 1600 4965 1615 4985
rect 1635 4965 1650 4985
rect 1600 4935 1650 4965
rect 1600 4915 1615 4935
rect 1635 4915 1650 4935
rect 1600 4885 1650 4915
rect 1600 4865 1615 4885
rect 1635 4865 1650 4885
rect 1600 4835 1650 4865
rect 1600 4815 1615 4835
rect 1635 4815 1650 4835
rect 1600 4785 1650 4815
rect 1600 4765 1615 4785
rect 1635 4765 1650 4785
rect 1600 4735 1650 4765
rect 1600 4715 1615 4735
rect 1635 4715 1650 4735
rect 1600 4685 1650 4715
rect 1600 4665 1615 4685
rect 1635 4665 1650 4685
rect 1600 4635 1650 4665
rect 1600 4615 1615 4635
rect 1635 4615 1650 4635
rect 1600 4600 1650 4615
rect 1750 5085 1800 5100
rect 1750 5065 1765 5085
rect 1785 5065 1800 5085
rect 1750 5035 1800 5065
rect 1750 5015 1765 5035
rect 1785 5015 1800 5035
rect 1750 4985 1800 5015
rect 1750 4965 1765 4985
rect 1785 4965 1800 4985
rect 1750 4935 1800 4965
rect 1750 4915 1765 4935
rect 1785 4915 1800 4935
rect 1750 4885 1800 4915
rect 1750 4865 1765 4885
rect 1785 4865 1800 4885
rect 1750 4835 1800 4865
rect 1750 4815 1765 4835
rect 1785 4815 1800 4835
rect 1750 4785 1800 4815
rect 1750 4765 1765 4785
rect 1785 4765 1800 4785
rect 1750 4735 1800 4765
rect 1750 4715 1765 4735
rect 1785 4715 1800 4735
rect 1750 4685 1800 4715
rect 1750 4665 1765 4685
rect 1785 4665 1800 4685
rect 1750 4635 1800 4665
rect 1750 4615 1765 4635
rect 1785 4615 1800 4635
rect 1750 4600 1800 4615
rect 1900 5085 1950 5100
rect 1900 5065 1915 5085
rect 1935 5065 1950 5085
rect 1900 5035 1950 5065
rect 1900 5015 1915 5035
rect 1935 5015 1950 5035
rect 1900 4985 1950 5015
rect 1900 4965 1915 4985
rect 1935 4965 1950 4985
rect 1900 4935 1950 4965
rect 1900 4915 1915 4935
rect 1935 4915 1950 4935
rect 1900 4885 1950 4915
rect 1900 4865 1915 4885
rect 1935 4865 1950 4885
rect 1900 4835 1950 4865
rect 1900 4815 1915 4835
rect 1935 4815 1950 4835
rect 1900 4785 1950 4815
rect 1900 4765 1915 4785
rect 1935 4765 1950 4785
rect 1900 4735 1950 4765
rect 1900 4715 1915 4735
rect 1935 4715 1950 4735
rect 1900 4685 1950 4715
rect 1900 4665 1915 4685
rect 1935 4665 1950 4685
rect 1900 4635 1950 4665
rect 1900 4615 1915 4635
rect 1935 4615 1950 4635
rect 1900 4600 1950 4615
rect 2050 5085 2100 5100
rect 2050 5065 2065 5085
rect 2085 5065 2100 5085
rect 2050 5035 2100 5065
rect 2050 5015 2065 5035
rect 2085 5015 2100 5035
rect 2050 4985 2100 5015
rect 2050 4965 2065 4985
rect 2085 4965 2100 4985
rect 2050 4935 2100 4965
rect 2050 4915 2065 4935
rect 2085 4915 2100 4935
rect 2050 4885 2100 4915
rect 2050 4865 2065 4885
rect 2085 4865 2100 4885
rect 2050 4835 2100 4865
rect 2050 4815 2065 4835
rect 2085 4815 2100 4835
rect 2050 4785 2100 4815
rect 2050 4765 2065 4785
rect 2085 4765 2100 4785
rect 2050 4735 2100 4765
rect 2050 4715 2065 4735
rect 2085 4715 2100 4735
rect 2050 4685 2100 4715
rect 2050 4665 2065 4685
rect 2085 4665 2100 4685
rect 2050 4635 2100 4665
rect 2050 4615 2065 4635
rect 2085 4615 2100 4635
rect 2050 4600 2100 4615
rect 2200 5085 2250 5100
rect 2200 5065 2215 5085
rect 2235 5065 2250 5085
rect 2200 5035 2250 5065
rect 2200 5015 2215 5035
rect 2235 5015 2250 5035
rect 2200 4985 2250 5015
rect 2200 4965 2215 4985
rect 2235 4965 2250 4985
rect 2200 4935 2250 4965
rect 2200 4915 2215 4935
rect 2235 4915 2250 4935
rect 2200 4885 2250 4915
rect 2200 4865 2215 4885
rect 2235 4865 2250 4885
rect 2200 4835 2250 4865
rect 2200 4815 2215 4835
rect 2235 4815 2250 4835
rect 2200 4785 2250 4815
rect 2200 4765 2215 4785
rect 2235 4765 2250 4785
rect 2200 4735 2250 4765
rect 2200 4715 2215 4735
rect 2235 4715 2250 4735
rect 2200 4685 2250 4715
rect 2200 4665 2215 4685
rect 2235 4665 2250 4685
rect 2200 4635 2250 4665
rect 2200 4615 2215 4635
rect 2235 4615 2250 4635
rect 2200 4600 2250 4615
rect 2350 5085 2400 5100
rect 2350 5065 2365 5085
rect 2385 5065 2400 5085
rect 2350 5035 2400 5065
rect 2350 5015 2365 5035
rect 2385 5015 2400 5035
rect 2350 4985 2400 5015
rect 2350 4965 2365 4985
rect 2385 4965 2400 4985
rect 2350 4935 2400 4965
rect 2350 4915 2365 4935
rect 2385 4915 2400 4935
rect 2350 4885 2400 4915
rect 2350 4865 2365 4885
rect 2385 4865 2400 4885
rect 2350 4835 2400 4865
rect 2350 4815 2365 4835
rect 2385 4815 2400 4835
rect 2350 4785 2400 4815
rect 2350 4765 2365 4785
rect 2385 4765 2400 4785
rect 2350 4735 2400 4765
rect 2350 4715 2365 4735
rect 2385 4715 2400 4735
rect 2350 4685 2400 4715
rect 2350 4665 2365 4685
rect 2385 4665 2400 4685
rect 2350 4635 2400 4665
rect 2350 4615 2365 4635
rect 2385 4615 2400 4635
rect 2350 4600 2400 4615
rect 2500 5085 2550 5100
rect 2500 5065 2515 5085
rect 2535 5065 2550 5085
rect 2500 5035 2550 5065
rect 2500 5015 2515 5035
rect 2535 5015 2550 5035
rect 2500 4985 2550 5015
rect 2500 4965 2515 4985
rect 2535 4965 2550 4985
rect 2500 4935 2550 4965
rect 2500 4915 2515 4935
rect 2535 4915 2550 4935
rect 2500 4885 2550 4915
rect 2500 4865 2515 4885
rect 2535 4865 2550 4885
rect 2500 4835 2550 4865
rect 2500 4815 2515 4835
rect 2535 4815 2550 4835
rect 2500 4785 2550 4815
rect 2500 4765 2515 4785
rect 2535 4765 2550 4785
rect 2500 4735 2550 4765
rect 2500 4715 2515 4735
rect 2535 4715 2550 4735
rect 2500 4685 2550 4715
rect 2500 4665 2515 4685
rect 2535 4665 2550 4685
rect 2500 4635 2550 4665
rect 2500 4615 2515 4635
rect 2535 4615 2550 4635
rect 2500 4600 2550 4615
rect 2650 5085 2700 5100
rect 2650 5065 2665 5085
rect 2685 5065 2700 5085
rect 2650 5035 2700 5065
rect 2650 5015 2665 5035
rect 2685 5015 2700 5035
rect 2650 4985 2700 5015
rect 2650 4965 2665 4985
rect 2685 4965 2700 4985
rect 2650 4935 2700 4965
rect 2650 4915 2665 4935
rect 2685 4915 2700 4935
rect 2650 4885 2700 4915
rect 2650 4865 2665 4885
rect 2685 4865 2700 4885
rect 2650 4835 2700 4865
rect 2650 4815 2665 4835
rect 2685 4815 2700 4835
rect 2650 4785 2700 4815
rect 2650 4765 2665 4785
rect 2685 4765 2700 4785
rect 2650 4735 2700 4765
rect 2650 4715 2665 4735
rect 2685 4715 2700 4735
rect 2650 4685 2700 4715
rect 2650 4665 2665 4685
rect 2685 4665 2700 4685
rect 2650 4635 2700 4665
rect 2650 4615 2665 4635
rect 2685 4615 2700 4635
rect 2650 4600 2700 4615
rect 2800 5085 2850 5100
rect 2800 5065 2815 5085
rect 2835 5065 2850 5085
rect 2800 5035 2850 5065
rect 2800 5015 2815 5035
rect 2835 5015 2850 5035
rect 2800 4985 2850 5015
rect 2800 4965 2815 4985
rect 2835 4965 2850 4985
rect 2800 4935 2850 4965
rect 2800 4915 2815 4935
rect 2835 4915 2850 4935
rect 2800 4885 2850 4915
rect 2800 4865 2815 4885
rect 2835 4865 2850 4885
rect 2800 4835 2850 4865
rect 2800 4815 2815 4835
rect 2835 4815 2850 4835
rect 2800 4785 2850 4815
rect 2800 4765 2815 4785
rect 2835 4765 2850 4785
rect 2800 4735 2850 4765
rect 2800 4715 2815 4735
rect 2835 4715 2850 4735
rect 2800 4685 2850 4715
rect 2800 4665 2815 4685
rect 2835 4665 2850 4685
rect 2800 4635 2850 4665
rect 2800 4615 2815 4635
rect 2835 4615 2850 4635
rect 2800 4600 2850 4615
rect 2950 5085 3000 5100
rect 2950 5065 2965 5085
rect 2985 5065 3000 5085
rect 2950 5035 3000 5065
rect 2950 5015 2965 5035
rect 2985 5015 3000 5035
rect 2950 4985 3000 5015
rect 2950 4965 2965 4985
rect 2985 4965 3000 4985
rect 2950 4935 3000 4965
rect 2950 4915 2965 4935
rect 2985 4915 3000 4935
rect 2950 4885 3000 4915
rect 2950 4865 2965 4885
rect 2985 4865 3000 4885
rect 2950 4835 3000 4865
rect 2950 4815 2965 4835
rect 2985 4815 3000 4835
rect 2950 4785 3000 4815
rect 2950 4765 2965 4785
rect 2985 4765 3000 4785
rect 2950 4735 3000 4765
rect 2950 4715 2965 4735
rect 2985 4715 3000 4735
rect 2950 4685 3000 4715
rect 2950 4665 2965 4685
rect 2985 4665 3000 4685
rect 2950 4635 3000 4665
rect 2950 4615 2965 4635
rect 2985 4615 3000 4635
rect 2950 4600 3000 4615
rect 3100 5085 3150 5100
rect 3100 5065 3115 5085
rect 3135 5065 3150 5085
rect 3100 5035 3150 5065
rect 3100 5015 3115 5035
rect 3135 5015 3150 5035
rect 3100 4985 3150 5015
rect 3100 4965 3115 4985
rect 3135 4965 3150 4985
rect 3100 4935 3150 4965
rect 3100 4915 3115 4935
rect 3135 4915 3150 4935
rect 3100 4885 3150 4915
rect 3100 4865 3115 4885
rect 3135 4865 3150 4885
rect 3100 4835 3150 4865
rect 3100 4815 3115 4835
rect 3135 4815 3150 4835
rect 3100 4785 3150 4815
rect 3100 4765 3115 4785
rect 3135 4765 3150 4785
rect 3100 4735 3150 4765
rect 3100 4715 3115 4735
rect 3135 4715 3150 4735
rect 3100 4685 3150 4715
rect 3100 4665 3115 4685
rect 3135 4665 3150 4685
rect 3100 4635 3150 4665
rect 3100 4615 3115 4635
rect 3135 4615 3150 4635
rect 3100 4600 3150 4615
rect 3250 5085 3300 5100
rect 3250 5065 3265 5085
rect 3285 5065 3300 5085
rect 3250 5035 3300 5065
rect 3250 5015 3265 5035
rect 3285 5015 3300 5035
rect 3250 4985 3300 5015
rect 3250 4965 3265 4985
rect 3285 4965 3300 4985
rect 3250 4935 3300 4965
rect 3250 4915 3265 4935
rect 3285 4915 3300 4935
rect 3250 4885 3300 4915
rect 3250 4865 3265 4885
rect 3285 4865 3300 4885
rect 3250 4835 3300 4865
rect 3250 4815 3265 4835
rect 3285 4815 3300 4835
rect 3250 4785 3300 4815
rect 3250 4765 3265 4785
rect 3285 4765 3300 4785
rect 3250 4735 3300 4765
rect 3250 4715 3265 4735
rect 3285 4715 3300 4735
rect 3250 4685 3300 4715
rect 3250 4665 3265 4685
rect 3285 4665 3300 4685
rect 3250 4635 3300 4665
rect 3250 4615 3265 4635
rect 3285 4615 3300 4635
rect 3250 4600 3300 4615
rect 3400 5085 3450 5100
rect 3400 5065 3415 5085
rect 3435 5065 3450 5085
rect 3400 5035 3450 5065
rect 3400 5015 3415 5035
rect 3435 5015 3450 5035
rect 3400 4985 3450 5015
rect 3400 4965 3415 4985
rect 3435 4965 3450 4985
rect 3400 4935 3450 4965
rect 3400 4915 3415 4935
rect 3435 4915 3450 4935
rect 3400 4885 3450 4915
rect 3400 4865 3415 4885
rect 3435 4865 3450 4885
rect 3400 4835 3450 4865
rect 3400 4815 3415 4835
rect 3435 4815 3450 4835
rect 3400 4785 3450 4815
rect 3400 4765 3415 4785
rect 3435 4765 3450 4785
rect 3400 4735 3450 4765
rect 3400 4715 3415 4735
rect 3435 4715 3450 4735
rect 3400 4685 3450 4715
rect 3400 4665 3415 4685
rect 3435 4665 3450 4685
rect 3400 4635 3450 4665
rect 3400 4615 3415 4635
rect 3435 4615 3450 4635
rect 3400 4600 3450 4615
rect 3550 5085 3600 5100
rect 3550 5065 3565 5085
rect 3585 5065 3600 5085
rect 3550 5035 3600 5065
rect 3550 5015 3565 5035
rect 3585 5015 3600 5035
rect 3550 4985 3600 5015
rect 3550 4965 3565 4985
rect 3585 4965 3600 4985
rect 3550 4935 3600 4965
rect 3550 4915 3565 4935
rect 3585 4915 3600 4935
rect 3550 4885 3600 4915
rect 3550 4865 3565 4885
rect 3585 4865 3600 4885
rect 3550 4835 3600 4865
rect 3550 4815 3565 4835
rect 3585 4815 3600 4835
rect 3550 4785 3600 4815
rect 3550 4765 3565 4785
rect 3585 4765 3600 4785
rect 3550 4735 3600 4765
rect 3550 4715 3565 4735
rect 3585 4715 3600 4735
rect 3550 4685 3600 4715
rect 3550 4665 3565 4685
rect 3585 4665 3600 4685
rect 3550 4635 3600 4665
rect 3550 4615 3565 4635
rect 3585 4615 3600 4635
rect 3550 4600 3600 4615
rect 4150 5085 4200 5100
rect 4150 5065 4165 5085
rect 4185 5065 4200 5085
rect 4150 5035 4200 5065
rect 4150 5015 4165 5035
rect 4185 5015 4200 5035
rect 4150 4985 4200 5015
rect 4150 4965 4165 4985
rect 4185 4965 4200 4985
rect 4150 4935 4200 4965
rect 4150 4915 4165 4935
rect 4185 4915 4200 4935
rect 4150 4885 4200 4915
rect 4150 4865 4165 4885
rect 4185 4865 4200 4885
rect 4150 4835 4200 4865
rect 4150 4815 4165 4835
rect 4185 4815 4200 4835
rect 4150 4785 4200 4815
rect 4150 4765 4165 4785
rect 4185 4765 4200 4785
rect 4150 4735 4200 4765
rect 4150 4715 4165 4735
rect 4185 4715 4200 4735
rect 4150 4685 4200 4715
rect 4150 4665 4165 4685
rect 4185 4665 4200 4685
rect 4150 4635 4200 4665
rect 4150 4615 4165 4635
rect 4185 4615 4200 4635
rect 4150 4600 4200 4615
rect 4750 5085 4800 5100
rect 4750 5065 4765 5085
rect 4785 5065 4800 5085
rect 4750 5035 4800 5065
rect 4750 5015 4765 5035
rect 4785 5015 4800 5035
rect 4750 4985 4800 5015
rect 4750 4965 4765 4985
rect 4785 4965 4800 4985
rect 4750 4935 4800 4965
rect 4750 4915 4765 4935
rect 4785 4915 4800 4935
rect 4750 4885 4800 4915
rect 4750 4865 4765 4885
rect 4785 4865 4800 4885
rect 4750 4835 4800 4865
rect 4750 4815 4765 4835
rect 4785 4815 4800 4835
rect 4750 4785 4800 4815
rect 4750 4765 4765 4785
rect 4785 4765 4800 4785
rect 4750 4735 4800 4765
rect 4750 4715 4765 4735
rect 4785 4715 4800 4735
rect 4750 4685 4800 4715
rect 4750 4665 4765 4685
rect 4785 4665 4800 4685
rect 4750 4635 4800 4665
rect 4750 4615 4765 4635
rect 4785 4615 4800 4635
rect 4750 4600 4800 4615
rect 4900 5085 4950 5100
rect 4900 5065 4915 5085
rect 4935 5065 4950 5085
rect 4900 5035 4950 5065
rect 4900 5015 4915 5035
rect 4935 5015 4950 5035
rect 4900 4985 4950 5015
rect 4900 4965 4915 4985
rect 4935 4965 4950 4985
rect 4900 4935 4950 4965
rect 4900 4915 4915 4935
rect 4935 4915 4950 4935
rect 4900 4885 4950 4915
rect 4900 4865 4915 4885
rect 4935 4865 4950 4885
rect 4900 4835 4950 4865
rect 4900 4815 4915 4835
rect 4935 4815 4950 4835
rect 4900 4785 4950 4815
rect 4900 4765 4915 4785
rect 4935 4765 4950 4785
rect 4900 4735 4950 4765
rect 4900 4715 4915 4735
rect 4935 4715 4950 4735
rect 4900 4685 4950 4715
rect 4900 4665 4915 4685
rect 4935 4665 4950 4685
rect 4900 4635 4950 4665
rect 4900 4615 4915 4635
rect 4935 4615 4950 4635
rect 4900 4600 4950 4615
rect 5050 5085 5100 5100
rect 5050 5065 5065 5085
rect 5085 5065 5100 5085
rect 5050 5035 5100 5065
rect 5050 5015 5065 5035
rect 5085 5015 5100 5035
rect 5050 4985 5100 5015
rect 5050 4965 5065 4985
rect 5085 4965 5100 4985
rect 5050 4935 5100 4965
rect 5050 4915 5065 4935
rect 5085 4915 5100 4935
rect 5050 4885 5100 4915
rect 5050 4865 5065 4885
rect 5085 4865 5100 4885
rect 5050 4835 5100 4865
rect 5050 4815 5065 4835
rect 5085 4815 5100 4835
rect 5050 4785 5100 4815
rect 5050 4765 5065 4785
rect 5085 4765 5100 4785
rect 5050 4735 5100 4765
rect 5050 4715 5065 4735
rect 5085 4715 5100 4735
rect 5050 4685 5100 4715
rect 5050 4665 5065 4685
rect 5085 4665 5100 4685
rect 5050 4635 5100 4665
rect 5050 4615 5065 4635
rect 5085 4615 5100 4635
rect 5050 4600 5100 4615
rect 5200 5085 5250 5100
rect 5200 5065 5215 5085
rect 5235 5065 5250 5085
rect 5200 5035 5250 5065
rect 5200 5015 5215 5035
rect 5235 5015 5250 5035
rect 5200 4985 5250 5015
rect 5200 4965 5215 4985
rect 5235 4965 5250 4985
rect 5200 4935 5250 4965
rect 5200 4915 5215 4935
rect 5235 4915 5250 4935
rect 5200 4885 5250 4915
rect 5200 4865 5215 4885
rect 5235 4865 5250 4885
rect 5200 4835 5250 4865
rect 5200 4815 5215 4835
rect 5235 4815 5250 4835
rect 5200 4785 5250 4815
rect 5200 4765 5215 4785
rect 5235 4765 5250 4785
rect 5200 4735 5250 4765
rect 5200 4715 5215 4735
rect 5235 4715 5250 4735
rect 5200 4685 5250 4715
rect 5200 4665 5215 4685
rect 5235 4665 5250 4685
rect 5200 4635 5250 4665
rect 5200 4615 5215 4635
rect 5235 4615 5250 4635
rect 5200 4600 5250 4615
rect 5350 5085 5400 5100
rect 5350 5065 5365 5085
rect 5385 5065 5400 5085
rect 5350 5035 5400 5065
rect 5350 5015 5365 5035
rect 5385 5015 5400 5035
rect 5350 4985 5400 5015
rect 5350 4965 5365 4985
rect 5385 4965 5400 4985
rect 5350 4935 5400 4965
rect 5350 4915 5365 4935
rect 5385 4915 5400 4935
rect 5350 4885 5400 4915
rect 5350 4865 5365 4885
rect 5385 4865 5400 4885
rect 5350 4835 5400 4865
rect 5350 4815 5365 4835
rect 5385 4815 5400 4835
rect 5350 4785 5400 4815
rect 5350 4765 5365 4785
rect 5385 4765 5400 4785
rect 5350 4735 5400 4765
rect 5350 4715 5365 4735
rect 5385 4715 5400 4735
rect 5350 4685 5400 4715
rect 5350 4665 5365 4685
rect 5385 4665 5400 4685
rect 5350 4635 5400 4665
rect 5350 4615 5365 4635
rect 5385 4615 5400 4635
rect 5350 4600 5400 4615
rect 5500 5085 5550 5100
rect 5500 5065 5515 5085
rect 5535 5065 5550 5085
rect 5500 5035 5550 5065
rect 5500 5015 5515 5035
rect 5535 5015 5550 5035
rect 5500 4985 5550 5015
rect 5500 4965 5515 4985
rect 5535 4965 5550 4985
rect 5500 4935 5550 4965
rect 5500 4915 5515 4935
rect 5535 4915 5550 4935
rect 5500 4885 5550 4915
rect 5500 4865 5515 4885
rect 5535 4865 5550 4885
rect 5500 4835 5550 4865
rect 5500 4815 5515 4835
rect 5535 4815 5550 4835
rect 5500 4785 5550 4815
rect 5500 4765 5515 4785
rect 5535 4765 5550 4785
rect 5500 4735 5550 4765
rect 5500 4715 5515 4735
rect 5535 4715 5550 4735
rect 5500 4685 5550 4715
rect 5500 4665 5515 4685
rect 5535 4665 5550 4685
rect 5500 4635 5550 4665
rect 5500 4615 5515 4635
rect 5535 4615 5550 4635
rect 5500 4600 5550 4615
rect 5650 5085 5700 5100
rect 5650 5065 5665 5085
rect 5685 5065 5700 5085
rect 5650 5035 5700 5065
rect 5650 5015 5665 5035
rect 5685 5015 5700 5035
rect 5650 4985 5700 5015
rect 5650 4965 5665 4985
rect 5685 4965 5700 4985
rect 5650 4935 5700 4965
rect 5650 4915 5665 4935
rect 5685 4915 5700 4935
rect 5650 4885 5700 4915
rect 5650 4865 5665 4885
rect 5685 4865 5700 4885
rect 5650 4835 5700 4865
rect 5650 4815 5665 4835
rect 5685 4815 5700 4835
rect 5650 4785 5700 4815
rect 5650 4765 5665 4785
rect 5685 4765 5700 4785
rect 5650 4735 5700 4765
rect 5650 4715 5665 4735
rect 5685 4715 5700 4735
rect 5650 4685 5700 4715
rect 5650 4665 5665 4685
rect 5685 4665 5700 4685
rect 5650 4635 5700 4665
rect 5650 4615 5665 4635
rect 5685 4615 5700 4635
rect 5650 4600 5700 4615
rect 5800 5085 5850 5100
rect 5800 5065 5815 5085
rect 5835 5065 5850 5085
rect 5800 5035 5850 5065
rect 5800 5015 5815 5035
rect 5835 5015 5850 5035
rect 5800 4985 5850 5015
rect 5800 4965 5815 4985
rect 5835 4965 5850 4985
rect 5800 4935 5850 4965
rect 5800 4915 5815 4935
rect 5835 4915 5850 4935
rect 5800 4885 5850 4915
rect 5800 4865 5815 4885
rect 5835 4865 5850 4885
rect 5800 4835 5850 4865
rect 5800 4815 5815 4835
rect 5835 4815 5850 4835
rect 5800 4785 5850 4815
rect 5800 4765 5815 4785
rect 5835 4765 5850 4785
rect 5800 4735 5850 4765
rect 5800 4715 5815 4735
rect 5835 4715 5850 4735
rect 5800 4685 5850 4715
rect 5800 4665 5815 4685
rect 5835 4665 5850 4685
rect 5800 4635 5850 4665
rect 5800 4615 5815 4635
rect 5835 4615 5850 4635
rect 5800 4600 5850 4615
rect 5950 5085 6000 5100
rect 5950 5065 5965 5085
rect 5985 5065 6000 5085
rect 5950 5035 6000 5065
rect 5950 5015 5965 5035
rect 5985 5015 6000 5035
rect 5950 4985 6000 5015
rect 5950 4965 5965 4985
rect 5985 4965 6000 4985
rect 5950 4935 6000 4965
rect 5950 4915 5965 4935
rect 5985 4915 6000 4935
rect 5950 4885 6000 4915
rect 5950 4865 5965 4885
rect 5985 4865 6000 4885
rect 5950 4835 6000 4865
rect 5950 4815 5965 4835
rect 5985 4815 6000 4835
rect 5950 4785 6000 4815
rect 5950 4765 5965 4785
rect 5985 4765 6000 4785
rect 5950 4735 6000 4765
rect 5950 4715 5965 4735
rect 5985 4715 6000 4735
rect 5950 4685 6000 4715
rect 5950 4665 5965 4685
rect 5985 4665 6000 4685
rect 5950 4635 6000 4665
rect 5950 4615 5965 4635
rect 5985 4615 6000 4635
rect 5950 4600 6000 4615
rect 6100 5085 6150 5100
rect 6100 5065 6115 5085
rect 6135 5065 6150 5085
rect 6100 5035 6150 5065
rect 6100 5015 6115 5035
rect 6135 5015 6150 5035
rect 6100 4985 6150 5015
rect 6100 4965 6115 4985
rect 6135 4965 6150 4985
rect 6100 4935 6150 4965
rect 6100 4915 6115 4935
rect 6135 4915 6150 4935
rect 6100 4885 6150 4915
rect 6100 4865 6115 4885
rect 6135 4865 6150 4885
rect 6100 4835 6150 4865
rect 6100 4815 6115 4835
rect 6135 4815 6150 4835
rect 6100 4785 6150 4815
rect 6100 4765 6115 4785
rect 6135 4765 6150 4785
rect 6100 4735 6150 4765
rect 6100 4715 6115 4735
rect 6135 4715 6150 4735
rect 6100 4685 6150 4715
rect 6100 4665 6115 4685
rect 6135 4665 6150 4685
rect 6100 4635 6150 4665
rect 6100 4615 6115 4635
rect 6135 4615 6150 4635
rect 6100 4600 6150 4615
rect 6250 5085 6300 5100
rect 6250 5065 6265 5085
rect 6285 5065 6300 5085
rect 6250 5035 6300 5065
rect 6250 5015 6265 5035
rect 6285 5015 6300 5035
rect 6250 4985 6300 5015
rect 6250 4965 6265 4985
rect 6285 4965 6300 4985
rect 6250 4935 6300 4965
rect 6250 4915 6265 4935
rect 6285 4915 6300 4935
rect 6250 4885 6300 4915
rect 6250 4865 6265 4885
rect 6285 4865 6300 4885
rect 6250 4835 6300 4865
rect 6250 4815 6265 4835
rect 6285 4815 6300 4835
rect 6250 4785 6300 4815
rect 6250 4765 6265 4785
rect 6285 4765 6300 4785
rect 6250 4735 6300 4765
rect 6250 4715 6265 4735
rect 6285 4715 6300 4735
rect 6250 4685 6300 4715
rect 6250 4665 6265 4685
rect 6285 4665 6300 4685
rect 6250 4635 6300 4665
rect 6250 4615 6265 4635
rect 6285 4615 6300 4635
rect 6250 4600 6300 4615
rect 6400 5085 6450 5100
rect 6400 5065 6415 5085
rect 6435 5065 6450 5085
rect 6400 5035 6450 5065
rect 6400 5015 6415 5035
rect 6435 5015 6450 5035
rect 6400 4985 6450 5015
rect 6400 4965 6415 4985
rect 6435 4965 6450 4985
rect 6400 4935 6450 4965
rect 6400 4915 6415 4935
rect 6435 4915 6450 4935
rect 6400 4885 6450 4915
rect 6400 4865 6415 4885
rect 6435 4865 6450 4885
rect 6400 4835 6450 4865
rect 6400 4815 6415 4835
rect 6435 4815 6450 4835
rect 6400 4785 6450 4815
rect 6400 4765 6415 4785
rect 6435 4765 6450 4785
rect 6400 4735 6450 4765
rect 6400 4715 6415 4735
rect 6435 4715 6450 4735
rect 6400 4685 6450 4715
rect 6400 4665 6415 4685
rect 6435 4665 6450 4685
rect 6400 4635 6450 4665
rect 6400 4615 6415 4635
rect 6435 4615 6450 4635
rect 6400 4600 6450 4615
rect 6550 5085 6600 5100
rect 6550 5065 6565 5085
rect 6585 5065 6600 5085
rect 6550 5035 6600 5065
rect 6550 5015 6565 5035
rect 6585 5015 6600 5035
rect 6550 4985 6600 5015
rect 6550 4965 6565 4985
rect 6585 4965 6600 4985
rect 6550 4935 6600 4965
rect 6550 4915 6565 4935
rect 6585 4915 6600 4935
rect 6550 4885 6600 4915
rect 6550 4865 6565 4885
rect 6585 4865 6600 4885
rect 6550 4835 6600 4865
rect 6550 4815 6565 4835
rect 6585 4815 6600 4835
rect 6550 4785 6600 4815
rect 6550 4765 6565 4785
rect 6585 4765 6600 4785
rect 6550 4735 6600 4765
rect 6550 4715 6565 4735
rect 6585 4715 6600 4735
rect 6550 4685 6600 4715
rect 6550 4665 6565 4685
rect 6585 4665 6600 4685
rect 6550 4635 6600 4665
rect 6550 4615 6565 4635
rect 6585 4615 6600 4635
rect 6550 4600 6600 4615
rect 6700 5085 6750 5100
rect 6700 5065 6715 5085
rect 6735 5065 6750 5085
rect 6700 5035 6750 5065
rect 6700 5015 6715 5035
rect 6735 5015 6750 5035
rect 6700 4985 6750 5015
rect 6700 4965 6715 4985
rect 6735 4965 6750 4985
rect 6700 4935 6750 4965
rect 6700 4915 6715 4935
rect 6735 4915 6750 4935
rect 6700 4885 6750 4915
rect 6700 4865 6715 4885
rect 6735 4865 6750 4885
rect 6700 4835 6750 4865
rect 6700 4815 6715 4835
rect 6735 4815 6750 4835
rect 6700 4785 6750 4815
rect 6700 4765 6715 4785
rect 6735 4765 6750 4785
rect 6700 4735 6750 4765
rect 6700 4715 6715 4735
rect 6735 4715 6750 4735
rect 6700 4685 6750 4715
rect 6700 4665 6715 4685
rect 6735 4665 6750 4685
rect 6700 4635 6750 4665
rect 6700 4615 6715 4635
rect 6735 4615 6750 4635
rect 6700 4600 6750 4615
rect 6850 5085 6900 5100
rect 6850 5065 6865 5085
rect 6885 5065 6900 5085
rect 6850 5035 6900 5065
rect 6850 5015 6865 5035
rect 6885 5015 6900 5035
rect 6850 4985 6900 5015
rect 6850 4965 6865 4985
rect 6885 4965 6900 4985
rect 6850 4935 6900 4965
rect 6850 4915 6865 4935
rect 6885 4915 6900 4935
rect 6850 4885 6900 4915
rect 6850 4865 6865 4885
rect 6885 4865 6900 4885
rect 6850 4835 6900 4865
rect 6850 4815 6865 4835
rect 6885 4815 6900 4835
rect 6850 4785 6900 4815
rect 6850 4765 6865 4785
rect 6885 4765 6900 4785
rect 6850 4735 6900 4765
rect 6850 4715 6865 4735
rect 6885 4715 6900 4735
rect 6850 4685 6900 4715
rect 6850 4665 6865 4685
rect 6885 4665 6900 4685
rect 6850 4635 6900 4665
rect 6850 4615 6865 4635
rect 6885 4615 6900 4635
rect 6850 4600 6900 4615
rect 7000 5085 7050 5100
rect 7000 5065 7015 5085
rect 7035 5065 7050 5085
rect 7000 5035 7050 5065
rect 7000 5015 7015 5035
rect 7035 5015 7050 5035
rect 7000 4985 7050 5015
rect 7000 4965 7015 4985
rect 7035 4965 7050 4985
rect 7000 4935 7050 4965
rect 7000 4915 7015 4935
rect 7035 4915 7050 4935
rect 7000 4885 7050 4915
rect 7000 4865 7015 4885
rect 7035 4865 7050 4885
rect 7000 4835 7050 4865
rect 7000 4815 7015 4835
rect 7035 4815 7050 4835
rect 7000 4785 7050 4815
rect 7000 4765 7015 4785
rect 7035 4765 7050 4785
rect 7000 4735 7050 4765
rect 7000 4715 7015 4735
rect 7035 4715 7050 4735
rect 7000 4685 7050 4715
rect 7000 4665 7015 4685
rect 7035 4665 7050 4685
rect 7000 4635 7050 4665
rect 7000 4615 7015 4635
rect 7035 4615 7050 4635
rect 7000 4600 7050 4615
rect 7150 5085 7200 5100
rect 7150 5065 7165 5085
rect 7185 5065 7200 5085
rect 7150 5035 7200 5065
rect 7150 5015 7165 5035
rect 7185 5015 7200 5035
rect 7150 4985 7200 5015
rect 7150 4965 7165 4985
rect 7185 4965 7200 4985
rect 7150 4935 7200 4965
rect 7150 4915 7165 4935
rect 7185 4915 7200 4935
rect 7150 4885 7200 4915
rect 7150 4865 7165 4885
rect 7185 4865 7200 4885
rect 7150 4835 7200 4865
rect 7150 4815 7165 4835
rect 7185 4815 7200 4835
rect 7150 4785 7200 4815
rect 7150 4765 7165 4785
rect 7185 4765 7200 4785
rect 7150 4735 7200 4765
rect 7150 4715 7165 4735
rect 7185 4715 7200 4735
rect 7150 4685 7200 4715
rect 7150 4665 7165 4685
rect 7185 4665 7200 4685
rect 7150 4635 7200 4665
rect 7150 4615 7165 4635
rect 7185 4615 7200 4635
rect 7150 4600 7200 4615
rect 7300 5085 7350 5100
rect 7300 5065 7315 5085
rect 7335 5065 7350 5085
rect 7300 5035 7350 5065
rect 7300 5015 7315 5035
rect 7335 5015 7350 5035
rect 7300 4985 7350 5015
rect 7300 4965 7315 4985
rect 7335 4965 7350 4985
rect 7300 4935 7350 4965
rect 7300 4915 7315 4935
rect 7335 4915 7350 4935
rect 7300 4885 7350 4915
rect 7300 4865 7315 4885
rect 7335 4865 7350 4885
rect 7300 4835 7350 4865
rect 7300 4815 7315 4835
rect 7335 4815 7350 4835
rect 7300 4785 7350 4815
rect 7300 4765 7315 4785
rect 7335 4765 7350 4785
rect 7300 4735 7350 4765
rect 7300 4715 7315 4735
rect 7335 4715 7350 4735
rect 7300 4685 7350 4715
rect 7300 4665 7315 4685
rect 7335 4665 7350 4685
rect 7300 4635 7350 4665
rect 7300 4615 7315 4635
rect 7335 4615 7350 4635
rect 7300 4600 7350 4615
rect 7450 5085 7500 5100
rect 7450 5065 7465 5085
rect 7485 5065 7500 5085
rect 7450 5035 7500 5065
rect 7450 5015 7465 5035
rect 7485 5015 7500 5035
rect 7450 4985 7500 5015
rect 7450 4965 7465 4985
rect 7485 4965 7500 4985
rect 7450 4935 7500 4965
rect 7450 4915 7465 4935
rect 7485 4915 7500 4935
rect 7450 4885 7500 4915
rect 7450 4865 7465 4885
rect 7485 4865 7500 4885
rect 7450 4835 7500 4865
rect 7450 4815 7465 4835
rect 7485 4815 7500 4835
rect 7450 4785 7500 4815
rect 7450 4765 7465 4785
rect 7485 4765 7500 4785
rect 7450 4735 7500 4765
rect 7450 4715 7465 4735
rect 7485 4715 7500 4735
rect 7450 4685 7500 4715
rect 7450 4665 7465 4685
rect 7485 4665 7500 4685
rect 7450 4635 7500 4665
rect 7450 4615 7465 4635
rect 7485 4615 7500 4635
rect 7450 4600 7500 4615
rect 7600 5085 7650 5100
rect 7600 5065 7615 5085
rect 7635 5065 7650 5085
rect 7600 5035 7650 5065
rect 7600 5015 7615 5035
rect 7635 5015 7650 5035
rect 7600 4985 7650 5015
rect 7600 4965 7615 4985
rect 7635 4965 7650 4985
rect 7600 4935 7650 4965
rect 7600 4915 7615 4935
rect 7635 4915 7650 4935
rect 7600 4885 7650 4915
rect 7600 4865 7615 4885
rect 7635 4865 7650 4885
rect 7600 4835 7650 4865
rect 7600 4815 7615 4835
rect 7635 4815 7650 4835
rect 7600 4785 7650 4815
rect 7600 4765 7615 4785
rect 7635 4765 7650 4785
rect 7600 4735 7650 4765
rect 7600 4715 7615 4735
rect 7635 4715 7650 4735
rect 7600 4685 7650 4715
rect 7600 4665 7615 4685
rect 7635 4665 7650 4685
rect 7600 4635 7650 4665
rect 7600 4615 7615 4635
rect 7635 4615 7650 4635
rect 7600 4600 7650 4615
rect 7750 5085 7800 5100
rect 7750 5065 7765 5085
rect 7785 5065 7800 5085
rect 7750 5035 7800 5065
rect 7750 5015 7765 5035
rect 7785 5015 7800 5035
rect 7750 4985 7800 5015
rect 7750 4965 7765 4985
rect 7785 4965 7800 4985
rect 7750 4935 7800 4965
rect 7750 4915 7765 4935
rect 7785 4915 7800 4935
rect 7750 4885 7800 4915
rect 7750 4865 7765 4885
rect 7785 4865 7800 4885
rect 7750 4835 7800 4865
rect 7750 4815 7765 4835
rect 7785 4815 7800 4835
rect 7750 4785 7800 4815
rect 7750 4765 7765 4785
rect 7785 4765 7800 4785
rect 7750 4735 7800 4765
rect 7750 4715 7765 4735
rect 7785 4715 7800 4735
rect 7750 4685 7800 4715
rect 7750 4665 7765 4685
rect 7785 4665 7800 4685
rect 7750 4635 7800 4665
rect 7750 4615 7765 4635
rect 7785 4615 7800 4635
rect 7750 4600 7800 4615
rect 8350 5085 8400 5100
rect 8350 5065 8365 5085
rect 8385 5065 8400 5085
rect 8350 5035 8400 5065
rect 8350 5015 8365 5035
rect 8385 5015 8400 5035
rect 8350 4985 8400 5015
rect 8350 4965 8365 4985
rect 8385 4965 8400 4985
rect 8350 4935 8400 4965
rect 8350 4915 8365 4935
rect 8385 4915 8400 4935
rect 8350 4885 8400 4915
rect 8350 4865 8365 4885
rect 8385 4865 8400 4885
rect 8350 4835 8400 4865
rect 8350 4815 8365 4835
rect 8385 4815 8400 4835
rect 8350 4785 8400 4815
rect 8350 4765 8365 4785
rect 8385 4765 8400 4785
rect 8350 4735 8400 4765
rect 8350 4715 8365 4735
rect 8385 4715 8400 4735
rect 8350 4685 8400 4715
rect 8350 4665 8365 4685
rect 8385 4665 8400 4685
rect 8350 4635 8400 4665
rect 8350 4615 8365 4635
rect 8385 4615 8400 4635
rect 8350 4600 8400 4615
rect 8500 5085 8550 5100
rect 8500 5065 8515 5085
rect 8535 5065 8550 5085
rect 8500 5035 8550 5065
rect 8500 5015 8515 5035
rect 8535 5015 8550 5035
rect 8500 4985 8550 5015
rect 8500 4965 8515 4985
rect 8535 4965 8550 4985
rect 8500 4935 8550 4965
rect 8500 4915 8515 4935
rect 8535 4915 8550 4935
rect 8500 4885 8550 4915
rect 8500 4865 8515 4885
rect 8535 4865 8550 4885
rect 8500 4835 8550 4865
rect 8500 4815 8515 4835
rect 8535 4815 8550 4835
rect 8500 4785 8550 4815
rect 8500 4765 8515 4785
rect 8535 4765 8550 4785
rect 8500 4735 8550 4765
rect 8500 4715 8515 4735
rect 8535 4715 8550 4735
rect 8500 4685 8550 4715
rect 8500 4665 8515 4685
rect 8535 4665 8550 4685
rect 8500 4635 8550 4665
rect 8500 4615 8515 4635
rect 8535 4615 8550 4635
rect 8500 4550 8550 4615
rect 8650 5085 8700 5100
rect 8650 5065 8665 5085
rect 8685 5065 8700 5085
rect 8650 5035 8700 5065
rect 8650 5015 8665 5035
rect 8685 5015 8700 5035
rect 8650 4985 8700 5015
rect 8650 4965 8665 4985
rect 8685 4965 8700 4985
rect 8650 4935 8700 4965
rect 8650 4915 8665 4935
rect 8685 4915 8700 4935
rect 8650 4885 8700 4915
rect 8650 4865 8665 4885
rect 8685 4865 8700 4885
rect 8650 4835 8700 4865
rect 8650 4815 8665 4835
rect 8685 4815 8700 4835
rect 8650 4785 8700 4815
rect 8650 4765 8665 4785
rect 8685 4765 8700 4785
rect 8650 4735 8700 4765
rect 8650 4715 8665 4735
rect 8685 4715 8700 4735
rect 8650 4685 8700 4715
rect 8650 4665 8665 4685
rect 8685 4665 8700 4685
rect 8650 4635 8700 4665
rect 8650 4615 8665 4635
rect 8685 4615 8700 4635
rect 8650 4600 8700 4615
rect 8800 5085 8850 5100
rect 8800 5065 8815 5085
rect 8835 5065 8850 5085
rect 8800 5035 8850 5065
rect 8800 5015 8815 5035
rect 8835 5015 8850 5035
rect 8800 4985 8850 5015
rect 8800 4965 8815 4985
rect 8835 4965 8850 4985
rect 8800 4935 8850 4965
rect 8800 4915 8815 4935
rect 8835 4915 8850 4935
rect 8800 4885 8850 4915
rect 8800 4865 8815 4885
rect 8835 4865 8850 4885
rect 8800 4835 8850 4865
rect 8800 4815 8815 4835
rect 8835 4815 8850 4835
rect 8800 4785 8850 4815
rect 8800 4765 8815 4785
rect 8835 4765 8850 4785
rect 8800 4735 8850 4765
rect 8800 4715 8815 4735
rect 8835 4715 8850 4735
rect 8800 4685 8850 4715
rect 8800 4665 8815 4685
rect 8835 4665 8850 4685
rect 8800 4635 8850 4665
rect 8800 4615 8815 4635
rect 8835 4615 8850 4635
rect 8800 4550 8850 4615
rect 8950 5085 9000 5100
rect 8950 5065 8965 5085
rect 8985 5065 9000 5085
rect 8950 5035 9000 5065
rect 8950 5015 8965 5035
rect 8985 5015 9000 5035
rect 8950 4985 9000 5015
rect 8950 4965 8965 4985
rect 8985 4965 9000 4985
rect 8950 4935 9000 4965
rect 8950 4915 8965 4935
rect 8985 4915 9000 4935
rect 8950 4885 9000 4915
rect 8950 4865 8965 4885
rect 8985 4865 9000 4885
rect 8950 4835 9000 4865
rect 8950 4815 8965 4835
rect 8985 4815 9000 4835
rect 8950 4785 9000 4815
rect 8950 4765 8965 4785
rect 8985 4765 9000 4785
rect 8950 4735 9000 4765
rect 8950 4715 8965 4735
rect 8985 4715 9000 4735
rect 8950 4685 9000 4715
rect 8950 4665 8965 4685
rect 8985 4665 9000 4685
rect 8950 4635 9000 4665
rect 8950 4615 8965 4635
rect 8985 4615 9000 4635
rect 8950 4600 9000 4615
rect 9100 5085 9150 5100
rect 9100 5065 9115 5085
rect 9135 5065 9150 5085
rect 9100 5035 9150 5065
rect 9100 5015 9115 5035
rect 9135 5015 9150 5035
rect 9100 4985 9150 5015
rect 9100 4965 9115 4985
rect 9135 4965 9150 4985
rect 9100 4935 9150 4965
rect 9100 4915 9115 4935
rect 9135 4915 9150 4935
rect 9100 4885 9150 4915
rect 9100 4865 9115 4885
rect 9135 4865 9150 4885
rect 9100 4835 9150 4865
rect 9100 4815 9115 4835
rect 9135 4815 9150 4835
rect 9100 4785 9150 4815
rect 9100 4765 9115 4785
rect 9135 4765 9150 4785
rect 9100 4735 9150 4765
rect 9100 4715 9115 4735
rect 9135 4715 9150 4735
rect 9100 4685 9150 4715
rect 9100 4665 9115 4685
rect 9135 4665 9150 4685
rect 9100 4635 9150 4665
rect 9100 4615 9115 4635
rect 9135 4615 9150 4635
rect 9100 4550 9150 4615
rect 9250 5085 9300 5100
rect 9250 5065 9265 5085
rect 9285 5065 9300 5085
rect 9250 5035 9300 5065
rect 9250 5015 9265 5035
rect 9285 5015 9300 5035
rect 9250 4985 9300 5015
rect 9250 4965 9265 4985
rect 9285 4965 9300 4985
rect 9250 4935 9300 4965
rect 9250 4915 9265 4935
rect 9285 4915 9300 4935
rect 9250 4885 9300 4915
rect 9250 4865 9265 4885
rect 9285 4865 9300 4885
rect 9250 4835 9300 4865
rect 9250 4815 9265 4835
rect 9285 4815 9300 4835
rect 9250 4785 9300 4815
rect 9250 4765 9265 4785
rect 9285 4765 9300 4785
rect 9250 4735 9300 4765
rect 9250 4715 9265 4735
rect 9285 4715 9300 4735
rect 9250 4685 9300 4715
rect 9250 4665 9265 4685
rect 9285 4665 9300 4685
rect 9250 4635 9300 4665
rect 9250 4615 9265 4635
rect 9285 4615 9300 4635
rect 9250 4600 9300 4615
rect 9400 5085 9450 5100
rect 9400 5065 9415 5085
rect 9435 5065 9450 5085
rect 9400 5035 9450 5065
rect 9400 5015 9415 5035
rect 9435 5015 9450 5035
rect 9400 4985 9450 5015
rect 9400 4965 9415 4985
rect 9435 4965 9450 4985
rect 9400 4935 9450 4965
rect 9400 4915 9415 4935
rect 9435 4915 9450 4935
rect 9400 4885 9450 4915
rect 9400 4865 9415 4885
rect 9435 4865 9450 4885
rect 9400 4835 9450 4865
rect 9400 4815 9415 4835
rect 9435 4815 9450 4835
rect 9400 4785 9450 4815
rect 9400 4765 9415 4785
rect 9435 4765 9450 4785
rect 9400 4735 9450 4765
rect 9400 4715 9415 4735
rect 9435 4715 9450 4735
rect 9400 4685 9450 4715
rect 9400 4665 9415 4685
rect 9435 4665 9450 4685
rect 9400 4635 9450 4665
rect 9400 4615 9415 4635
rect 9435 4615 9450 4635
rect 9400 4550 9450 4615
rect 9550 5085 9600 5100
rect 9550 5065 9565 5085
rect 9585 5065 9600 5085
rect 9550 5035 9600 5065
rect 9550 5015 9565 5035
rect 9585 5015 9600 5035
rect 9550 4985 9600 5015
rect 9550 4965 9565 4985
rect 9585 4965 9600 4985
rect 9550 4935 9600 4965
rect 9550 4915 9565 4935
rect 9585 4915 9600 4935
rect 9550 4885 9600 4915
rect 9550 4865 9565 4885
rect 9585 4865 9600 4885
rect 9550 4835 9600 4865
rect 9550 4815 9565 4835
rect 9585 4815 9600 4835
rect 9550 4785 9600 4815
rect 9550 4765 9565 4785
rect 9585 4765 9600 4785
rect 9550 4735 9600 4765
rect 9550 4715 9565 4735
rect 9585 4715 9600 4735
rect 9550 4685 9600 4715
rect 9550 4665 9565 4685
rect 9585 4665 9600 4685
rect 9550 4635 9600 4665
rect 9550 4615 9565 4635
rect 9585 4615 9600 4635
rect 9550 4600 9600 4615
rect 9700 5085 9750 5100
rect 9700 5065 9715 5085
rect 9735 5065 9750 5085
rect 9700 5035 9750 5065
rect 9700 5015 9715 5035
rect 9735 5015 9750 5035
rect 9700 4985 9750 5015
rect 9700 4965 9715 4985
rect 9735 4965 9750 4985
rect 9700 4935 9750 4965
rect 9700 4915 9715 4935
rect 9735 4915 9750 4935
rect 9700 4885 9750 4915
rect 9700 4865 9715 4885
rect 9735 4865 9750 4885
rect 9700 4835 9750 4865
rect 9700 4815 9715 4835
rect 9735 4815 9750 4835
rect 9700 4785 9750 4815
rect 9700 4765 9715 4785
rect 9735 4765 9750 4785
rect 9700 4735 9750 4765
rect 9700 4715 9715 4735
rect 9735 4715 9750 4735
rect 9700 4685 9750 4715
rect 9700 4665 9715 4685
rect 9735 4665 9750 4685
rect 9700 4635 9750 4665
rect 9700 4615 9715 4635
rect 9735 4615 9750 4635
rect 9700 4550 9750 4615
rect 9850 5085 9900 5100
rect 9850 5065 9865 5085
rect 9885 5065 9900 5085
rect 9850 5035 9900 5065
rect 9850 5015 9865 5035
rect 9885 5015 9900 5035
rect 9850 4985 9900 5015
rect 9850 4965 9865 4985
rect 9885 4965 9900 4985
rect 9850 4935 9900 4965
rect 9850 4915 9865 4935
rect 9885 4915 9900 4935
rect 9850 4885 9900 4915
rect 9850 4865 9865 4885
rect 9885 4865 9900 4885
rect 9850 4835 9900 4865
rect 9850 4815 9865 4835
rect 9885 4815 9900 4835
rect 9850 4785 9900 4815
rect 9850 4765 9865 4785
rect 9885 4765 9900 4785
rect 9850 4735 9900 4765
rect 9850 4715 9865 4735
rect 9885 4715 9900 4735
rect 9850 4685 9900 4715
rect 9850 4665 9865 4685
rect 9885 4665 9900 4685
rect 9850 4635 9900 4665
rect 9850 4615 9865 4635
rect 9885 4615 9900 4635
rect 9850 4600 9900 4615
rect 10000 5085 10050 5100
rect 10000 5065 10015 5085
rect 10035 5065 10050 5085
rect 10000 5035 10050 5065
rect 10000 5015 10015 5035
rect 10035 5015 10050 5035
rect 10000 4985 10050 5015
rect 10000 4965 10015 4985
rect 10035 4965 10050 4985
rect 10000 4935 10050 4965
rect 10000 4915 10015 4935
rect 10035 4915 10050 4935
rect 10000 4885 10050 4915
rect 10000 4865 10015 4885
rect 10035 4865 10050 4885
rect 10000 4835 10050 4865
rect 10000 4815 10015 4835
rect 10035 4815 10050 4835
rect 10000 4785 10050 4815
rect 10000 4765 10015 4785
rect 10035 4765 10050 4785
rect 10000 4735 10050 4765
rect 10000 4715 10015 4735
rect 10035 4715 10050 4735
rect 10000 4685 10050 4715
rect 10000 4665 10015 4685
rect 10035 4665 10050 4685
rect 10000 4635 10050 4665
rect 10000 4615 10015 4635
rect 10035 4615 10050 4635
rect 10000 4550 10050 4615
rect 10150 5085 10200 5100
rect 10150 5065 10165 5085
rect 10185 5065 10200 5085
rect 10150 5035 10200 5065
rect 10150 5015 10165 5035
rect 10185 5015 10200 5035
rect 10150 4985 10200 5015
rect 10150 4965 10165 4985
rect 10185 4965 10200 4985
rect 10150 4935 10200 4965
rect 10150 4915 10165 4935
rect 10185 4915 10200 4935
rect 10150 4885 10200 4915
rect 10150 4865 10165 4885
rect 10185 4865 10200 4885
rect 10150 4835 10200 4865
rect 10150 4815 10165 4835
rect 10185 4815 10200 4835
rect 10150 4785 10200 4815
rect 10150 4765 10165 4785
rect 10185 4765 10200 4785
rect 10150 4735 10200 4765
rect 10150 4715 10165 4735
rect 10185 4715 10200 4735
rect 10150 4685 10200 4715
rect 10150 4665 10165 4685
rect 10185 4665 10200 4685
rect 10150 4635 10200 4665
rect 10150 4615 10165 4635
rect 10185 4615 10200 4635
rect 10150 4600 10200 4615
rect 10300 5085 10350 5100
rect 10300 5065 10315 5085
rect 10335 5065 10350 5085
rect 10300 5035 10350 5065
rect 10300 5015 10315 5035
rect 10335 5015 10350 5035
rect 10300 4985 10350 5015
rect 10300 4965 10315 4985
rect 10335 4965 10350 4985
rect 10300 4935 10350 4965
rect 10300 4915 10315 4935
rect 10335 4915 10350 4935
rect 10300 4885 10350 4915
rect 10300 4865 10315 4885
rect 10335 4865 10350 4885
rect 10300 4835 10350 4865
rect 10300 4815 10315 4835
rect 10335 4815 10350 4835
rect 10300 4785 10350 4815
rect 10300 4765 10315 4785
rect 10335 4765 10350 4785
rect 10300 4735 10350 4765
rect 10300 4715 10315 4735
rect 10335 4715 10350 4735
rect 10300 4685 10350 4715
rect 10300 4665 10315 4685
rect 10335 4665 10350 4685
rect 10300 4635 10350 4665
rect 10300 4615 10315 4635
rect 10335 4615 10350 4635
rect 10300 4550 10350 4615
rect 10450 5085 10500 5100
rect 10450 5065 10465 5085
rect 10485 5065 10500 5085
rect 10450 5035 10500 5065
rect 10450 5015 10465 5035
rect 10485 5015 10500 5035
rect 10450 4985 10500 5015
rect 10450 4965 10465 4985
rect 10485 4965 10500 4985
rect 10450 4935 10500 4965
rect 10450 4915 10465 4935
rect 10485 4915 10500 4935
rect 10450 4885 10500 4915
rect 10450 4865 10465 4885
rect 10485 4865 10500 4885
rect 10450 4835 10500 4865
rect 10450 4815 10465 4835
rect 10485 4815 10500 4835
rect 10450 4785 10500 4815
rect 10450 4765 10465 4785
rect 10485 4765 10500 4785
rect 10450 4735 10500 4765
rect 10450 4715 10465 4735
rect 10485 4715 10500 4735
rect 10450 4685 10500 4715
rect 10450 4665 10465 4685
rect 10485 4665 10500 4685
rect 10450 4635 10500 4665
rect 10450 4615 10465 4635
rect 10485 4615 10500 4635
rect 10450 4600 10500 4615
rect 10600 5085 10650 5100
rect 10600 5065 10615 5085
rect 10635 5065 10650 5085
rect 10600 5035 10650 5065
rect 10600 5015 10615 5035
rect 10635 5015 10650 5035
rect 10600 4985 10650 5015
rect 10600 4965 10615 4985
rect 10635 4965 10650 4985
rect 10600 4935 10650 4965
rect 10600 4915 10615 4935
rect 10635 4915 10650 4935
rect 10600 4885 10650 4915
rect 10600 4865 10615 4885
rect 10635 4865 10650 4885
rect 10600 4835 10650 4865
rect 10600 4815 10615 4835
rect 10635 4815 10650 4835
rect 10600 4785 10650 4815
rect 10600 4765 10615 4785
rect 10635 4765 10650 4785
rect 10600 4735 10650 4765
rect 10600 4715 10615 4735
rect 10635 4715 10650 4735
rect 10600 4685 10650 4715
rect 10600 4665 10615 4685
rect 10635 4665 10650 4685
rect 10600 4635 10650 4665
rect 10600 4615 10615 4635
rect 10635 4615 10650 4635
rect 10600 4550 10650 4615
rect 10750 5085 10800 5100
rect 10750 5065 10765 5085
rect 10785 5065 10800 5085
rect 10750 5035 10800 5065
rect 10750 5015 10765 5035
rect 10785 5015 10800 5035
rect 10750 4985 10800 5015
rect 10750 4965 10765 4985
rect 10785 4965 10800 4985
rect 10750 4935 10800 4965
rect 10750 4915 10765 4935
rect 10785 4915 10800 4935
rect 10750 4885 10800 4915
rect 10750 4865 10765 4885
rect 10785 4865 10800 4885
rect 10750 4835 10800 4865
rect 10750 4815 10765 4835
rect 10785 4815 10800 4835
rect 10750 4785 10800 4815
rect 10750 4765 10765 4785
rect 10785 4765 10800 4785
rect 10750 4735 10800 4765
rect 10750 4715 10765 4735
rect 10785 4715 10800 4735
rect 10750 4685 10800 4715
rect 10750 4665 10765 4685
rect 10785 4665 10800 4685
rect 10750 4635 10800 4665
rect 10750 4615 10765 4635
rect 10785 4615 10800 4635
rect 10750 4600 10800 4615
rect 11350 5085 11400 5100
rect 11350 5065 11365 5085
rect 11385 5065 11400 5085
rect 11350 5035 11400 5065
rect 11350 5015 11365 5035
rect 11385 5015 11400 5035
rect 11350 4985 11400 5015
rect 11350 4965 11365 4985
rect 11385 4965 11400 4985
rect 11350 4935 11400 4965
rect 11350 4915 11365 4935
rect 11385 4915 11400 4935
rect 11350 4885 11400 4915
rect 11350 4865 11365 4885
rect 11385 4865 11400 4885
rect 11350 4835 11400 4865
rect 11350 4815 11365 4835
rect 11385 4815 11400 4835
rect 11350 4785 11400 4815
rect 11350 4765 11365 4785
rect 11385 4765 11400 4785
rect 11350 4735 11400 4765
rect 11350 4715 11365 4735
rect 11385 4715 11400 4735
rect 11350 4685 11400 4715
rect 11350 4665 11365 4685
rect 11385 4665 11400 4685
rect 11350 4635 11400 4665
rect 11350 4615 11365 4635
rect 11385 4615 11400 4635
rect 11350 4600 11400 4615
rect 11950 5085 12000 5100
rect 11950 5065 11965 5085
rect 11985 5065 12000 5085
rect 11950 5035 12000 5065
rect 11950 5015 11965 5035
rect 11985 5015 12000 5035
rect 11950 4985 12000 5015
rect 11950 4965 11965 4985
rect 11985 4965 12000 4985
rect 11950 4935 12000 4965
rect 11950 4915 11965 4935
rect 11985 4915 12000 4935
rect 11950 4885 12000 4915
rect 11950 4865 11965 4885
rect 11985 4865 12000 4885
rect 11950 4835 12000 4865
rect 11950 4815 11965 4835
rect 11985 4815 12000 4835
rect 11950 4785 12000 4815
rect 11950 4765 11965 4785
rect 11985 4765 12000 4785
rect 11950 4735 12000 4765
rect 11950 4715 11965 4735
rect 11985 4715 12000 4735
rect 11950 4685 12000 4715
rect 11950 4665 11965 4685
rect 11985 4665 12000 4685
rect 11950 4635 12000 4665
rect 11950 4615 11965 4635
rect 11985 4615 12000 4635
rect 11950 4600 12000 4615
rect 12550 5085 12600 5100
rect 12550 5065 12565 5085
rect 12585 5065 12600 5085
rect 12550 5035 12600 5065
rect 12550 5015 12565 5035
rect 12585 5015 12600 5035
rect 12550 4985 12600 5015
rect 12550 4965 12565 4985
rect 12585 4965 12600 4985
rect 12550 4935 12600 4965
rect 12550 4915 12565 4935
rect 12585 4915 12600 4935
rect 12550 4885 12600 4915
rect 12550 4865 12565 4885
rect 12585 4865 12600 4885
rect 12550 4835 12600 4865
rect 12550 4815 12565 4835
rect 12585 4815 12600 4835
rect 12550 4785 12600 4815
rect 12550 4765 12565 4785
rect 12585 4765 12600 4785
rect 12550 4735 12600 4765
rect 12550 4715 12565 4735
rect 12585 4715 12600 4735
rect 12550 4685 12600 4715
rect 12550 4665 12565 4685
rect 12585 4665 12600 4685
rect 12550 4635 12600 4665
rect 12550 4615 12565 4635
rect 12585 4615 12600 4635
rect 12550 4600 12600 4615
rect 13150 5085 13200 5100
rect 13150 5065 13165 5085
rect 13185 5065 13200 5085
rect 13150 5035 13200 5065
rect 13150 5015 13165 5035
rect 13185 5015 13200 5035
rect 13150 4985 13200 5015
rect 13150 4965 13165 4985
rect 13185 4965 13200 4985
rect 13150 4935 13200 4965
rect 13150 4915 13165 4935
rect 13185 4915 13200 4935
rect 13150 4885 13200 4915
rect 13150 4865 13165 4885
rect 13185 4865 13200 4885
rect 13150 4835 13200 4865
rect 13150 4815 13165 4835
rect 13185 4815 13200 4835
rect 13150 4785 13200 4815
rect 13150 4765 13165 4785
rect 13185 4765 13200 4785
rect 13150 4735 13200 4765
rect 13150 4715 13165 4735
rect 13185 4715 13200 4735
rect 13150 4685 13200 4715
rect 13150 4665 13165 4685
rect 13185 4665 13200 4685
rect 13150 4635 13200 4665
rect 13150 4615 13165 4635
rect 13185 4615 13200 4635
rect 13150 4600 13200 4615
rect 13750 5085 13800 5100
rect 13750 5065 13765 5085
rect 13785 5065 13800 5085
rect 13750 5035 13800 5065
rect 13750 5015 13765 5035
rect 13785 5015 13800 5035
rect 13750 4985 13800 5015
rect 13750 4965 13765 4985
rect 13785 4965 13800 4985
rect 13750 4935 13800 4965
rect 13750 4915 13765 4935
rect 13785 4915 13800 4935
rect 13750 4885 13800 4915
rect 13750 4865 13765 4885
rect 13785 4865 13800 4885
rect 13750 4835 13800 4865
rect 13750 4815 13765 4835
rect 13785 4815 13800 4835
rect 13750 4785 13800 4815
rect 13750 4765 13765 4785
rect 13785 4765 13800 4785
rect 13750 4735 13800 4765
rect 13750 4715 13765 4735
rect 13785 4715 13800 4735
rect 13750 4685 13800 4715
rect 13750 4665 13765 4685
rect 13785 4665 13800 4685
rect 13750 4635 13800 4665
rect 13750 4615 13765 4635
rect 13785 4615 13800 4635
rect 13750 4600 13800 4615
rect 14350 5085 14400 5100
rect 14350 5065 14365 5085
rect 14385 5065 14400 5085
rect 14350 5035 14400 5065
rect 14350 5015 14365 5035
rect 14385 5015 14400 5035
rect 14350 4985 14400 5015
rect 14350 4965 14365 4985
rect 14385 4965 14400 4985
rect 14350 4935 14400 4965
rect 14350 4915 14365 4935
rect 14385 4915 14400 4935
rect 14350 4885 14400 4915
rect 14350 4865 14365 4885
rect 14385 4865 14400 4885
rect 14350 4835 14400 4865
rect 14350 4815 14365 4835
rect 14385 4815 14400 4835
rect 14350 4785 14400 4815
rect 14350 4765 14365 4785
rect 14385 4765 14400 4785
rect 14350 4735 14400 4765
rect 14350 4715 14365 4735
rect 14385 4715 14400 4735
rect 14350 4685 14400 4715
rect 14350 4665 14365 4685
rect 14385 4665 14400 4685
rect 14350 4635 14400 4665
rect 14350 4615 14365 4635
rect 14385 4615 14400 4635
rect 14350 4600 14400 4615
rect 14950 5085 15000 5100
rect 14950 5065 14965 5085
rect 14985 5065 15000 5085
rect 14950 5035 15000 5065
rect 14950 5015 14965 5035
rect 14985 5015 15000 5035
rect 14950 4985 15000 5015
rect 14950 4965 14965 4985
rect 14985 4965 15000 4985
rect 14950 4935 15000 4965
rect 14950 4915 14965 4935
rect 14985 4915 15000 4935
rect 14950 4885 15000 4915
rect 14950 4865 14965 4885
rect 14985 4865 15000 4885
rect 14950 4835 15000 4865
rect 14950 4815 14965 4835
rect 14985 4815 15000 4835
rect 14950 4785 15000 4815
rect 14950 4765 14965 4785
rect 14985 4765 15000 4785
rect 14950 4735 15000 4765
rect 14950 4715 14965 4735
rect 14985 4715 15000 4735
rect 14950 4685 15000 4715
rect 14950 4665 14965 4685
rect 14985 4665 15000 4685
rect 14950 4635 15000 4665
rect 14950 4615 14965 4635
rect 14985 4615 15000 4635
rect 14950 4600 15000 4615
rect 15550 5085 15600 5100
rect 15550 5065 15565 5085
rect 15585 5065 15600 5085
rect 15550 5035 15600 5065
rect 15550 5015 15565 5035
rect 15585 5015 15600 5035
rect 15550 4985 15600 5015
rect 15550 4965 15565 4985
rect 15585 4965 15600 4985
rect 15550 4935 15600 4965
rect 15550 4915 15565 4935
rect 15585 4915 15600 4935
rect 15550 4885 15600 4915
rect 15550 4865 15565 4885
rect 15585 4865 15600 4885
rect 15550 4835 15600 4865
rect 15550 4815 15565 4835
rect 15585 4815 15600 4835
rect 15550 4785 15600 4815
rect 15550 4765 15565 4785
rect 15585 4765 15600 4785
rect 15550 4735 15600 4765
rect 15550 4715 15565 4735
rect 15585 4715 15600 4735
rect 15550 4685 15600 4715
rect 15550 4665 15565 4685
rect 15585 4665 15600 4685
rect 15550 4635 15600 4665
rect 15550 4615 15565 4635
rect 15585 4615 15600 4635
rect 15550 4600 15600 4615
rect 16150 5085 16200 5100
rect 16150 5065 16165 5085
rect 16185 5065 16200 5085
rect 16150 5035 16200 5065
rect 16150 5015 16165 5035
rect 16185 5015 16200 5035
rect 16150 4985 16200 5015
rect 16150 4965 16165 4985
rect 16185 4965 16200 4985
rect 16150 4935 16200 4965
rect 16150 4915 16165 4935
rect 16185 4915 16200 4935
rect 16150 4885 16200 4915
rect 16150 4865 16165 4885
rect 16185 4865 16200 4885
rect 16150 4835 16200 4865
rect 16150 4815 16165 4835
rect 16185 4815 16200 4835
rect 16150 4785 16200 4815
rect 16150 4765 16165 4785
rect 16185 4765 16200 4785
rect 16150 4735 16200 4765
rect 16150 4715 16165 4735
rect 16185 4715 16200 4735
rect 16150 4685 16200 4715
rect 16150 4665 16165 4685
rect 16185 4665 16200 4685
rect 16150 4635 16200 4665
rect 16150 4615 16165 4635
rect 16185 4615 16200 4635
rect 16150 4600 16200 4615
rect 16300 5085 16350 5100
rect 16300 5065 16315 5085
rect 16335 5065 16350 5085
rect 16300 5035 16350 5065
rect 16300 5015 16315 5035
rect 16335 5015 16350 5035
rect 16300 4985 16350 5015
rect 16300 4965 16315 4985
rect 16335 4965 16350 4985
rect 16300 4935 16350 4965
rect 16300 4915 16315 4935
rect 16335 4915 16350 4935
rect 16300 4885 16350 4915
rect 16300 4865 16315 4885
rect 16335 4865 16350 4885
rect 16300 4835 16350 4865
rect 16300 4815 16315 4835
rect 16335 4815 16350 4835
rect 16300 4785 16350 4815
rect 16300 4765 16315 4785
rect 16335 4765 16350 4785
rect 16300 4735 16350 4765
rect 16300 4715 16315 4735
rect 16335 4715 16350 4735
rect 16300 4685 16350 4715
rect 16300 4665 16315 4685
rect 16335 4665 16350 4685
rect 16300 4635 16350 4665
rect 16300 4615 16315 4635
rect 16335 4615 16350 4635
rect 16300 4600 16350 4615
rect 16450 5085 16500 5100
rect 16450 5065 16465 5085
rect 16485 5065 16500 5085
rect 16450 5035 16500 5065
rect 16450 5015 16465 5035
rect 16485 5015 16500 5035
rect 16450 4985 16500 5015
rect 16450 4965 16465 4985
rect 16485 4965 16500 4985
rect 16450 4935 16500 4965
rect 16450 4915 16465 4935
rect 16485 4915 16500 4935
rect 16450 4885 16500 4915
rect 16450 4865 16465 4885
rect 16485 4865 16500 4885
rect 16450 4835 16500 4865
rect 16450 4815 16465 4835
rect 16485 4815 16500 4835
rect 16450 4785 16500 4815
rect 16450 4765 16465 4785
rect 16485 4765 16500 4785
rect 16450 4735 16500 4765
rect 16450 4715 16465 4735
rect 16485 4715 16500 4735
rect 16450 4685 16500 4715
rect 16450 4665 16465 4685
rect 16485 4665 16500 4685
rect 16450 4635 16500 4665
rect 16450 4615 16465 4635
rect 16485 4615 16500 4635
rect 16450 4600 16500 4615
rect 16600 5085 16650 5100
rect 16600 5065 16615 5085
rect 16635 5065 16650 5085
rect 16600 5035 16650 5065
rect 16600 5015 16615 5035
rect 16635 5015 16650 5035
rect 16600 4985 16650 5015
rect 16600 4965 16615 4985
rect 16635 4965 16650 4985
rect 16600 4935 16650 4965
rect 16600 4915 16615 4935
rect 16635 4915 16650 4935
rect 16600 4885 16650 4915
rect 16600 4865 16615 4885
rect 16635 4865 16650 4885
rect 16600 4835 16650 4865
rect 16600 4815 16615 4835
rect 16635 4815 16650 4835
rect 16600 4785 16650 4815
rect 16600 4765 16615 4785
rect 16635 4765 16650 4785
rect 16600 4735 16650 4765
rect 16600 4715 16615 4735
rect 16635 4715 16650 4735
rect 16600 4685 16650 4715
rect 16600 4665 16615 4685
rect 16635 4665 16650 4685
rect 16600 4635 16650 4665
rect 16600 4615 16615 4635
rect 16635 4615 16650 4635
rect 16600 4600 16650 4615
rect 16750 5085 16800 5100
rect 16750 5065 16765 5085
rect 16785 5065 16800 5085
rect 16750 5035 16800 5065
rect 16750 5015 16765 5035
rect 16785 5015 16800 5035
rect 16750 4985 16800 5015
rect 16750 4965 16765 4985
rect 16785 4965 16800 4985
rect 16750 4935 16800 4965
rect 16750 4915 16765 4935
rect 16785 4915 16800 4935
rect 16750 4885 16800 4915
rect 16750 4865 16765 4885
rect 16785 4865 16800 4885
rect 16750 4835 16800 4865
rect 16750 4815 16765 4835
rect 16785 4815 16800 4835
rect 16750 4785 16800 4815
rect 16750 4765 16765 4785
rect 16785 4765 16800 4785
rect 16750 4735 16800 4765
rect 16750 4715 16765 4735
rect 16785 4715 16800 4735
rect 16750 4685 16800 4715
rect 16750 4665 16765 4685
rect 16785 4665 16800 4685
rect 16750 4635 16800 4665
rect 16750 4615 16765 4635
rect 16785 4615 16800 4635
rect 16750 4600 16800 4615
rect 16900 5085 16950 5100
rect 16900 5065 16915 5085
rect 16935 5065 16950 5085
rect 16900 5035 16950 5065
rect 16900 5015 16915 5035
rect 16935 5015 16950 5035
rect 16900 4985 16950 5015
rect 16900 4965 16915 4985
rect 16935 4965 16950 4985
rect 16900 4935 16950 4965
rect 16900 4915 16915 4935
rect 16935 4915 16950 4935
rect 16900 4885 16950 4915
rect 16900 4865 16915 4885
rect 16935 4865 16950 4885
rect 16900 4835 16950 4865
rect 16900 4815 16915 4835
rect 16935 4815 16950 4835
rect 16900 4785 16950 4815
rect 16900 4765 16915 4785
rect 16935 4765 16950 4785
rect 16900 4735 16950 4765
rect 16900 4715 16915 4735
rect 16935 4715 16950 4735
rect 16900 4685 16950 4715
rect 16900 4665 16915 4685
rect 16935 4665 16950 4685
rect 16900 4635 16950 4665
rect 16900 4615 16915 4635
rect 16935 4615 16950 4635
rect 16900 4600 16950 4615
rect 17050 5085 17100 5100
rect 17050 5065 17065 5085
rect 17085 5065 17100 5085
rect 17050 5035 17100 5065
rect 17050 5015 17065 5035
rect 17085 5015 17100 5035
rect 17050 4985 17100 5015
rect 17050 4965 17065 4985
rect 17085 4965 17100 4985
rect 17050 4935 17100 4965
rect 17050 4915 17065 4935
rect 17085 4915 17100 4935
rect 17050 4885 17100 4915
rect 17050 4865 17065 4885
rect 17085 4865 17100 4885
rect 17050 4835 17100 4865
rect 17050 4815 17065 4835
rect 17085 4815 17100 4835
rect 17050 4785 17100 4815
rect 17050 4765 17065 4785
rect 17085 4765 17100 4785
rect 17050 4735 17100 4765
rect 17050 4715 17065 4735
rect 17085 4715 17100 4735
rect 17050 4685 17100 4715
rect 17050 4665 17065 4685
rect 17085 4665 17100 4685
rect 17050 4635 17100 4665
rect 17050 4615 17065 4635
rect 17085 4615 17100 4635
rect 17050 4600 17100 4615
rect 17200 5085 17250 5100
rect 17200 5065 17215 5085
rect 17235 5065 17250 5085
rect 17200 5035 17250 5065
rect 17200 5015 17215 5035
rect 17235 5015 17250 5035
rect 17200 4985 17250 5015
rect 17200 4965 17215 4985
rect 17235 4965 17250 4985
rect 17200 4935 17250 4965
rect 17200 4915 17215 4935
rect 17235 4915 17250 4935
rect 17200 4885 17250 4915
rect 17200 4865 17215 4885
rect 17235 4865 17250 4885
rect 17200 4835 17250 4865
rect 17200 4815 17215 4835
rect 17235 4815 17250 4835
rect 17200 4785 17250 4815
rect 17200 4765 17215 4785
rect 17235 4765 17250 4785
rect 17200 4735 17250 4765
rect 17200 4715 17215 4735
rect 17235 4715 17250 4735
rect 17200 4685 17250 4715
rect 17200 4665 17215 4685
rect 17235 4665 17250 4685
rect 17200 4635 17250 4665
rect 17200 4615 17215 4635
rect 17235 4615 17250 4635
rect 17200 4600 17250 4615
rect 17350 5085 17400 5100
rect 17350 5065 17365 5085
rect 17385 5065 17400 5085
rect 17350 5035 17400 5065
rect 17350 5015 17365 5035
rect 17385 5015 17400 5035
rect 17350 4985 17400 5015
rect 17350 4965 17365 4985
rect 17385 4965 17400 4985
rect 17350 4935 17400 4965
rect 17350 4915 17365 4935
rect 17385 4915 17400 4935
rect 17350 4885 17400 4915
rect 17350 4865 17365 4885
rect 17385 4865 17400 4885
rect 17350 4835 17400 4865
rect 17350 4815 17365 4835
rect 17385 4815 17400 4835
rect 17350 4785 17400 4815
rect 17350 4765 17365 4785
rect 17385 4765 17400 4785
rect 17350 4735 17400 4765
rect 17350 4715 17365 4735
rect 17385 4715 17400 4735
rect 17350 4685 17400 4715
rect 17350 4665 17365 4685
rect 17385 4665 17400 4685
rect 17350 4635 17400 4665
rect 17350 4615 17365 4635
rect 17385 4615 17400 4635
rect 17350 4600 17400 4615
rect 17950 5085 18000 5100
rect 17950 5065 17965 5085
rect 17985 5065 18000 5085
rect 17950 5035 18000 5065
rect 17950 5015 17965 5035
rect 17985 5015 18000 5035
rect 17950 4985 18000 5015
rect 17950 4965 17965 4985
rect 17985 4965 18000 4985
rect 17950 4935 18000 4965
rect 17950 4915 17965 4935
rect 17985 4915 18000 4935
rect 17950 4885 18000 4915
rect 17950 4865 17965 4885
rect 17985 4865 18000 4885
rect 17950 4835 18000 4865
rect 17950 4815 17965 4835
rect 17985 4815 18000 4835
rect 17950 4785 18000 4815
rect 17950 4765 17965 4785
rect 17985 4765 18000 4785
rect 17950 4735 18000 4765
rect 17950 4715 17965 4735
rect 17985 4715 18000 4735
rect 17950 4685 18000 4715
rect 17950 4665 17965 4685
rect 17985 4665 18000 4685
rect 17950 4635 18000 4665
rect 17950 4615 17965 4635
rect 17985 4615 18000 4635
rect 17950 4600 18000 4615
rect 18550 5085 18600 5100
rect 18550 5065 18565 5085
rect 18585 5065 18600 5085
rect 18550 5035 18600 5065
rect 18550 5015 18565 5035
rect 18585 5015 18600 5035
rect 18550 4985 18600 5015
rect 18550 4965 18565 4985
rect 18585 4965 18600 4985
rect 18550 4935 18600 4965
rect 18550 4915 18565 4935
rect 18585 4915 18600 4935
rect 18550 4885 18600 4915
rect 18550 4865 18565 4885
rect 18585 4865 18600 4885
rect 18550 4835 18600 4865
rect 18550 4815 18565 4835
rect 18585 4815 18600 4835
rect 18550 4785 18600 4815
rect 18550 4765 18565 4785
rect 18585 4765 18600 4785
rect 18550 4735 18600 4765
rect 18550 4715 18565 4735
rect 18585 4715 18600 4735
rect 18550 4685 18600 4715
rect 18550 4665 18565 4685
rect 18585 4665 18600 4685
rect 18550 4635 18600 4665
rect 18550 4615 18565 4635
rect 18585 4615 18600 4635
rect 18550 4600 18600 4615
rect 18700 5085 18750 5100
rect 18700 5065 18715 5085
rect 18735 5065 18750 5085
rect 18700 5035 18750 5065
rect 18700 5015 18715 5035
rect 18735 5015 18750 5035
rect 18700 4985 18750 5015
rect 18700 4965 18715 4985
rect 18735 4965 18750 4985
rect 18700 4935 18750 4965
rect 18700 4915 18715 4935
rect 18735 4915 18750 4935
rect 18700 4885 18750 4915
rect 18700 4865 18715 4885
rect 18735 4865 18750 4885
rect 18700 4835 18750 4865
rect 18700 4815 18715 4835
rect 18735 4815 18750 4835
rect 18700 4785 18750 4815
rect 18700 4765 18715 4785
rect 18735 4765 18750 4785
rect 18700 4735 18750 4765
rect 18700 4715 18715 4735
rect 18735 4715 18750 4735
rect 18700 4685 18750 4715
rect 18700 4665 18715 4685
rect 18735 4665 18750 4685
rect 18700 4635 18750 4665
rect 18700 4615 18715 4635
rect 18735 4615 18750 4635
rect 18700 4600 18750 4615
rect 18850 5085 18900 5100
rect 18850 5065 18865 5085
rect 18885 5065 18900 5085
rect 18850 5035 18900 5065
rect 18850 5015 18865 5035
rect 18885 5015 18900 5035
rect 18850 4985 18900 5015
rect 18850 4965 18865 4985
rect 18885 4965 18900 4985
rect 18850 4935 18900 4965
rect 18850 4915 18865 4935
rect 18885 4915 18900 4935
rect 18850 4885 18900 4915
rect 18850 4865 18865 4885
rect 18885 4865 18900 4885
rect 18850 4835 18900 4865
rect 18850 4815 18865 4835
rect 18885 4815 18900 4835
rect 18850 4785 18900 4815
rect 18850 4765 18865 4785
rect 18885 4765 18900 4785
rect 18850 4735 18900 4765
rect 18850 4715 18865 4735
rect 18885 4715 18900 4735
rect 18850 4685 18900 4715
rect 18850 4665 18865 4685
rect 18885 4665 18900 4685
rect 18850 4635 18900 4665
rect 18850 4615 18865 4635
rect 18885 4615 18900 4635
rect 18850 4600 18900 4615
rect 19000 5085 19050 5100
rect 19000 5065 19015 5085
rect 19035 5065 19050 5085
rect 19000 5035 19050 5065
rect 19000 5015 19015 5035
rect 19035 5015 19050 5035
rect 19000 4985 19050 5015
rect 19000 4965 19015 4985
rect 19035 4965 19050 4985
rect 19000 4935 19050 4965
rect 19000 4915 19015 4935
rect 19035 4915 19050 4935
rect 19000 4885 19050 4915
rect 19000 4865 19015 4885
rect 19035 4865 19050 4885
rect 19000 4835 19050 4865
rect 19000 4815 19015 4835
rect 19035 4815 19050 4835
rect 19000 4785 19050 4815
rect 19000 4765 19015 4785
rect 19035 4765 19050 4785
rect 19000 4735 19050 4765
rect 19000 4715 19015 4735
rect 19035 4715 19050 4735
rect 19000 4685 19050 4715
rect 19000 4665 19015 4685
rect 19035 4665 19050 4685
rect 19000 4635 19050 4665
rect 19000 4615 19015 4635
rect 19035 4615 19050 4635
rect 19000 4600 19050 4615
rect 19150 5085 19200 5100
rect 19150 5065 19165 5085
rect 19185 5065 19200 5085
rect 19150 5035 19200 5065
rect 19150 5015 19165 5035
rect 19185 5015 19200 5035
rect 19150 4985 19200 5015
rect 19150 4965 19165 4985
rect 19185 4965 19200 4985
rect 19150 4935 19200 4965
rect 19150 4915 19165 4935
rect 19185 4915 19200 4935
rect 19150 4885 19200 4915
rect 19150 4865 19165 4885
rect 19185 4865 19200 4885
rect 19150 4835 19200 4865
rect 19150 4815 19165 4835
rect 19185 4815 19200 4835
rect 19150 4785 19200 4815
rect 19150 4765 19165 4785
rect 19185 4765 19200 4785
rect 19150 4735 19200 4765
rect 19150 4715 19165 4735
rect 19185 4715 19200 4735
rect 19150 4685 19200 4715
rect 19150 4665 19165 4685
rect 19185 4665 19200 4685
rect 19150 4635 19200 4665
rect 19150 4615 19165 4635
rect 19185 4615 19200 4635
rect 19150 4600 19200 4615
rect 19300 5085 19350 5100
rect 19300 5065 19315 5085
rect 19335 5065 19350 5085
rect 19300 5035 19350 5065
rect 19300 5015 19315 5035
rect 19335 5015 19350 5035
rect 19300 4985 19350 5015
rect 19300 4965 19315 4985
rect 19335 4965 19350 4985
rect 19300 4935 19350 4965
rect 19300 4915 19315 4935
rect 19335 4915 19350 4935
rect 19300 4885 19350 4915
rect 19300 4865 19315 4885
rect 19335 4865 19350 4885
rect 19300 4835 19350 4865
rect 19300 4815 19315 4835
rect 19335 4815 19350 4835
rect 19300 4785 19350 4815
rect 19300 4765 19315 4785
rect 19335 4765 19350 4785
rect 19300 4735 19350 4765
rect 19300 4715 19315 4735
rect 19335 4715 19350 4735
rect 19300 4685 19350 4715
rect 19300 4665 19315 4685
rect 19335 4665 19350 4685
rect 19300 4635 19350 4665
rect 19300 4615 19315 4635
rect 19335 4615 19350 4635
rect 19300 4600 19350 4615
rect 19450 5085 19500 5100
rect 19450 5065 19465 5085
rect 19485 5065 19500 5085
rect 19450 5035 19500 5065
rect 19450 5015 19465 5035
rect 19485 5015 19500 5035
rect 19450 4985 19500 5015
rect 19450 4965 19465 4985
rect 19485 4965 19500 4985
rect 19450 4935 19500 4965
rect 19450 4915 19465 4935
rect 19485 4915 19500 4935
rect 19450 4885 19500 4915
rect 19450 4865 19465 4885
rect 19485 4865 19500 4885
rect 19450 4835 19500 4865
rect 19450 4815 19465 4835
rect 19485 4815 19500 4835
rect 19450 4785 19500 4815
rect 19450 4765 19465 4785
rect 19485 4765 19500 4785
rect 19450 4735 19500 4765
rect 19450 4715 19465 4735
rect 19485 4715 19500 4735
rect 19450 4685 19500 4715
rect 19450 4665 19465 4685
rect 19485 4665 19500 4685
rect 19450 4635 19500 4665
rect 19450 4615 19465 4635
rect 19485 4615 19500 4635
rect 19450 4600 19500 4615
rect 19600 5085 19650 5100
rect 19600 5065 19615 5085
rect 19635 5065 19650 5085
rect 19600 5035 19650 5065
rect 19600 5015 19615 5035
rect 19635 5015 19650 5035
rect 19600 4985 19650 5015
rect 19600 4965 19615 4985
rect 19635 4965 19650 4985
rect 19600 4935 19650 4965
rect 19600 4915 19615 4935
rect 19635 4915 19650 4935
rect 19600 4885 19650 4915
rect 19600 4865 19615 4885
rect 19635 4865 19650 4885
rect 19600 4835 19650 4865
rect 19600 4815 19615 4835
rect 19635 4815 19650 4835
rect 19600 4785 19650 4815
rect 19600 4765 19615 4785
rect 19635 4765 19650 4785
rect 19600 4735 19650 4765
rect 19600 4715 19615 4735
rect 19635 4715 19650 4735
rect 19600 4685 19650 4715
rect 19600 4665 19615 4685
rect 19635 4665 19650 4685
rect 19600 4635 19650 4665
rect 19600 4615 19615 4635
rect 19635 4615 19650 4635
rect 19600 4600 19650 4615
rect 19750 5085 19800 5100
rect 19750 5065 19765 5085
rect 19785 5065 19800 5085
rect 19750 5035 19800 5065
rect 19750 5015 19765 5035
rect 19785 5015 19800 5035
rect 19750 4985 19800 5015
rect 19750 4965 19765 4985
rect 19785 4965 19800 4985
rect 19750 4935 19800 4965
rect 19750 4915 19765 4935
rect 19785 4915 19800 4935
rect 19750 4885 19800 4915
rect 19750 4865 19765 4885
rect 19785 4865 19800 4885
rect 19750 4835 19800 4865
rect 19750 4815 19765 4835
rect 19785 4815 19800 4835
rect 19750 4785 19800 4815
rect 19750 4765 19765 4785
rect 19785 4765 19800 4785
rect 19750 4735 19800 4765
rect 19750 4715 19765 4735
rect 19785 4715 19800 4735
rect 19750 4685 19800 4715
rect 19750 4665 19765 4685
rect 19785 4665 19800 4685
rect 19750 4635 19800 4665
rect 19750 4615 19765 4635
rect 19785 4615 19800 4635
rect 19750 4600 19800 4615
rect 20350 5085 20400 5100
rect 20350 5065 20365 5085
rect 20385 5065 20400 5085
rect 20350 5035 20400 5065
rect 20350 5015 20365 5035
rect 20385 5015 20400 5035
rect 20350 4985 20400 5015
rect 20350 4965 20365 4985
rect 20385 4965 20400 4985
rect 20350 4935 20400 4965
rect 20350 4915 20365 4935
rect 20385 4915 20400 4935
rect 20350 4885 20400 4915
rect 20350 4865 20365 4885
rect 20385 4865 20400 4885
rect 20350 4835 20400 4865
rect 20350 4815 20365 4835
rect 20385 4815 20400 4835
rect 20350 4785 20400 4815
rect 20350 4765 20365 4785
rect 20385 4765 20400 4785
rect 20350 4735 20400 4765
rect 20350 4715 20365 4735
rect 20385 4715 20400 4735
rect 20350 4685 20400 4715
rect 20350 4665 20365 4685
rect 20385 4665 20400 4685
rect 20350 4635 20400 4665
rect 20350 4615 20365 4635
rect 20385 4615 20400 4635
rect 20350 4600 20400 4615
rect -600 4535 -350 4550
rect -600 4515 -585 4535
rect -565 4515 -535 4535
rect -515 4515 -485 4535
rect -465 4515 -435 4535
rect -415 4515 -385 4535
rect -365 4515 -350 4535
rect -600 4500 -350 4515
rect -300 4535 -50 4550
rect -300 4515 -285 4535
rect -265 4515 -235 4535
rect -215 4515 -185 4535
rect -165 4515 -135 4535
rect -115 4515 -85 4535
rect -65 4515 -50 4535
rect -300 4500 -50 4515
rect 0 4535 250 4550
rect 0 4515 15 4535
rect 35 4515 65 4535
rect 85 4515 115 4535
rect 135 4515 165 4535
rect 185 4515 215 4535
rect 235 4515 250 4535
rect 0 4500 250 4515
rect 300 4535 550 4550
rect 300 4515 315 4535
rect 335 4515 365 4535
rect 385 4515 415 4535
rect 435 4515 465 4535
rect 485 4515 515 4535
rect 535 4515 550 4535
rect 300 4500 550 4515
rect 600 4535 850 4550
rect 600 4515 615 4535
rect 635 4515 665 4535
rect 685 4515 715 4535
rect 735 4515 765 4535
rect 785 4515 815 4535
rect 835 4515 850 4535
rect 600 4500 850 4515
rect 900 4535 1150 4550
rect 900 4515 915 4535
rect 935 4515 965 4535
rect 985 4515 1015 4535
rect 1035 4515 1065 4535
rect 1085 4515 1115 4535
rect 1135 4515 1150 4535
rect 900 4500 1150 4515
rect 1200 4535 1450 4550
rect 1200 4515 1215 4535
rect 1235 4515 1265 4535
rect 1285 4515 1315 4535
rect 1335 4515 1365 4535
rect 1385 4515 1415 4535
rect 1435 4515 1450 4535
rect 1200 4500 1450 4515
rect 1500 4535 1750 4550
rect 1500 4515 1515 4535
rect 1535 4515 1565 4535
rect 1585 4515 1615 4535
rect 1635 4515 1665 4535
rect 1685 4515 1715 4535
rect 1735 4515 1750 4535
rect 1500 4500 1750 4515
rect 1800 4535 2050 4550
rect 1800 4515 1815 4535
rect 1835 4515 1865 4535
rect 1885 4515 1915 4535
rect 1935 4515 1965 4535
rect 1985 4515 2015 4535
rect 2035 4515 2050 4535
rect 1800 4500 2050 4515
rect 2100 4535 2350 4550
rect 2100 4515 2115 4535
rect 2135 4515 2165 4535
rect 2185 4515 2215 4535
rect 2235 4515 2265 4535
rect 2285 4515 2315 4535
rect 2335 4515 2350 4535
rect 2100 4500 2350 4515
rect 2400 4535 2650 4550
rect 2400 4515 2415 4535
rect 2435 4515 2465 4535
rect 2485 4515 2515 4535
rect 2535 4515 2565 4535
rect 2585 4515 2615 4535
rect 2635 4515 2650 4535
rect 2400 4500 2650 4515
rect 2700 4535 2950 4550
rect 2700 4515 2715 4535
rect 2735 4515 2765 4535
rect 2785 4515 2815 4535
rect 2835 4515 2865 4535
rect 2885 4515 2915 4535
rect 2935 4515 2950 4535
rect 2700 4500 2950 4515
rect 3000 4535 3250 4550
rect 3000 4515 3015 4535
rect 3035 4515 3065 4535
rect 3085 4515 3115 4535
rect 3135 4515 3165 4535
rect 3185 4515 3215 4535
rect 3235 4515 3250 4535
rect 3000 4500 3250 4515
rect 3300 4535 3550 4550
rect 3300 4515 3315 4535
rect 3335 4515 3365 4535
rect 3385 4515 3415 4535
rect 3435 4515 3465 4535
rect 3485 4515 3515 4535
rect 3535 4515 3550 4535
rect 3300 4500 3550 4515
rect 3600 4535 3850 4550
rect 3600 4515 3615 4535
rect 3635 4515 3665 4535
rect 3685 4515 3715 4535
rect 3735 4515 3765 4535
rect 3785 4515 3815 4535
rect 3835 4515 3850 4535
rect 3600 4500 3850 4515
rect 3900 4535 4150 4550
rect 3900 4515 3915 4535
rect 3935 4515 3965 4535
rect 3985 4515 4015 4535
rect 4035 4515 4065 4535
rect 4085 4515 4115 4535
rect 4135 4515 4150 4535
rect 3900 4500 4150 4515
rect 4200 4535 4450 4550
rect 4200 4515 4215 4535
rect 4235 4515 4265 4535
rect 4285 4515 4315 4535
rect 4335 4515 4365 4535
rect 4385 4515 4415 4535
rect 4435 4515 4450 4535
rect 4200 4500 4450 4515
rect 4500 4535 4750 4550
rect 4500 4515 4515 4535
rect 4535 4515 4565 4535
rect 4585 4515 4615 4535
rect 4635 4515 4665 4535
rect 4685 4515 4715 4535
rect 4735 4515 4750 4535
rect 4500 4500 4750 4515
rect 4800 4535 5050 4550
rect 4800 4515 4815 4535
rect 4835 4515 4865 4535
rect 4885 4515 4915 4535
rect 4935 4515 4965 4535
rect 4985 4515 5015 4535
rect 5035 4515 5050 4535
rect 4800 4500 5050 4515
rect 5100 4535 5350 4550
rect 5100 4515 5115 4535
rect 5135 4515 5165 4535
rect 5185 4515 5215 4535
rect 5235 4515 5265 4535
rect 5285 4515 5315 4535
rect 5335 4515 5350 4535
rect 5100 4500 5350 4515
rect 5400 4535 5650 4550
rect 5400 4515 5415 4535
rect 5435 4515 5465 4535
rect 5485 4515 5515 4535
rect 5535 4515 5565 4535
rect 5585 4515 5615 4535
rect 5635 4515 5650 4535
rect 5400 4500 5650 4515
rect 5700 4535 5950 4550
rect 5700 4515 5715 4535
rect 5735 4515 5765 4535
rect 5785 4515 5815 4535
rect 5835 4515 5865 4535
rect 5885 4515 5915 4535
rect 5935 4515 5950 4535
rect 5700 4500 5950 4515
rect 6000 4535 6250 4550
rect 6000 4515 6015 4535
rect 6035 4515 6065 4535
rect 6085 4515 6115 4535
rect 6135 4515 6165 4535
rect 6185 4515 6215 4535
rect 6235 4515 6250 4535
rect 6000 4500 6250 4515
rect 6300 4535 6550 4550
rect 6300 4515 6315 4535
rect 6335 4515 6365 4535
rect 6385 4515 6415 4535
rect 6435 4515 6465 4535
rect 6485 4515 6515 4535
rect 6535 4515 6550 4535
rect 6300 4500 6550 4515
rect 6600 4535 6850 4550
rect 6600 4515 6615 4535
rect 6635 4515 6665 4535
rect 6685 4515 6715 4535
rect 6735 4515 6765 4535
rect 6785 4515 6815 4535
rect 6835 4515 6850 4535
rect 6600 4500 6850 4515
rect 6900 4535 7150 4550
rect 6900 4515 6915 4535
rect 6935 4515 6965 4535
rect 6985 4515 7015 4535
rect 7035 4515 7065 4535
rect 7085 4515 7115 4535
rect 7135 4515 7150 4535
rect 6900 4500 7150 4515
rect 7200 4535 7450 4550
rect 7200 4515 7215 4535
rect 7235 4515 7265 4535
rect 7285 4515 7315 4535
rect 7335 4515 7365 4535
rect 7385 4515 7415 4535
rect 7435 4515 7450 4535
rect 7200 4500 7450 4515
rect 7500 4535 7750 4550
rect 7500 4515 7515 4535
rect 7535 4515 7565 4535
rect 7585 4515 7615 4535
rect 7635 4515 7665 4535
rect 7685 4515 7715 4535
rect 7735 4515 7750 4535
rect 7500 4500 7750 4515
rect 7800 4535 8050 4550
rect 7800 4515 7815 4535
rect 7835 4515 7865 4535
rect 7885 4515 7915 4535
rect 7935 4515 7965 4535
rect 7985 4515 8015 4535
rect 8035 4515 8050 4535
rect 7800 4500 8050 4515
rect 8100 4535 8350 4550
rect 8100 4515 8115 4535
rect 8135 4515 8165 4535
rect 8185 4515 8215 4535
rect 8235 4515 8265 4535
rect 8285 4515 8315 4535
rect 8335 4515 8350 4535
rect 8100 4500 8350 4515
rect 8400 4535 10750 4550
rect 8400 4515 8415 4535
rect 8435 4515 8465 4535
rect 8485 4515 8515 4535
rect 8535 4515 8565 4535
rect 8585 4515 8615 4535
rect 8635 4515 8715 4535
rect 8735 4515 8765 4535
rect 8785 4515 8815 4535
rect 8835 4515 8865 4535
rect 8885 4515 8915 4535
rect 8935 4515 9015 4535
rect 9035 4515 9065 4535
rect 9085 4515 9115 4535
rect 9135 4515 9165 4535
rect 9185 4515 9215 4535
rect 9235 4515 9315 4535
rect 9335 4515 9365 4535
rect 9385 4515 9415 4535
rect 9435 4515 9465 4535
rect 9485 4515 9515 4535
rect 9535 4515 9615 4535
rect 9635 4515 9665 4535
rect 9685 4515 9715 4535
rect 9735 4515 9765 4535
rect 9785 4515 9815 4535
rect 9835 4515 9915 4535
rect 9935 4515 9965 4535
rect 9985 4515 10015 4535
rect 10035 4515 10065 4535
rect 10085 4515 10115 4535
rect 10135 4515 10215 4535
rect 10235 4515 10265 4535
rect 10285 4515 10315 4535
rect 10335 4515 10365 4535
rect 10385 4515 10415 4535
rect 10435 4515 10515 4535
rect 10535 4515 10565 4535
rect 10585 4515 10615 4535
rect 10635 4515 10665 4535
rect 10685 4515 10715 4535
rect 10735 4515 10750 4535
rect 8400 4500 10750 4515
rect 10800 4535 11050 4550
rect 10800 4515 10815 4535
rect 10835 4515 10865 4535
rect 10885 4515 10915 4535
rect 10935 4515 10965 4535
rect 10985 4515 11015 4535
rect 11035 4515 11050 4535
rect 10800 4500 11050 4515
rect 11100 4535 11350 4550
rect 11100 4515 11115 4535
rect 11135 4515 11165 4535
rect 11185 4515 11215 4535
rect 11235 4515 11265 4535
rect 11285 4515 11315 4535
rect 11335 4515 11350 4535
rect 11100 4500 11350 4515
rect 11400 4535 11650 4550
rect 11400 4515 11415 4535
rect 11435 4515 11465 4535
rect 11485 4515 11515 4535
rect 11535 4515 11565 4535
rect 11585 4515 11615 4535
rect 11635 4515 11650 4535
rect 11400 4500 11650 4515
rect 11700 4535 11950 4550
rect 11700 4515 11715 4535
rect 11735 4515 11765 4535
rect 11785 4515 11815 4535
rect 11835 4515 11865 4535
rect 11885 4515 11915 4535
rect 11935 4515 11950 4535
rect 11700 4500 11950 4515
rect 12000 4535 12250 4550
rect 12000 4515 12015 4535
rect 12035 4515 12065 4535
rect 12085 4515 12115 4535
rect 12135 4515 12165 4535
rect 12185 4515 12215 4535
rect 12235 4515 12250 4535
rect 12000 4500 12250 4515
rect 12300 4535 12550 4550
rect 12300 4515 12315 4535
rect 12335 4515 12365 4535
rect 12385 4515 12415 4535
rect 12435 4515 12465 4535
rect 12485 4515 12515 4535
rect 12535 4515 12550 4535
rect 12300 4500 12550 4515
rect 12600 4535 12850 4550
rect 12600 4515 12615 4535
rect 12635 4515 12665 4535
rect 12685 4515 12715 4535
rect 12735 4515 12765 4535
rect 12785 4515 12815 4535
rect 12835 4515 12850 4535
rect 12600 4500 12850 4515
rect 12900 4535 13150 4550
rect 12900 4515 12915 4535
rect 12935 4515 12965 4535
rect 12985 4515 13015 4535
rect 13035 4515 13065 4535
rect 13085 4515 13115 4535
rect 13135 4515 13150 4535
rect 12900 4500 13150 4515
rect 13200 4535 13450 4550
rect 13200 4515 13215 4535
rect 13235 4515 13265 4535
rect 13285 4515 13315 4535
rect 13335 4515 13365 4535
rect 13385 4515 13415 4535
rect 13435 4515 13450 4535
rect 13200 4500 13450 4515
rect 13500 4535 13750 4550
rect 13500 4515 13515 4535
rect 13535 4515 13565 4535
rect 13585 4515 13615 4535
rect 13635 4515 13665 4535
rect 13685 4515 13715 4535
rect 13735 4515 13750 4535
rect 13500 4500 13750 4515
rect 13800 4535 14050 4550
rect 13800 4515 13815 4535
rect 13835 4515 13865 4535
rect 13885 4515 13915 4535
rect 13935 4515 13965 4535
rect 13985 4515 14015 4535
rect 14035 4515 14050 4535
rect 13800 4500 14050 4515
rect 14100 4535 14350 4550
rect 14100 4515 14115 4535
rect 14135 4515 14165 4535
rect 14185 4515 14215 4535
rect 14235 4515 14265 4535
rect 14285 4515 14315 4535
rect 14335 4515 14350 4535
rect 14100 4500 14350 4515
rect 14400 4535 14650 4550
rect 14400 4515 14415 4535
rect 14435 4515 14465 4535
rect 14485 4515 14515 4535
rect 14535 4515 14565 4535
rect 14585 4515 14615 4535
rect 14635 4515 14650 4535
rect 14400 4500 14650 4515
rect 14700 4535 14950 4550
rect 14700 4515 14715 4535
rect 14735 4515 14765 4535
rect 14785 4515 14815 4535
rect 14835 4515 14865 4535
rect 14885 4515 14915 4535
rect 14935 4515 14950 4535
rect 14700 4500 14950 4515
rect 15000 4535 15250 4550
rect 15000 4515 15015 4535
rect 15035 4515 15065 4535
rect 15085 4515 15115 4535
rect 15135 4515 15165 4535
rect 15185 4515 15215 4535
rect 15235 4515 15250 4535
rect 15000 4500 15250 4515
rect 15300 4535 15550 4550
rect 15300 4515 15315 4535
rect 15335 4515 15365 4535
rect 15385 4515 15415 4535
rect 15435 4515 15465 4535
rect 15485 4515 15515 4535
rect 15535 4515 15550 4535
rect 15300 4500 15550 4515
rect 15600 4535 15850 4550
rect 15600 4515 15615 4535
rect 15635 4515 15665 4535
rect 15685 4515 15715 4535
rect 15735 4515 15765 4535
rect 15785 4515 15815 4535
rect 15835 4515 15850 4535
rect 15600 4500 15850 4515
rect 15900 4535 16150 4550
rect 15900 4515 15915 4535
rect 15935 4515 15965 4535
rect 15985 4515 16015 4535
rect 16035 4515 16065 4535
rect 16085 4515 16115 4535
rect 16135 4515 16150 4535
rect 15900 4500 16150 4515
rect 16200 4535 16450 4550
rect 16200 4515 16215 4535
rect 16235 4515 16265 4535
rect 16285 4515 16315 4535
rect 16335 4515 16365 4535
rect 16385 4515 16415 4535
rect 16435 4515 16450 4535
rect 16200 4500 16450 4515
rect 16500 4535 16750 4550
rect 16500 4515 16515 4535
rect 16535 4515 16565 4535
rect 16585 4515 16615 4535
rect 16635 4515 16665 4535
rect 16685 4515 16715 4535
rect 16735 4515 16750 4535
rect 16500 4500 16750 4515
rect 16800 4535 17050 4550
rect 16800 4515 16815 4535
rect 16835 4515 16865 4535
rect 16885 4515 16915 4535
rect 16935 4515 16965 4535
rect 16985 4515 17015 4535
rect 17035 4515 17050 4535
rect 16800 4500 17050 4515
rect 17100 4535 17350 4550
rect 17100 4515 17115 4535
rect 17135 4515 17165 4535
rect 17185 4515 17215 4535
rect 17235 4515 17265 4535
rect 17285 4515 17315 4535
rect 17335 4515 17350 4535
rect 17100 4500 17350 4515
rect 17400 4535 17650 4550
rect 17400 4515 17415 4535
rect 17435 4515 17465 4535
rect 17485 4515 17515 4535
rect 17535 4515 17565 4535
rect 17585 4515 17615 4535
rect 17635 4515 17650 4535
rect 17400 4500 17650 4515
rect 17700 4535 17950 4550
rect 17700 4515 17715 4535
rect 17735 4515 17765 4535
rect 17785 4515 17815 4535
rect 17835 4515 17865 4535
rect 17885 4515 17915 4535
rect 17935 4515 17950 4535
rect 17700 4500 17950 4515
rect 18000 4535 18250 4550
rect 18000 4515 18015 4535
rect 18035 4515 18065 4535
rect 18085 4515 18115 4535
rect 18135 4515 18165 4535
rect 18185 4515 18215 4535
rect 18235 4515 18250 4535
rect 18000 4500 18250 4515
rect 18300 4535 18550 4550
rect 18300 4515 18315 4535
rect 18335 4515 18365 4535
rect 18385 4515 18415 4535
rect 18435 4515 18465 4535
rect 18485 4515 18515 4535
rect 18535 4515 18550 4535
rect 18300 4500 18550 4515
rect 18600 4535 18850 4550
rect 18600 4515 18615 4535
rect 18635 4515 18665 4535
rect 18685 4515 18715 4535
rect 18735 4515 18765 4535
rect 18785 4515 18815 4535
rect 18835 4515 18850 4535
rect 18600 4500 18850 4515
rect 18900 4535 19150 4550
rect 18900 4515 18915 4535
rect 18935 4515 18965 4535
rect 18985 4515 19015 4535
rect 19035 4515 19065 4535
rect 19085 4515 19115 4535
rect 19135 4515 19150 4535
rect 18900 4500 19150 4515
rect 19200 4535 19450 4550
rect 19200 4515 19215 4535
rect 19235 4515 19265 4535
rect 19285 4515 19315 4535
rect 19335 4515 19365 4535
rect 19385 4515 19415 4535
rect 19435 4515 19450 4535
rect 19200 4500 19450 4515
rect 19500 4535 19750 4550
rect 19500 4515 19515 4535
rect 19535 4515 19565 4535
rect 19585 4515 19615 4535
rect 19635 4515 19665 4535
rect 19685 4515 19715 4535
rect 19735 4515 19750 4535
rect 19500 4500 19750 4515
rect 19800 4535 20050 4550
rect 19800 4515 19815 4535
rect 19835 4515 19865 4535
rect 19885 4515 19915 4535
rect 19935 4515 19965 4535
rect 19985 4515 20015 4535
rect 20035 4515 20050 4535
rect 19800 4500 20050 4515
rect 20100 4535 20350 4550
rect 20100 4515 20115 4535
rect 20135 4515 20165 4535
rect 20185 4515 20215 4535
rect 20235 4515 20265 4535
rect 20285 4515 20315 4535
rect 20335 4515 20350 4535
rect 20100 4500 20350 4515
rect -650 4435 -600 4450
rect -650 4415 -635 4435
rect -615 4415 -600 4435
rect -650 4385 -600 4415
rect -650 4365 -635 4385
rect -615 4365 -600 4385
rect -650 4335 -600 4365
rect -650 4315 -635 4335
rect -615 4315 -600 4335
rect -650 4285 -600 4315
rect -650 4265 -635 4285
rect -615 4265 -600 4285
rect -650 4235 -600 4265
rect -650 4215 -635 4235
rect -615 4215 -600 4235
rect -650 4185 -600 4215
rect -650 4165 -635 4185
rect -615 4165 -600 4185
rect -650 4135 -600 4165
rect -650 4115 -635 4135
rect -615 4115 -600 4135
rect -650 4085 -600 4115
rect -650 4065 -635 4085
rect -615 4065 -600 4085
rect -650 4035 -600 4065
rect -650 4015 -635 4035
rect -615 4015 -600 4035
rect -650 3985 -600 4015
rect -650 3965 -635 3985
rect -615 3965 -600 3985
rect -650 3950 -600 3965
rect -500 4435 -450 4450
rect -500 4415 -485 4435
rect -465 4415 -450 4435
rect -500 4385 -450 4415
rect -500 4365 -485 4385
rect -465 4365 -450 4385
rect -500 4335 -450 4365
rect -500 4315 -485 4335
rect -465 4315 -450 4335
rect -500 4285 -450 4315
rect -500 4265 -485 4285
rect -465 4265 -450 4285
rect -500 4235 -450 4265
rect -500 4215 -485 4235
rect -465 4215 -450 4235
rect -500 4185 -450 4215
rect -500 4165 -485 4185
rect -465 4165 -450 4185
rect -500 4135 -450 4165
rect -500 4115 -485 4135
rect -465 4115 -450 4135
rect -500 4085 -450 4115
rect -500 4065 -485 4085
rect -465 4065 -450 4085
rect -500 4035 -450 4065
rect -500 4015 -485 4035
rect -465 4015 -450 4035
rect -500 3985 -450 4015
rect -500 3965 -485 3985
rect -465 3965 -450 3985
rect -500 3950 -450 3965
rect -350 4435 -300 4450
rect -350 4415 -335 4435
rect -315 4415 -300 4435
rect -350 4385 -300 4415
rect -350 4365 -335 4385
rect -315 4365 -300 4385
rect -350 4335 -300 4365
rect -350 4315 -335 4335
rect -315 4315 -300 4335
rect -350 4285 -300 4315
rect -350 4265 -335 4285
rect -315 4265 -300 4285
rect -350 4235 -300 4265
rect -350 4215 -335 4235
rect -315 4215 -300 4235
rect -350 4185 -300 4215
rect -350 4165 -335 4185
rect -315 4165 -300 4185
rect -350 4135 -300 4165
rect -350 4115 -335 4135
rect -315 4115 -300 4135
rect -350 4085 -300 4115
rect -350 4065 -335 4085
rect -315 4065 -300 4085
rect -350 4035 -300 4065
rect -350 4015 -335 4035
rect -315 4015 -300 4035
rect -350 3985 -300 4015
rect -350 3965 -335 3985
rect -315 3965 -300 3985
rect -350 3950 -300 3965
rect -200 4435 -150 4450
rect -200 4415 -185 4435
rect -165 4415 -150 4435
rect -200 4385 -150 4415
rect -200 4365 -185 4385
rect -165 4365 -150 4385
rect -200 4335 -150 4365
rect -200 4315 -185 4335
rect -165 4315 -150 4335
rect -200 4285 -150 4315
rect -200 4265 -185 4285
rect -165 4265 -150 4285
rect -200 4235 -150 4265
rect -200 4215 -185 4235
rect -165 4215 -150 4235
rect -200 4185 -150 4215
rect -200 4165 -185 4185
rect -165 4165 -150 4185
rect -200 4135 -150 4165
rect -200 4115 -185 4135
rect -165 4115 -150 4135
rect -200 4085 -150 4115
rect -200 4065 -185 4085
rect -165 4065 -150 4085
rect -200 4035 -150 4065
rect -200 4015 -185 4035
rect -165 4015 -150 4035
rect -200 3985 -150 4015
rect -200 3965 -185 3985
rect -165 3965 -150 3985
rect -200 3950 -150 3965
rect -50 4435 0 4450
rect -50 4415 -35 4435
rect -15 4415 0 4435
rect -50 4385 0 4415
rect -50 4365 -35 4385
rect -15 4365 0 4385
rect -50 4335 0 4365
rect -50 4315 -35 4335
rect -15 4315 0 4335
rect -50 4285 0 4315
rect -50 4265 -35 4285
rect -15 4265 0 4285
rect -50 4235 0 4265
rect -50 4215 -35 4235
rect -15 4215 0 4235
rect -50 4185 0 4215
rect -50 4165 -35 4185
rect -15 4165 0 4185
rect -50 4135 0 4165
rect -50 4115 -35 4135
rect -15 4115 0 4135
rect -50 4085 0 4115
rect -50 4065 -35 4085
rect -15 4065 0 4085
rect -50 4035 0 4065
rect -50 4015 -35 4035
rect -15 4015 0 4035
rect -50 3985 0 4015
rect -50 3965 -35 3985
rect -15 3965 0 3985
rect -50 3950 0 3965
rect 550 4435 600 4450
rect 550 4415 565 4435
rect 585 4415 600 4435
rect 550 4385 600 4415
rect 550 4365 565 4385
rect 585 4365 600 4385
rect 550 4335 600 4365
rect 550 4315 565 4335
rect 585 4315 600 4335
rect 550 4285 600 4315
rect 550 4265 565 4285
rect 585 4265 600 4285
rect 550 4235 600 4265
rect 550 4215 565 4235
rect 585 4215 600 4235
rect 550 4185 600 4215
rect 550 4165 565 4185
rect 585 4165 600 4185
rect 550 4135 600 4165
rect 550 4115 565 4135
rect 585 4115 600 4135
rect 550 4085 600 4115
rect 550 4065 565 4085
rect 585 4065 600 4085
rect 550 4035 600 4065
rect 550 4015 565 4035
rect 585 4015 600 4035
rect 550 3985 600 4015
rect 550 3965 565 3985
rect 585 3965 600 3985
rect 550 3950 600 3965
rect 700 4435 750 4450
rect 700 4415 715 4435
rect 735 4415 750 4435
rect 700 4385 750 4415
rect 700 4365 715 4385
rect 735 4365 750 4385
rect 700 4335 750 4365
rect 700 4315 715 4335
rect 735 4315 750 4335
rect 700 4285 750 4315
rect 700 4265 715 4285
rect 735 4265 750 4285
rect 700 4235 750 4265
rect 700 4215 715 4235
rect 735 4215 750 4235
rect 700 4185 750 4215
rect 700 4165 715 4185
rect 735 4165 750 4185
rect 700 4135 750 4165
rect 700 4115 715 4135
rect 735 4115 750 4135
rect 700 4085 750 4115
rect 700 4065 715 4085
rect 735 4065 750 4085
rect 700 4035 750 4065
rect 700 4015 715 4035
rect 735 4015 750 4035
rect 700 3985 750 4015
rect 700 3965 715 3985
rect 735 3965 750 3985
rect 700 3950 750 3965
rect 850 4435 900 4450
rect 850 4415 865 4435
rect 885 4415 900 4435
rect 850 4385 900 4415
rect 850 4365 865 4385
rect 885 4365 900 4385
rect 850 4335 900 4365
rect 850 4315 865 4335
rect 885 4315 900 4335
rect 850 4285 900 4315
rect 850 4265 865 4285
rect 885 4265 900 4285
rect 850 4235 900 4265
rect 850 4215 865 4235
rect 885 4215 900 4235
rect 850 4185 900 4215
rect 850 4165 865 4185
rect 885 4165 900 4185
rect 850 4135 900 4165
rect 850 4115 865 4135
rect 885 4115 900 4135
rect 850 4085 900 4115
rect 850 4065 865 4085
rect 885 4065 900 4085
rect 850 4035 900 4065
rect 850 4015 865 4035
rect 885 4015 900 4035
rect 850 3985 900 4015
rect 850 3965 865 3985
rect 885 3965 900 3985
rect 850 3950 900 3965
rect 1000 4435 1050 4450
rect 1000 4415 1015 4435
rect 1035 4415 1050 4435
rect 1000 4385 1050 4415
rect 1000 4365 1015 4385
rect 1035 4365 1050 4385
rect 1000 4335 1050 4365
rect 1000 4315 1015 4335
rect 1035 4315 1050 4335
rect 1000 4285 1050 4315
rect 1000 4265 1015 4285
rect 1035 4265 1050 4285
rect 1000 4235 1050 4265
rect 1000 4215 1015 4235
rect 1035 4215 1050 4235
rect 1000 4185 1050 4215
rect 1000 4165 1015 4185
rect 1035 4165 1050 4185
rect 1000 4135 1050 4165
rect 1000 4115 1015 4135
rect 1035 4115 1050 4135
rect 1000 4085 1050 4115
rect 1000 4065 1015 4085
rect 1035 4065 1050 4085
rect 1000 4035 1050 4065
rect 1000 4015 1015 4035
rect 1035 4015 1050 4035
rect 1000 3985 1050 4015
rect 1000 3965 1015 3985
rect 1035 3965 1050 3985
rect 1000 3950 1050 3965
rect 1150 4435 1200 4450
rect 1150 4415 1165 4435
rect 1185 4415 1200 4435
rect 1150 4385 1200 4415
rect 1150 4365 1165 4385
rect 1185 4365 1200 4385
rect 1150 4335 1200 4365
rect 1150 4315 1165 4335
rect 1185 4315 1200 4335
rect 1150 4285 1200 4315
rect 1150 4265 1165 4285
rect 1185 4265 1200 4285
rect 1150 4235 1200 4265
rect 1150 4215 1165 4235
rect 1185 4215 1200 4235
rect 1150 4185 1200 4215
rect 1150 4165 1165 4185
rect 1185 4165 1200 4185
rect 1150 4135 1200 4165
rect 1150 4115 1165 4135
rect 1185 4115 1200 4135
rect 1150 4085 1200 4115
rect 1150 4065 1165 4085
rect 1185 4065 1200 4085
rect 1150 4035 1200 4065
rect 1150 4015 1165 4035
rect 1185 4015 1200 4035
rect 1150 3985 1200 4015
rect 1150 3965 1165 3985
rect 1185 3965 1200 3985
rect 1150 3950 1200 3965
rect 1300 4435 1350 4450
rect 1300 4415 1315 4435
rect 1335 4415 1350 4435
rect 1300 4385 1350 4415
rect 1300 4365 1315 4385
rect 1335 4365 1350 4385
rect 1300 4335 1350 4365
rect 1300 4315 1315 4335
rect 1335 4315 1350 4335
rect 1300 4285 1350 4315
rect 1300 4265 1315 4285
rect 1335 4265 1350 4285
rect 1300 4235 1350 4265
rect 1300 4215 1315 4235
rect 1335 4215 1350 4235
rect 1300 4185 1350 4215
rect 1300 4165 1315 4185
rect 1335 4165 1350 4185
rect 1300 4135 1350 4165
rect 1300 4115 1315 4135
rect 1335 4115 1350 4135
rect 1300 4085 1350 4115
rect 1300 4065 1315 4085
rect 1335 4065 1350 4085
rect 1300 4035 1350 4065
rect 1300 4015 1315 4035
rect 1335 4015 1350 4035
rect 1300 3985 1350 4015
rect 1300 3965 1315 3985
rect 1335 3965 1350 3985
rect 1300 3950 1350 3965
rect 1450 4435 1500 4450
rect 1450 4415 1465 4435
rect 1485 4415 1500 4435
rect 1450 4385 1500 4415
rect 1450 4365 1465 4385
rect 1485 4365 1500 4385
rect 1450 4335 1500 4365
rect 1450 4315 1465 4335
rect 1485 4315 1500 4335
rect 1450 4285 1500 4315
rect 1450 4265 1465 4285
rect 1485 4265 1500 4285
rect 1450 4235 1500 4265
rect 1450 4215 1465 4235
rect 1485 4215 1500 4235
rect 1450 4185 1500 4215
rect 1450 4165 1465 4185
rect 1485 4165 1500 4185
rect 1450 4135 1500 4165
rect 1450 4115 1465 4135
rect 1485 4115 1500 4135
rect 1450 4085 1500 4115
rect 1450 4065 1465 4085
rect 1485 4065 1500 4085
rect 1450 4035 1500 4065
rect 1450 4015 1465 4035
rect 1485 4015 1500 4035
rect 1450 3985 1500 4015
rect 1450 3965 1465 3985
rect 1485 3965 1500 3985
rect 1450 3950 1500 3965
rect 1600 4435 1650 4450
rect 1600 4415 1615 4435
rect 1635 4415 1650 4435
rect 1600 4385 1650 4415
rect 1600 4365 1615 4385
rect 1635 4365 1650 4385
rect 1600 4335 1650 4365
rect 1600 4315 1615 4335
rect 1635 4315 1650 4335
rect 1600 4285 1650 4315
rect 1600 4265 1615 4285
rect 1635 4265 1650 4285
rect 1600 4235 1650 4265
rect 1600 4215 1615 4235
rect 1635 4215 1650 4235
rect 1600 4185 1650 4215
rect 1600 4165 1615 4185
rect 1635 4165 1650 4185
rect 1600 4135 1650 4165
rect 1600 4115 1615 4135
rect 1635 4115 1650 4135
rect 1600 4085 1650 4115
rect 1600 4065 1615 4085
rect 1635 4065 1650 4085
rect 1600 4035 1650 4065
rect 1600 4015 1615 4035
rect 1635 4015 1650 4035
rect 1600 3985 1650 4015
rect 1600 3965 1615 3985
rect 1635 3965 1650 3985
rect 1600 3950 1650 3965
rect 1750 4435 1800 4450
rect 1750 4415 1765 4435
rect 1785 4415 1800 4435
rect 1750 4385 1800 4415
rect 1750 4365 1765 4385
rect 1785 4365 1800 4385
rect 1750 4335 1800 4365
rect 1750 4315 1765 4335
rect 1785 4315 1800 4335
rect 1750 4285 1800 4315
rect 1750 4265 1765 4285
rect 1785 4265 1800 4285
rect 1750 4235 1800 4265
rect 1750 4215 1765 4235
rect 1785 4215 1800 4235
rect 1750 4185 1800 4215
rect 1750 4165 1765 4185
rect 1785 4165 1800 4185
rect 1750 4135 1800 4165
rect 1750 4115 1765 4135
rect 1785 4115 1800 4135
rect 1750 4085 1800 4115
rect 1750 4065 1765 4085
rect 1785 4065 1800 4085
rect 1750 4035 1800 4065
rect 1750 4015 1765 4035
rect 1785 4015 1800 4035
rect 1750 3985 1800 4015
rect 1750 3965 1765 3985
rect 1785 3965 1800 3985
rect 1750 3950 1800 3965
rect 1900 4435 1950 4450
rect 1900 4415 1915 4435
rect 1935 4415 1950 4435
rect 1900 4385 1950 4415
rect 1900 4365 1915 4385
rect 1935 4365 1950 4385
rect 1900 4335 1950 4365
rect 1900 4315 1915 4335
rect 1935 4315 1950 4335
rect 1900 4285 1950 4315
rect 1900 4265 1915 4285
rect 1935 4265 1950 4285
rect 1900 4235 1950 4265
rect 1900 4215 1915 4235
rect 1935 4215 1950 4235
rect 1900 4185 1950 4215
rect 1900 4165 1915 4185
rect 1935 4165 1950 4185
rect 1900 4135 1950 4165
rect 1900 4115 1915 4135
rect 1935 4115 1950 4135
rect 1900 4085 1950 4115
rect 1900 4065 1915 4085
rect 1935 4065 1950 4085
rect 1900 4035 1950 4065
rect 1900 4015 1915 4035
rect 1935 4015 1950 4035
rect 1900 3985 1950 4015
rect 1900 3965 1915 3985
rect 1935 3965 1950 3985
rect 1900 3950 1950 3965
rect 2050 4435 2100 4450
rect 2050 4415 2065 4435
rect 2085 4415 2100 4435
rect 2050 4385 2100 4415
rect 2050 4365 2065 4385
rect 2085 4365 2100 4385
rect 2050 4335 2100 4365
rect 2050 4315 2065 4335
rect 2085 4315 2100 4335
rect 2050 4285 2100 4315
rect 2050 4265 2065 4285
rect 2085 4265 2100 4285
rect 2050 4235 2100 4265
rect 2050 4215 2065 4235
rect 2085 4215 2100 4235
rect 2050 4185 2100 4215
rect 2050 4165 2065 4185
rect 2085 4165 2100 4185
rect 2050 4135 2100 4165
rect 2050 4115 2065 4135
rect 2085 4115 2100 4135
rect 2050 4085 2100 4115
rect 2050 4065 2065 4085
rect 2085 4065 2100 4085
rect 2050 4035 2100 4065
rect 2050 4015 2065 4035
rect 2085 4015 2100 4035
rect 2050 3985 2100 4015
rect 2050 3965 2065 3985
rect 2085 3965 2100 3985
rect 2050 3950 2100 3965
rect 2200 4435 2250 4450
rect 2200 4415 2215 4435
rect 2235 4415 2250 4435
rect 2200 4385 2250 4415
rect 2200 4365 2215 4385
rect 2235 4365 2250 4385
rect 2200 4335 2250 4365
rect 2200 4315 2215 4335
rect 2235 4315 2250 4335
rect 2200 4285 2250 4315
rect 2200 4265 2215 4285
rect 2235 4265 2250 4285
rect 2200 4235 2250 4265
rect 2200 4215 2215 4235
rect 2235 4215 2250 4235
rect 2200 4185 2250 4215
rect 2200 4165 2215 4185
rect 2235 4165 2250 4185
rect 2200 4135 2250 4165
rect 2200 4115 2215 4135
rect 2235 4115 2250 4135
rect 2200 4085 2250 4115
rect 2200 4065 2215 4085
rect 2235 4065 2250 4085
rect 2200 4035 2250 4065
rect 2200 4015 2215 4035
rect 2235 4015 2250 4035
rect 2200 3985 2250 4015
rect 2200 3965 2215 3985
rect 2235 3965 2250 3985
rect 2200 3950 2250 3965
rect 2350 4435 2400 4450
rect 2350 4415 2365 4435
rect 2385 4415 2400 4435
rect 2350 4385 2400 4415
rect 2350 4365 2365 4385
rect 2385 4365 2400 4385
rect 2350 4335 2400 4365
rect 2350 4315 2365 4335
rect 2385 4315 2400 4335
rect 2350 4285 2400 4315
rect 2350 4265 2365 4285
rect 2385 4265 2400 4285
rect 2350 4235 2400 4265
rect 2350 4215 2365 4235
rect 2385 4215 2400 4235
rect 2350 4185 2400 4215
rect 2350 4165 2365 4185
rect 2385 4165 2400 4185
rect 2350 4135 2400 4165
rect 2350 4115 2365 4135
rect 2385 4115 2400 4135
rect 2350 4085 2400 4115
rect 2350 4065 2365 4085
rect 2385 4065 2400 4085
rect 2350 4035 2400 4065
rect 2350 4015 2365 4035
rect 2385 4015 2400 4035
rect 2350 3985 2400 4015
rect 2350 3965 2365 3985
rect 2385 3965 2400 3985
rect 2350 3950 2400 3965
rect 2500 4435 2550 4450
rect 2500 4415 2515 4435
rect 2535 4415 2550 4435
rect 2500 4385 2550 4415
rect 2500 4365 2515 4385
rect 2535 4365 2550 4385
rect 2500 4335 2550 4365
rect 2500 4315 2515 4335
rect 2535 4315 2550 4335
rect 2500 4285 2550 4315
rect 2500 4265 2515 4285
rect 2535 4265 2550 4285
rect 2500 4235 2550 4265
rect 2500 4215 2515 4235
rect 2535 4215 2550 4235
rect 2500 4185 2550 4215
rect 2500 4165 2515 4185
rect 2535 4165 2550 4185
rect 2500 4135 2550 4165
rect 2500 4115 2515 4135
rect 2535 4115 2550 4135
rect 2500 4085 2550 4115
rect 2500 4065 2515 4085
rect 2535 4065 2550 4085
rect 2500 4035 2550 4065
rect 2500 4015 2515 4035
rect 2535 4015 2550 4035
rect 2500 3985 2550 4015
rect 2500 3965 2515 3985
rect 2535 3965 2550 3985
rect 2500 3950 2550 3965
rect 2650 4435 2700 4450
rect 2650 4415 2665 4435
rect 2685 4415 2700 4435
rect 2650 4385 2700 4415
rect 2650 4365 2665 4385
rect 2685 4365 2700 4385
rect 2650 4335 2700 4365
rect 2650 4315 2665 4335
rect 2685 4315 2700 4335
rect 2650 4285 2700 4315
rect 2650 4265 2665 4285
rect 2685 4265 2700 4285
rect 2650 4235 2700 4265
rect 2650 4215 2665 4235
rect 2685 4215 2700 4235
rect 2650 4185 2700 4215
rect 2650 4165 2665 4185
rect 2685 4165 2700 4185
rect 2650 4135 2700 4165
rect 2650 4115 2665 4135
rect 2685 4115 2700 4135
rect 2650 4085 2700 4115
rect 2650 4065 2665 4085
rect 2685 4065 2700 4085
rect 2650 4035 2700 4065
rect 2650 4015 2665 4035
rect 2685 4015 2700 4035
rect 2650 3985 2700 4015
rect 2650 3965 2665 3985
rect 2685 3965 2700 3985
rect 2650 3950 2700 3965
rect 2800 4435 2850 4450
rect 2800 4415 2815 4435
rect 2835 4415 2850 4435
rect 2800 4385 2850 4415
rect 2800 4365 2815 4385
rect 2835 4365 2850 4385
rect 2800 4335 2850 4365
rect 2800 4315 2815 4335
rect 2835 4315 2850 4335
rect 2800 4285 2850 4315
rect 2800 4265 2815 4285
rect 2835 4265 2850 4285
rect 2800 4235 2850 4265
rect 2800 4215 2815 4235
rect 2835 4215 2850 4235
rect 2800 4185 2850 4215
rect 2800 4165 2815 4185
rect 2835 4165 2850 4185
rect 2800 4135 2850 4165
rect 2800 4115 2815 4135
rect 2835 4115 2850 4135
rect 2800 4085 2850 4115
rect 2800 4065 2815 4085
rect 2835 4065 2850 4085
rect 2800 4035 2850 4065
rect 2800 4015 2815 4035
rect 2835 4015 2850 4035
rect 2800 3985 2850 4015
rect 2800 3965 2815 3985
rect 2835 3965 2850 3985
rect 2800 3950 2850 3965
rect 2950 4435 3000 4450
rect 2950 4415 2965 4435
rect 2985 4415 3000 4435
rect 2950 4385 3000 4415
rect 2950 4365 2965 4385
rect 2985 4365 3000 4385
rect 2950 4335 3000 4365
rect 2950 4315 2965 4335
rect 2985 4315 3000 4335
rect 2950 4285 3000 4315
rect 2950 4265 2965 4285
rect 2985 4265 3000 4285
rect 2950 4235 3000 4265
rect 2950 4215 2965 4235
rect 2985 4215 3000 4235
rect 2950 4185 3000 4215
rect 2950 4165 2965 4185
rect 2985 4165 3000 4185
rect 2950 4135 3000 4165
rect 2950 4115 2965 4135
rect 2985 4115 3000 4135
rect 2950 4085 3000 4115
rect 2950 4065 2965 4085
rect 2985 4065 3000 4085
rect 2950 4035 3000 4065
rect 2950 4015 2965 4035
rect 2985 4015 3000 4035
rect 2950 3985 3000 4015
rect 2950 3965 2965 3985
rect 2985 3965 3000 3985
rect 2950 3950 3000 3965
rect 3100 4435 3150 4450
rect 3100 4415 3115 4435
rect 3135 4415 3150 4435
rect 3100 4385 3150 4415
rect 3100 4365 3115 4385
rect 3135 4365 3150 4385
rect 3100 4335 3150 4365
rect 3100 4315 3115 4335
rect 3135 4315 3150 4335
rect 3100 4285 3150 4315
rect 3100 4265 3115 4285
rect 3135 4265 3150 4285
rect 3100 4235 3150 4265
rect 3100 4215 3115 4235
rect 3135 4215 3150 4235
rect 3100 4185 3150 4215
rect 3100 4165 3115 4185
rect 3135 4165 3150 4185
rect 3100 4135 3150 4165
rect 3100 4115 3115 4135
rect 3135 4115 3150 4135
rect 3100 4085 3150 4115
rect 3100 4065 3115 4085
rect 3135 4065 3150 4085
rect 3100 4035 3150 4065
rect 3100 4015 3115 4035
rect 3135 4015 3150 4035
rect 3100 3985 3150 4015
rect 3100 3965 3115 3985
rect 3135 3965 3150 3985
rect 3100 3950 3150 3965
rect 3250 4435 3300 4450
rect 3250 4415 3265 4435
rect 3285 4415 3300 4435
rect 3250 4385 3300 4415
rect 3250 4365 3265 4385
rect 3285 4365 3300 4385
rect 3250 4335 3300 4365
rect 3250 4315 3265 4335
rect 3285 4315 3300 4335
rect 3250 4285 3300 4315
rect 3250 4265 3265 4285
rect 3285 4265 3300 4285
rect 3250 4235 3300 4265
rect 3250 4215 3265 4235
rect 3285 4215 3300 4235
rect 3250 4185 3300 4215
rect 3250 4165 3265 4185
rect 3285 4165 3300 4185
rect 3250 4135 3300 4165
rect 3250 4115 3265 4135
rect 3285 4115 3300 4135
rect 3250 4085 3300 4115
rect 3250 4065 3265 4085
rect 3285 4065 3300 4085
rect 3250 4035 3300 4065
rect 3250 4015 3265 4035
rect 3285 4015 3300 4035
rect 3250 3985 3300 4015
rect 3250 3965 3265 3985
rect 3285 3965 3300 3985
rect 3250 3950 3300 3965
rect 3400 4435 3450 4450
rect 3400 4415 3415 4435
rect 3435 4415 3450 4435
rect 3400 4385 3450 4415
rect 3400 4365 3415 4385
rect 3435 4365 3450 4385
rect 3400 4335 3450 4365
rect 3400 4315 3415 4335
rect 3435 4315 3450 4335
rect 3400 4285 3450 4315
rect 3400 4265 3415 4285
rect 3435 4265 3450 4285
rect 3400 4235 3450 4265
rect 3400 4215 3415 4235
rect 3435 4215 3450 4235
rect 3400 4185 3450 4215
rect 3400 4165 3415 4185
rect 3435 4165 3450 4185
rect 3400 4135 3450 4165
rect 3400 4115 3415 4135
rect 3435 4115 3450 4135
rect 3400 4085 3450 4115
rect 3400 4065 3415 4085
rect 3435 4065 3450 4085
rect 3400 4035 3450 4065
rect 3400 4015 3415 4035
rect 3435 4015 3450 4035
rect 3400 3985 3450 4015
rect 3400 3965 3415 3985
rect 3435 3965 3450 3985
rect 3400 3950 3450 3965
rect 3550 4435 3600 4450
rect 3550 4415 3565 4435
rect 3585 4415 3600 4435
rect 3550 4385 3600 4415
rect 3550 4365 3565 4385
rect 3585 4365 3600 4385
rect 3550 4335 3600 4365
rect 3550 4315 3565 4335
rect 3585 4315 3600 4335
rect 3550 4285 3600 4315
rect 3550 4265 3565 4285
rect 3585 4265 3600 4285
rect 3550 4235 3600 4265
rect 3550 4215 3565 4235
rect 3585 4215 3600 4235
rect 3550 4185 3600 4215
rect 3550 4165 3565 4185
rect 3585 4165 3600 4185
rect 3550 4135 3600 4165
rect 3550 4115 3565 4135
rect 3585 4115 3600 4135
rect 3550 4085 3600 4115
rect 3550 4065 3565 4085
rect 3585 4065 3600 4085
rect 3550 4035 3600 4065
rect 3550 4015 3565 4035
rect 3585 4015 3600 4035
rect 3550 3985 3600 4015
rect 3550 3965 3565 3985
rect 3585 3965 3600 3985
rect 3550 3950 3600 3965
rect 4150 4435 4200 4450
rect 4150 4415 4165 4435
rect 4185 4415 4200 4435
rect 4150 4385 4200 4415
rect 4150 4365 4165 4385
rect 4185 4365 4200 4385
rect 4150 4335 4200 4365
rect 4150 4315 4165 4335
rect 4185 4315 4200 4335
rect 4150 4285 4200 4315
rect 4150 4265 4165 4285
rect 4185 4265 4200 4285
rect 4150 4235 4200 4265
rect 4150 4215 4165 4235
rect 4185 4215 4200 4235
rect 4150 4185 4200 4215
rect 4150 4165 4165 4185
rect 4185 4165 4200 4185
rect 4150 4135 4200 4165
rect 4150 4115 4165 4135
rect 4185 4115 4200 4135
rect 4150 4085 4200 4115
rect 4150 4065 4165 4085
rect 4185 4065 4200 4085
rect 4150 4035 4200 4065
rect 4150 4015 4165 4035
rect 4185 4015 4200 4035
rect 4150 3985 4200 4015
rect 4150 3965 4165 3985
rect 4185 3965 4200 3985
rect 4150 3950 4200 3965
rect 4750 4435 4800 4450
rect 4750 4415 4765 4435
rect 4785 4415 4800 4435
rect 4750 4385 4800 4415
rect 4750 4365 4765 4385
rect 4785 4365 4800 4385
rect 4750 4335 4800 4365
rect 4750 4315 4765 4335
rect 4785 4315 4800 4335
rect 4750 4285 4800 4315
rect 4750 4265 4765 4285
rect 4785 4265 4800 4285
rect 4750 4235 4800 4265
rect 4750 4215 4765 4235
rect 4785 4215 4800 4235
rect 4750 4185 4800 4215
rect 4750 4165 4765 4185
rect 4785 4165 4800 4185
rect 4750 4135 4800 4165
rect 4750 4115 4765 4135
rect 4785 4115 4800 4135
rect 4750 4085 4800 4115
rect 4750 4065 4765 4085
rect 4785 4065 4800 4085
rect 4750 4035 4800 4065
rect 4750 4015 4765 4035
rect 4785 4015 4800 4035
rect 4750 3985 4800 4015
rect 4750 3965 4765 3985
rect 4785 3965 4800 3985
rect 4750 3950 4800 3965
rect 4900 4435 4950 4450
rect 4900 4415 4915 4435
rect 4935 4415 4950 4435
rect 4900 4385 4950 4415
rect 4900 4365 4915 4385
rect 4935 4365 4950 4385
rect 4900 4335 4950 4365
rect 4900 4315 4915 4335
rect 4935 4315 4950 4335
rect 4900 4285 4950 4315
rect 4900 4265 4915 4285
rect 4935 4265 4950 4285
rect 4900 4235 4950 4265
rect 4900 4215 4915 4235
rect 4935 4215 4950 4235
rect 4900 4185 4950 4215
rect 4900 4165 4915 4185
rect 4935 4165 4950 4185
rect 4900 4135 4950 4165
rect 4900 4115 4915 4135
rect 4935 4115 4950 4135
rect 4900 4085 4950 4115
rect 4900 4065 4915 4085
rect 4935 4065 4950 4085
rect 4900 4035 4950 4065
rect 4900 4015 4915 4035
rect 4935 4015 4950 4035
rect 4900 3985 4950 4015
rect 4900 3965 4915 3985
rect 4935 3965 4950 3985
rect 4900 3950 4950 3965
rect 5050 4435 5100 4450
rect 5050 4415 5065 4435
rect 5085 4415 5100 4435
rect 5050 4385 5100 4415
rect 5050 4365 5065 4385
rect 5085 4365 5100 4385
rect 5050 4335 5100 4365
rect 5050 4315 5065 4335
rect 5085 4315 5100 4335
rect 5050 4285 5100 4315
rect 5050 4265 5065 4285
rect 5085 4265 5100 4285
rect 5050 4235 5100 4265
rect 5050 4215 5065 4235
rect 5085 4215 5100 4235
rect 5050 4185 5100 4215
rect 5050 4165 5065 4185
rect 5085 4165 5100 4185
rect 5050 4135 5100 4165
rect 5050 4115 5065 4135
rect 5085 4115 5100 4135
rect 5050 4085 5100 4115
rect 5050 4065 5065 4085
rect 5085 4065 5100 4085
rect 5050 4035 5100 4065
rect 5050 4015 5065 4035
rect 5085 4015 5100 4035
rect 5050 3985 5100 4015
rect 5050 3965 5065 3985
rect 5085 3965 5100 3985
rect 5050 3950 5100 3965
rect 5200 4435 5250 4450
rect 5200 4415 5215 4435
rect 5235 4415 5250 4435
rect 5200 4385 5250 4415
rect 5200 4365 5215 4385
rect 5235 4365 5250 4385
rect 5200 4335 5250 4365
rect 5200 4315 5215 4335
rect 5235 4315 5250 4335
rect 5200 4285 5250 4315
rect 5200 4265 5215 4285
rect 5235 4265 5250 4285
rect 5200 4235 5250 4265
rect 5200 4215 5215 4235
rect 5235 4215 5250 4235
rect 5200 4185 5250 4215
rect 5200 4165 5215 4185
rect 5235 4165 5250 4185
rect 5200 4135 5250 4165
rect 5200 4115 5215 4135
rect 5235 4115 5250 4135
rect 5200 4085 5250 4115
rect 5200 4065 5215 4085
rect 5235 4065 5250 4085
rect 5200 4035 5250 4065
rect 5200 4015 5215 4035
rect 5235 4015 5250 4035
rect 5200 3985 5250 4015
rect 5200 3965 5215 3985
rect 5235 3965 5250 3985
rect 5200 3950 5250 3965
rect 5350 4435 5400 4450
rect 5350 4415 5365 4435
rect 5385 4415 5400 4435
rect 5350 4385 5400 4415
rect 5350 4365 5365 4385
rect 5385 4365 5400 4385
rect 5350 4335 5400 4365
rect 5350 4315 5365 4335
rect 5385 4315 5400 4335
rect 5350 4285 5400 4315
rect 5350 4265 5365 4285
rect 5385 4265 5400 4285
rect 5350 4235 5400 4265
rect 5350 4215 5365 4235
rect 5385 4215 5400 4235
rect 5350 4185 5400 4215
rect 5350 4165 5365 4185
rect 5385 4165 5400 4185
rect 5350 4135 5400 4165
rect 5350 4115 5365 4135
rect 5385 4115 5400 4135
rect 5350 4085 5400 4115
rect 5350 4065 5365 4085
rect 5385 4065 5400 4085
rect 5350 4035 5400 4065
rect 5350 4015 5365 4035
rect 5385 4015 5400 4035
rect 5350 3985 5400 4015
rect 5350 3965 5365 3985
rect 5385 3965 5400 3985
rect 5350 3950 5400 3965
rect 5500 4435 5550 4450
rect 5500 4415 5515 4435
rect 5535 4415 5550 4435
rect 5500 4385 5550 4415
rect 5500 4365 5515 4385
rect 5535 4365 5550 4385
rect 5500 4335 5550 4365
rect 5500 4315 5515 4335
rect 5535 4315 5550 4335
rect 5500 4285 5550 4315
rect 5500 4265 5515 4285
rect 5535 4265 5550 4285
rect 5500 4235 5550 4265
rect 5500 4215 5515 4235
rect 5535 4215 5550 4235
rect 5500 4185 5550 4215
rect 5500 4165 5515 4185
rect 5535 4165 5550 4185
rect 5500 4135 5550 4165
rect 5500 4115 5515 4135
rect 5535 4115 5550 4135
rect 5500 4085 5550 4115
rect 5500 4065 5515 4085
rect 5535 4065 5550 4085
rect 5500 4035 5550 4065
rect 5500 4015 5515 4035
rect 5535 4015 5550 4035
rect 5500 3985 5550 4015
rect 5500 3965 5515 3985
rect 5535 3965 5550 3985
rect 5500 3950 5550 3965
rect 5650 4435 5700 4450
rect 5650 4415 5665 4435
rect 5685 4415 5700 4435
rect 5650 4385 5700 4415
rect 5650 4365 5665 4385
rect 5685 4365 5700 4385
rect 5650 4335 5700 4365
rect 5650 4315 5665 4335
rect 5685 4315 5700 4335
rect 5650 4285 5700 4315
rect 5650 4265 5665 4285
rect 5685 4265 5700 4285
rect 5650 4235 5700 4265
rect 5650 4215 5665 4235
rect 5685 4215 5700 4235
rect 5650 4185 5700 4215
rect 5650 4165 5665 4185
rect 5685 4165 5700 4185
rect 5650 4135 5700 4165
rect 5650 4115 5665 4135
rect 5685 4115 5700 4135
rect 5650 4085 5700 4115
rect 5650 4065 5665 4085
rect 5685 4065 5700 4085
rect 5650 4035 5700 4065
rect 5650 4015 5665 4035
rect 5685 4015 5700 4035
rect 5650 3985 5700 4015
rect 5650 3965 5665 3985
rect 5685 3965 5700 3985
rect 5650 3950 5700 3965
rect 5800 4435 5850 4450
rect 5800 4415 5815 4435
rect 5835 4415 5850 4435
rect 5800 4385 5850 4415
rect 5800 4365 5815 4385
rect 5835 4365 5850 4385
rect 5800 4335 5850 4365
rect 5800 4315 5815 4335
rect 5835 4315 5850 4335
rect 5800 4285 5850 4315
rect 5800 4265 5815 4285
rect 5835 4265 5850 4285
rect 5800 4235 5850 4265
rect 5800 4215 5815 4235
rect 5835 4215 5850 4235
rect 5800 4185 5850 4215
rect 5800 4165 5815 4185
rect 5835 4165 5850 4185
rect 5800 4135 5850 4165
rect 5800 4115 5815 4135
rect 5835 4115 5850 4135
rect 5800 4085 5850 4115
rect 5800 4065 5815 4085
rect 5835 4065 5850 4085
rect 5800 4035 5850 4065
rect 5800 4015 5815 4035
rect 5835 4015 5850 4035
rect 5800 3985 5850 4015
rect 5800 3965 5815 3985
rect 5835 3965 5850 3985
rect 5800 3950 5850 3965
rect 5950 4435 6000 4450
rect 5950 4415 5965 4435
rect 5985 4415 6000 4435
rect 5950 4385 6000 4415
rect 5950 4365 5965 4385
rect 5985 4365 6000 4385
rect 5950 4335 6000 4365
rect 5950 4315 5965 4335
rect 5985 4315 6000 4335
rect 5950 4285 6000 4315
rect 5950 4265 5965 4285
rect 5985 4265 6000 4285
rect 5950 4235 6000 4265
rect 5950 4215 5965 4235
rect 5985 4215 6000 4235
rect 5950 4185 6000 4215
rect 5950 4165 5965 4185
rect 5985 4165 6000 4185
rect 5950 4135 6000 4165
rect 5950 4115 5965 4135
rect 5985 4115 6000 4135
rect 5950 4085 6000 4115
rect 5950 4065 5965 4085
rect 5985 4065 6000 4085
rect 5950 4035 6000 4065
rect 5950 4015 5965 4035
rect 5985 4015 6000 4035
rect 5950 3985 6000 4015
rect 5950 3965 5965 3985
rect 5985 3965 6000 3985
rect 5950 3950 6000 3965
rect 6100 4435 6150 4450
rect 6100 4415 6115 4435
rect 6135 4415 6150 4435
rect 6100 4385 6150 4415
rect 6100 4365 6115 4385
rect 6135 4365 6150 4385
rect 6100 4335 6150 4365
rect 6100 4315 6115 4335
rect 6135 4315 6150 4335
rect 6100 4285 6150 4315
rect 6100 4265 6115 4285
rect 6135 4265 6150 4285
rect 6100 4235 6150 4265
rect 6100 4215 6115 4235
rect 6135 4215 6150 4235
rect 6100 4185 6150 4215
rect 6100 4165 6115 4185
rect 6135 4165 6150 4185
rect 6100 4135 6150 4165
rect 6100 4115 6115 4135
rect 6135 4115 6150 4135
rect 6100 4085 6150 4115
rect 6100 4065 6115 4085
rect 6135 4065 6150 4085
rect 6100 4035 6150 4065
rect 6100 4015 6115 4035
rect 6135 4015 6150 4035
rect 6100 3985 6150 4015
rect 6100 3965 6115 3985
rect 6135 3965 6150 3985
rect 6100 3950 6150 3965
rect 6250 4435 6300 4450
rect 6250 4415 6265 4435
rect 6285 4415 6300 4435
rect 6250 4385 6300 4415
rect 6250 4365 6265 4385
rect 6285 4365 6300 4385
rect 6250 4335 6300 4365
rect 6250 4315 6265 4335
rect 6285 4315 6300 4335
rect 6250 4285 6300 4315
rect 6250 4265 6265 4285
rect 6285 4265 6300 4285
rect 6250 4235 6300 4265
rect 6250 4215 6265 4235
rect 6285 4215 6300 4235
rect 6250 4185 6300 4215
rect 6250 4165 6265 4185
rect 6285 4165 6300 4185
rect 6250 4135 6300 4165
rect 6250 4115 6265 4135
rect 6285 4115 6300 4135
rect 6250 4085 6300 4115
rect 6250 4065 6265 4085
rect 6285 4065 6300 4085
rect 6250 4035 6300 4065
rect 6250 4015 6265 4035
rect 6285 4015 6300 4035
rect 6250 3985 6300 4015
rect 6250 3965 6265 3985
rect 6285 3965 6300 3985
rect 6250 3950 6300 3965
rect 6400 4435 6450 4450
rect 6400 4415 6415 4435
rect 6435 4415 6450 4435
rect 6400 4385 6450 4415
rect 6400 4365 6415 4385
rect 6435 4365 6450 4385
rect 6400 4335 6450 4365
rect 6400 4315 6415 4335
rect 6435 4315 6450 4335
rect 6400 4285 6450 4315
rect 6400 4265 6415 4285
rect 6435 4265 6450 4285
rect 6400 4235 6450 4265
rect 6400 4215 6415 4235
rect 6435 4215 6450 4235
rect 6400 4185 6450 4215
rect 6400 4165 6415 4185
rect 6435 4165 6450 4185
rect 6400 4135 6450 4165
rect 6400 4115 6415 4135
rect 6435 4115 6450 4135
rect 6400 4085 6450 4115
rect 6400 4065 6415 4085
rect 6435 4065 6450 4085
rect 6400 4035 6450 4065
rect 6400 4015 6415 4035
rect 6435 4015 6450 4035
rect 6400 3985 6450 4015
rect 6400 3965 6415 3985
rect 6435 3965 6450 3985
rect 6400 3950 6450 3965
rect 6550 4435 6600 4450
rect 6550 4415 6565 4435
rect 6585 4415 6600 4435
rect 6550 4385 6600 4415
rect 6550 4365 6565 4385
rect 6585 4365 6600 4385
rect 6550 4335 6600 4365
rect 6550 4315 6565 4335
rect 6585 4315 6600 4335
rect 6550 4285 6600 4315
rect 6550 4265 6565 4285
rect 6585 4265 6600 4285
rect 6550 4235 6600 4265
rect 6550 4215 6565 4235
rect 6585 4215 6600 4235
rect 6550 4185 6600 4215
rect 6550 4165 6565 4185
rect 6585 4165 6600 4185
rect 6550 4135 6600 4165
rect 6550 4115 6565 4135
rect 6585 4115 6600 4135
rect 6550 4085 6600 4115
rect 6550 4065 6565 4085
rect 6585 4065 6600 4085
rect 6550 4035 6600 4065
rect 6550 4015 6565 4035
rect 6585 4015 6600 4035
rect 6550 3985 6600 4015
rect 6550 3965 6565 3985
rect 6585 3965 6600 3985
rect 6550 3950 6600 3965
rect 6700 4435 6750 4450
rect 6700 4415 6715 4435
rect 6735 4415 6750 4435
rect 6700 4385 6750 4415
rect 6700 4365 6715 4385
rect 6735 4365 6750 4385
rect 6700 4335 6750 4365
rect 6700 4315 6715 4335
rect 6735 4315 6750 4335
rect 6700 4285 6750 4315
rect 6700 4265 6715 4285
rect 6735 4265 6750 4285
rect 6700 4235 6750 4265
rect 6700 4215 6715 4235
rect 6735 4215 6750 4235
rect 6700 4185 6750 4215
rect 6700 4165 6715 4185
rect 6735 4165 6750 4185
rect 6700 4135 6750 4165
rect 6700 4115 6715 4135
rect 6735 4115 6750 4135
rect 6700 4085 6750 4115
rect 6700 4065 6715 4085
rect 6735 4065 6750 4085
rect 6700 4035 6750 4065
rect 6700 4015 6715 4035
rect 6735 4015 6750 4035
rect 6700 3985 6750 4015
rect 6700 3965 6715 3985
rect 6735 3965 6750 3985
rect 6700 3950 6750 3965
rect 6850 4435 6900 4450
rect 6850 4415 6865 4435
rect 6885 4415 6900 4435
rect 6850 4385 6900 4415
rect 6850 4365 6865 4385
rect 6885 4365 6900 4385
rect 6850 4335 6900 4365
rect 6850 4315 6865 4335
rect 6885 4315 6900 4335
rect 6850 4285 6900 4315
rect 6850 4265 6865 4285
rect 6885 4265 6900 4285
rect 6850 4235 6900 4265
rect 6850 4215 6865 4235
rect 6885 4215 6900 4235
rect 6850 4185 6900 4215
rect 6850 4165 6865 4185
rect 6885 4165 6900 4185
rect 6850 4135 6900 4165
rect 6850 4115 6865 4135
rect 6885 4115 6900 4135
rect 6850 4085 6900 4115
rect 6850 4065 6865 4085
rect 6885 4065 6900 4085
rect 6850 4035 6900 4065
rect 6850 4015 6865 4035
rect 6885 4015 6900 4035
rect 6850 3985 6900 4015
rect 6850 3965 6865 3985
rect 6885 3965 6900 3985
rect 6850 3950 6900 3965
rect 7000 4435 7050 4450
rect 7000 4415 7015 4435
rect 7035 4415 7050 4435
rect 7000 4385 7050 4415
rect 7000 4365 7015 4385
rect 7035 4365 7050 4385
rect 7000 4335 7050 4365
rect 7000 4315 7015 4335
rect 7035 4315 7050 4335
rect 7000 4285 7050 4315
rect 7000 4265 7015 4285
rect 7035 4265 7050 4285
rect 7000 4235 7050 4265
rect 7000 4215 7015 4235
rect 7035 4215 7050 4235
rect 7000 4185 7050 4215
rect 7000 4165 7015 4185
rect 7035 4165 7050 4185
rect 7000 4135 7050 4165
rect 7000 4115 7015 4135
rect 7035 4115 7050 4135
rect 7000 4085 7050 4115
rect 7000 4065 7015 4085
rect 7035 4065 7050 4085
rect 7000 4035 7050 4065
rect 7000 4015 7015 4035
rect 7035 4015 7050 4035
rect 7000 3985 7050 4015
rect 7000 3965 7015 3985
rect 7035 3965 7050 3985
rect 7000 3950 7050 3965
rect 7150 4435 7200 4450
rect 7150 4415 7165 4435
rect 7185 4415 7200 4435
rect 7150 4385 7200 4415
rect 7150 4365 7165 4385
rect 7185 4365 7200 4385
rect 7150 4335 7200 4365
rect 7150 4315 7165 4335
rect 7185 4315 7200 4335
rect 7150 4285 7200 4315
rect 7150 4265 7165 4285
rect 7185 4265 7200 4285
rect 7150 4235 7200 4265
rect 7150 4215 7165 4235
rect 7185 4215 7200 4235
rect 7150 4185 7200 4215
rect 7150 4165 7165 4185
rect 7185 4165 7200 4185
rect 7150 4135 7200 4165
rect 7150 4115 7165 4135
rect 7185 4115 7200 4135
rect 7150 4085 7200 4115
rect 7150 4065 7165 4085
rect 7185 4065 7200 4085
rect 7150 4035 7200 4065
rect 7150 4015 7165 4035
rect 7185 4015 7200 4035
rect 7150 3985 7200 4015
rect 7150 3965 7165 3985
rect 7185 3965 7200 3985
rect 7150 3950 7200 3965
rect 7300 4435 7350 4450
rect 7300 4415 7315 4435
rect 7335 4415 7350 4435
rect 7300 4385 7350 4415
rect 7300 4365 7315 4385
rect 7335 4365 7350 4385
rect 7300 4335 7350 4365
rect 7300 4315 7315 4335
rect 7335 4315 7350 4335
rect 7300 4285 7350 4315
rect 7300 4265 7315 4285
rect 7335 4265 7350 4285
rect 7300 4235 7350 4265
rect 7300 4215 7315 4235
rect 7335 4215 7350 4235
rect 7300 4185 7350 4215
rect 7300 4165 7315 4185
rect 7335 4165 7350 4185
rect 7300 4135 7350 4165
rect 7300 4115 7315 4135
rect 7335 4115 7350 4135
rect 7300 4085 7350 4115
rect 7300 4065 7315 4085
rect 7335 4065 7350 4085
rect 7300 4035 7350 4065
rect 7300 4015 7315 4035
rect 7335 4015 7350 4035
rect 7300 3985 7350 4015
rect 7300 3965 7315 3985
rect 7335 3965 7350 3985
rect 7300 3950 7350 3965
rect 7450 4435 7500 4450
rect 7450 4415 7465 4435
rect 7485 4415 7500 4435
rect 7450 4385 7500 4415
rect 7450 4365 7465 4385
rect 7485 4365 7500 4385
rect 7450 4335 7500 4365
rect 7450 4315 7465 4335
rect 7485 4315 7500 4335
rect 7450 4285 7500 4315
rect 7450 4265 7465 4285
rect 7485 4265 7500 4285
rect 7450 4235 7500 4265
rect 7450 4215 7465 4235
rect 7485 4215 7500 4235
rect 7450 4185 7500 4215
rect 7450 4165 7465 4185
rect 7485 4165 7500 4185
rect 7450 4135 7500 4165
rect 7450 4115 7465 4135
rect 7485 4115 7500 4135
rect 7450 4085 7500 4115
rect 7450 4065 7465 4085
rect 7485 4065 7500 4085
rect 7450 4035 7500 4065
rect 7450 4015 7465 4035
rect 7485 4015 7500 4035
rect 7450 3985 7500 4015
rect 7450 3965 7465 3985
rect 7485 3965 7500 3985
rect 7450 3950 7500 3965
rect 7600 4435 7650 4450
rect 7600 4415 7615 4435
rect 7635 4415 7650 4435
rect 7600 4385 7650 4415
rect 7600 4365 7615 4385
rect 7635 4365 7650 4385
rect 7600 4335 7650 4365
rect 7600 4315 7615 4335
rect 7635 4315 7650 4335
rect 7600 4285 7650 4315
rect 7600 4265 7615 4285
rect 7635 4265 7650 4285
rect 7600 4235 7650 4265
rect 7600 4215 7615 4235
rect 7635 4215 7650 4235
rect 7600 4185 7650 4215
rect 7600 4165 7615 4185
rect 7635 4165 7650 4185
rect 7600 4135 7650 4165
rect 7600 4115 7615 4135
rect 7635 4115 7650 4135
rect 7600 4085 7650 4115
rect 7600 4065 7615 4085
rect 7635 4065 7650 4085
rect 7600 4035 7650 4065
rect 7600 4015 7615 4035
rect 7635 4015 7650 4035
rect 7600 3985 7650 4015
rect 7600 3965 7615 3985
rect 7635 3965 7650 3985
rect 7600 3950 7650 3965
rect 7750 4435 7800 4450
rect 7750 4415 7765 4435
rect 7785 4415 7800 4435
rect 7750 4385 7800 4415
rect 7750 4365 7765 4385
rect 7785 4365 7800 4385
rect 7750 4335 7800 4365
rect 7750 4315 7765 4335
rect 7785 4315 7800 4335
rect 7750 4285 7800 4315
rect 7750 4265 7765 4285
rect 7785 4265 7800 4285
rect 7750 4235 7800 4265
rect 7750 4215 7765 4235
rect 7785 4215 7800 4235
rect 7750 4185 7800 4215
rect 7750 4165 7765 4185
rect 7785 4165 7800 4185
rect 7750 4135 7800 4165
rect 7750 4115 7765 4135
rect 7785 4115 7800 4135
rect 7750 4085 7800 4115
rect 7750 4065 7765 4085
rect 7785 4065 7800 4085
rect 7750 4035 7800 4065
rect 7750 4015 7765 4035
rect 7785 4015 7800 4035
rect 7750 3985 7800 4015
rect 7750 3965 7765 3985
rect 7785 3965 7800 3985
rect 7750 3950 7800 3965
rect 8350 4435 8400 4450
rect 8350 4415 8365 4435
rect 8385 4415 8400 4435
rect 8350 4385 8400 4415
rect 8350 4365 8365 4385
rect 8385 4365 8400 4385
rect 8350 4335 8400 4365
rect 8350 4315 8365 4335
rect 8385 4315 8400 4335
rect 8350 4285 8400 4315
rect 8350 4265 8365 4285
rect 8385 4265 8400 4285
rect 8350 4235 8400 4265
rect 8350 4215 8365 4235
rect 8385 4215 8400 4235
rect 8350 4185 8400 4215
rect 8350 4165 8365 4185
rect 8385 4165 8400 4185
rect 8350 4135 8400 4165
rect 8350 4115 8365 4135
rect 8385 4115 8400 4135
rect 8350 4085 8400 4115
rect 8350 4065 8365 4085
rect 8385 4065 8400 4085
rect 8350 4035 8400 4065
rect 8350 4015 8365 4035
rect 8385 4015 8400 4035
rect 8350 3985 8400 4015
rect 8350 3965 8365 3985
rect 8385 3965 8400 3985
rect 8350 3950 8400 3965
rect 8500 4435 8550 4500
rect 8500 4415 8515 4435
rect 8535 4415 8550 4435
rect 8500 4385 8550 4415
rect 8500 4365 8515 4385
rect 8535 4365 8550 4385
rect 8500 4335 8550 4365
rect 8500 4315 8515 4335
rect 8535 4315 8550 4335
rect 8500 4285 8550 4315
rect 8500 4265 8515 4285
rect 8535 4265 8550 4285
rect 8500 4235 8550 4265
rect 8500 4215 8515 4235
rect 8535 4215 8550 4235
rect 8500 4185 8550 4215
rect 8500 4165 8515 4185
rect 8535 4165 8550 4185
rect 8500 4135 8550 4165
rect 8500 4115 8515 4135
rect 8535 4115 8550 4135
rect 8500 4085 8550 4115
rect 8500 4065 8515 4085
rect 8535 4065 8550 4085
rect 8500 4035 8550 4065
rect 8500 4015 8515 4035
rect 8535 4015 8550 4035
rect 8500 3985 8550 4015
rect 8500 3965 8515 3985
rect 8535 3965 8550 3985
rect 8500 3950 8550 3965
rect 8650 4435 8700 4450
rect 8650 4415 8665 4435
rect 8685 4415 8700 4435
rect 8650 4385 8700 4415
rect 8650 4365 8665 4385
rect 8685 4365 8700 4385
rect 8650 4335 8700 4365
rect 8650 4315 8665 4335
rect 8685 4315 8700 4335
rect 8650 4285 8700 4315
rect 8650 4265 8665 4285
rect 8685 4265 8700 4285
rect 8650 4235 8700 4265
rect 8650 4215 8665 4235
rect 8685 4215 8700 4235
rect 8650 4185 8700 4215
rect 8650 4165 8665 4185
rect 8685 4165 8700 4185
rect 8650 4135 8700 4165
rect 8650 4115 8665 4135
rect 8685 4115 8700 4135
rect 8650 4085 8700 4115
rect 8650 4065 8665 4085
rect 8685 4065 8700 4085
rect 8650 4035 8700 4065
rect 8650 4015 8665 4035
rect 8685 4015 8700 4035
rect 8650 3985 8700 4015
rect 8650 3965 8665 3985
rect 8685 3965 8700 3985
rect 8650 3950 8700 3965
rect 8800 4435 8850 4500
rect 8800 4415 8815 4435
rect 8835 4415 8850 4435
rect 8800 4385 8850 4415
rect 8800 4365 8815 4385
rect 8835 4365 8850 4385
rect 8800 4335 8850 4365
rect 8800 4315 8815 4335
rect 8835 4315 8850 4335
rect 8800 4285 8850 4315
rect 8800 4265 8815 4285
rect 8835 4265 8850 4285
rect 8800 4235 8850 4265
rect 8800 4215 8815 4235
rect 8835 4215 8850 4235
rect 8800 4185 8850 4215
rect 8800 4165 8815 4185
rect 8835 4165 8850 4185
rect 8800 4135 8850 4165
rect 8800 4115 8815 4135
rect 8835 4115 8850 4135
rect 8800 4085 8850 4115
rect 8800 4065 8815 4085
rect 8835 4065 8850 4085
rect 8800 4035 8850 4065
rect 8800 4015 8815 4035
rect 8835 4015 8850 4035
rect 8800 3985 8850 4015
rect 8800 3965 8815 3985
rect 8835 3965 8850 3985
rect 8800 3950 8850 3965
rect 8950 4435 9000 4450
rect 8950 4415 8965 4435
rect 8985 4415 9000 4435
rect 8950 4385 9000 4415
rect 8950 4365 8965 4385
rect 8985 4365 9000 4385
rect 8950 4335 9000 4365
rect 8950 4315 8965 4335
rect 8985 4315 9000 4335
rect 8950 4285 9000 4315
rect 8950 4265 8965 4285
rect 8985 4265 9000 4285
rect 8950 4235 9000 4265
rect 8950 4215 8965 4235
rect 8985 4215 9000 4235
rect 8950 4185 9000 4215
rect 8950 4165 8965 4185
rect 8985 4165 9000 4185
rect 8950 4135 9000 4165
rect 8950 4115 8965 4135
rect 8985 4115 9000 4135
rect 8950 4085 9000 4115
rect 8950 4065 8965 4085
rect 8985 4065 9000 4085
rect 8950 4035 9000 4065
rect 8950 4015 8965 4035
rect 8985 4015 9000 4035
rect 8950 3985 9000 4015
rect 8950 3965 8965 3985
rect 8985 3965 9000 3985
rect 8950 3950 9000 3965
rect 9100 4435 9150 4500
rect 9100 4415 9115 4435
rect 9135 4415 9150 4435
rect 9100 4385 9150 4415
rect 9100 4365 9115 4385
rect 9135 4365 9150 4385
rect 9100 4335 9150 4365
rect 9100 4315 9115 4335
rect 9135 4315 9150 4335
rect 9100 4285 9150 4315
rect 9100 4265 9115 4285
rect 9135 4265 9150 4285
rect 9100 4235 9150 4265
rect 9100 4215 9115 4235
rect 9135 4215 9150 4235
rect 9100 4185 9150 4215
rect 9100 4165 9115 4185
rect 9135 4165 9150 4185
rect 9100 4135 9150 4165
rect 9100 4115 9115 4135
rect 9135 4115 9150 4135
rect 9100 4085 9150 4115
rect 9100 4065 9115 4085
rect 9135 4065 9150 4085
rect 9100 4035 9150 4065
rect 9100 4015 9115 4035
rect 9135 4015 9150 4035
rect 9100 3985 9150 4015
rect 9100 3965 9115 3985
rect 9135 3965 9150 3985
rect 9100 3950 9150 3965
rect 9250 4435 9300 4450
rect 9250 4415 9265 4435
rect 9285 4415 9300 4435
rect 9250 4385 9300 4415
rect 9250 4365 9265 4385
rect 9285 4365 9300 4385
rect 9250 4335 9300 4365
rect 9250 4315 9265 4335
rect 9285 4315 9300 4335
rect 9250 4285 9300 4315
rect 9250 4265 9265 4285
rect 9285 4265 9300 4285
rect 9250 4235 9300 4265
rect 9250 4215 9265 4235
rect 9285 4215 9300 4235
rect 9250 4185 9300 4215
rect 9250 4165 9265 4185
rect 9285 4165 9300 4185
rect 9250 4135 9300 4165
rect 9250 4115 9265 4135
rect 9285 4115 9300 4135
rect 9250 4085 9300 4115
rect 9250 4065 9265 4085
rect 9285 4065 9300 4085
rect 9250 4035 9300 4065
rect 9250 4015 9265 4035
rect 9285 4015 9300 4035
rect 9250 3985 9300 4015
rect 9250 3965 9265 3985
rect 9285 3965 9300 3985
rect 9250 3950 9300 3965
rect 9400 4435 9450 4500
rect 9400 4415 9415 4435
rect 9435 4415 9450 4435
rect 9400 4385 9450 4415
rect 9400 4365 9415 4385
rect 9435 4365 9450 4385
rect 9400 4335 9450 4365
rect 9400 4315 9415 4335
rect 9435 4315 9450 4335
rect 9400 4285 9450 4315
rect 9400 4265 9415 4285
rect 9435 4265 9450 4285
rect 9400 4235 9450 4265
rect 9400 4215 9415 4235
rect 9435 4215 9450 4235
rect 9400 4185 9450 4215
rect 9400 4165 9415 4185
rect 9435 4165 9450 4185
rect 9400 4135 9450 4165
rect 9400 4115 9415 4135
rect 9435 4115 9450 4135
rect 9400 4085 9450 4115
rect 9400 4065 9415 4085
rect 9435 4065 9450 4085
rect 9400 4035 9450 4065
rect 9400 4015 9415 4035
rect 9435 4015 9450 4035
rect 9400 3985 9450 4015
rect 9400 3965 9415 3985
rect 9435 3965 9450 3985
rect 9400 3950 9450 3965
rect 9550 4435 9600 4450
rect 9550 4415 9565 4435
rect 9585 4415 9600 4435
rect 9550 4385 9600 4415
rect 9550 4365 9565 4385
rect 9585 4365 9600 4385
rect 9550 4335 9600 4365
rect 9550 4315 9565 4335
rect 9585 4315 9600 4335
rect 9550 4285 9600 4315
rect 9550 4265 9565 4285
rect 9585 4265 9600 4285
rect 9550 4235 9600 4265
rect 9550 4215 9565 4235
rect 9585 4215 9600 4235
rect 9550 4185 9600 4215
rect 9550 4165 9565 4185
rect 9585 4165 9600 4185
rect 9550 4135 9600 4165
rect 9550 4115 9565 4135
rect 9585 4115 9600 4135
rect 9550 4085 9600 4115
rect 9550 4065 9565 4085
rect 9585 4065 9600 4085
rect 9550 4035 9600 4065
rect 9550 4015 9565 4035
rect 9585 4015 9600 4035
rect 9550 3985 9600 4015
rect 9550 3965 9565 3985
rect 9585 3965 9600 3985
rect 9550 3950 9600 3965
rect 9700 4435 9750 4500
rect 9700 4415 9715 4435
rect 9735 4415 9750 4435
rect 9700 4385 9750 4415
rect 9700 4365 9715 4385
rect 9735 4365 9750 4385
rect 9700 4335 9750 4365
rect 9700 4315 9715 4335
rect 9735 4315 9750 4335
rect 9700 4285 9750 4315
rect 9700 4265 9715 4285
rect 9735 4265 9750 4285
rect 9700 4235 9750 4265
rect 9700 4215 9715 4235
rect 9735 4215 9750 4235
rect 9700 4185 9750 4215
rect 9700 4165 9715 4185
rect 9735 4165 9750 4185
rect 9700 4135 9750 4165
rect 9700 4115 9715 4135
rect 9735 4115 9750 4135
rect 9700 4085 9750 4115
rect 9700 4065 9715 4085
rect 9735 4065 9750 4085
rect 9700 4035 9750 4065
rect 9700 4015 9715 4035
rect 9735 4015 9750 4035
rect 9700 3985 9750 4015
rect 9700 3965 9715 3985
rect 9735 3965 9750 3985
rect 9700 3950 9750 3965
rect 9850 4435 9900 4450
rect 9850 4415 9865 4435
rect 9885 4415 9900 4435
rect 9850 4385 9900 4415
rect 9850 4365 9865 4385
rect 9885 4365 9900 4385
rect 9850 4335 9900 4365
rect 9850 4315 9865 4335
rect 9885 4315 9900 4335
rect 9850 4285 9900 4315
rect 9850 4265 9865 4285
rect 9885 4265 9900 4285
rect 9850 4235 9900 4265
rect 9850 4215 9865 4235
rect 9885 4215 9900 4235
rect 9850 4185 9900 4215
rect 9850 4165 9865 4185
rect 9885 4165 9900 4185
rect 9850 4135 9900 4165
rect 9850 4115 9865 4135
rect 9885 4115 9900 4135
rect 9850 4085 9900 4115
rect 9850 4065 9865 4085
rect 9885 4065 9900 4085
rect 9850 4035 9900 4065
rect 9850 4015 9865 4035
rect 9885 4015 9900 4035
rect 9850 3985 9900 4015
rect 9850 3965 9865 3985
rect 9885 3965 9900 3985
rect 9850 3950 9900 3965
rect 10000 4435 10050 4500
rect 10000 4415 10015 4435
rect 10035 4415 10050 4435
rect 10000 4385 10050 4415
rect 10000 4365 10015 4385
rect 10035 4365 10050 4385
rect 10000 4335 10050 4365
rect 10000 4315 10015 4335
rect 10035 4315 10050 4335
rect 10000 4285 10050 4315
rect 10000 4265 10015 4285
rect 10035 4265 10050 4285
rect 10000 4235 10050 4265
rect 10000 4215 10015 4235
rect 10035 4215 10050 4235
rect 10000 4185 10050 4215
rect 10000 4165 10015 4185
rect 10035 4165 10050 4185
rect 10000 4135 10050 4165
rect 10000 4115 10015 4135
rect 10035 4115 10050 4135
rect 10000 4085 10050 4115
rect 10000 4065 10015 4085
rect 10035 4065 10050 4085
rect 10000 4035 10050 4065
rect 10000 4015 10015 4035
rect 10035 4015 10050 4035
rect 10000 3985 10050 4015
rect 10000 3965 10015 3985
rect 10035 3965 10050 3985
rect 10000 3950 10050 3965
rect 10150 4435 10200 4450
rect 10150 4415 10165 4435
rect 10185 4415 10200 4435
rect 10150 4385 10200 4415
rect 10150 4365 10165 4385
rect 10185 4365 10200 4385
rect 10150 4335 10200 4365
rect 10150 4315 10165 4335
rect 10185 4315 10200 4335
rect 10150 4285 10200 4315
rect 10150 4265 10165 4285
rect 10185 4265 10200 4285
rect 10150 4235 10200 4265
rect 10150 4215 10165 4235
rect 10185 4215 10200 4235
rect 10150 4185 10200 4215
rect 10150 4165 10165 4185
rect 10185 4165 10200 4185
rect 10150 4135 10200 4165
rect 10150 4115 10165 4135
rect 10185 4115 10200 4135
rect 10150 4085 10200 4115
rect 10150 4065 10165 4085
rect 10185 4065 10200 4085
rect 10150 4035 10200 4065
rect 10150 4015 10165 4035
rect 10185 4015 10200 4035
rect 10150 3985 10200 4015
rect 10150 3965 10165 3985
rect 10185 3965 10200 3985
rect 10150 3950 10200 3965
rect 10300 4435 10350 4500
rect 10300 4415 10315 4435
rect 10335 4415 10350 4435
rect 10300 4385 10350 4415
rect 10300 4365 10315 4385
rect 10335 4365 10350 4385
rect 10300 4335 10350 4365
rect 10300 4315 10315 4335
rect 10335 4315 10350 4335
rect 10300 4285 10350 4315
rect 10300 4265 10315 4285
rect 10335 4265 10350 4285
rect 10300 4235 10350 4265
rect 10300 4215 10315 4235
rect 10335 4215 10350 4235
rect 10300 4185 10350 4215
rect 10300 4165 10315 4185
rect 10335 4165 10350 4185
rect 10300 4135 10350 4165
rect 10300 4115 10315 4135
rect 10335 4115 10350 4135
rect 10300 4085 10350 4115
rect 10300 4065 10315 4085
rect 10335 4065 10350 4085
rect 10300 4035 10350 4065
rect 10300 4015 10315 4035
rect 10335 4015 10350 4035
rect 10300 3985 10350 4015
rect 10300 3965 10315 3985
rect 10335 3965 10350 3985
rect 10300 3950 10350 3965
rect 10450 4435 10500 4450
rect 10450 4415 10465 4435
rect 10485 4415 10500 4435
rect 10450 4385 10500 4415
rect 10450 4365 10465 4385
rect 10485 4365 10500 4385
rect 10450 4335 10500 4365
rect 10450 4315 10465 4335
rect 10485 4315 10500 4335
rect 10450 4285 10500 4315
rect 10450 4265 10465 4285
rect 10485 4265 10500 4285
rect 10450 4235 10500 4265
rect 10450 4215 10465 4235
rect 10485 4215 10500 4235
rect 10450 4185 10500 4215
rect 10450 4165 10465 4185
rect 10485 4165 10500 4185
rect 10450 4135 10500 4165
rect 10450 4115 10465 4135
rect 10485 4115 10500 4135
rect 10450 4085 10500 4115
rect 10450 4065 10465 4085
rect 10485 4065 10500 4085
rect 10450 4035 10500 4065
rect 10450 4015 10465 4035
rect 10485 4015 10500 4035
rect 10450 3985 10500 4015
rect 10450 3965 10465 3985
rect 10485 3965 10500 3985
rect 10450 3950 10500 3965
rect 10600 4435 10650 4500
rect 10600 4415 10615 4435
rect 10635 4415 10650 4435
rect 10600 4385 10650 4415
rect 10600 4365 10615 4385
rect 10635 4365 10650 4385
rect 10600 4335 10650 4365
rect 10600 4315 10615 4335
rect 10635 4315 10650 4335
rect 10600 4285 10650 4315
rect 10600 4265 10615 4285
rect 10635 4265 10650 4285
rect 10600 4235 10650 4265
rect 10600 4215 10615 4235
rect 10635 4215 10650 4235
rect 10600 4185 10650 4215
rect 10600 4165 10615 4185
rect 10635 4165 10650 4185
rect 10600 4135 10650 4165
rect 10600 4115 10615 4135
rect 10635 4115 10650 4135
rect 10600 4085 10650 4115
rect 10600 4065 10615 4085
rect 10635 4065 10650 4085
rect 10600 4035 10650 4065
rect 10600 4015 10615 4035
rect 10635 4015 10650 4035
rect 10600 3985 10650 4015
rect 10600 3965 10615 3985
rect 10635 3965 10650 3985
rect 10600 3950 10650 3965
rect 10750 4435 10800 4450
rect 10750 4415 10765 4435
rect 10785 4415 10800 4435
rect 10750 4385 10800 4415
rect 10750 4365 10765 4385
rect 10785 4365 10800 4385
rect 10750 4335 10800 4365
rect 10750 4315 10765 4335
rect 10785 4315 10800 4335
rect 10750 4285 10800 4315
rect 10750 4265 10765 4285
rect 10785 4265 10800 4285
rect 10750 4235 10800 4265
rect 10750 4215 10765 4235
rect 10785 4215 10800 4235
rect 10750 4185 10800 4215
rect 10750 4165 10765 4185
rect 10785 4165 10800 4185
rect 10750 4135 10800 4165
rect 10750 4115 10765 4135
rect 10785 4115 10800 4135
rect 10750 4085 10800 4115
rect 10750 4065 10765 4085
rect 10785 4065 10800 4085
rect 10750 4035 10800 4065
rect 10750 4015 10765 4035
rect 10785 4015 10800 4035
rect 10750 3985 10800 4015
rect 10750 3965 10765 3985
rect 10785 3965 10800 3985
rect 10750 3950 10800 3965
rect 11350 4435 11400 4450
rect 11350 4415 11365 4435
rect 11385 4415 11400 4435
rect 11350 4385 11400 4415
rect 11350 4365 11365 4385
rect 11385 4365 11400 4385
rect 11350 4335 11400 4365
rect 11350 4315 11365 4335
rect 11385 4315 11400 4335
rect 11350 4285 11400 4315
rect 11350 4265 11365 4285
rect 11385 4265 11400 4285
rect 11350 4235 11400 4265
rect 11350 4215 11365 4235
rect 11385 4215 11400 4235
rect 11350 4185 11400 4215
rect 11350 4165 11365 4185
rect 11385 4165 11400 4185
rect 11350 4135 11400 4165
rect 11350 4115 11365 4135
rect 11385 4115 11400 4135
rect 11350 4085 11400 4115
rect 11350 4065 11365 4085
rect 11385 4065 11400 4085
rect 11350 4035 11400 4065
rect 11350 4015 11365 4035
rect 11385 4015 11400 4035
rect 11350 3985 11400 4015
rect 11350 3965 11365 3985
rect 11385 3965 11400 3985
rect 11350 3950 11400 3965
rect 11950 4435 12000 4450
rect 11950 4415 11965 4435
rect 11985 4415 12000 4435
rect 11950 4385 12000 4415
rect 11950 4365 11965 4385
rect 11985 4365 12000 4385
rect 11950 4335 12000 4365
rect 11950 4315 11965 4335
rect 11985 4315 12000 4335
rect 11950 4285 12000 4315
rect 11950 4265 11965 4285
rect 11985 4265 12000 4285
rect 11950 4235 12000 4265
rect 11950 4215 11965 4235
rect 11985 4215 12000 4235
rect 11950 4185 12000 4215
rect 11950 4165 11965 4185
rect 11985 4165 12000 4185
rect 11950 4135 12000 4165
rect 11950 4115 11965 4135
rect 11985 4115 12000 4135
rect 11950 4085 12000 4115
rect 11950 4065 11965 4085
rect 11985 4065 12000 4085
rect 11950 4035 12000 4065
rect 11950 4015 11965 4035
rect 11985 4015 12000 4035
rect 11950 3985 12000 4015
rect 11950 3965 11965 3985
rect 11985 3965 12000 3985
rect 11950 3950 12000 3965
rect 12550 4435 12600 4450
rect 12550 4415 12565 4435
rect 12585 4415 12600 4435
rect 12550 4385 12600 4415
rect 12550 4365 12565 4385
rect 12585 4365 12600 4385
rect 12550 4335 12600 4365
rect 12550 4315 12565 4335
rect 12585 4315 12600 4335
rect 12550 4285 12600 4315
rect 12550 4265 12565 4285
rect 12585 4265 12600 4285
rect 12550 4235 12600 4265
rect 12550 4215 12565 4235
rect 12585 4215 12600 4235
rect 12550 4185 12600 4215
rect 12550 4165 12565 4185
rect 12585 4165 12600 4185
rect 12550 4135 12600 4165
rect 12550 4115 12565 4135
rect 12585 4115 12600 4135
rect 12550 4085 12600 4115
rect 12550 4065 12565 4085
rect 12585 4065 12600 4085
rect 12550 4035 12600 4065
rect 12550 4015 12565 4035
rect 12585 4015 12600 4035
rect 12550 3985 12600 4015
rect 12550 3965 12565 3985
rect 12585 3965 12600 3985
rect 12550 3950 12600 3965
rect 13150 4435 13200 4450
rect 13150 4415 13165 4435
rect 13185 4415 13200 4435
rect 13150 4385 13200 4415
rect 13150 4365 13165 4385
rect 13185 4365 13200 4385
rect 13150 4335 13200 4365
rect 13150 4315 13165 4335
rect 13185 4315 13200 4335
rect 13150 4285 13200 4315
rect 13150 4265 13165 4285
rect 13185 4265 13200 4285
rect 13150 4235 13200 4265
rect 13150 4215 13165 4235
rect 13185 4215 13200 4235
rect 13150 4185 13200 4215
rect 13150 4165 13165 4185
rect 13185 4165 13200 4185
rect 13150 4135 13200 4165
rect 13150 4115 13165 4135
rect 13185 4115 13200 4135
rect 13150 4085 13200 4115
rect 13150 4065 13165 4085
rect 13185 4065 13200 4085
rect 13150 4035 13200 4065
rect 13150 4015 13165 4035
rect 13185 4015 13200 4035
rect 13150 3985 13200 4015
rect 13150 3965 13165 3985
rect 13185 3965 13200 3985
rect 13150 3950 13200 3965
rect 13750 4435 13800 4450
rect 13750 4415 13765 4435
rect 13785 4415 13800 4435
rect 13750 4385 13800 4415
rect 13750 4365 13765 4385
rect 13785 4365 13800 4385
rect 13750 4335 13800 4365
rect 13750 4315 13765 4335
rect 13785 4315 13800 4335
rect 13750 4285 13800 4315
rect 13750 4265 13765 4285
rect 13785 4265 13800 4285
rect 13750 4235 13800 4265
rect 13750 4215 13765 4235
rect 13785 4215 13800 4235
rect 13750 4185 13800 4215
rect 13750 4165 13765 4185
rect 13785 4165 13800 4185
rect 13750 4135 13800 4165
rect 13750 4115 13765 4135
rect 13785 4115 13800 4135
rect 13750 4085 13800 4115
rect 13750 4065 13765 4085
rect 13785 4065 13800 4085
rect 13750 4035 13800 4065
rect 13750 4015 13765 4035
rect 13785 4015 13800 4035
rect 13750 3985 13800 4015
rect 13750 3965 13765 3985
rect 13785 3965 13800 3985
rect 13750 3950 13800 3965
rect 14350 4435 14400 4450
rect 14350 4415 14365 4435
rect 14385 4415 14400 4435
rect 14350 4385 14400 4415
rect 14350 4365 14365 4385
rect 14385 4365 14400 4385
rect 14350 4335 14400 4365
rect 14350 4315 14365 4335
rect 14385 4315 14400 4335
rect 14350 4285 14400 4315
rect 14350 4265 14365 4285
rect 14385 4265 14400 4285
rect 14350 4235 14400 4265
rect 14350 4215 14365 4235
rect 14385 4215 14400 4235
rect 14350 4185 14400 4215
rect 14350 4165 14365 4185
rect 14385 4165 14400 4185
rect 14350 4135 14400 4165
rect 14350 4115 14365 4135
rect 14385 4115 14400 4135
rect 14350 4085 14400 4115
rect 14350 4065 14365 4085
rect 14385 4065 14400 4085
rect 14350 4035 14400 4065
rect 14350 4015 14365 4035
rect 14385 4015 14400 4035
rect 14350 3985 14400 4015
rect 14350 3965 14365 3985
rect 14385 3965 14400 3985
rect 14350 3950 14400 3965
rect 14950 4435 15000 4450
rect 14950 4415 14965 4435
rect 14985 4415 15000 4435
rect 14950 4385 15000 4415
rect 14950 4365 14965 4385
rect 14985 4365 15000 4385
rect 14950 4335 15000 4365
rect 14950 4315 14965 4335
rect 14985 4315 15000 4335
rect 14950 4285 15000 4315
rect 14950 4265 14965 4285
rect 14985 4265 15000 4285
rect 14950 4235 15000 4265
rect 14950 4215 14965 4235
rect 14985 4215 15000 4235
rect 14950 4185 15000 4215
rect 14950 4165 14965 4185
rect 14985 4165 15000 4185
rect 14950 4135 15000 4165
rect 14950 4115 14965 4135
rect 14985 4115 15000 4135
rect 14950 4085 15000 4115
rect 14950 4065 14965 4085
rect 14985 4065 15000 4085
rect 14950 4035 15000 4065
rect 14950 4015 14965 4035
rect 14985 4015 15000 4035
rect 14950 3985 15000 4015
rect 14950 3965 14965 3985
rect 14985 3965 15000 3985
rect 14950 3950 15000 3965
rect 15550 4435 15600 4450
rect 15550 4415 15565 4435
rect 15585 4415 15600 4435
rect 15550 4385 15600 4415
rect 15550 4365 15565 4385
rect 15585 4365 15600 4385
rect 15550 4335 15600 4365
rect 15550 4315 15565 4335
rect 15585 4315 15600 4335
rect 15550 4285 15600 4315
rect 15550 4265 15565 4285
rect 15585 4265 15600 4285
rect 15550 4235 15600 4265
rect 15550 4215 15565 4235
rect 15585 4215 15600 4235
rect 15550 4185 15600 4215
rect 15550 4165 15565 4185
rect 15585 4165 15600 4185
rect 15550 4135 15600 4165
rect 15550 4115 15565 4135
rect 15585 4115 15600 4135
rect 15550 4085 15600 4115
rect 15550 4065 15565 4085
rect 15585 4065 15600 4085
rect 15550 4035 15600 4065
rect 15550 4015 15565 4035
rect 15585 4015 15600 4035
rect 15550 3985 15600 4015
rect 15550 3965 15565 3985
rect 15585 3965 15600 3985
rect 15550 3950 15600 3965
rect 16150 4435 16200 4450
rect 16150 4415 16165 4435
rect 16185 4415 16200 4435
rect 16150 4385 16200 4415
rect 16150 4365 16165 4385
rect 16185 4365 16200 4385
rect 16150 4335 16200 4365
rect 16150 4315 16165 4335
rect 16185 4315 16200 4335
rect 16150 4285 16200 4315
rect 16150 4265 16165 4285
rect 16185 4265 16200 4285
rect 16150 4235 16200 4265
rect 16150 4215 16165 4235
rect 16185 4215 16200 4235
rect 16150 4185 16200 4215
rect 16150 4165 16165 4185
rect 16185 4165 16200 4185
rect 16150 4135 16200 4165
rect 16150 4115 16165 4135
rect 16185 4115 16200 4135
rect 16150 4085 16200 4115
rect 16150 4065 16165 4085
rect 16185 4065 16200 4085
rect 16150 4035 16200 4065
rect 16150 4015 16165 4035
rect 16185 4015 16200 4035
rect 16150 3985 16200 4015
rect 16150 3965 16165 3985
rect 16185 3965 16200 3985
rect 16150 3950 16200 3965
rect 16300 4435 16350 4450
rect 16300 4415 16315 4435
rect 16335 4415 16350 4435
rect 16300 4385 16350 4415
rect 16300 4365 16315 4385
rect 16335 4365 16350 4385
rect 16300 4335 16350 4365
rect 16300 4315 16315 4335
rect 16335 4315 16350 4335
rect 16300 4285 16350 4315
rect 16300 4265 16315 4285
rect 16335 4265 16350 4285
rect 16300 4235 16350 4265
rect 16300 4215 16315 4235
rect 16335 4215 16350 4235
rect 16300 4185 16350 4215
rect 16300 4165 16315 4185
rect 16335 4165 16350 4185
rect 16300 4135 16350 4165
rect 16300 4115 16315 4135
rect 16335 4115 16350 4135
rect 16300 4085 16350 4115
rect 16300 4065 16315 4085
rect 16335 4065 16350 4085
rect 16300 4035 16350 4065
rect 16300 4015 16315 4035
rect 16335 4015 16350 4035
rect 16300 3985 16350 4015
rect 16300 3965 16315 3985
rect 16335 3965 16350 3985
rect 16300 3950 16350 3965
rect 16450 4435 16500 4450
rect 16450 4415 16465 4435
rect 16485 4415 16500 4435
rect 16450 4385 16500 4415
rect 16450 4365 16465 4385
rect 16485 4365 16500 4385
rect 16450 4335 16500 4365
rect 16450 4315 16465 4335
rect 16485 4315 16500 4335
rect 16450 4285 16500 4315
rect 16450 4265 16465 4285
rect 16485 4265 16500 4285
rect 16450 4235 16500 4265
rect 16450 4215 16465 4235
rect 16485 4215 16500 4235
rect 16450 4185 16500 4215
rect 16450 4165 16465 4185
rect 16485 4165 16500 4185
rect 16450 4135 16500 4165
rect 16450 4115 16465 4135
rect 16485 4115 16500 4135
rect 16450 4085 16500 4115
rect 16450 4065 16465 4085
rect 16485 4065 16500 4085
rect 16450 4035 16500 4065
rect 16450 4015 16465 4035
rect 16485 4015 16500 4035
rect 16450 3985 16500 4015
rect 16450 3965 16465 3985
rect 16485 3965 16500 3985
rect 16450 3950 16500 3965
rect 16600 4435 16650 4450
rect 16600 4415 16615 4435
rect 16635 4415 16650 4435
rect 16600 4385 16650 4415
rect 16600 4365 16615 4385
rect 16635 4365 16650 4385
rect 16600 4335 16650 4365
rect 16600 4315 16615 4335
rect 16635 4315 16650 4335
rect 16600 4285 16650 4315
rect 16600 4265 16615 4285
rect 16635 4265 16650 4285
rect 16600 4235 16650 4265
rect 16600 4215 16615 4235
rect 16635 4215 16650 4235
rect 16600 4185 16650 4215
rect 16600 4165 16615 4185
rect 16635 4165 16650 4185
rect 16600 4135 16650 4165
rect 16600 4115 16615 4135
rect 16635 4115 16650 4135
rect 16600 4085 16650 4115
rect 16600 4065 16615 4085
rect 16635 4065 16650 4085
rect 16600 4035 16650 4065
rect 16600 4015 16615 4035
rect 16635 4015 16650 4035
rect 16600 3985 16650 4015
rect 16600 3965 16615 3985
rect 16635 3965 16650 3985
rect 16600 3950 16650 3965
rect 16750 4435 16800 4450
rect 16750 4415 16765 4435
rect 16785 4415 16800 4435
rect 16750 4385 16800 4415
rect 16750 4365 16765 4385
rect 16785 4365 16800 4385
rect 16750 4335 16800 4365
rect 16750 4315 16765 4335
rect 16785 4315 16800 4335
rect 16750 4285 16800 4315
rect 16750 4265 16765 4285
rect 16785 4265 16800 4285
rect 16750 4235 16800 4265
rect 16750 4215 16765 4235
rect 16785 4215 16800 4235
rect 16750 4185 16800 4215
rect 16750 4165 16765 4185
rect 16785 4165 16800 4185
rect 16750 4135 16800 4165
rect 16750 4115 16765 4135
rect 16785 4115 16800 4135
rect 16750 4085 16800 4115
rect 16750 4065 16765 4085
rect 16785 4065 16800 4085
rect 16750 4035 16800 4065
rect 16750 4015 16765 4035
rect 16785 4015 16800 4035
rect 16750 3985 16800 4015
rect 16750 3965 16765 3985
rect 16785 3965 16800 3985
rect 16750 3950 16800 3965
rect 16900 4435 16950 4450
rect 16900 4415 16915 4435
rect 16935 4415 16950 4435
rect 16900 4385 16950 4415
rect 16900 4365 16915 4385
rect 16935 4365 16950 4385
rect 16900 4335 16950 4365
rect 16900 4315 16915 4335
rect 16935 4315 16950 4335
rect 16900 4285 16950 4315
rect 16900 4265 16915 4285
rect 16935 4265 16950 4285
rect 16900 4235 16950 4265
rect 16900 4215 16915 4235
rect 16935 4215 16950 4235
rect 16900 4185 16950 4215
rect 16900 4165 16915 4185
rect 16935 4165 16950 4185
rect 16900 4135 16950 4165
rect 16900 4115 16915 4135
rect 16935 4115 16950 4135
rect 16900 4085 16950 4115
rect 16900 4065 16915 4085
rect 16935 4065 16950 4085
rect 16900 4035 16950 4065
rect 16900 4015 16915 4035
rect 16935 4015 16950 4035
rect 16900 3985 16950 4015
rect 16900 3965 16915 3985
rect 16935 3965 16950 3985
rect 16900 3950 16950 3965
rect 17050 4435 17100 4450
rect 17050 4415 17065 4435
rect 17085 4415 17100 4435
rect 17050 4385 17100 4415
rect 17050 4365 17065 4385
rect 17085 4365 17100 4385
rect 17050 4335 17100 4365
rect 17050 4315 17065 4335
rect 17085 4315 17100 4335
rect 17050 4285 17100 4315
rect 17050 4265 17065 4285
rect 17085 4265 17100 4285
rect 17050 4235 17100 4265
rect 17050 4215 17065 4235
rect 17085 4215 17100 4235
rect 17050 4185 17100 4215
rect 17050 4165 17065 4185
rect 17085 4165 17100 4185
rect 17050 4135 17100 4165
rect 17050 4115 17065 4135
rect 17085 4115 17100 4135
rect 17050 4085 17100 4115
rect 17050 4065 17065 4085
rect 17085 4065 17100 4085
rect 17050 4035 17100 4065
rect 17050 4015 17065 4035
rect 17085 4015 17100 4035
rect 17050 3985 17100 4015
rect 17050 3965 17065 3985
rect 17085 3965 17100 3985
rect 17050 3950 17100 3965
rect 17200 4435 17250 4450
rect 17200 4415 17215 4435
rect 17235 4415 17250 4435
rect 17200 4385 17250 4415
rect 17200 4365 17215 4385
rect 17235 4365 17250 4385
rect 17200 4335 17250 4365
rect 17200 4315 17215 4335
rect 17235 4315 17250 4335
rect 17200 4285 17250 4315
rect 17200 4265 17215 4285
rect 17235 4265 17250 4285
rect 17200 4235 17250 4265
rect 17200 4215 17215 4235
rect 17235 4215 17250 4235
rect 17200 4185 17250 4215
rect 17200 4165 17215 4185
rect 17235 4165 17250 4185
rect 17200 4135 17250 4165
rect 17200 4115 17215 4135
rect 17235 4115 17250 4135
rect 17200 4085 17250 4115
rect 17200 4065 17215 4085
rect 17235 4065 17250 4085
rect 17200 4035 17250 4065
rect 17200 4015 17215 4035
rect 17235 4015 17250 4035
rect 17200 3985 17250 4015
rect 17200 3965 17215 3985
rect 17235 3965 17250 3985
rect 17200 3950 17250 3965
rect 17350 4435 17400 4450
rect 17350 4415 17365 4435
rect 17385 4415 17400 4435
rect 17350 4385 17400 4415
rect 17350 4365 17365 4385
rect 17385 4365 17400 4385
rect 17350 4335 17400 4365
rect 17350 4315 17365 4335
rect 17385 4315 17400 4335
rect 17350 4285 17400 4315
rect 17350 4265 17365 4285
rect 17385 4265 17400 4285
rect 17350 4235 17400 4265
rect 17350 4215 17365 4235
rect 17385 4215 17400 4235
rect 17350 4185 17400 4215
rect 17350 4165 17365 4185
rect 17385 4165 17400 4185
rect 17350 4135 17400 4165
rect 17350 4115 17365 4135
rect 17385 4115 17400 4135
rect 17350 4085 17400 4115
rect 17350 4065 17365 4085
rect 17385 4065 17400 4085
rect 17350 4035 17400 4065
rect 17350 4015 17365 4035
rect 17385 4015 17400 4035
rect 17350 3985 17400 4015
rect 17350 3965 17365 3985
rect 17385 3965 17400 3985
rect 17350 3950 17400 3965
rect 17950 4435 18000 4450
rect 17950 4415 17965 4435
rect 17985 4415 18000 4435
rect 17950 4385 18000 4415
rect 17950 4365 17965 4385
rect 17985 4365 18000 4385
rect 17950 4335 18000 4365
rect 17950 4315 17965 4335
rect 17985 4315 18000 4335
rect 17950 4285 18000 4315
rect 17950 4265 17965 4285
rect 17985 4265 18000 4285
rect 17950 4235 18000 4265
rect 17950 4215 17965 4235
rect 17985 4215 18000 4235
rect 17950 4185 18000 4215
rect 17950 4165 17965 4185
rect 17985 4165 18000 4185
rect 17950 4135 18000 4165
rect 17950 4115 17965 4135
rect 17985 4115 18000 4135
rect 17950 4085 18000 4115
rect 17950 4065 17965 4085
rect 17985 4065 18000 4085
rect 17950 4035 18000 4065
rect 17950 4015 17965 4035
rect 17985 4015 18000 4035
rect 17950 3985 18000 4015
rect 17950 3965 17965 3985
rect 17985 3965 18000 3985
rect 17950 3950 18000 3965
rect 18550 4435 18600 4450
rect 18550 4415 18565 4435
rect 18585 4415 18600 4435
rect 18550 4385 18600 4415
rect 18550 4365 18565 4385
rect 18585 4365 18600 4385
rect 18550 4335 18600 4365
rect 18550 4315 18565 4335
rect 18585 4315 18600 4335
rect 18550 4285 18600 4315
rect 18550 4265 18565 4285
rect 18585 4265 18600 4285
rect 18550 4235 18600 4265
rect 18550 4215 18565 4235
rect 18585 4215 18600 4235
rect 18550 4185 18600 4215
rect 18550 4165 18565 4185
rect 18585 4165 18600 4185
rect 18550 4135 18600 4165
rect 18550 4115 18565 4135
rect 18585 4115 18600 4135
rect 18550 4085 18600 4115
rect 18550 4065 18565 4085
rect 18585 4065 18600 4085
rect 18550 4035 18600 4065
rect 18550 4015 18565 4035
rect 18585 4015 18600 4035
rect 18550 3985 18600 4015
rect 18550 3965 18565 3985
rect 18585 3965 18600 3985
rect 18550 3950 18600 3965
rect 18700 4435 18750 4450
rect 18700 4415 18715 4435
rect 18735 4415 18750 4435
rect 18700 4385 18750 4415
rect 18700 4365 18715 4385
rect 18735 4365 18750 4385
rect 18700 4335 18750 4365
rect 18700 4315 18715 4335
rect 18735 4315 18750 4335
rect 18700 4285 18750 4315
rect 18700 4265 18715 4285
rect 18735 4265 18750 4285
rect 18700 4235 18750 4265
rect 18700 4215 18715 4235
rect 18735 4215 18750 4235
rect 18700 4185 18750 4215
rect 18700 4165 18715 4185
rect 18735 4165 18750 4185
rect 18700 4135 18750 4165
rect 18700 4115 18715 4135
rect 18735 4115 18750 4135
rect 18700 4085 18750 4115
rect 18700 4065 18715 4085
rect 18735 4065 18750 4085
rect 18700 4035 18750 4065
rect 18700 4015 18715 4035
rect 18735 4015 18750 4035
rect 18700 3985 18750 4015
rect 18700 3965 18715 3985
rect 18735 3965 18750 3985
rect 18700 3950 18750 3965
rect 18850 4435 18900 4450
rect 18850 4415 18865 4435
rect 18885 4415 18900 4435
rect 18850 4385 18900 4415
rect 18850 4365 18865 4385
rect 18885 4365 18900 4385
rect 18850 4335 18900 4365
rect 18850 4315 18865 4335
rect 18885 4315 18900 4335
rect 18850 4285 18900 4315
rect 18850 4265 18865 4285
rect 18885 4265 18900 4285
rect 18850 4235 18900 4265
rect 18850 4215 18865 4235
rect 18885 4215 18900 4235
rect 18850 4185 18900 4215
rect 18850 4165 18865 4185
rect 18885 4165 18900 4185
rect 18850 4135 18900 4165
rect 18850 4115 18865 4135
rect 18885 4115 18900 4135
rect 18850 4085 18900 4115
rect 18850 4065 18865 4085
rect 18885 4065 18900 4085
rect 18850 4035 18900 4065
rect 18850 4015 18865 4035
rect 18885 4015 18900 4035
rect 18850 3985 18900 4015
rect 18850 3965 18865 3985
rect 18885 3965 18900 3985
rect 18850 3950 18900 3965
rect 19000 4435 19050 4450
rect 19000 4415 19015 4435
rect 19035 4415 19050 4435
rect 19000 4385 19050 4415
rect 19000 4365 19015 4385
rect 19035 4365 19050 4385
rect 19000 4335 19050 4365
rect 19000 4315 19015 4335
rect 19035 4315 19050 4335
rect 19000 4285 19050 4315
rect 19000 4265 19015 4285
rect 19035 4265 19050 4285
rect 19000 4235 19050 4265
rect 19000 4215 19015 4235
rect 19035 4215 19050 4235
rect 19000 4185 19050 4215
rect 19000 4165 19015 4185
rect 19035 4165 19050 4185
rect 19000 4135 19050 4165
rect 19000 4115 19015 4135
rect 19035 4115 19050 4135
rect 19000 4085 19050 4115
rect 19000 4065 19015 4085
rect 19035 4065 19050 4085
rect 19000 4035 19050 4065
rect 19000 4015 19015 4035
rect 19035 4015 19050 4035
rect 19000 3985 19050 4015
rect 19000 3965 19015 3985
rect 19035 3965 19050 3985
rect 19000 3950 19050 3965
rect 19150 4435 19200 4450
rect 19150 4415 19165 4435
rect 19185 4415 19200 4435
rect 19150 4385 19200 4415
rect 19150 4365 19165 4385
rect 19185 4365 19200 4385
rect 19150 4335 19200 4365
rect 19150 4315 19165 4335
rect 19185 4315 19200 4335
rect 19150 4285 19200 4315
rect 19150 4265 19165 4285
rect 19185 4265 19200 4285
rect 19150 4235 19200 4265
rect 19150 4215 19165 4235
rect 19185 4215 19200 4235
rect 19150 4185 19200 4215
rect 19150 4165 19165 4185
rect 19185 4165 19200 4185
rect 19150 4135 19200 4165
rect 19150 4115 19165 4135
rect 19185 4115 19200 4135
rect 19150 4085 19200 4115
rect 19150 4065 19165 4085
rect 19185 4065 19200 4085
rect 19150 4035 19200 4065
rect 19150 4015 19165 4035
rect 19185 4015 19200 4035
rect 19150 3985 19200 4015
rect 19150 3965 19165 3985
rect 19185 3965 19200 3985
rect 19150 3950 19200 3965
rect 19300 4435 19350 4450
rect 19300 4415 19315 4435
rect 19335 4415 19350 4435
rect 19300 4385 19350 4415
rect 19300 4365 19315 4385
rect 19335 4365 19350 4385
rect 19300 4335 19350 4365
rect 19300 4315 19315 4335
rect 19335 4315 19350 4335
rect 19300 4285 19350 4315
rect 19300 4265 19315 4285
rect 19335 4265 19350 4285
rect 19300 4235 19350 4265
rect 19300 4215 19315 4235
rect 19335 4215 19350 4235
rect 19300 4185 19350 4215
rect 19300 4165 19315 4185
rect 19335 4165 19350 4185
rect 19300 4135 19350 4165
rect 19300 4115 19315 4135
rect 19335 4115 19350 4135
rect 19300 4085 19350 4115
rect 19300 4065 19315 4085
rect 19335 4065 19350 4085
rect 19300 4035 19350 4065
rect 19300 4015 19315 4035
rect 19335 4015 19350 4035
rect 19300 3985 19350 4015
rect 19300 3965 19315 3985
rect 19335 3965 19350 3985
rect 19300 3950 19350 3965
rect 19450 4435 19500 4450
rect 19450 4415 19465 4435
rect 19485 4415 19500 4435
rect 19450 4385 19500 4415
rect 19450 4365 19465 4385
rect 19485 4365 19500 4385
rect 19450 4335 19500 4365
rect 19450 4315 19465 4335
rect 19485 4315 19500 4335
rect 19450 4285 19500 4315
rect 19450 4265 19465 4285
rect 19485 4265 19500 4285
rect 19450 4235 19500 4265
rect 19450 4215 19465 4235
rect 19485 4215 19500 4235
rect 19450 4185 19500 4215
rect 19450 4165 19465 4185
rect 19485 4165 19500 4185
rect 19450 4135 19500 4165
rect 19450 4115 19465 4135
rect 19485 4115 19500 4135
rect 19450 4085 19500 4115
rect 19450 4065 19465 4085
rect 19485 4065 19500 4085
rect 19450 4035 19500 4065
rect 19450 4015 19465 4035
rect 19485 4015 19500 4035
rect 19450 3985 19500 4015
rect 19450 3965 19465 3985
rect 19485 3965 19500 3985
rect 19450 3950 19500 3965
rect 19600 4435 19650 4450
rect 19600 4415 19615 4435
rect 19635 4415 19650 4435
rect 19600 4385 19650 4415
rect 19600 4365 19615 4385
rect 19635 4365 19650 4385
rect 19600 4335 19650 4365
rect 19600 4315 19615 4335
rect 19635 4315 19650 4335
rect 19600 4285 19650 4315
rect 19600 4265 19615 4285
rect 19635 4265 19650 4285
rect 19600 4235 19650 4265
rect 19600 4215 19615 4235
rect 19635 4215 19650 4235
rect 19600 4185 19650 4215
rect 19600 4165 19615 4185
rect 19635 4165 19650 4185
rect 19600 4135 19650 4165
rect 19600 4115 19615 4135
rect 19635 4115 19650 4135
rect 19600 4085 19650 4115
rect 19600 4065 19615 4085
rect 19635 4065 19650 4085
rect 19600 4035 19650 4065
rect 19600 4015 19615 4035
rect 19635 4015 19650 4035
rect 19600 3985 19650 4015
rect 19600 3965 19615 3985
rect 19635 3965 19650 3985
rect 19600 3950 19650 3965
rect 19750 4435 19800 4450
rect 19750 4415 19765 4435
rect 19785 4415 19800 4435
rect 19750 4385 19800 4415
rect 19750 4365 19765 4385
rect 19785 4365 19800 4385
rect 19750 4335 19800 4365
rect 19750 4315 19765 4335
rect 19785 4315 19800 4335
rect 19750 4285 19800 4315
rect 19750 4265 19765 4285
rect 19785 4265 19800 4285
rect 19750 4235 19800 4265
rect 19750 4215 19765 4235
rect 19785 4215 19800 4235
rect 19750 4185 19800 4215
rect 19750 4165 19765 4185
rect 19785 4165 19800 4185
rect 19750 4135 19800 4165
rect 19750 4115 19765 4135
rect 19785 4115 19800 4135
rect 19750 4085 19800 4115
rect 19750 4065 19765 4085
rect 19785 4065 19800 4085
rect 19750 4035 19800 4065
rect 19750 4015 19765 4035
rect 19785 4015 19800 4035
rect 19750 3985 19800 4015
rect 19750 3965 19765 3985
rect 19785 3965 19800 3985
rect 19750 3950 19800 3965
rect 20350 4435 20400 4450
rect 20350 4415 20365 4435
rect 20385 4415 20400 4435
rect 20350 4385 20400 4415
rect 20350 4365 20365 4385
rect 20385 4365 20400 4385
rect 20350 4335 20400 4365
rect 20350 4315 20365 4335
rect 20385 4315 20400 4335
rect 20350 4285 20400 4315
rect 20350 4265 20365 4285
rect 20385 4265 20400 4285
rect 20350 4235 20400 4265
rect 20350 4215 20365 4235
rect 20385 4215 20400 4235
rect 20350 4185 20400 4215
rect 20350 4165 20365 4185
rect 20385 4165 20400 4185
rect 20350 4135 20400 4165
rect 20350 4115 20365 4135
rect 20385 4115 20400 4135
rect 20350 4085 20400 4115
rect 20350 4065 20365 4085
rect 20385 4065 20400 4085
rect 20350 4035 20400 4065
rect 20350 4015 20365 4035
rect 20385 4015 20400 4035
rect 20350 3985 20400 4015
rect 20350 3965 20365 3985
rect 20385 3965 20400 3985
rect 20350 3950 20400 3965
rect -650 3885 20400 3900
rect -650 3865 -635 3885
rect -615 3865 -585 3885
rect -565 3865 -535 3885
rect -515 3865 -485 3885
rect -465 3865 -435 3885
rect -415 3865 -385 3885
rect -365 3865 -335 3885
rect -315 3865 -285 3885
rect -265 3865 -235 3885
rect -215 3865 -185 3885
rect -165 3865 -135 3885
rect -115 3865 -85 3885
rect -65 3865 -35 3885
rect -15 3865 15 3885
rect 35 3865 65 3885
rect 85 3865 115 3885
rect 135 3865 165 3885
rect 185 3865 215 3885
rect 235 3865 265 3885
rect 285 3865 315 3885
rect 335 3865 365 3885
rect 385 3865 415 3885
rect 435 3865 465 3885
rect 485 3865 515 3885
rect 535 3865 565 3885
rect 585 3865 615 3885
rect 635 3865 665 3885
rect 685 3865 715 3885
rect 735 3865 765 3885
rect 785 3865 815 3885
rect 835 3865 865 3885
rect 885 3865 915 3885
rect 935 3865 965 3885
rect 985 3865 1015 3885
rect 1035 3865 1065 3885
rect 1085 3865 1115 3885
rect 1135 3865 1165 3885
rect 1185 3865 1215 3885
rect 1235 3865 1265 3885
rect 1285 3865 1315 3885
rect 1335 3865 1365 3885
rect 1385 3865 1415 3885
rect 1435 3865 1465 3885
rect 1485 3865 1515 3885
rect 1535 3865 1565 3885
rect 1585 3865 1615 3885
rect 1635 3865 1665 3885
rect 1685 3865 1715 3885
rect 1735 3865 1765 3885
rect 1785 3865 1815 3885
rect 1835 3865 1865 3885
rect 1885 3865 1915 3885
rect 1935 3865 1965 3885
rect 1985 3865 2015 3885
rect 2035 3865 2065 3885
rect 2085 3865 2115 3885
rect 2135 3865 2165 3885
rect 2185 3865 2215 3885
rect 2235 3865 2265 3885
rect 2285 3865 2315 3885
rect 2335 3865 2365 3885
rect 2385 3865 2415 3885
rect 2435 3865 2465 3885
rect 2485 3865 2515 3885
rect 2535 3865 2565 3885
rect 2585 3865 2615 3885
rect 2635 3865 2665 3885
rect 2685 3865 2715 3885
rect 2735 3865 2765 3885
rect 2785 3865 2815 3885
rect 2835 3865 2865 3885
rect 2885 3865 2915 3885
rect 2935 3865 2965 3885
rect 2985 3865 3015 3885
rect 3035 3865 3065 3885
rect 3085 3865 3115 3885
rect 3135 3865 3165 3885
rect 3185 3865 3215 3885
rect 3235 3865 3265 3885
rect 3285 3865 3315 3885
rect 3335 3865 3365 3885
rect 3385 3865 3415 3885
rect 3435 3865 3465 3885
rect 3485 3865 3515 3885
rect 3535 3865 3565 3885
rect 3585 3865 3615 3885
rect 3635 3865 3665 3885
rect 3685 3865 3715 3885
rect 3735 3865 3765 3885
rect 3785 3865 3815 3885
rect 3835 3865 3865 3885
rect 3885 3865 3915 3885
rect 3935 3865 3965 3885
rect 3985 3865 4015 3885
rect 4035 3865 4065 3885
rect 4085 3865 4115 3885
rect 4135 3865 4165 3885
rect 4185 3865 4215 3885
rect 4235 3865 4265 3885
rect 4285 3865 4315 3885
rect 4335 3865 4365 3885
rect 4385 3865 4415 3885
rect 4435 3865 4465 3885
rect 4485 3865 4515 3885
rect 4535 3865 4565 3885
rect 4585 3865 4615 3885
rect 4635 3865 4665 3885
rect 4685 3865 4715 3885
rect 4735 3865 4765 3885
rect 4785 3865 4815 3885
rect 4835 3865 4865 3885
rect 4885 3865 4915 3885
rect 4935 3865 4965 3885
rect 4985 3865 5015 3885
rect 5035 3865 5065 3885
rect 5085 3865 5115 3885
rect 5135 3865 5165 3885
rect 5185 3865 5215 3885
rect 5235 3865 5265 3885
rect 5285 3865 5315 3885
rect 5335 3865 5365 3885
rect 5385 3865 5415 3885
rect 5435 3865 5465 3885
rect 5485 3865 5515 3885
rect 5535 3865 5565 3885
rect 5585 3865 5615 3885
rect 5635 3865 5665 3885
rect 5685 3865 5715 3885
rect 5735 3865 5765 3885
rect 5785 3865 5815 3885
rect 5835 3865 5865 3885
rect 5885 3865 5915 3885
rect 5935 3865 5965 3885
rect 5985 3865 6015 3885
rect 6035 3865 6065 3885
rect 6085 3865 6115 3885
rect 6135 3865 6165 3885
rect 6185 3865 6215 3885
rect 6235 3865 6265 3885
rect 6285 3865 6315 3885
rect 6335 3865 6365 3885
rect 6385 3865 6415 3885
rect 6435 3865 6465 3885
rect 6485 3865 6515 3885
rect 6535 3865 6565 3885
rect 6585 3865 6615 3885
rect 6635 3865 6665 3885
rect 6685 3865 6715 3885
rect 6735 3865 6765 3885
rect 6785 3865 6815 3885
rect 6835 3865 6865 3885
rect 6885 3865 6915 3885
rect 6935 3865 6965 3885
rect 6985 3865 7015 3885
rect 7035 3865 7065 3885
rect 7085 3865 7115 3885
rect 7135 3865 7165 3885
rect 7185 3865 7215 3885
rect 7235 3865 7265 3885
rect 7285 3865 7315 3885
rect 7335 3865 7365 3885
rect 7385 3865 7415 3885
rect 7435 3865 7465 3885
rect 7485 3865 7515 3885
rect 7535 3865 7565 3885
rect 7585 3865 7615 3885
rect 7635 3865 7665 3885
rect 7685 3865 7715 3885
rect 7735 3865 7765 3885
rect 7785 3865 7815 3885
rect 7835 3865 7865 3885
rect 7885 3865 7915 3885
rect 7935 3865 7965 3885
rect 7985 3865 8015 3885
rect 8035 3865 8065 3885
rect 8085 3865 8115 3885
rect 8135 3865 8165 3885
rect 8185 3865 8215 3885
rect 8235 3865 8265 3885
rect 8285 3865 8315 3885
rect 8335 3865 8365 3885
rect 8385 3865 8415 3885
rect 8435 3865 8465 3885
rect 8485 3865 8515 3885
rect 8535 3865 8565 3885
rect 8585 3865 8615 3885
rect 8635 3865 8665 3885
rect 8685 3865 8715 3885
rect 8735 3865 8765 3885
rect 8785 3865 8815 3885
rect 8835 3865 8865 3885
rect 8885 3865 8915 3885
rect 8935 3865 8965 3885
rect 8985 3865 9015 3885
rect 9035 3865 9065 3885
rect 9085 3865 9115 3885
rect 9135 3865 9165 3885
rect 9185 3865 9215 3885
rect 9235 3865 9265 3885
rect 9285 3865 9315 3885
rect 9335 3865 9365 3885
rect 9385 3865 9415 3885
rect 9435 3865 9465 3885
rect 9485 3865 9515 3885
rect 9535 3865 9565 3885
rect 9585 3865 9615 3885
rect 9635 3865 9665 3885
rect 9685 3865 9715 3885
rect 9735 3865 9765 3885
rect 9785 3865 9815 3885
rect 9835 3865 9865 3885
rect 9885 3865 9915 3885
rect 9935 3865 9965 3885
rect 9985 3865 10015 3885
rect 10035 3865 10065 3885
rect 10085 3865 10115 3885
rect 10135 3865 10165 3885
rect 10185 3865 10215 3885
rect 10235 3865 10265 3885
rect 10285 3865 10315 3885
rect 10335 3865 10365 3885
rect 10385 3865 10415 3885
rect 10435 3865 10465 3885
rect 10485 3865 10515 3885
rect 10535 3865 10565 3885
rect 10585 3865 10615 3885
rect 10635 3865 10665 3885
rect 10685 3865 10715 3885
rect 10735 3865 10765 3885
rect 10785 3865 10815 3885
rect 10835 3865 10865 3885
rect 10885 3865 10915 3885
rect 10935 3865 10965 3885
rect 10985 3865 11015 3885
rect 11035 3865 11065 3885
rect 11085 3865 11115 3885
rect 11135 3865 11165 3885
rect 11185 3865 11215 3885
rect 11235 3865 11265 3885
rect 11285 3865 11315 3885
rect 11335 3865 11365 3885
rect 11385 3865 11415 3885
rect 11435 3865 11465 3885
rect 11485 3865 11515 3885
rect 11535 3865 11565 3885
rect 11585 3865 11615 3885
rect 11635 3865 11665 3885
rect 11685 3865 11715 3885
rect 11735 3865 11765 3885
rect 11785 3865 11815 3885
rect 11835 3865 11865 3885
rect 11885 3865 11915 3885
rect 11935 3865 11965 3885
rect 11985 3865 12015 3885
rect 12035 3865 12065 3885
rect 12085 3865 12115 3885
rect 12135 3865 12165 3885
rect 12185 3865 12215 3885
rect 12235 3865 12265 3885
rect 12285 3865 12315 3885
rect 12335 3865 12365 3885
rect 12385 3865 12415 3885
rect 12435 3865 12465 3885
rect 12485 3865 12515 3885
rect 12535 3865 12565 3885
rect 12585 3865 12615 3885
rect 12635 3865 12665 3885
rect 12685 3865 12715 3885
rect 12735 3865 12765 3885
rect 12785 3865 12815 3885
rect 12835 3865 12865 3885
rect 12885 3865 12915 3885
rect 12935 3865 12965 3885
rect 12985 3865 13015 3885
rect 13035 3865 13065 3885
rect 13085 3865 13115 3885
rect 13135 3865 13165 3885
rect 13185 3865 13215 3885
rect 13235 3865 13265 3885
rect 13285 3865 13315 3885
rect 13335 3865 13365 3885
rect 13385 3865 13415 3885
rect 13435 3865 13465 3885
rect 13485 3865 13515 3885
rect 13535 3865 13565 3885
rect 13585 3865 13615 3885
rect 13635 3865 13665 3885
rect 13685 3865 13715 3885
rect 13735 3865 13765 3885
rect 13785 3865 13815 3885
rect 13835 3865 13865 3885
rect 13885 3865 13915 3885
rect 13935 3865 13965 3885
rect 13985 3865 14015 3885
rect 14035 3865 14065 3885
rect 14085 3865 14115 3885
rect 14135 3865 14165 3885
rect 14185 3865 14215 3885
rect 14235 3865 14265 3885
rect 14285 3865 14315 3885
rect 14335 3865 14365 3885
rect 14385 3865 14415 3885
rect 14435 3865 14465 3885
rect 14485 3865 14515 3885
rect 14535 3865 14565 3885
rect 14585 3865 14615 3885
rect 14635 3865 14665 3885
rect 14685 3865 14715 3885
rect 14735 3865 14765 3885
rect 14785 3865 14815 3885
rect 14835 3865 14865 3885
rect 14885 3865 14915 3885
rect 14935 3865 14965 3885
rect 14985 3865 15015 3885
rect 15035 3865 15065 3885
rect 15085 3865 15115 3885
rect 15135 3865 15165 3885
rect 15185 3865 15215 3885
rect 15235 3865 15265 3885
rect 15285 3865 15315 3885
rect 15335 3865 15365 3885
rect 15385 3865 15415 3885
rect 15435 3865 15465 3885
rect 15485 3865 15515 3885
rect 15535 3865 15565 3885
rect 15585 3865 15615 3885
rect 15635 3865 15665 3885
rect 15685 3865 15715 3885
rect 15735 3865 15765 3885
rect 15785 3865 15815 3885
rect 15835 3865 15865 3885
rect 15885 3865 15915 3885
rect 15935 3865 15965 3885
rect 15985 3865 16015 3885
rect 16035 3865 16065 3885
rect 16085 3865 16115 3885
rect 16135 3865 16165 3885
rect 16185 3865 16215 3885
rect 16235 3865 16265 3885
rect 16285 3865 16315 3885
rect 16335 3865 16365 3885
rect 16385 3865 16415 3885
rect 16435 3865 16465 3885
rect 16485 3865 16515 3885
rect 16535 3865 16565 3885
rect 16585 3865 16615 3885
rect 16635 3865 16665 3885
rect 16685 3865 16715 3885
rect 16735 3865 16765 3885
rect 16785 3865 16815 3885
rect 16835 3865 16865 3885
rect 16885 3865 16915 3885
rect 16935 3865 16965 3885
rect 16985 3865 17015 3885
rect 17035 3865 17065 3885
rect 17085 3865 17115 3885
rect 17135 3865 17165 3885
rect 17185 3865 17215 3885
rect 17235 3865 17265 3885
rect 17285 3865 17315 3885
rect 17335 3865 17365 3885
rect 17385 3865 17415 3885
rect 17435 3865 17465 3885
rect 17485 3865 17515 3885
rect 17535 3865 17565 3885
rect 17585 3865 17615 3885
rect 17635 3865 17665 3885
rect 17685 3865 17715 3885
rect 17735 3865 17765 3885
rect 17785 3865 17815 3885
rect 17835 3865 17865 3885
rect 17885 3865 17915 3885
rect 17935 3865 17965 3885
rect 17985 3865 18015 3885
rect 18035 3865 18065 3885
rect 18085 3865 18115 3885
rect 18135 3865 18165 3885
rect 18185 3865 18215 3885
rect 18235 3865 18265 3885
rect 18285 3865 18315 3885
rect 18335 3865 18365 3885
rect 18385 3865 18415 3885
rect 18435 3865 18465 3885
rect 18485 3865 18515 3885
rect 18535 3865 18565 3885
rect 18585 3865 18615 3885
rect 18635 3865 18665 3885
rect 18685 3865 18715 3885
rect 18735 3865 18765 3885
rect 18785 3865 18815 3885
rect 18835 3865 18865 3885
rect 18885 3865 18915 3885
rect 18935 3865 18965 3885
rect 18985 3865 19015 3885
rect 19035 3865 19065 3885
rect 19085 3865 19115 3885
rect 19135 3865 19165 3885
rect 19185 3865 19215 3885
rect 19235 3865 19265 3885
rect 19285 3865 19315 3885
rect 19335 3865 19365 3885
rect 19385 3865 19415 3885
rect 19435 3865 19465 3885
rect 19485 3865 19515 3885
rect 19535 3865 19565 3885
rect 19585 3865 19615 3885
rect 19635 3865 19665 3885
rect 19685 3865 19715 3885
rect 19735 3865 19765 3885
rect 19785 3865 19815 3885
rect 19835 3865 19865 3885
rect 19885 3865 19915 3885
rect 19935 3865 19965 3885
rect 19985 3865 20015 3885
rect 20035 3865 20065 3885
rect 20085 3865 20115 3885
rect 20135 3865 20165 3885
rect 20185 3865 20215 3885
rect 20235 3865 20265 3885
rect 20285 3865 20315 3885
rect 20335 3865 20365 3885
rect 20385 3865 20400 3885
rect -650 3850 20400 3865
rect -650 3785 -600 3800
rect -650 3765 -635 3785
rect -615 3765 -600 3785
rect -650 3735 -600 3765
rect -650 3715 -635 3735
rect -615 3715 -600 3735
rect -650 3685 -600 3715
rect -650 3665 -635 3685
rect -615 3665 -600 3685
rect -650 3635 -600 3665
rect -650 3615 -635 3635
rect -615 3615 -600 3635
rect -650 3585 -600 3615
rect -650 3565 -635 3585
rect -615 3565 -600 3585
rect -650 3535 -600 3565
rect -650 3515 -635 3535
rect -615 3515 -600 3535
rect -650 3485 -600 3515
rect -650 3465 -635 3485
rect -615 3465 -600 3485
rect -650 3435 -600 3465
rect -650 3415 -635 3435
rect -615 3415 -600 3435
rect -650 3385 -600 3415
rect -650 3365 -635 3385
rect -615 3365 -600 3385
rect -650 3335 -600 3365
rect -650 3315 -635 3335
rect -615 3315 -600 3335
rect -650 3300 -600 3315
rect -500 3785 -450 3800
rect -500 3765 -485 3785
rect -465 3765 -450 3785
rect -500 3735 -450 3765
rect -500 3715 -485 3735
rect -465 3715 -450 3735
rect -500 3685 -450 3715
rect -500 3665 -485 3685
rect -465 3665 -450 3685
rect -500 3635 -450 3665
rect -500 3615 -485 3635
rect -465 3615 -450 3635
rect -500 3585 -450 3615
rect -500 3565 -485 3585
rect -465 3565 -450 3585
rect -500 3535 -450 3565
rect -500 3515 -485 3535
rect -465 3515 -450 3535
rect -500 3485 -450 3515
rect -500 3465 -485 3485
rect -465 3465 -450 3485
rect -500 3435 -450 3465
rect -500 3415 -485 3435
rect -465 3415 -450 3435
rect -500 3385 -450 3415
rect -500 3365 -485 3385
rect -465 3365 -450 3385
rect -500 3335 -450 3365
rect -500 3315 -485 3335
rect -465 3315 -450 3335
rect -500 3300 -450 3315
rect -350 3785 -300 3800
rect -350 3765 -335 3785
rect -315 3765 -300 3785
rect -350 3735 -300 3765
rect -350 3715 -335 3735
rect -315 3715 -300 3735
rect -350 3685 -300 3715
rect -350 3665 -335 3685
rect -315 3665 -300 3685
rect -350 3635 -300 3665
rect -350 3615 -335 3635
rect -315 3615 -300 3635
rect -350 3585 -300 3615
rect -350 3565 -335 3585
rect -315 3565 -300 3585
rect -350 3535 -300 3565
rect -350 3515 -335 3535
rect -315 3515 -300 3535
rect -350 3485 -300 3515
rect -350 3465 -335 3485
rect -315 3465 -300 3485
rect -350 3435 -300 3465
rect -350 3415 -335 3435
rect -315 3415 -300 3435
rect -350 3385 -300 3415
rect -350 3365 -335 3385
rect -315 3365 -300 3385
rect -350 3335 -300 3365
rect -350 3315 -335 3335
rect -315 3315 -300 3335
rect -350 3300 -300 3315
rect -200 3785 -150 3800
rect -200 3765 -185 3785
rect -165 3765 -150 3785
rect -200 3735 -150 3765
rect -200 3715 -185 3735
rect -165 3715 -150 3735
rect -200 3685 -150 3715
rect -200 3665 -185 3685
rect -165 3665 -150 3685
rect -200 3635 -150 3665
rect -200 3615 -185 3635
rect -165 3615 -150 3635
rect -200 3585 -150 3615
rect -200 3565 -185 3585
rect -165 3565 -150 3585
rect -200 3535 -150 3565
rect -200 3515 -185 3535
rect -165 3515 -150 3535
rect -200 3485 -150 3515
rect -200 3465 -185 3485
rect -165 3465 -150 3485
rect -200 3435 -150 3465
rect -200 3415 -185 3435
rect -165 3415 -150 3435
rect -200 3385 -150 3415
rect -200 3365 -185 3385
rect -165 3365 -150 3385
rect -200 3335 -150 3365
rect -200 3315 -185 3335
rect -165 3315 -150 3335
rect -200 3300 -150 3315
rect -50 3785 0 3800
rect -50 3765 -35 3785
rect -15 3765 0 3785
rect -50 3735 0 3765
rect -50 3715 -35 3735
rect -15 3715 0 3735
rect -50 3685 0 3715
rect -50 3665 -35 3685
rect -15 3665 0 3685
rect -50 3635 0 3665
rect -50 3615 -35 3635
rect -15 3615 0 3635
rect -50 3585 0 3615
rect -50 3565 -35 3585
rect -15 3565 0 3585
rect -50 3535 0 3565
rect -50 3515 -35 3535
rect -15 3515 0 3535
rect -50 3485 0 3515
rect -50 3465 -35 3485
rect -15 3465 0 3485
rect -50 3435 0 3465
rect -50 3415 -35 3435
rect -15 3415 0 3435
rect -50 3385 0 3415
rect -50 3365 -35 3385
rect -15 3365 0 3385
rect -50 3335 0 3365
rect -50 3315 -35 3335
rect -15 3315 0 3335
rect -50 3300 0 3315
rect 550 3785 600 3800
rect 550 3765 565 3785
rect 585 3765 600 3785
rect 550 3735 600 3765
rect 550 3715 565 3735
rect 585 3715 600 3735
rect 550 3685 600 3715
rect 550 3665 565 3685
rect 585 3665 600 3685
rect 550 3635 600 3665
rect 550 3615 565 3635
rect 585 3615 600 3635
rect 550 3585 600 3615
rect 550 3565 565 3585
rect 585 3565 600 3585
rect 550 3535 600 3565
rect 550 3515 565 3535
rect 585 3515 600 3535
rect 550 3485 600 3515
rect 550 3465 565 3485
rect 585 3465 600 3485
rect 550 3435 600 3465
rect 550 3415 565 3435
rect 585 3415 600 3435
rect 550 3385 600 3415
rect 550 3365 565 3385
rect 585 3365 600 3385
rect 550 3335 600 3365
rect 550 3315 565 3335
rect 585 3315 600 3335
rect 550 3300 600 3315
rect 700 3785 750 3800
rect 700 3765 715 3785
rect 735 3765 750 3785
rect 700 3735 750 3765
rect 700 3715 715 3735
rect 735 3715 750 3735
rect 700 3685 750 3715
rect 700 3665 715 3685
rect 735 3665 750 3685
rect 700 3635 750 3665
rect 700 3615 715 3635
rect 735 3615 750 3635
rect 700 3585 750 3615
rect 700 3565 715 3585
rect 735 3565 750 3585
rect 700 3535 750 3565
rect 700 3515 715 3535
rect 735 3515 750 3535
rect 700 3485 750 3515
rect 700 3465 715 3485
rect 735 3465 750 3485
rect 700 3435 750 3465
rect 700 3415 715 3435
rect 735 3415 750 3435
rect 700 3385 750 3415
rect 700 3365 715 3385
rect 735 3365 750 3385
rect 700 3335 750 3365
rect 700 3315 715 3335
rect 735 3315 750 3335
rect 700 3300 750 3315
rect 850 3785 900 3800
rect 850 3765 865 3785
rect 885 3765 900 3785
rect 850 3735 900 3765
rect 850 3715 865 3735
rect 885 3715 900 3735
rect 850 3685 900 3715
rect 850 3665 865 3685
rect 885 3665 900 3685
rect 850 3635 900 3665
rect 850 3615 865 3635
rect 885 3615 900 3635
rect 850 3585 900 3615
rect 850 3565 865 3585
rect 885 3565 900 3585
rect 850 3535 900 3565
rect 850 3515 865 3535
rect 885 3515 900 3535
rect 850 3485 900 3515
rect 850 3465 865 3485
rect 885 3465 900 3485
rect 850 3435 900 3465
rect 850 3415 865 3435
rect 885 3415 900 3435
rect 850 3385 900 3415
rect 850 3365 865 3385
rect 885 3365 900 3385
rect 850 3335 900 3365
rect 850 3315 865 3335
rect 885 3315 900 3335
rect 850 3300 900 3315
rect 1000 3785 1050 3800
rect 1000 3765 1015 3785
rect 1035 3765 1050 3785
rect 1000 3735 1050 3765
rect 1000 3715 1015 3735
rect 1035 3715 1050 3735
rect 1000 3685 1050 3715
rect 1000 3665 1015 3685
rect 1035 3665 1050 3685
rect 1000 3635 1050 3665
rect 1000 3615 1015 3635
rect 1035 3615 1050 3635
rect 1000 3585 1050 3615
rect 1000 3565 1015 3585
rect 1035 3565 1050 3585
rect 1000 3535 1050 3565
rect 1000 3515 1015 3535
rect 1035 3515 1050 3535
rect 1000 3485 1050 3515
rect 1000 3465 1015 3485
rect 1035 3465 1050 3485
rect 1000 3435 1050 3465
rect 1000 3415 1015 3435
rect 1035 3415 1050 3435
rect 1000 3385 1050 3415
rect 1000 3365 1015 3385
rect 1035 3365 1050 3385
rect 1000 3335 1050 3365
rect 1000 3315 1015 3335
rect 1035 3315 1050 3335
rect 1000 3300 1050 3315
rect 1150 3785 1200 3800
rect 1150 3765 1165 3785
rect 1185 3765 1200 3785
rect 1150 3735 1200 3765
rect 1150 3715 1165 3735
rect 1185 3715 1200 3735
rect 1150 3685 1200 3715
rect 1150 3665 1165 3685
rect 1185 3665 1200 3685
rect 1150 3635 1200 3665
rect 1150 3615 1165 3635
rect 1185 3615 1200 3635
rect 1150 3585 1200 3615
rect 1150 3565 1165 3585
rect 1185 3565 1200 3585
rect 1150 3535 1200 3565
rect 1150 3515 1165 3535
rect 1185 3515 1200 3535
rect 1150 3485 1200 3515
rect 1150 3465 1165 3485
rect 1185 3465 1200 3485
rect 1150 3435 1200 3465
rect 1150 3415 1165 3435
rect 1185 3415 1200 3435
rect 1150 3385 1200 3415
rect 1150 3365 1165 3385
rect 1185 3365 1200 3385
rect 1150 3335 1200 3365
rect 1150 3315 1165 3335
rect 1185 3315 1200 3335
rect 1150 3300 1200 3315
rect 1300 3785 1350 3800
rect 1300 3765 1315 3785
rect 1335 3765 1350 3785
rect 1300 3735 1350 3765
rect 1300 3715 1315 3735
rect 1335 3715 1350 3735
rect 1300 3685 1350 3715
rect 1300 3665 1315 3685
rect 1335 3665 1350 3685
rect 1300 3635 1350 3665
rect 1300 3615 1315 3635
rect 1335 3615 1350 3635
rect 1300 3585 1350 3615
rect 1300 3565 1315 3585
rect 1335 3565 1350 3585
rect 1300 3535 1350 3565
rect 1300 3515 1315 3535
rect 1335 3515 1350 3535
rect 1300 3485 1350 3515
rect 1300 3465 1315 3485
rect 1335 3465 1350 3485
rect 1300 3435 1350 3465
rect 1300 3415 1315 3435
rect 1335 3415 1350 3435
rect 1300 3385 1350 3415
rect 1300 3365 1315 3385
rect 1335 3365 1350 3385
rect 1300 3335 1350 3365
rect 1300 3315 1315 3335
rect 1335 3315 1350 3335
rect 1300 3300 1350 3315
rect 1450 3785 1500 3800
rect 1450 3765 1465 3785
rect 1485 3765 1500 3785
rect 1450 3735 1500 3765
rect 1450 3715 1465 3735
rect 1485 3715 1500 3735
rect 1450 3685 1500 3715
rect 1450 3665 1465 3685
rect 1485 3665 1500 3685
rect 1450 3635 1500 3665
rect 1450 3615 1465 3635
rect 1485 3615 1500 3635
rect 1450 3585 1500 3615
rect 1450 3565 1465 3585
rect 1485 3565 1500 3585
rect 1450 3535 1500 3565
rect 1450 3515 1465 3535
rect 1485 3515 1500 3535
rect 1450 3485 1500 3515
rect 1450 3465 1465 3485
rect 1485 3465 1500 3485
rect 1450 3435 1500 3465
rect 1450 3415 1465 3435
rect 1485 3415 1500 3435
rect 1450 3385 1500 3415
rect 1450 3365 1465 3385
rect 1485 3365 1500 3385
rect 1450 3335 1500 3365
rect 1450 3315 1465 3335
rect 1485 3315 1500 3335
rect 1450 3300 1500 3315
rect 1600 3785 1650 3800
rect 1600 3765 1615 3785
rect 1635 3765 1650 3785
rect 1600 3735 1650 3765
rect 1600 3715 1615 3735
rect 1635 3715 1650 3735
rect 1600 3685 1650 3715
rect 1600 3665 1615 3685
rect 1635 3665 1650 3685
rect 1600 3635 1650 3665
rect 1600 3615 1615 3635
rect 1635 3615 1650 3635
rect 1600 3585 1650 3615
rect 1600 3565 1615 3585
rect 1635 3565 1650 3585
rect 1600 3535 1650 3565
rect 1600 3515 1615 3535
rect 1635 3515 1650 3535
rect 1600 3485 1650 3515
rect 1600 3465 1615 3485
rect 1635 3465 1650 3485
rect 1600 3435 1650 3465
rect 1600 3415 1615 3435
rect 1635 3415 1650 3435
rect 1600 3385 1650 3415
rect 1600 3365 1615 3385
rect 1635 3365 1650 3385
rect 1600 3335 1650 3365
rect 1600 3315 1615 3335
rect 1635 3315 1650 3335
rect 1600 3300 1650 3315
rect 1750 3785 1800 3800
rect 1750 3765 1765 3785
rect 1785 3765 1800 3785
rect 1750 3735 1800 3765
rect 1750 3715 1765 3735
rect 1785 3715 1800 3735
rect 1750 3685 1800 3715
rect 1750 3665 1765 3685
rect 1785 3665 1800 3685
rect 1750 3635 1800 3665
rect 1750 3615 1765 3635
rect 1785 3615 1800 3635
rect 1750 3585 1800 3615
rect 1750 3565 1765 3585
rect 1785 3565 1800 3585
rect 1750 3535 1800 3565
rect 1750 3515 1765 3535
rect 1785 3515 1800 3535
rect 1750 3485 1800 3515
rect 1750 3465 1765 3485
rect 1785 3465 1800 3485
rect 1750 3435 1800 3465
rect 1750 3415 1765 3435
rect 1785 3415 1800 3435
rect 1750 3385 1800 3415
rect 1750 3365 1765 3385
rect 1785 3365 1800 3385
rect 1750 3335 1800 3365
rect 1750 3315 1765 3335
rect 1785 3315 1800 3335
rect 1750 3300 1800 3315
rect 1900 3785 1950 3800
rect 1900 3765 1915 3785
rect 1935 3765 1950 3785
rect 1900 3735 1950 3765
rect 1900 3715 1915 3735
rect 1935 3715 1950 3735
rect 1900 3685 1950 3715
rect 1900 3665 1915 3685
rect 1935 3665 1950 3685
rect 1900 3635 1950 3665
rect 1900 3615 1915 3635
rect 1935 3615 1950 3635
rect 1900 3585 1950 3615
rect 1900 3565 1915 3585
rect 1935 3565 1950 3585
rect 1900 3535 1950 3565
rect 1900 3515 1915 3535
rect 1935 3515 1950 3535
rect 1900 3485 1950 3515
rect 1900 3465 1915 3485
rect 1935 3465 1950 3485
rect 1900 3435 1950 3465
rect 1900 3415 1915 3435
rect 1935 3415 1950 3435
rect 1900 3385 1950 3415
rect 1900 3365 1915 3385
rect 1935 3365 1950 3385
rect 1900 3335 1950 3365
rect 1900 3315 1915 3335
rect 1935 3315 1950 3335
rect 1900 3300 1950 3315
rect 2050 3785 2100 3800
rect 2050 3765 2065 3785
rect 2085 3765 2100 3785
rect 2050 3735 2100 3765
rect 2050 3715 2065 3735
rect 2085 3715 2100 3735
rect 2050 3685 2100 3715
rect 2050 3665 2065 3685
rect 2085 3665 2100 3685
rect 2050 3635 2100 3665
rect 2050 3615 2065 3635
rect 2085 3615 2100 3635
rect 2050 3585 2100 3615
rect 2050 3565 2065 3585
rect 2085 3565 2100 3585
rect 2050 3535 2100 3565
rect 2050 3515 2065 3535
rect 2085 3515 2100 3535
rect 2050 3485 2100 3515
rect 2050 3465 2065 3485
rect 2085 3465 2100 3485
rect 2050 3435 2100 3465
rect 2050 3415 2065 3435
rect 2085 3415 2100 3435
rect 2050 3385 2100 3415
rect 2050 3365 2065 3385
rect 2085 3365 2100 3385
rect 2050 3335 2100 3365
rect 2050 3315 2065 3335
rect 2085 3315 2100 3335
rect 2050 3300 2100 3315
rect 2200 3785 2250 3800
rect 2200 3765 2215 3785
rect 2235 3765 2250 3785
rect 2200 3735 2250 3765
rect 2200 3715 2215 3735
rect 2235 3715 2250 3735
rect 2200 3685 2250 3715
rect 2200 3665 2215 3685
rect 2235 3665 2250 3685
rect 2200 3635 2250 3665
rect 2200 3615 2215 3635
rect 2235 3615 2250 3635
rect 2200 3585 2250 3615
rect 2200 3565 2215 3585
rect 2235 3565 2250 3585
rect 2200 3535 2250 3565
rect 2200 3515 2215 3535
rect 2235 3515 2250 3535
rect 2200 3485 2250 3515
rect 2200 3465 2215 3485
rect 2235 3465 2250 3485
rect 2200 3435 2250 3465
rect 2200 3415 2215 3435
rect 2235 3415 2250 3435
rect 2200 3385 2250 3415
rect 2200 3365 2215 3385
rect 2235 3365 2250 3385
rect 2200 3335 2250 3365
rect 2200 3315 2215 3335
rect 2235 3315 2250 3335
rect 2200 3300 2250 3315
rect 2350 3785 2400 3800
rect 2350 3765 2365 3785
rect 2385 3765 2400 3785
rect 2350 3735 2400 3765
rect 2350 3715 2365 3735
rect 2385 3715 2400 3735
rect 2350 3685 2400 3715
rect 2350 3665 2365 3685
rect 2385 3665 2400 3685
rect 2350 3635 2400 3665
rect 2350 3615 2365 3635
rect 2385 3615 2400 3635
rect 2350 3585 2400 3615
rect 2350 3565 2365 3585
rect 2385 3565 2400 3585
rect 2350 3535 2400 3565
rect 2350 3515 2365 3535
rect 2385 3515 2400 3535
rect 2350 3485 2400 3515
rect 2350 3465 2365 3485
rect 2385 3465 2400 3485
rect 2350 3435 2400 3465
rect 2350 3415 2365 3435
rect 2385 3415 2400 3435
rect 2350 3385 2400 3415
rect 2350 3365 2365 3385
rect 2385 3365 2400 3385
rect 2350 3335 2400 3365
rect 2350 3315 2365 3335
rect 2385 3315 2400 3335
rect 2350 3300 2400 3315
rect 2500 3785 2550 3800
rect 2500 3765 2515 3785
rect 2535 3765 2550 3785
rect 2500 3735 2550 3765
rect 2500 3715 2515 3735
rect 2535 3715 2550 3735
rect 2500 3685 2550 3715
rect 2500 3665 2515 3685
rect 2535 3665 2550 3685
rect 2500 3635 2550 3665
rect 2500 3615 2515 3635
rect 2535 3615 2550 3635
rect 2500 3585 2550 3615
rect 2500 3565 2515 3585
rect 2535 3565 2550 3585
rect 2500 3535 2550 3565
rect 2500 3515 2515 3535
rect 2535 3515 2550 3535
rect 2500 3485 2550 3515
rect 2500 3465 2515 3485
rect 2535 3465 2550 3485
rect 2500 3435 2550 3465
rect 2500 3415 2515 3435
rect 2535 3415 2550 3435
rect 2500 3385 2550 3415
rect 2500 3365 2515 3385
rect 2535 3365 2550 3385
rect 2500 3335 2550 3365
rect 2500 3315 2515 3335
rect 2535 3315 2550 3335
rect 2500 3300 2550 3315
rect 2650 3785 2700 3800
rect 2650 3765 2665 3785
rect 2685 3765 2700 3785
rect 2650 3735 2700 3765
rect 2650 3715 2665 3735
rect 2685 3715 2700 3735
rect 2650 3685 2700 3715
rect 2650 3665 2665 3685
rect 2685 3665 2700 3685
rect 2650 3635 2700 3665
rect 2650 3615 2665 3635
rect 2685 3615 2700 3635
rect 2650 3585 2700 3615
rect 2650 3565 2665 3585
rect 2685 3565 2700 3585
rect 2650 3535 2700 3565
rect 2650 3515 2665 3535
rect 2685 3515 2700 3535
rect 2650 3485 2700 3515
rect 2650 3465 2665 3485
rect 2685 3465 2700 3485
rect 2650 3435 2700 3465
rect 2650 3415 2665 3435
rect 2685 3415 2700 3435
rect 2650 3385 2700 3415
rect 2650 3365 2665 3385
rect 2685 3365 2700 3385
rect 2650 3335 2700 3365
rect 2650 3315 2665 3335
rect 2685 3315 2700 3335
rect 2650 3300 2700 3315
rect 2800 3785 2850 3800
rect 2800 3765 2815 3785
rect 2835 3765 2850 3785
rect 2800 3735 2850 3765
rect 2800 3715 2815 3735
rect 2835 3715 2850 3735
rect 2800 3685 2850 3715
rect 2800 3665 2815 3685
rect 2835 3665 2850 3685
rect 2800 3635 2850 3665
rect 2800 3615 2815 3635
rect 2835 3615 2850 3635
rect 2800 3585 2850 3615
rect 2800 3565 2815 3585
rect 2835 3565 2850 3585
rect 2800 3535 2850 3565
rect 2800 3515 2815 3535
rect 2835 3515 2850 3535
rect 2800 3485 2850 3515
rect 2800 3465 2815 3485
rect 2835 3465 2850 3485
rect 2800 3435 2850 3465
rect 2800 3415 2815 3435
rect 2835 3415 2850 3435
rect 2800 3385 2850 3415
rect 2800 3365 2815 3385
rect 2835 3365 2850 3385
rect 2800 3335 2850 3365
rect 2800 3315 2815 3335
rect 2835 3315 2850 3335
rect 2800 3300 2850 3315
rect 2950 3785 3000 3800
rect 2950 3765 2965 3785
rect 2985 3765 3000 3785
rect 2950 3735 3000 3765
rect 2950 3715 2965 3735
rect 2985 3715 3000 3735
rect 2950 3685 3000 3715
rect 2950 3665 2965 3685
rect 2985 3665 3000 3685
rect 2950 3635 3000 3665
rect 2950 3615 2965 3635
rect 2985 3615 3000 3635
rect 2950 3585 3000 3615
rect 2950 3565 2965 3585
rect 2985 3565 3000 3585
rect 2950 3535 3000 3565
rect 2950 3515 2965 3535
rect 2985 3515 3000 3535
rect 2950 3485 3000 3515
rect 2950 3465 2965 3485
rect 2985 3465 3000 3485
rect 2950 3435 3000 3465
rect 2950 3415 2965 3435
rect 2985 3415 3000 3435
rect 2950 3385 3000 3415
rect 2950 3365 2965 3385
rect 2985 3365 3000 3385
rect 2950 3335 3000 3365
rect 2950 3315 2965 3335
rect 2985 3315 3000 3335
rect 2950 3300 3000 3315
rect 3100 3785 3150 3800
rect 3100 3765 3115 3785
rect 3135 3765 3150 3785
rect 3100 3735 3150 3765
rect 3100 3715 3115 3735
rect 3135 3715 3150 3735
rect 3100 3685 3150 3715
rect 3100 3665 3115 3685
rect 3135 3665 3150 3685
rect 3100 3635 3150 3665
rect 3100 3615 3115 3635
rect 3135 3615 3150 3635
rect 3100 3585 3150 3615
rect 3100 3565 3115 3585
rect 3135 3565 3150 3585
rect 3100 3535 3150 3565
rect 3100 3515 3115 3535
rect 3135 3515 3150 3535
rect 3100 3485 3150 3515
rect 3100 3465 3115 3485
rect 3135 3465 3150 3485
rect 3100 3435 3150 3465
rect 3100 3415 3115 3435
rect 3135 3415 3150 3435
rect 3100 3385 3150 3415
rect 3100 3365 3115 3385
rect 3135 3365 3150 3385
rect 3100 3335 3150 3365
rect 3100 3315 3115 3335
rect 3135 3315 3150 3335
rect 3100 3300 3150 3315
rect 3250 3785 3300 3800
rect 3250 3765 3265 3785
rect 3285 3765 3300 3785
rect 3250 3735 3300 3765
rect 3250 3715 3265 3735
rect 3285 3715 3300 3735
rect 3250 3685 3300 3715
rect 3250 3665 3265 3685
rect 3285 3665 3300 3685
rect 3250 3635 3300 3665
rect 3250 3615 3265 3635
rect 3285 3615 3300 3635
rect 3250 3585 3300 3615
rect 3250 3565 3265 3585
rect 3285 3565 3300 3585
rect 3250 3535 3300 3565
rect 3250 3515 3265 3535
rect 3285 3515 3300 3535
rect 3250 3485 3300 3515
rect 3250 3465 3265 3485
rect 3285 3465 3300 3485
rect 3250 3435 3300 3465
rect 3250 3415 3265 3435
rect 3285 3415 3300 3435
rect 3250 3385 3300 3415
rect 3250 3365 3265 3385
rect 3285 3365 3300 3385
rect 3250 3335 3300 3365
rect 3250 3315 3265 3335
rect 3285 3315 3300 3335
rect 3250 3300 3300 3315
rect 3400 3785 3450 3800
rect 3400 3765 3415 3785
rect 3435 3765 3450 3785
rect 3400 3735 3450 3765
rect 3400 3715 3415 3735
rect 3435 3715 3450 3735
rect 3400 3685 3450 3715
rect 3400 3665 3415 3685
rect 3435 3665 3450 3685
rect 3400 3635 3450 3665
rect 3400 3615 3415 3635
rect 3435 3615 3450 3635
rect 3400 3585 3450 3615
rect 3400 3565 3415 3585
rect 3435 3565 3450 3585
rect 3400 3535 3450 3565
rect 3400 3515 3415 3535
rect 3435 3515 3450 3535
rect 3400 3485 3450 3515
rect 3400 3465 3415 3485
rect 3435 3465 3450 3485
rect 3400 3435 3450 3465
rect 3400 3415 3415 3435
rect 3435 3415 3450 3435
rect 3400 3385 3450 3415
rect 3400 3365 3415 3385
rect 3435 3365 3450 3385
rect 3400 3335 3450 3365
rect 3400 3315 3415 3335
rect 3435 3315 3450 3335
rect 3400 3300 3450 3315
rect 3550 3785 3600 3800
rect 3550 3765 3565 3785
rect 3585 3765 3600 3785
rect 3550 3735 3600 3765
rect 3550 3715 3565 3735
rect 3585 3715 3600 3735
rect 3550 3685 3600 3715
rect 3550 3665 3565 3685
rect 3585 3665 3600 3685
rect 3550 3635 3600 3665
rect 3550 3615 3565 3635
rect 3585 3615 3600 3635
rect 3550 3585 3600 3615
rect 3550 3565 3565 3585
rect 3585 3565 3600 3585
rect 3550 3535 3600 3565
rect 3550 3515 3565 3535
rect 3585 3515 3600 3535
rect 3550 3485 3600 3515
rect 3550 3465 3565 3485
rect 3585 3465 3600 3485
rect 3550 3435 3600 3465
rect 3550 3415 3565 3435
rect 3585 3415 3600 3435
rect 3550 3385 3600 3415
rect 3550 3365 3565 3385
rect 3585 3365 3600 3385
rect 3550 3335 3600 3365
rect 3550 3315 3565 3335
rect 3585 3315 3600 3335
rect 3550 3300 3600 3315
rect 4150 3785 4200 3800
rect 4150 3765 4165 3785
rect 4185 3765 4200 3785
rect 4150 3735 4200 3765
rect 4150 3715 4165 3735
rect 4185 3715 4200 3735
rect 4150 3685 4200 3715
rect 4150 3665 4165 3685
rect 4185 3665 4200 3685
rect 4150 3635 4200 3665
rect 4150 3615 4165 3635
rect 4185 3615 4200 3635
rect 4150 3585 4200 3615
rect 4150 3565 4165 3585
rect 4185 3565 4200 3585
rect 4150 3535 4200 3565
rect 4150 3515 4165 3535
rect 4185 3515 4200 3535
rect 4150 3485 4200 3515
rect 4150 3465 4165 3485
rect 4185 3465 4200 3485
rect 4150 3435 4200 3465
rect 4150 3415 4165 3435
rect 4185 3415 4200 3435
rect 4150 3385 4200 3415
rect 4150 3365 4165 3385
rect 4185 3365 4200 3385
rect 4150 3335 4200 3365
rect 4150 3315 4165 3335
rect 4185 3315 4200 3335
rect 4150 3300 4200 3315
rect 4750 3785 4800 3800
rect 4750 3765 4765 3785
rect 4785 3765 4800 3785
rect 4750 3735 4800 3765
rect 4750 3715 4765 3735
rect 4785 3715 4800 3735
rect 4750 3685 4800 3715
rect 4750 3665 4765 3685
rect 4785 3665 4800 3685
rect 4750 3635 4800 3665
rect 4750 3615 4765 3635
rect 4785 3615 4800 3635
rect 4750 3585 4800 3615
rect 4750 3565 4765 3585
rect 4785 3565 4800 3585
rect 4750 3535 4800 3565
rect 4750 3515 4765 3535
rect 4785 3515 4800 3535
rect 4750 3485 4800 3515
rect 4750 3465 4765 3485
rect 4785 3465 4800 3485
rect 4750 3435 4800 3465
rect 4750 3415 4765 3435
rect 4785 3415 4800 3435
rect 4750 3385 4800 3415
rect 4750 3365 4765 3385
rect 4785 3365 4800 3385
rect 4750 3335 4800 3365
rect 4750 3315 4765 3335
rect 4785 3315 4800 3335
rect 4750 3300 4800 3315
rect 4900 3785 4950 3800
rect 4900 3765 4915 3785
rect 4935 3765 4950 3785
rect 4900 3735 4950 3765
rect 4900 3715 4915 3735
rect 4935 3715 4950 3735
rect 4900 3685 4950 3715
rect 4900 3665 4915 3685
rect 4935 3665 4950 3685
rect 4900 3635 4950 3665
rect 4900 3615 4915 3635
rect 4935 3615 4950 3635
rect 4900 3585 4950 3615
rect 4900 3565 4915 3585
rect 4935 3565 4950 3585
rect 4900 3535 4950 3565
rect 4900 3515 4915 3535
rect 4935 3515 4950 3535
rect 4900 3485 4950 3515
rect 4900 3465 4915 3485
rect 4935 3465 4950 3485
rect 4900 3435 4950 3465
rect 4900 3415 4915 3435
rect 4935 3415 4950 3435
rect 4900 3385 4950 3415
rect 4900 3365 4915 3385
rect 4935 3365 4950 3385
rect 4900 3335 4950 3365
rect 4900 3315 4915 3335
rect 4935 3315 4950 3335
rect 4900 3300 4950 3315
rect 5050 3785 5100 3800
rect 5050 3765 5065 3785
rect 5085 3765 5100 3785
rect 5050 3735 5100 3765
rect 5050 3715 5065 3735
rect 5085 3715 5100 3735
rect 5050 3685 5100 3715
rect 5050 3665 5065 3685
rect 5085 3665 5100 3685
rect 5050 3635 5100 3665
rect 5050 3615 5065 3635
rect 5085 3615 5100 3635
rect 5050 3585 5100 3615
rect 5050 3565 5065 3585
rect 5085 3565 5100 3585
rect 5050 3535 5100 3565
rect 5050 3515 5065 3535
rect 5085 3515 5100 3535
rect 5050 3485 5100 3515
rect 5050 3465 5065 3485
rect 5085 3465 5100 3485
rect 5050 3435 5100 3465
rect 5050 3415 5065 3435
rect 5085 3415 5100 3435
rect 5050 3385 5100 3415
rect 5050 3365 5065 3385
rect 5085 3365 5100 3385
rect 5050 3335 5100 3365
rect 5050 3315 5065 3335
rect 5085 3315 5100 3335
rect 5050 3300 5100 3315
rect 5200 3785 5250 3800
rect 5200 3765 5215 3785
rect 5235 3765 5250 3785
rect 5200 3735 5250 3765
rect 5200 3715 5215 3735
rect 5235 3715 5250 3735
rect 5200 3685 5250 3715
rect 5200 3665 5215 3685
rect 5235 3665 5250 3685
rect 5200 3635 5250 3665
rect 5200 3615 5215 3635
rect 5235 3615 5250 3635
rect 5200 3585 5250 3615
rect 5200 3565 5215 3585
rect 5235 3565 5250 3585
rect 5200 3535 5250 3565
rect 5200 3515 5215 3535
rect 5235 3515 5250 3535
rect 5200 3485 5250 3515
rect 5200 3465 5215 3485
rect 5235 3465 5250 3485
rect 5200 3435 5250 3465
rect 5200 3415 5215 3435
rect 5235 3415 5250 3435
rect 5200 3385 5250 3415
rect 5200 3365 5215 3385
rect 5235 3365 5250 3385
rect 5200 3335 5250 3365
rect 5200 3315 5215 3335
rect 5235 3315 5250 3335
rect 5200 3300 5250 3315
rect 5350 3785 5400 3800
rect 5350 3765 5365 3785
rect 5385 3765 5400 3785
rect 5350 3735 5400 3765
rect 5350 3715 5365 3735
rect 5385 3715 5400 3735
rect 5350 3685 5400 3715
rect 5350 3665 5365 3685
rect 5385 3665 5400 3685
rect 5350 3635 5400 3665
rect 5350 3615 5365 3635
rect 5385 3615 5400 3635
rect 5350 3585 5400 3615
rect 5350 3565 5365 3585
rect 5385 3565 5400 3585
rect 5350 3535 5400 3565
rect 5350 3515 5365 3535
rect 5385 3515 5400 3535
rect 5350 3485 5400 3515
rect 5350 3465 5365 3485
rect 5385 3465 5400 3485
rect 5350 3435 5400 3465
rect 5350 3415 5365 3435
rect 5385 3415 5400 3435
rect 5350 3385 5400 3415
rect 5350 3365 5365 3385
rect 5385 3365 5400 3385
rect 5350 3335 5400 3365
rect 5350 3315 5365 3335
rect 5385 3315 5400 3335
rect 5350 3300 5400 3315
rect 5500 3785 5550 3800
rect 5500 3765 5515 3785
rect 5535 3765 5550 3785
rect 5500 3735 5550 3765
rect 5500 3715 5515 3735
rect 5535 3715 5550 3735
rect 5500 3685 5550 3715
rect 5500 3665 5515 3685
rect 5535 3665 5550 3685
rect 5500 3635 5550 3665
rect 5500 3615 5515 3635
rect 5535 3615 5550 3635
rect 5500 3585 5550 3615
rect 5500 3565 5515 3585
rect 5535 3565 5550 3585
rect 5500 3535 5550 3565
rect 5500 3515 5515 3535
rect 5535 3515 5550 3535
rect 5500 3485 5550 3515
rect 5500 3465 5515 3485
rect 5535 3465 5550 3485
rect 5500 3435 5550 3465
rect 5500 3415 5515 3435
rect 5535 3415 5550 3435
rect 5500 3385 5550 3415
rect 5500 3365 5515 3385
rect 5535 3365 5550 3385
rect 5500 3335 5550 3365
rect 5500 3315 5515 3335
rect 5535 3315 5550 3335
rect 5500 3300 5550 3315
rect 5650 3785 5700 3800
rect 5650 3765 5665 3785
rect 5685 3765 5700 3785
rect 5650 3735 5700 3765
rect 5650 3715 5665 3735
rect 5685 3715 5700 3735
rect 5650 3685 5700 3715
rect 5650 3665 5665 3685
rect 5685 3665 5700 3685
rect 5650 3635 5700 3665
rect 5650 3615 5665 3635
rect 5685 3615 5700 3635
rect 5650 3585 5700 3615
rect 5650 3565 5665 3585
rect 5685 3565 5700 3585
rect 5650 3535 5700 3565
rect 5650 3515 5665 3535
rect 5685 3515 5700 3535
rect 5650 3485 5700 3515
rect 5650 3465 5665 3485
rect 5685 3465 5700 3485
rect 5650 3435 5700 3465
rect 5650 3415 5665 3435
rect 5685 3415 5700 3435
rect 5650 3385 5700 3415
rect 5650 3365 5665 3385
rect 5685 3365 5700 3385
rect 5650 3335 5700 3365
rect 5650 3315 5665 3335
rect 5685 3315 5700 3335
rect 5650 3300 5700 3315
rect 5800 3785 5850 3800
rect 5800 3765 5815 3785
rect 5835 3765 5850 3785
rect 5800 3735 5850 3765
rect 5800 3715 5815 3735
rect 5835 3715 5850 3735
rect 5800 3685 5850 3715
rect 5800 3665 5815 3685
rect 5835 3665 5850 3685
rect 5800 3635 5850 3665
rect 5800 3615 5815 3635
rect 5835 3615 5850 3635
rect 5800 3585 5850 3615
rect 5800 3565 5815 3585
rect 5835 3565 5850 3585
rect 5800 3535 5850 3565
rect 5800 3515 5815 3535
rect 5835 3515 5850 3535
rect 5800 3485 5850 3515
rect 5800 3465 5815 3485
rect 5835 3465 5850 3485
rect 5800 3435 5850 3465
rect 5800 3415 5815 3435
rect 5835 3415 5850 3435
rect 5800 3385 5850 3415
rect 5800 3365 5815 3385
rect 5835 3365 5850 3385
rect 5800 3335 5850 3365
rect 5800 3315 5815 3335
rect 5835 3315 5850 3335
rect 5800 3300 5850 3315
rect 5950 3785 6000 3800
rect 5950 3765 5965 3785
rect 5985 3765 6000 3785
rect 5950 3735 6000 3765
rect 5950 3715 5965 3735
rect 5985 3715 6000 3735
rect 5950 3685 6000 3715
rect 5950 3665 5965 3685
rect 5985 3665 6000 3685
rect 5950 3635 6000 3665
rect 5950 3615 5965 3635
rect 5985 3615 6000 3635
rect 5950 3585 6000 3615
rect 5950 3565 5965 3585
rect 5985 3565 6000 3585
rect 5950 3535 6000 3565
rect 5950 3515 5965 3535
rect 5985 3515 6000 3535
rect 5950 3485 6000 3515
rect 5950 3465 5965 3485
rect 5985 3465 6000 3485
rect 5950 3435 6000 3465
rect 5950 3415 5965 3435
rect 5985 3415 6000 3435
rect 5950 3385 6000 3415
rect 5950 3365 5965 3385
rect 5985 3365 6000 3385
rect 5950 3335 6000 3365
rect 5950 3315 5965 3335
rect 5985 3315 6000 3335
rect 5950 3300 6000 3315
rect 6100 3785 6150 3800
rect 6100 3765 6115 3785
rect 6135 3765 6150 3785
rect 6100 3735 6150 3765
rect 6100 3715 6115 3735
rect 6135 3715 6150 3735
rect 6100 3685 6150 3715
rect 6100 3665 6115 3685
rect 6135 3665 6150 3685
rect 6100 3635 6150 3665
rect 6100 3615 6115 3635
rect 6135 3615 6150 3635
rect 6100 3585 6150 3615
rect 6100 3565 6115 3585
rect 6135 3565 6150 3585
rect 6100 3535 6150 3565
rect 6100 3515 6115 3535
rect 6135 3515 6150 3535
rect 6100 3485 6150 3515
rect 6100 3465 6115 3485
rect 6135 3465 6150 3485
rect 6100 3435 6150 3465
rect 6100 3415 6115 3435
rect 6135 3415 6150 3435
rect 6100 3385 6150 3415
rect 6100 3365 6115 3385
rect 6135 3365 6150 3385
rect 6100 3335 6150 3365
rect 6100 3315 6115 3335
rect 6135 3315 6150 3335
rect 6100 3300 6150 3315
rect 6250 3785 6300 3800
rect 6250 3765 6265 3785
rect 6285 3765 6300 3785
rect 6250 3735 6300 3765
rect 6250 3715 6265 3735
rect 6285 3715 6300 3735
rect 6250 3685 6300 3715
rect 6250 3665 6265 3685
rect 6285 3665 6300 3685
rect 6250 3635 6300 3665
rect 6250 3615 6265 3635
rect 6285 3615 6300 3635
rect 6250 3585 6300 3615
rect 6250 3565 6265 3585
rect 6285 3565 6300 3585
rect 6250 3535 6300 3565
rect 6250 3515 6265 3535
rect 6285 3515 6300 3535
rect 6250 3485 6300 3515
rect 6250 3465 6265 3485
rect 6285 3465 6300 3485
rect 6250 3435 6300 3465
rect 6250 3415 6265 3435
rect 6285 3415 6300 3435
rect 6250 3385 6300 3415
rect 6250 3365 6265 3385
rect 6285 3365 6300 3385
rect 6250 3335 6300 3365
rect 6250 3315 6265 3335
rect 6285 3315 6300 3335
rect 6250 3300 6300 3315
rect 6400 3785 6450 3800
rect 6400 3765 6415 3785
rect 6435 3765 6450 3785
rect 6400 3735 6450 3765
rect 6400 3715 6415 3735
rect 6435 3715 6450 3735
rect 6400 3685 6450 3715
rect 6400 3665 6415 3685
rect 6435 3665 6450 3685
rect 6400 3635 6450 3665
rect 6400 3615 6415 3635
rect 6435 3615 6450 3635
rect 6400 3585 6450 3615
rect 6400 3565 6415 3585
rect 6435 3565 6450 3585
rect 6400 3535 6450 3565
rect 6400 3515 6415 3535
rect 6435 3515 6450 3535
rect 6400 3485 6450 3515
rect 6400 3465 6415 3485
rect 6435 3465 6450 3485
rect 6400 3435 6450 3465
rect 6400 3415 6415 3435
rect 6435 3415 6450 3435
rect 6400 3385 6450 3415
rect 6400 3365 6415 3385
rect 6435 3365 6450 3385
rect 6400 3335 6450 3365
rect 6400 3315 6415 3335
rect 6435 3315 6450 3335
rect 6400 3300 6450 3315
rect 6550 3785 6600 3800
rect 6550 3765 6565 3785
rect 6585 3765 6600 3785
rect 6550 3735 6600 3765
rect 6550 3715 6565 3735
rect 6585 3715 6600 3735
rect 6550 3685 6600 3715
rect 6550 3665 6565 3685
rect 6585 3665 6600 3685
rect 6550 3635 6600 3665
rect 6550 3615 6565 3635
rect 6585 3615 6600 3635
rect 6550 3585 6600 3615
rect 6550 3565 6565 3585
rect 6585 3565 6600 3585
rect 6550 3535 6600 3565
rect 6550 3515 6565 3535
rect 6585 3515 6600 3535
rect 6550 3485 6600 3515
rect 6550 3465 6565 3485
rect 6585 3465 6600 3485
rect 6550 3435 6600 3465
rect 6550 3415 6565 3435
rect 6585 3415 6600 3435
rect 6550 3385 6600 3415
rect 6550 3365 6565 3385
rect 6585 3365 6600 3385
rect 6550 3335 6600 3365
rect 6550 3315 6565 3335
rect 6585 3315 6600 3335
rect 6550 3300 6600 3315
rect 6700 3785 6750 3800
rect 6700 3765 6715 3785
rect 6735 3765 6750 3785
rect 6700 3735 6750 3765
rect 6700 3715 6715 3735
rect 6735 3715 6750 3735
rect 6700 3685 6750 3715
rect 6700 3665 6715 3685
rect 6735 3665 6750 3685
rect 6700 3635 6750 3665
rect 6700 3615 6715 3635
rect 6735 3615 6750 3635
rect 6700 3585 6750 3615
rect 6700 3565 6715 3585
rect 6735 3565 6750 3585
rect 6700 3535 6750 3565
rect 6700 3515 6715 3535
rect 6735 3515 6750 3535
rect 6700 3485 6750 3515
rect 6700 3465 6715 3485
rect 6735 3465 6750 3485
rect 6700 3435 6750 3465
rect 6700 3415 6715 3435
rect 6735 3415 6750 3435
rect 6700 3385 6750 3415
rect 6700 3365 6715 3385
rect 6735 3365 6750 3385
rect 6700 3335 6750 3365
rect 6700 3315 6715 3335
rect 6735 3315 6750 3335
rect 6700 3300 6750 3315
rect 6850 3785 6900 3800
rect 6850 3765 6865 3785
rect 6885 3765 6900 3785
rect 6850 3735 6900 3765
rect 6850 3715 6865 3735
rect 6885 3715 6900 3735
rect 6850 3685 6900 3715
rect 6850 3665 6865 3685
rect 6885 3665 6900 3685
rect 6850 3635 6900 3665
rect 6850 3615 6865 3635
rect 6885 3615 6900 3635
rect 6850 3585 6900 3615
rect 6850 3565 6865 3585
rect 6885 3565 6900 3585
rect 6850 3535 6900 3565
rect 6850 3515 6865 3535
rect 6885 3515 6900 3535
rect 6850 3485 6900 3515
rect 6850 3465 6865 3485
rect 6885 3465 6900 3485
rect 6850 3435 6900 3465
rect 6850 3415 6865 3435
rect 6885 3415 6900 3435
rect 6850 3385 6900 3415
rect 6850 3365 6865 3385
rect 6885 3365 6900 3385
rect 6850 3335 6900 3365
rect 6850 3315 6865 3335
rect 6885 3315 6900 3335
rect 6850 3300 6900 3315
rect 7000 3785 7050 3800
rect 7000 3765 7015 3785
rect 7035 3765 7050 3785
rect 7000 3735 7050 3765
rect 7000 3715 7015 3735
rect 7035 3715 7050 3735
rect 7000 3685 7050 3715
rect 7000 3665 7015 3685
rect 7035 3665 7050 3685
rect 7000 3635 7050 3665
rect 7000 3615 7015 3635
rect 7035 3615 7050 3635
rect 7000 3585 7050 3615
rect 7000 3565 7015 3585
rect 7035 3565 7050 3585
rect 7000 3535 7050 3565
rect 7000 3515 7015 3535
rect 7035 3515 7050 3535
rect 7000 3485 7050 3515
rect 7000 3465 7015 3485
rect 7035 3465 7050 3485
rect 7000 3435 7050 3465
rect 7000 3415 7015 3435
rect 7035 3415 7050 3435
rect 7000 3385 7050 3415
rect 7000 3365 7015 3385
rect 7035 3365 7050 3385
rect 7000 3335 7050 3365
rect 7000 3315 7015 3335
rect 7035 3315 7050 3335
rect 7000 3300 7050 3315
rect 7150 3785 7200 3800
rect 7150 3765 7165 3785
rect 7185 3765 7200 3785
rect 7150 3735 7200 3765
rect 7150 3715 7165 3735
rect 7185 3715 7200 3735
rect 7150 3685 7200 3715
rect 7150 3665 7165 3685
rect 7185 3665 7200 3685
rect 7150 3635 7200 3665
rect 7150 3615 7165 3635
rect 7185 3615 7200 3635
rect 7150 3585 7200 3615
rect 7150 3565 7165 3585
rect 7185 3565 7200 3585
rect 7150 3535 7200 3565
rect 7150 3515 7165 3535
rect 7185 3515 7200 3535
rect 7150 3485 7200 3515
rect 7150 3465 7165 3485
rect 7185 3465 7200 3485
rect 7150 3435 7200 3465
rect 7150 3415 7165 3435
rect 7185 3415 7200 3435
rect 7150 3385 7200 3415
rect 7150 3365 7165 3385
rect 7185 3365 7200 3385
rect 7150 3335 7200 3365
rect 7150 3315 7165 3335
rect 7185 3315 7200 3335
rect 7150 3300 7200 3315
rect 7300 3785 7350 3800
rect 7300 3765 7315 3785
rect 7335 3765 7350 3785
rect 7300 3735 7350 3765
rect 7300 3715 7315 3735
rect 7335 3715 7350 3735
rect 7300 3685 7350 3715
rect 7300 3665 7315 3685
rect 7335 3665 7350 3685
rect 7300 3635 7350 3665
rect 7300 3615 7315 3635
rect 7335 3615 7350 3635
rect 7300 3585 7350 3615
rect 7300 3565 7315 3585
rect 7335 3565 7350 3585
rect 7300 3535 7350 3565
rect 7300 3515 7315 3535
rect 7335 3515 7350 3535
rect 7300 3485 7350 3515
rect 7300 3465 7315 3485
rect 7335 3465 7350 3485
rect 7300 3435 7350 3465
rect 7300 3415 7315 3435
rect 7335 3415 7350 3435
rect 7300 3385 7350 3415
rect 7300 3365 7315 3385
rect 7335 3365 7350 3385
rect 7300 3335 7350 3365
rect 7300 3315 7315 3335
rect 7335 3315 7350 3335
rect 7300 3300 7350 3315
rect 7450 3785 7500 3800
rect 7450 3765 7465 3785
rect 7485 3765 7500 3785
rect 7450 3735 7500 3765
rect 7450 3715 7465 3735
rect 7485 3715 7500 3735
rect 7450 3685 7500 3715
rect 7450 3665 7465 3685
rect 7485 3665 7500 3685
rect 7450 3635 7500 3665
rect 7450 3615 7465 3635
rect 7485 3615 7500 3635
rect 7450 3585 7500 3615
rect 7450 3565 7465 3585
rect 7485 3565 7500 3585
rect 7450 3535 7500 3565
rect 7450 3515 7465 3535
rect 7485 3515 7500 3535
rect 7450 3485 7500 3515
rect 7450 3465 7465 3485
rect 7485 3465 7500 3485
rect 7450 3435 7500 3465
rect 7450 3415 7465 3435
rect 7485 3415 7500 3435
rect 7450 3385 7500 3415
rect 7450 3365 7465 3385
rect 7485 3365 7500 3385
rect 7450 3335 7500 3365
rect 7450 3315 7465 3335
rect 7485 3315 7500 3335
rect 7450 3300 7500 3315
rect 7600 3785 7650 3800
rect 7600 3765 7615 3785
rect 7635 3765 7650 3785
rect 7600 3735 7650 3765
rect 7600 3715 7615 3735
rect 7635 3715 7650 3735
rect 7600 3685 7650 3715
rect 7600 3665 7615 3685
rect 7635 3665 7650 3685
rect 7600 3635 7650 3665
rect 7600 3615 7615 3635
rect 7635 3615 7650 3635
rect 7600 3585 7650 3615
rect 7600 3565 7615 3585
rect 7635 3565 7650 3585
rect 7600 3535 7650 3565
rect 7600 3515 7615 3535
rect 7635 3515 7650 3535
rect 7600 3485 7650 3515
rect 7600 3465 7615 3485
rect 7635 3465 7650 3485
rect 7600 3435 7650 3465
rect 7600 3415 7615 3435
rect 7635 3415 7650 3435
rect 7600 3385 7650 3415
rect 7600 3365 7615 3385
rect 7635 3365 7650 3385
rect 7600 3335 7650 3365
rect 7600 3315 7615 3335
rect 7635 3315 7650 3335
rect 7600 3300 7650 3315
rect 7750 3785 7800 3800
rect 7750 3765 7765 3785
rect 7785 3765 7800 3785
rect 7750 3735 7800 3765
rect 7750 3715 7765 3735
rect 7785 3715 7800 3735
rect 7750 3685 7800 3715
rect 7750 3665 7765 3685
rect 7785 3665 7800 3685
rect 7750 3635 7800 3665
rect 7750 3615 7765 3635
rect 7785 3615 7800 3635
rect 7750 3585 7800 3615
rect 7750 3565 7765 3585
rect 7785 3565 7800 3585
rect 7750 3535 7800 3565
rect 7750 3515 7765 3535
rect 7785 3515 7800 3535
rect 7750 3485 7800 3515
rect 7750 3465 7765 3485
rect 7785 3465 7800 3485
rect 7750 3435 7800 3465
rect 7750 3415 7765 3435
rect 7785 3415 7800 3435
rect 7750 3385 7800 3415
rect 7750 3365 7765 3385
rect 7785 3365 7800 3385
rect 7750 3335 7800 3365
rect 7750 3315 7765 3335
rect 7785 3315 7800 3335
rect 7750 3300 7800 3315
rect 8350 3785 8400 3800
rect 8350 3765 8365 3785
rect 8385 3765 8400 3785
rect 8350 3735 8400 3765
rect 8350 3715 8365 3735
rect 8385 3715 8400 3735
rect 8350 3685 8400 3715
rect 8350 3665 8365 3685
rect 8385 3665 8400 3685
rect 8350 3635 8400 3665
rect 8350 3615 8365 3635
rect 8385 3615 8400 3635
rect 8350 3585 8400 3615
rect 8350 3565 8365 3585
rect 8385 3565 8400 3585
rect 8350 3535 8400 3565
rect 8350 3515 8365 3535
rect 8385 3515 8400 3535
rect 8350 3485 8400 3515
rect 8350 3465 8365 3485
rect 8385 3465 8400 3485
rect 8350 3435 8400 3465
rect 8350 3415 8365 3435
rect 8385 3415 8400 3435
rect 8350 3385 8400 3415
rect 8350 3365 8365 3385
rect 8385 3365 8400 3385
rect 8350 3335 8400 3365
rect 8350 3315 8365 3335
rect 8385 3315 8400 3335
rect 8350 3300 8400 3315
rect 8500 3785 8550 3800
rect 8500 3765 8515 3785
rect 8535 3765 8550 3785
rect 8500 3735 8550 3765
rect 8500 3715 8515 3735
rect 8535 3715 8550 3735
rect 8500 3685 8550 3715
rect 8500 3665 8515 3685
rect 8535 3665 8550 3685
rect 8500 3635 8550 3665
rect 8500 3615 8515 3635
rect 8535 3615 8550 3635
rect 8500 3585 8550 3615
rect 8500 3565 8515 3585
rect 8535 3565 8550 3585
rect 8500 3535 8550 3565
rect 8500 3515 8515 3535
rect 8535 3515 8550 3535
rect 8500 3485 8550 3515
rect 8500 3465 8515 3485
rect 8535 3465 8550 3485
rect 8500 3435 8550 3465
rect 8500 3415 8515 3435
rect 8535 3415 8550 3435
rect 8500 3385 8550 3415
rect 8500 3365 8515 3385
rect 8535 3365 8550 3385
rect 8500 3335 8550 3365
rect 8500 3315 8515 3335
rect 8535 3315 8550 3335
rect 8500 3250 8550 3315
rect 8650 3785 8700 3800
rect 8650 3765 8665 3785
rect 8685 3765 8700 3785
rect 8650 3735 8700 3765
rect 8650 3715 8665 3735
rect 8685 3715 8700 3735
rect 8650 3685 8700 3715
rect 8650 3665 8665 3685
rect 8685 3665 8700 3685
rect 8650 3635 8700 3665
rect 8650 3615 8665 3635
rect 8685 3615 8700 3635
rect 8650 3585 8700 3615
rect 8650 3565 8665 3585
rect 8685 3565 8700 3585
rect 8650 3535 8700 3565
rect 8650 3515 8665 3535
rect 8685 3515 8700 3535
rect 8650 3485 8700 3515
rect 8650 3465 8665 3485
rect 8685 3465 8700 3485
rect 8650 3435 8700 3465
rect 8650 3415 8665 3435
rect 8685 3415 8700 3435
rect 8650 3385 8700 3415
rect 8650 3365 8665 3385
rect 8685 3365 8700 3385
rect 8650 3335 8700 3365
rect 8650 3315 8665 3335
rect 8685 3315 8700 3335
rect 8650 3300 8700 3315
rect 8800 3785 8850 3800
rect 8800 3765 8815 3785
rect 8835 3765 8850 3785
rect 8800 3735 8850 3765
rect 8800 3715 8815 3735
rect 8835 3715 8850 3735
rect 8800 3685 8850 3715
rect 8800 3665 8815 3685
rect 8835 3665 8850 3685
rect 8800 3635 8850 3665
rect 8800 3615 8815 3635
rect 8835 3615 8850 3635
rect 8800 3585 8850 3615
rect 8800 3565 8815 3585
rect 8835 3565 8850 3585
rect 8800 3535 8850 3565
rect 8800 3515 8815 3535
rect 8835 3515 8850 3535
rect 8800 3485 8850 3515
rect 8800 3465 8815 3485
rect 8835 3465 8850 3485
rect 8800 3435 8850 3465
rect 8800 3415 8815 3435
rect 8835 3415 8850 3435
rect 8800 3385 8850 3415
rect 8800 3365 8815 3385
rect 8835 3365 8850 3385
rect 8800 3335 8850 3365
rect 8800 3315 8815 3335
rect 8835 3315 8850 3335
rect 8800 3250 8850 3315
rect 8950 3785 9000 3800
rect 8950 3765 8965 3785
rect 8985 3765 9000 3785
rect 8950 3735 9000 3765
rect 8950 3715 8965 3735
rect 8985 3715 9000 3735
rect 8950 3685 9000 3715
rect 8950 3665 8965 3685
rect 8985 3665 9000 3685
rect 8950 3635 9000 3665
rect 8950 3615 8965 3635
rect 8985 3615 9000 3635
rect 8950 3585 9000 3615
rect 8950 3565 8965 3585
rect 8985 3565 9000 3585
rect 8950 3535 9000 3565
rect 8950 3515 8965 3535
rect 8985 3515 9000 3535
rect 8950 3485 9000 3515
rect 8950 3465 8965 3485
rect 8985 3465 9000 3485
rect 8950 3435 9000 3465
rect 8950 3415 8965 3435
rect 8985 3415 9000 3435
rect 8950 3385 9000 3415
rect 8950 3365 8965 3385
rect 8985 3365 9000 3385
rect 8950 3335 9000 3365
rect 8950 3315 8965 3335
rect 8985 3315 9000 3335
rect 8950 3300 9000 3315
rect 9100 3785 9150 3800
rect 9100 3765 9115 3785
rect 9135 3765 9150 3785
rect 9100 3735 9150 3765
rect 9100 3715 9115 3735
rect 9135 3715 9150 3735
rect 9100 3685 9150 3715
rect 9100 3665 9115 3685
rect 9135 3665 9150 3685
rect 9100 3635 9150 3665
rect 9100 3615 9115 3635
rect 9135 3615 9150 3635
rect 9100 3585 9150 3615
rect 9100 3565 9115 3585
rect 9135 3565 9150 3585
rect 9100 3535 9150 3565
rect 9100 3515 9115 3535
rect 9135 3515 9150 3535
rect 9100 3485 9150 3515
rect 9100 3465 9115 3485
rect 9135 3465 9150 3485
rect 9100 3435 9150 3465
rect 9100 3415 9115 3435
rect 9135 3415 9150 3435
rect 9100 3385 9150 3415
rect 9100 3365 9115 3385
rect 9135 3365 9150 3385
rect 9100 3335 9150 3365
rect 9100 3315 9115 3335
rect 9135 3315 9150 3335
rect 9100 3250 9150 3315
rect 9250 3785 9300 3800
rect 9250 3765 9265 3785
rect 9285 3765 9300 3785
rect 9250 3735 9300 3765
rect 9250 3715 9265 3735
rect 9285 3715 9300 3735
rect 9250 3685 9300 3715
rect 9250 3665 9265 3685
rect 9285 3665 9300 3685
rect 9250 3635 9300 3665
rect 9250 3615 9265 3635
rect 9285 3615 9300 3635
rect 9250 3585 9300 3615
rect 9250 3565 9265 3585
rect 9285 3565 9300 3585
rect 9250 3535 9300 3565
rect 9250 3515 9265 3535
rect 9285 3515 9300 3535
rect 9250 3485 9300 3515
rect 9250 3465 9265 3485
rect 9285 3465 9300 3485
rect 9250 3435 9300 3465
rect 9250 3415 9265 3435
rect 9285 3415 9300 3435
rect 9250 3385 9300 3415
rect 9250 3365 9265 3385
rect 9285 3365 9300 3385
rect 9250 3335 9300 3365
rect 9250 3315 9265 3335
rect 9285 3315 9300 3335
rect 9250 3300 9300 3315
rect 9400 3785 9450 3800
rect 9400 3765 9415 3785
rect 9435 3765 9450 3785
rect 9400 3735 9450 3765
rect 9400 3715 9415 3735
rect 9435 3715 9450 3735
rect 9400 3685 9450 3715
rect 9400 3665 9415 3685
rect 9435 3665 9450 3685
rect 9400 3635 9450 3665
rect 9400 3615 9415 3635
rect 9435 3615 9450 3635
rect 9400 3585 9450 3615
rect 9400 3565 9415 3585
rect 9435 3565 9450 3585
rect 9400 3535 9450 3565
rect 9400 3515 9415 3535
rect 9435 3515 9450 3535
rect 9400 3485 9450 3515
rect 9400 3465 9415 3485
rect 9435 3465 9450 3485
rect 9400 3435 9450 3465
rect 9400 3415 9415 3435
rect 9435 3415 9450 3435
rect 9400 3385 9450 3415
rect 9400 3365 9415 3385
rect 9435 3365 9450 3385
rect 9400 3335 9450 3365
rect 9400 3315 9415 3335
rect 9435 3315 9450 3335
rect 9400 3250 9450 3315
rect 9550 3785 9600 3800
rect 9550 3765 9565 3785
rect 9585 3765 9600 3785
rect 9550 3735 9600 3765
rect 9550 3715 9565 3735
rect 9585 3715 9600 3735
rect 9550 3685 9600 3715
rect 9550 3665 9565 3685
rect 9585 3665 9600 3685
rect 9550 3635 9600 3665
rect 9550 3615 9565 3635
rect 9585 3615 9600 3635
rect 9550 3585 9600 3615
rect 9550 3565 9565 3585
rect 9585 3565 9600 3585
rect 9550 3535 9600 3565
rect 9550 3515 9565 3535
rect 9585 3515 9600 3535
rect 9550 3485 9600 3515
rect 9550 3465 9565 3485
rect 9585 3465 9600 3485
rect 9550 3435 9600 3465
rect 9550 3415 9565 3435
rect 9585 3415 9600 3435
rect 9550 3385 9600 3415
rect 9550 3365 9565 3385
rect 9585 3365 9600 3385
rect 9550 3335 9600 3365
rect 9550 3315 9565 3335
rect 9585 3315 9600 3335
rect 9550 3300 9600 3315
rect 9700 3785 9750 3800
rect 9700 3765 9715 3785
rect 9735 3765 9750 3785
rect 9700 3735 9750 3765
rect 9700 3715 9715 3735
rect 9735 3715 9750 3735
rect 9700 3685 9750 3715
rect 9700 3665 9715 3685
rect 9735 3665 9750 3685
rect 9700 3635 9750 3665
rect 9700 3615 9715 3635
rect 9735 3615 9750 3635
rect 9700 3585 9750 3615
rect 9700 3565 9715 3585
rect 9735 3565 9750 3585
rect 9700 3535 9750 3565
rect 9700 3515 9715 3535
rect 9735 3515 9750 3535
rect 9700 3485 9750 3515
rect 9700 3465 9715 3485
rect 9735 3465 9750 3485
rect 9700 3435 9750 3465
rect 9700 3415 9715 3435
rect 9735 3415 9750 3435
rect 9700 3385 9750 3415
rect 9700 3365 9715 3385
rect 9735 3365 9750 3385
rect 9700 3335 9750 3365
rect 9700 3315 9715 3335
rect 9735 3315 9750 3335
rect 9700 3250 9750 3315
rect 9850 3785 9900 3800
rect 9850 3765 9865 3785
rect 9885 3765 9900 3785
rect 9850 3735 9900 3765
rect 9850 3715 9865 3735
rect 9885 3715 9900 3735
rect 9850 3685 9900 3715
rect 9850 3665 9865 3685
rect 9885 3665 9900 3685
rect 9850 3635 9900 3665
rect 9850 3615 9865 3635
rect 9885 3615 9900 3635
rect 9850 3585 9900 3615
rect 9850 3565 9865 3585
rect 9885 3565 9900 3585
rect 9850 3535 9900 3565
rect 9850 3515 9865 3535
rect 9885 3515 9900 3535
rect 9850 3485 9900 3515
rect 9850 3465 9865 3485
rect 9885 3465 9900 3485
rect 9850 3435 9900 3465
rect 9850 3415 9865 3435
rect 9885 3415 9900 3435
rect 9850 3385 9900 3415
rect 9850 3365 9865 3385
rect 9885 3365 9900 3385
rect 9850 3335 9900 3365
rect 9850 3315 9865 3335
rect 9885 3315 9900 3335
rect 9850 3300 9900 3315
rect 10000 3785 10050 3800
rect 10000 3765 10015 3785
rect 10035 3765 10050 3785
rect 10000 3735 10050 3765
rect 10000 3715 10015 3735
rect 10035 3715 10050 3735
rect 10000 3685 10050 3715
rect 10000 3665 10015 3685
rect 10035 3665 10050 3685
rect 10000 3635 10050 3665
rect 10000 3615 10015 3635
rect 10035 3615 10050 3635
rect 10000 3585 10050 3615
rect 10000 3565 10015 3585
rect 10035 3565 10050 3585
rect 10000 3535 10050 3565
rect 10000 3515 10015 3535
rect 10035 3515 10050 3535
rect 10000 3485 10050 3515
rect 10000 3465 10015 3485
rect 10035 3465 10050 3485
rect 10000 3435 10050 3465
rect 10000 3415 10015 3435
rect 10035 3415 10050 3435
rect 10000 3385 10050 3415
rect 10000 3365 10015 3385
rect 10035 3365 10050 3385
rect 10000 3335 10050 3365
rect 10000 3315 10015 3335
rect 10035 3315 10050 3335
rect 10000 3250 10050 3315
rect 10150 3785 10200 3800
rect 10150 3765 10165 3785
rect 10185 3765 10200 3785
rect 10150 3735 10200 3765
rect 10150 3715 10165 3735
rect 10185 3715 10200 3735
rect 10150 3685 10200 3715
rect 10150 3665 10165 3685
rect 10185 3665 10200 3685
rect 10150 3635 10200 3665
rect 10150 3615 10165 3635
rect 10185 3615 10200 3635
rect 10150 3585 10200 3615
rect 10150 3565 10165 3585
rect 10185 3565 10200 3585
rect 10150 3535 10200 3565
rect 10150 3515 10165 3535
rect 10185 3515 10200 3535
rect 10150 3485 10200 3515
rect 10150 3465 10165 3485
rect 10185 3465 10200 3485
rect 10150 3435 10200 3465
rect 10150 3415 10165 3435
rect 10185 3415 10200 3435
rect 10150 3385 10200 3415
rect 10150 3365 10165 3385
rect 10185 3365 10200 3385
rect 10150 3335 10200 3365
rect 10150 3315 10165 3335
rect 10185 3315 10200 3335
rect 10150 3300 10200 3315
rect 10300 3785 10350 3800
rect 10300 3765 10315 3785
rect 10335 3765 10350 3785
rect 10300 3735 10350 3765
rect 10300 3715 10315 3735
rect 10335 3715 10350 3735
rect 10300 3685 10350 3715
rect 10300 3665 10315 3685
rect 10335 3665 10350 3685
rect 10300 3635 10350 3665
rect 10300 3615 10315 3635
rect 10335 3615 10350 3635
rect 10300 3585 10350 3615
rect 10300 3565 10315 3585
rect 10335 3565 10350 3585
rect 10300 3535 10350 3565
rect 10300 3515 10315 3535
rect 10335 3515 10350 3535
rect 10300 3485 10350 3515
rect 10300 3465 10315 3485
rect 10335 3465 10350 3485
rect 10300 3435 10350 3465
rect 10300 3415 10315 3435
rect 10335 3415 10350 3435
rect 10300 3385 10350 3415
rect 10300 3365 10315 3385
rect 10335 3365 10350 3385
rect 10300 3335 10350 3365
rect 10300 3315 10315 3335
rect 10335 3315 10350 3335
rect 10300 3250 10350 3315
rect 10450 3785 10500 3800
rect 10450 3765 10465 3785
rect 10485 3765 10500 3785
rect 10450 3735 10500 3765
rect 10450 3715 10465 3735
rect 10485 3715 10500 3735
rect 10450 3685 10500 3715
rect 10450 3665 10465 3685
rect 10485 3665 10500 3685
rect 10450 3635 10500 3665
rect 10450 3615 10465 3635
rect 10485 3615 10500 3635
rect 10450 3585 10500 3615
rect 10450 3565 10465 3585
rect 10485 3565 10500 3585
rect 10450 3535 10500 3565
rect 10450 3515 10465 3535
rect 10485 3515 10500 3535
rect 10450 3485 10500 3515
rect 10450 3465 10465 3485
rect 10485 3465 10500 3485
rect 10450 3435 10500 3465
rect 10450 3415 10465 3435
rect 10485 3415 10500 3435
rect 10450 3385 10500 3415
rect 10450 3365 10465 3385
rect 10485 3365 10500 3385
rect 10450 3335 10500 3365
rect 10450 3315 10465 3335
rect 10485 3315 10500 3335
rect 10450 3300 10500 3315
rect 10600 3785 10650 3800
rect 10600 3765 10615 3785
rect 10635 3765 10650 3785
rect 10600 3735 10650 3765
rect 10600 3715 10615 3735
rect 10635 3715 10650 3735
rect 10600 3685 10650 3715
rect 10600 3665 10615 3685
rect 10635 3665 10650 3685
rect 10600 3635 10650 3665
rect 10600 3615 10615 3635
rect 10635 3615 10650 3635
rect 10600 3585 10650 3615
rect 10600 3565 10615 3585
rect 10635 3565 10650 3585
rect 10600 3535 10650 3565
rect 10600 3515 10615 3535
rect 10635 3515 10650 3535
rect 10600 3485 10650 3515
rect 10600 3465 10615 3485
rect 10635 3465 10650 3485
rect 10600 3435 10650 3465
rect 10600 3415 10615 3435
rect 10635 3415 10650 3435
rect 10600 3385 10650 3415
rect 10600 3365 10615 3385
rect 10635 3365 10650 3385
rect 10600 3335 10650 3365
rect 10600 3315 10615 3335
rect 10635 3315 10650 3335
rect 10600 3250 10650 3315
rect 10750 3785 10800 3800
rect 10750 3765 10765 3785
rect 10785 3765 10800 3785
rect 10750 3735 10800 3765
rect 10750 3715 10765 3735
rect 10785 3715 10800 3735
rect 10750 3685 10800 3715
rect 10750 3665 10765 3685
rect 10785 3665 10800 3685
rect 10750 3635 10800 3665
rect 10750 3615 10765 3635
rect 10785 3615 10800 3635
rect 10750 3585 10800 3615
rect 10750 3565 10765 3585
rect 10785 3565 10800 3585
rect 10750 3535 10800 3565
rect 10750 3515 10765 3535
rect 10785 3515 10800 3535
rect 10750 3485 10800 3515
rect 10750 3465 10765 3485
rect 10785 3465 10800 3485
rect 10750 3435 10800 3465
rect 10750 3415 10765 3435
rect 10785 3415 10800 3435
rect 10750 3385 10800 3415
rect 10750 3365 10765 3385
rect 10785 3365 10800 3385
rect 10750 3335 10800 3365
rect 10750 3315 10765 3335
rect 10785 3315 10800 3335
rect 10750 3300 10800 3315
rect 11350 3785 11400 3800
rect 11350 3765 11365 3785
rect 11385 3765 11400 3785
rect 11350 3735 11400 3765
rect 11350 3715 11365 3735
rect 11385 3715 11400 3735
rect 11350 3685 11400 3715
rect 11350 3665 11365 3685
rect 11385 3665 11400 3685
rect 11350 3635 11400 3665
rect 11350 3615 11365 3635
rect 11385 3615 11400 3635
rect 11350 3585 11400 3615
rect 11350 3565 11365 3585
rect 11385 3565 11400 3585
rect 11350 3535 11400 3565
rect 11350 3515 11365 3535
rect 11385 3515 11400 3535
rect 11350 3485 11400 3515
rect 11350 3465 11365 3485
rect 11385 3465 11400 3485
rect 11350 3435 11400 3465
rect 11350 3415 11365 3435
rect 11385 3415 11400 3435
rect 11350 3385 11400 3415
rect 11350 3365 11365 3385
rect 11385 3365 11400 3385
rect 11350 3335 11400 3365
rect 11350 3315 11365 3335
rect 11385 3315 11400 3335
rect 11350 3300 11400 3315
rect 11950 3785 12000 3800
rect 11950 3765 11965 3785
rect 11985 3765 12000 3785
rect 11950 3735 12000 3765
rect 11950 3715 11965 3735
rect 11985 3715 12000 3735
rect 11950 3685 12000 3715
rect 11950 3665 11965 3685
rect 11985 3665 12000 3685
rect 11950 3635 12000 3665
rect 11950 3615 11965 3635
rect 11985 3615 12000 3635
rect 11950 3585 12000 3615
rect 11950 3565 11965 3585
rect 11985 3565 12000 3585
rect 11950 3535 12000 3565
rect 11950 3515 11965 3535
rect 11985 3515 12000 3535
rect 11950 3485 12000 3515
rect 11950 3465 11965 3485
rect 11985 3465 12000 3485
rect 11950 3435 12000 3465
rect 11950 3415 11965 3435
rect 11985 3415 12000 3435
rect 11950 3385 12000 3415
rect 11950 3365 11965 3385
rect 11985 3365 12000 3385
rect 11950 3335 12000 3365
rect 11950 3315 11965 3335
rect 11985 3315 12000 3335
rect 11950 3300 12000 3315
rect 12550 3785 12600 3800
rect 12550 3765 12565 3785
rect 12585 3765 12600 3785
rect 12550 3735 12600 3765
rect 12550 3715 12565 3735
rect 12585 3715 12600 3735
rect 12550 3685 12600 3715
rect 12550 3665 12565 3685
rect 12585 3665 12600 3685
rect 12550 3635 12600 3665
rect 12550 3615 12565 3635
rect 12585 3615 12600 3635
rect 12550 3585 12600 3615
rect 12550 3565 12565 3585
rect 12585 3565 12600 3585
rect 12550 3535 12600 3565
rect 12550 3515 12565 3535
rect 12585 3515 12600 3535
rect 12550 3485 12600 3515
rect 12550 3465 12565 3485
rect 12585 3465 12600 3485
rect 12550 3435 12600 3465
rect 12550 3415 12565 3435
rect 12585 3415 12600 3435
rect 12550 3385 12600 3415
rect 12550 3365 12565 3385
rect 12585 3365 12600 3385
rect 12550 3335 12600 3365
rect 12550 3315 12565 3335
rect 12585 3315 12600 3335
rect 12550 3300 12600 3315
rect 13150 3785 13200 3800
rect 13150 3765 13165 3785
rect 13185 3765 13200 3785
rect 13150 3735 13200 3765
rect 13150 3715 13165 3735
rect 13185 3715 13200 3735
rect 13150 3685 13200 3715
rect 13150 3665 13165 3685
rect 13185 3665 13200 3685
rect 13150 3635 13200 3665
rect 13150 3615 13165 3635
rect 13185 3615 13200 3635
rect 13150 3585 13200 3615
rect 13150 3565 13165 3585
rect 13185 3565 13200 3585
rect 13150 3535 13200 3565
rect 13150 3515 13165 3535
rect 13185 3515 13200 3535
rect 13150 3485 13200 3515
rect 13150 3465 13165 3485
rect 13185 3465 13200 3485
rect 13150 3435 13200 3465
rect 13150 3415 13165 3435
rect 13185 3415 13200 3435
rect 13150 3385 13200 3415
rect 13150 3365 13165 3385
rect 13185 3365 13200 3385
rect 13150 3335 13200 3365
rect 13150 3315 13165 3335
rect 13185 3315 13200 3335
rect 13150 3300 13200 3315
rect 13750 3785 13800 3800
rect 13750 3765 13765 3785
rect 13785 3765 13800 3785
rect 13750 3735 13800 3765
rect 13750 3715 13765 3735
rect 13785 3715 13800 3735
rect 13750 3685 13800 3715
rect 13750 3665 13765 3685
rect 13785 3665 13800 3685
rect 13750 3635 13800 3665
rect 13750 3615 13765 3635
rect 13785 3615 13800 3635
rect 13750 3585 13800 3615
rect 13750 3565 13765 3585
rect 13785 3565 13800 3585
rect 13750 3535 13800 3565
rect 13750 3515 13765 3535
rect 13785 3515 13800 3535
rect 13750 3485 13800 3515
rect 13750 3465 13765 3485
rect 13785 3465 13800 3485
rect 13750 3435 13800 3465
rect 13750 3415 13765 3435
rect 13785 3415 13800 3435
rect 13750 3385 13800 3415
rect 13750 3365 13765 3385
rect 13785 3365 13800 3385
rect 13750 3335 13800 3365
rect 13750 3315 13765 3335
rect 13785 3315 13800 3335
rect 13750 3300 13800 3315
rect 14350 3785 14400 3800
rect 14350 3765 14365 3785
rect 14385 3765 14400 3785
rect 14350 3735 14400 3765
rect 14350 3715 14365 3735
rect 14385 3715 14400 3735
rect 14350 3685 14400 3715
rect 14350 3665 14365 3685
rect 14385 3665 14400 3685
rect 14350 3635 14400 3665
rect 14350 3615 14365 3635
rect 14385 3615 14400 3635
rect 14350 3585 14400 3615
rect 14350 3565 14365 3585
rect 14385 3565 14400 3585
rect 14350 3535 14400 3565
rect 14350 3515 14365 3535
rect 14385 3515 14400 3535
rect 14350 3485 14400 3515
rect 14350 3465 14365 3485
rect 14385 3465 14400 3485
rect 14350 3435 14400 3465
rect 14350 3415 14365 3435
rect 14385 3415 14400 3435
rect 14350 3385 14400 3415
rect 14350 3365 14365 3385
rect 14385 3365 14400 3385
rect 14350 3335 14400 3365
rect 14350 3315 14365 3335
rect 14385 3315 14400 3335
rect 14350 3300 14400 3315
rect 14950 3785 15000 3800
rect 14950 3765 14965 3785
rect 14985 3765 15000 3785
rect 14950 3735 15000 3765
rect 14950 3715 14965 3735
rect 14985 3715 15000 3735
rect 14950 3685 15000 3715
rect 14950 3665 14965 3685
rect 14985 3665 15000 3685
rect 14950 3635 15000 3665
rect 14950 3615 14965 3635
rect 14985 3615 15000 3635
rect 14950 3585 15000 3615
rect 14950 3565 14965 3585
rect 14985 3565 15000 3585
rect 14950 3535 15000 3565
rect 14950 3515 14965 3535
rect 14985 3515 15000 3535
rect 14950 3485 15000 3515
rect 14950 3465 14965 3485
rect 14985 3465 15000 3485
rect 14950 3435 15000 3465
rect 14950 3415 14965 3435
rect 14985 3415 15000 3435
rect 14950 3385 15000 3415
rect 14950 3365 14965 3385
rect 14985 3365 15000 3385
rect 14950 3335 15000 3365
rect 14950 3315 14965 3335
rect 14985 3315 15000 3335
rect 14950 3300 15000 3315
rect 15550 3785 15600 3800
rect 15550 3765 15565 3785
rect 15585 3765 15600 3785
rect 15550 3735 15600 3765
rect 15550 3715 15565 3735
rect 15585 3715 15600 3735
rect 15550 3685 15600 3715
rect 15550 3665 15565 3685
rect 15585 3665 15600 3685
rect 15550 3635 15600 3665
rect 15550 3615 15565 3635
rect 15585 3615 15600 3635
rect 15550 3585 15600 3615
rect 15550 3565 15565 3585
rect 15585 3565 15600 3585
rect 15550 3535 15600 3565
rect 15550 3515 15565 3535
rect 15585 3515 15600 3535
rect 15550 3485 15600 3515
rect 15550 3465 15565 3485
rect 15585 3465 15600 3485
rect 15550 3435 15600 3465
rect 15550 3415 15565 3435
rect 15585 3415 15600 3435
rect 15550 3385 15600 3415
rect 15550 3365 15565 3385
rect 15585 3365 15600 3385
rect 15550 3335 15600 3365
rect 15550 3315 15565 3335
rect 15585 3315 15600 3335
rect 15550 3300 15600 3315
rect 16150 3785 16200 3800
rect 16150 3765 16165 3785
rect 16185 3765 16200 3785
rect 16150 3735 16200 3765
rect 16150 3715 16165 3735
rect 16185 3715 16200 3735
rect 16150 3685 16200 3715
rect 16150 3665 16165 3685
rect 16185 3665 16200 3685
rect 16150 3635 16200 3665
rect 16150 3615 16165 3635
rect 16185 3615 16200 3635
rect 16150 3585 16200 3615
rect 16150 3565 16165 3585
rect 16185 3565 16200 3585
rect 16150 3535 16200 3565
rect 16150 3515 16165 3535
rect 16185 3515 16200 3535
rect 16150 3485 16200 3515
rect 16150 3465 16165 3485
rect 16185 3465 16200 3485
rect 16150 3435 16200 3465
rect 16150 3415 16165 3435
rect 16185 3415 16200 3435
rect 16150 3385 16200 3415
rect 16150 3365 16165 3385
rect 16185 3365 16200 3385
rect 16150 3335 16200 3365
rect 16150 3315 16165 3335
rect 16185 3315 16200 3335
rect 16150 3300 16200 3315
rect 16300 3785 16350 3800
rect 16300 3765 16315 3785
rect 16335 3765 16350 3785
rect 16300 3735 16350 3765
rect 16300 3715 16315 3735
rect 16335 3715 16350 3735
rect 16300 3685 16350 3715
rect 16300 3665 16315 3685
rect 16335 3665 16350 3685
rect 16300 3635 16350 3665
rect 16300 3615 16315 3635
rect 16335 3615 16350 3635
rect 16300 3585 16350 3615
rect 16300 3565 16315 3585
rect 16335 3565 16350 3585
rect 16300 3535 16350 3565
rect 16300 3515 16315 3535
rect 16335 3515 16350 3535
rect 16300 3485 16350 3515
rect 16300 3465 16315 3485
rect 16335 3465 16350 3485
rect 16300 3435 16350 3465
rect 16300 3415 16315 3435
rect 16335 3415 16350 3435
rect 16300 3385 16350 3415
rect 16300 3365 16315 3385
rect 16335 3365 16350 3385
rect 16300 3335 16350 3365
rect 16300 3315 16315 3335
rect 16335 3315 16350 3335
rect 16300 3300 16350 3315
rect 16450 3785 16500 3800
rect 16450 3765 16465 3785
rect 16485 3765 16500 3785
rect 16450 3735 16500 3765
rect 16450 3715 16465 3735
rect 16485 3715 16500 3735
rect 16450 3685 16500 3715
rect 16450 3665 16465 3685
rect 16485 3665 16500 3685
rect 16450 3635 16500 3665
rect 16450 3615 16465 3635
rect 16485 3615 16500 3635
rect 16450 3585 16500 3615
rect 16450 3565 16465 3585
rect 16485 3565 16500 3585
rect 16450 3535 16500 3565
rect 16450 3515 16465 3535
rect 16485 3515 16500 3535
rect 16450 3485 16500 3515
rect 16450 3465 16465 3485
rect 16485 3465 16500 3485
rect 16450 3435 16500 3465
rect 16450 3415 16465 3435
rect 16485 3415 16500 3435
rect 16450 3385 16500 3415
rect 16450 3365 16465 3385
rect 16485 3365 16500 3385
rect 16450 3335 16500 3365
rect 16450 3315 16465 3335
rect 16485 3315 16500 3335
rect 16450 3300 16500 3315
rect 16600 3785 16650 3800
rect 16600 3765 16615 3785
rect 16635 3765 16650 3785
rect 16600 3735 16650 3765
rect 16600 3715 16615 3735
rect 16635 3715 16650 3735
rect 16600 3685 16650 3715
rect 16600 3665 16615 3685
rect 16635 3665 16650 3685
rect 16600 3635 16650 3665
rect 16600 3615 16615 3635
rect 16635 3615 16650 3635
rect 16600 3585 16650 3615
rect 16600 3565 16615 3585
rect 16635 3565 16650 3585
rect 16600 3535 16650 3565
rect 16600 3515 16615 3535
rect 16635 3515 16650 3535
rect 16600 3485 16650 3515
rect 16600 3465 16615 3485
rect 16635 3465 16650 3485
rect 16600 3435 16650 3465
rect 16600 3415 16615 3435
rect 16635 3415 16650 3435
rect 16600 3385 16650 3415
rect 16600 3365 16615 3385
rect 16635 3365 16650 3385
rect 16600 3335 16650 3365
rect 16600 3315 16615 3335
rect 16635 3315 16650 3335
rect 16600 3300 16650 3315
rect 16750 3785 16800 3800
rect 16750 3765 16765 3785
rect 16785 3765 16800 3785
rect 16750 3735 16800 3765
rect 16750 3715 16765 3735
rect 16785 3715 16800 3735
rect 16750 3685 16800 3715
rect 16750 3665 16765 3685
rect 16785 3665 16800 3685
rect 16750 3635 16800 3665
rect 16750 3615 16765 3635
rect 16785 3615 16800 3635
rect 16750 3585 16800 3615
rect 16750 3565 16765 3585
rect 16785 3565 16800 3585
rect 16750 3535 16800 3565
rect 16750 3515 16765 3535
rect 16785 3515 16800 3535
rect 16750 3485 16800 3515
rect 16750 3465 16765 3485
rect 16785 3465 16800 3485
rect 16750 3435 16800 3465
rect 16750 3415 16765 3435
rect 16785 3415 16800 3435
rect 16750 3385 16800 3415
rect 16750 3365 16765 3385
rect 16785 3365 16800 3385
rect 16750 3335 16800 3365
rect 16750 3315 16765 3335
rect 16785 3315 16800 3335
rect 16750 3300 16800 3315
rect 16900 3785 16950 3800
rect 16900 3765 16915 3785
rect 16935 3765 16950 3785
rect 16900 3735 16950 3765
rect 16900 3715 16915 3735
rect 16935 3715 16950 3735
rect 16900 3685 16950 3715
rect 16900 3665 16915 3685
rect 16935 3665 16950 3685
rect 16900 3635 16950 3665
rect 16900 3615 16915 3635
rect 16935 3615 16950 3635
rect 16900 3585 16950 3615
rect 16900 3565 16915 3585
rect 16935 3565 16950 3585
rect 16900 3535 16950 3565
rect 16900 3515 16915 3535
rect 16935 3515 16950 3535
rect 16900 3485 16950 3515
rect 16900 3465 16915 3485
rect 16935 3465 16950 3485
rect 16900 3435 16950 3465
rect 16900 3415 16915 3435
rect 16935 3415 16950 3435
rect 16900 3385 16950 3415
rect 16900 3365 16915 3385
rect 16935 3365 16950 3385
rect 16900 3335 16950 3365
rect 16900 3315 16915 3335
rect 16935 3315 16950 3335
rect 16900 3300 16950 3315
rect 17050 3785 17100 3800
rect 17050 3765 17065 3785
rect 17085 3765 17100 3785
rect 17050 3735 17100 3765
rect 17050 3715 17065 3735
rect 17085 3715 17100 3735
rect 17050 3685 17100 3715
rect 17050 3665 17065 3685
rect 17085 3665 17100 3685
rect 17050 3635 17100 3665
rect 17050 3615 17065 3635
rect 17085 3615 17100 3635
rect 17050 3585 17100 3615
rect 17050 3565 17065 3585
rect 17085 3565 17100 3585
rect 17050 3535 17100 3565
rect 17050 3515 17065 3535
rect 17085 3515 17100 3535
rect 17050 3485 17100 3515
rect 17050 3465 17065 3485
rect 17085 3465 17100 3485
rect 17050 3435 17100 3465
rect 17050 3415 17065 3435
rect 17085 3415 17100 3435
rect 17050 3385 17100 3415
rect 17050 3365 17065 3385
rect 17085 3365 17100 3385
rect 17050 3335 17100 3365
rect 17050 3315 17065 3335
rect 17085 3315 17100 3335
rect 17050 3300 17100 3315
rect 17200 3785 17250 3800
rect 17200 3765 17215 3785
rect 17235 3765 17250 3785
rect 17200 3735 17250 3765
rect 17200 3715 17215 3735
rect 17235 3715 17250 3735
rect 17200 3685 17250 3715
rect 17200 3665 17215 3685
rect 17235 3665 17250 3685
rect 17200 3635 17250 3665
rect 17200 3615 17215 3635
rect 17235 3615 17250 3635
rect 17200 3585 17250 3615
rect 17200 3565 17215 3585
rect 17235 3565 17250 3585
rect 17200 3535 17250 3565
rect 17200 3515 17215 3535
rect 17235 3515 17250 3535
rect 17200 3485 17250 3515
rect 17200 3465 17215 3485
rect 17235 3465 17250 3485
rect 17200 3435 17250 3465
rect 17200 3415 17215 3435
rect 17235 3415 17250 3435
rect 17200 3385 17250 3415
rect 17200 3365 17215 3385
rect 17235 3365 17250 3385
rect 17200 3335 17250 3365
rect 17200 3315 17215 3335
rect 17235 3315 17250 3335
rect 17200 3300 17250 3315
rect 17350 3785 17400 3800
rect 17350 3765 17365 3785
rect 17385 3765 17400 3785
rect 17350 3735 17400 3765
rect 17350 3715 17365 3735
rect 17385 3715 17400 3735
rect 17350 3685 17400 3715
rect 17350 3665 17365 3685
rect 17385 3665 17400 3685
rect 17350 3635 17400 3665
rect 17350 3615 17365 3635
rect 17385 3615 17400 3635
rect 17350 3585 17400 3615
rect 17350 3565 17365 3585
rect 17385 3565 17400 3585
rect 17350 3535 17400 3565
rect 17350 3515 17365 3535
rect 17385 3515 17400 3535
rect 17350 3485 17400 3515
rect 17350 3465 17365 3485
rect 17385 3465 17400 3485
rect 17350 3435 17400 3465
rect 17350 3415 17365 3435
rect 17385 3415 17400 3435
rect 17350 3385 17400 3415
rect 17350 3365 17365 3385
rect 17385 3365 17400 3385
rect 17350 3335 17400 3365
rect 17350 3315 17365 3335
rect 17385 3315 17400 3335
rect 17350 3300 17400 3315
rect 17950 3785 18000 3800
rect 17950 3765 17965 3785
rect 17985 3765 18000 3785
rect 17950 3735 18000 3765
rect 17950 3715 17965 3735
rect 17985 3715 18000 3735
rect 17950 3685 18000 3715
rect 17950 3665 17965 3685
rect 17985 3665 18000 3685
rect 17950 3635 18000 3665
rect 17950 3615 17965 3635
rect 17985 3615 18000 3635
rect 17950 3585 18000 3615
rect 17950 3565 17965 3585
rect 17985 3565 18000 3585
rect 17950 3535 18000 3565
rect 17950 3515 17965 3535
rect 17985 3515 18000 3535
rect 17950 3485 18000 3515
rect 17950 3465 17965 3485
rect 17985 3465 18000 3485
rect 17950 3435 18000 3465
rect 17950 3415 17965 3435
rect 17985 3415 18000 3435
rect 17950 3385 18000 3415
rect 17950 3365 17965 3385
rect 17985 3365 18000 3385
rect 17950 3335 18000 3365
rect 17950 3315 17965 3335
rect 17985 3315 18000 3335
rect 17950 3300 18000 3315
rect 18550 3785 18600 3800
rect 18550 3765 18565 3785
rect 18585 3765 18600 3785
rect 18550 3735 18600 3765
rect 18550 3715 18565 3735
rect 18585 3715 18600 3735
rect 18550 3685 18600 3715
rect 18550 3665 18565 3685
rect 18585 3665 18600 3685
rect 18550 3635 18600 3665
rect 18550 3615 18565 3635
rect 18585 3615 18600 3635
rect 18550 3585 18600 3615
rect 18550 3565 18565 3585
rect 18585 3565 18600 3585
rect 18550 3535 18600 3565
rect 18550 3515 18565 3535
rect 18585 3515 18600 3535
rect 18550 3485 18600 3515
rect 18550 3465 18565 3485
rect 18585 3465 18600 3485
rect 18550 3435 18600 3465
rect 18550 3415 18565 3435
rect 18585 3415 18600 3435
rect 18550 3385 18600 3415
rect 18550 3365 18565 3385
rect 18585 3365 18600 3385
rect 18550 3335 18600 3365
rect 18550 3315 18565 3335
rect 18585 3315 18600 3335
rect 18550 3300 18600 3315
rect 18700 3785 18750 3800
rect 18700 3765 18715 3785
rect 18735 3765 18750 3785
rect 18700 3735 18750 3765
rect 18700 3715 18715 3735
rect 18735 3715 18750 3735
rect 18700 3685 18750 3715
rect 18700 3665 18715 3685
rect 18735 3665 18750 3685
rect 18700 3635 18750 3665
rect 18700 3615 18715 3635
rect 18735 3615 18750 3635
rect 18700 3585 18750 3615
rect 18700 3565 18715 3585
rect 18735 3565 18750 3585
rect 18700 3535 18750 3565
rect 18700 3515 18715 3535
rect 18735 3515 18750 3535
rect 18700 3485 18750 3515
rect 18700 3465 18715 3485
rect 18735 3465 18750 3485
rect 18700 3435 18750 3465
rect 18700 3415 18715 3435
rect 18735 3415 18750 3435
rect 18700 3385 18750 3415
rect 18700 3365 18715 3385
rect 18735 3365 18750 3385
rect 18700 3335 18750 3365
rect 18700 3315 18715 3335
rect 18735 3315 18750 3335
rect 18700 3300 18750 3315
rect 18850 3785 18900 3800
rect 18850 3765 18865 3785
rect 18885 3765 18900 3785
rect 18850 3735 18900 3765
rect 18850 3715 18865 3735
rect 18885 3715 18900 3735
rect 18850 3685 18900 3715
rect 18850 3665 18865 3685
rect 18885 3665 18900 3685
rect 18850 3635 18900 3665
rect 18850 3615 18865 3635
rect 18885 3615 18900 3635
rect 18850 3585 18900 3615
rect 18850 3565 18865 3585
rect 18885 3565 18900 3585
rect 18850 3535 18900 3565
rect 18850 3515 18865 3535
rect 18885 3515 18900 3535
rect 18850 3485 18900 3515
rect 18850 3465 18865 3485
rect 18885 3465 18900 3485
rect 18850 3435 18900 3465
rect 18850 3415 18865 3435
rect 18885 3415 18900 3435
rect 18850 3385 18900 3415
rect 18850 3365 18865 3385
rect 18885 3365 18900 3385
rect 18850 3335 18900 3365
rect 18850 3315 18865 3335
rect 18885 3315 18900 3335
rect 18850 3300 18900 3315
rect 19000 3785 19050 3800
rect 19000 3765 19015 3785
rect 19035 3765 19050 3785
rect 19000 3735 19050 3765
rect 19000 3715 19015 3735
rect 19035 3715 19050 3735
rect 19000 3685 19050 3715
rect 19000 3665 19015 3685
rect 19035 3665 19050 3685
rect 19000 3635 19050 3665
rect 19000 3615 19015 3635
rect 19035 3615 19050 3635
rect 19000 3585 19050 3615
rect 19000 3565 19015 3585
rect 19035 3565 19050 3585
rect 19000 3535 19050 3565
rect 19000 3515 19015 3535
rect 19035 3515 19050 3535
rect 19000 3485 19050 3515
rect 19000 3465 19015 3485
rect 19035 3465 19050 3485
rect 19000 3435 19050 3465
rect 19000 3415 19015 3435
rect 19035 3415 19050 3435
rect 19000 3385 19050 3415
rect 19000 3365 19015 3385
rect 19035 3365 19050 3385
rect 19000 3335 19050 3365
rect 19000 3315 19015 3335
rect 19035 3315 19050 3335
rect 19000 3300 19050 3315
rect 19150 3785 19200 3800
rect 19150 3765 19165 3785
rect 19185 3765 19200 3785
rect 19150 3735 19200 3765
rect 19150 3715 19165 3735
rect 19185 3715 19200 3735
rect 19150 3685 19200 3715
rect 19150 3665 19165 3685
rect 19185 3665 19200 3685
rect 19150 3635 19200 3665
rect 19150 3615 19165 3635
rect 19185 3615 19200 3635
rect 19150 3585 19200 3615
rect 19150 3565 19165 3585
rect 19185 3565 19200 3585
rect 19150 3535 19200 3565
rect 19150 3515 19165 3535
rect 19185 3515 19200 3535
rect 19150 3485 19200 3515
rect 19150 3465 19165 3485
rect 19185 3465 19200 3485
rect 19150 3435 19200 3465
rect 19150 3415 19165 3435
rect 19185 3415 19200 3435
rect 19150 3385 19200 3415
rect 19150 3365 19165 3385
rect 19185 3365 19200 3385
rect 19150 3335 19200 3365
rect 19150 3315 19165 3335
rect 19185 3315 19200 3335
rect 19150 3300 19200 3315
rect 19300 3785 19350 3800
rect 19300 3765 19315 3785
rect 19335 3765 19350 3785
rect 19300 3735 19350 3765
rect 19300 3715 19315 3735
rect 19335 3715 19350 3735
rect 19300 3685 19350 3715
rect 19300 3665 19315 3685
rect 19335 3665 19350 3685
rect 19300 3635 19350 3665
rect 19300 3615 19315 3635
rect 19335 3615 19350 3635
rect 19300 3585 19350 3615
rect 19300 3565 19315 3585
rect 19335 3565 19350 3585
rect 19300 3535 19350 3565
rect 19300 3515 19315 3535
rect 19335 3515 19350 3535
rect 19300 3485 19350 3515
rect 19300 3465 19315 3485
rect 19335 3465 19350 3485
rect 19300 3435 19350 3465
rect 19300 3415 19315 3435
rect 19335 3415 19350 3435
rect 19300 3385 19350 3415
rect 19300 3365 19315 3385
rect 19335 3365 19350 3385
rect 19300 3335 19350 3365
rect 19300 3315 19315 3335
rect 19335 3315 19350 3335
rect 19300 3300 19350 3315
rect 19450 3785 19500 3800
rect 19450 3765 19465 3785
rect 19485 3765 19500 3785
rect 19450 3735 19500 3765
rect 19450 3715 19465 3735
rect 19485 3715 19500 3735
rect 19450 3685 19500 3715
rect 19450 3665 19465 3685
rect 19485 3665 19500 3685
rect 19450 3635 19500 3665
rect 19450 3615 19465 3635
rect 19485 3615 19500 3635
rect 19450 3585 19500 3615
rect 19450 3565 19465 3585
rect 19485 3565 19500 3585
rect 19450 3535 19500 3565
rect 19450 3515 19465 3535
rect 19485 3515 19500 3535
rect 19450 3485 19500 3515
rect 19450 3465 19465 3485
rect 19485 3465 19500 3485
rect 19450 3435 19500 3465
rect 19450 3415 19465 3435
rect 19485 3415 19500 3435
rect 19450 3385 19500 3415
rect 19450 3365 19465 3385
rect 19485 3365 19500 3385
rect 19450 3335 19500 3365
rect 19450 3315 19465 3335
rect 19485 3315 19500 3335
rect 19450 3300 19500 3315
rect 19600 3785 19650 3800
rect 19600 3765 19615 3785
rect 19635 3765 19650 3785
rect 19600 3735 19650 3765
rect 19600 3715 19615 3735
rect 19635 3715 19650 3735
rect 19600 3685 19650 3715
rect 19600 3665 19615 3685
rect 19635 3665 19650 3685
rect 19600 3635 19650 3665
rect 19600 3615 19615 3635
rect 19635 3615 19650 3635
rect 19600 3585 19650 3615
rect 19600 3565 19615 3585
rect 19635 3565 19650 3585
rect 19600 3535 19650 3565
rect 19600 3515 19615 3535
rect 19635 3515 19650 3535
rect 19600 3485 19650 3515
rect 19600 3465 19615 3485
rect 19635 3465 19650 3485
rect 19600 3435 19650 3465
rect 19600 3415 19615 3435
rect 19635 3415 19650 3435
rect 19600 3385 19650 3415
rect 19600 3365 19615 3385
rect 19635 3365 19650 3385
rect 19600 3335 19650 3365
rect 19600 3315 19615 3335
rect 19635 3315 19650 3335
rect 19600 3300 19650 3315
rect 19750 3785 19800 3800
rect 19750 3765 19765 3785
rect 19785 3765 19800 3785
rect 19750 3735 19800 3765
rect 19750 3715 19765 3735
rect 19785 3715 19800 3735
rect 19750 3685 19800 3715
rect 19750 3665 19765 3685
rect 19785 3665 19800 3685
rect 19750 3635 19800 3665
rect 19750 3615 19765 3635
rect 19785 3615 19800 3635
rect 19750 3585 19800 3615
rect 19750 3565 19765 3585
rect 19785 3565 19800 3585
rect 19750 3535 19800 3565
rect 19750 3515 19765 3535
rect 19785 3515 19800 3535
rect 19750 3485 19800 3515
rect 19750 3465 19765 3485
rect 19785 3465 19800 3485
rect 19750 3435 19800 3465
rect 19750 3415 19765 3435
rect 19785 3415 19800 3435
rect 19750 3385 19800 3415
rect 19750 3365 19765 3385
rect 19785 3365 19800 3385
rect 19750 3335 19800 3365
rect 19750 3315 19765 3335
rect 19785 3315 19800 3335
rect 19750 3300 19800 3315
rect 20350 3785 20400 3800
rect 20350 3765 20365 3785
rect 20385 3765 20400 3785
rect 20350 3735 20400 3765
rect 20350 3715 20365 3735
rect 20385 3715 20400 3735
rect 20350 3685 20400 3715
rect 20350 3665 20365 3685
rect 20385 3665 20400 3685
rect 20350 3635 20400 3665
rect 20350 3615 20365 3635
rect 20385 3615 20400 3635
rect 20350 3585 20400 3615
rect 20350 3565 20365 3585
rect 20385 3565 20400 3585
rect 20350 3535 20400 3565
rect 20350 3515 20365 3535
rect 20385 3515 20400 3535
rect 20350 3485 20400 3515
rect 20350 3465 20365 3485
rect 20385 3465 20400 3485
rect 20350 3435 20400 3465
rect 20350 3415 20365 3435
rect 20385 3415 20400 3435
rect 20350 3385 20400 3415
rect 20350 3365 20365 3385
rect 20385 3365 20400 3385
rect 20350 3335 20400 3365
rect 20350 3315 20365 3335
rect 20385 3315 20400 3335
rect 20350 3300 20400 3315
rect -600 3235 -350 3250
rect -600 3215 -585 3235
rect -565 3215 -535 3235
rect -515 3215 -485 3235
rect -465 3215 -435 3235
rect -415 3215 -385 3235
rect -365 3215 -350 3235
rect -600 3200 -350 3215
rect -300 3235 -50 3250
rect -300 3215 -285 3235
rect -265 3215 -235 3235
rect -215 3215 -185 3235
rect -165 3215 -135 3235
rect -115 3215 -85 3235
rect -65 3215 -50 3235
rect -300 3200 -50 3215
rect 0 3235 250 3250
rect 0 3215 15 3235
rect 35 3215 65 3235
rect 85 3215 115 3235
rect 135 3215 165 3235
rect 185 3215 215 3235
rect 235 3215 250 3235
rect 0 3200 250 3215
rect 300 3235 550 3250
rect 300 3215 315 3235
rect 335 3215 365 3235
rect 385 3215 415 3235
rect 435 3215 465 3235
rect 485 3215 515 3235
rect 535 3215 550 3235
rect 300 3200 550 3215
rect 600 3235 850 3250
rect 600 3215 615 3235
rect 635 3215 665 3235
rect 685 3215 715 3235
rect 735 3215 765 3235
rect 785 3215 815 3235
rect 835 3215 850 3235
rect 600 3200 850 3215
rect 900 3235 1150 3250
rect 900 3215 915 3235
rect 935 3215 965 3235
rect 985 3215 1015 3235
rect 1035 3215 1065 3235
rect 1085 3215 1115 3235
rect 1135 3215 1150 3235
rect 900 3200 1150 3215
rect 1200 3235 1450 3250
rect 1200 3215 1215 3235
rect 1235 3215 1265 3235
rect 1285 3215 1315 3235
rect 1335 3215 1365 3235
rect 1385 3215 1415 3235
rect 1435 3215 1450 3235
rect 1200 3200 1450 3215
rect 1500 3235 1750 3250
rect 1500 3215 1515 3235
rect 1535 3215 1565 3235
rect 1585 3215 1615 3235
rect 1635 3215 1665 3235
rect 1685 3215 1715 3235
rect 1735 3215 1750 3235
rect 1500 3200 1750 3215
rect 1800 3235 2050 3250
rect 1800 3215 1815 3235
rect 1835 3215 1865 3235
rect 1885 3215 1915 3235
rect 1935 3215 1965 3235
rect 1985 3215 2015 3235
rect 2035 3215 2050 3235
rect 1800 3200 2050 3215
rect 2100 3235 2350 3250
rect 2100 3215 2115 3235
rect 2135 3215 2165 3235
rect 2185 3215 2215 3235
rect 2235 3215 2265 3235
rect 2285 3215 2315 3235
rect 2335 3215 2350 3235
rect 2100 3200 2350 3215
rect 2400 3235 2650 3250
rect 2400 3215 2415 3235
rect 2435 3215 2465 3235
rect 2485 3215 2515 3235
rect 2535 3215 2565 3235
rect 2585 3215 2615 3235
rect 2635 3215 2650 3235
rect 2400 3200 2650 3215
rect 2700 3235 2950 3250
rect 2700 3215 2715 3235
rect 2735 3215 2765 3235
rect 2785 3215 2815 3235
rect 2835 3215 2865 3235
rect 2885 3215 2915 3235
rect 2935 3215 2950 3235
rect 2700 3200 2950 3215
rect 3000 3235 3250 3250
rect 3000 3215 3015 3235
rect 3035 3215 3065 3235
rect 3085 3215 3115 3235
rect 3135 3215 3165 3235
rect 3185 3215 3215 3235
rect 3235 3215 3250 3235
rect 3000 3200 3250 3215
rect 3300 3235 3550 3250
rect 3300 3215 3315 3235
rect 3335 3215 3365 3235
rect 3385 3215 3415 3235
rect 3435 3215 3465 3235
rect 3485 3215 3515 3235
rect 3535 3215 3550 3235
rect 3300 3200 3550 3215
rect 3600 3235 3850 3250
rect 3600 3215 3615 3235
rect 3635 3215 3665 3235
rect 3685 3215 3715 3235
rect 3735 3215 3765 3235
rect 3785 3215 3815 3235
rect 3835 3215 3850 3235
rect 3600 3200 3850 3215
rect 3900 3235 4150 3250
rect 3900 3215 3915 3235
rect 3935 3215 3965 3235
rect 3985 3215 4015 3235
rect 4035 3215 4065 3235
rect 4085 3215 4115 3235
rect 4135 3215 4150 3235
rect 3900 3200 4150 3215
rect 4200 3235 4450 3250
rect 4200 3215 4215 3235
rect 4235 3215 4265 3235
rect 4285 3215 4315 3235
rect 4335 3215 4365 3235
rect 4385 3215 4415 3235
rect 4435 3215 4450 3235
rect 4200 3200 4450 3215
rect 4500 3235 4750 3250
rect 4500 3215 4515 3235
rect 4535 3215 4565 3235
rect 4585 3215 4615 3235
rect 4635 3215 4665 3235
rect 4685 3215 4715 3235
rect 4735 3215 4750 3235
rect 4500 3200 4750 3215
rect 4800 3235 5050 3250
rect 4800 3215 4815 3235
rect 4835 3215 4865 3235
rect 4885 3215 4915 3235
rect 4935 3215 4965 3235
rect 4985 3215 5015 3235
rect 5035 3215 5050 3235
rect 4800 3200 5050 3215
rect 5100 3235 5350 3250
rect 5100 3215 5115 3235
rect 5135 3215 5165 3235
rect 5185 3215 5215 3235
rect 5235 3215 5265 3235
rect 5285 3215 5315 3235
rect 5335 3215 5350 3235
rect 5100 3200 5350 3215
rect 5400 3235 5650 3250
rect 5400 3215 5415 3235
rect 5435 3215 5465 3235
rect 5485 3215 5515 3235
rect 5535 3215 5565 3235
rect 5585 3215 5615 3235
rect 5635 3215 5650 3235
rect 5400 3200 5650 3215
rect 5700 3235 5950 3250
rect 5700 3215 5715 3235
rect 5735 3215 5765 3235
rect 5785 3215 5815 3235
rect 5835 3215 5865 3235
rect 5885 3215 5915 3235
rect 5935 3215 5950 3235
rect 5700 3200 5950 3215
rect 6000 3235 6250 3250
rect 6000 3215 6015 3235
rect 6035 3215 6065 3235
rect 6085 3215 6115 3235
rect 6135 3215 6165 3235
rect 6185 3215 6215 3235
rect 6235 3215 6250 3235
rect 6000 3200 6250 3215
rect 6300 3235 6550 3250
rect 6300 3215 6315 3235
rect 6335 3215 6365 3235
rect 6385 3215 6415 3235
rect 6435 3215 6465 3235
rect 6485 3215 6515 3235
rect 6535 3215 6550 3235
rect 6300 3200 6550 3215
rect 6600 3235 6850 3250
rect 6600 3215 6615 3235
rect 6635 3215 6665 3235
rect 6685 3215 6715 3235
rect 6735 3215 6765 3235
rect 6785 3215 6815 3235
rect 6835 3215 6850 3235
rect 6600 3200 6850 3215
rect 6900 3235 7150 3250
rect 6900 3215 6915 3235
rect 6935 3215 6965 3235
rect 6985 3215 7015 3235
rect 7035 3215 7065 3235
rect 7085 3215 7115 3235
rect 7135 3215 7150 3235
rect 6900 3200 7150 3215
rect 7200 3235 7450 3250
rect 7200 3215 7215 3235
rect 7235 3215 7265 3235
rect 7285 3215 7315 3235
rect 7335 3215 7365 3235
rect 7385 3215 7415 3235
rect 7435 3215 7450 3235
rect 7200 3200 7450 3215
rect 7500 3235 7750 3250
rect 7500 3215 7515 3235
rect 7535 3215 7565 3235
rect 7585 3215 7615 3235
rect 7635 3215 7665 3235
rect 7685 3215 7715 3235
rect 7735 3215 7750 3235
rect 7500 3200 7750 3215
rect 7800 3235 8050 3250
rect 7800 3215 7815 3235
rect 7835 3215 7865 3235
rect 7885 3215 7915 3235
rect 7935 3215 7965 3235
rect 7985 3215 8015 3235
rect 8035 3215 8050 3235
rect 7800 3200 8050 3215
rect 8100 3235 8350 3250
rect 8100 3215 8115 3235
rect 8135 3215 8165 3235
rect 8185 3215 8215 3235
rect 8235 3215 8265 3235
rect 8285 3215 8315 3235
rect 8335 3215 8350 3235
rect 8100 3200 8350 3215
rect 8400 3235 10750 3250
rect 8400 3215 8415 3235
rect 8435 3215 8465 3235
rect 8485 3215 8515 3235
rect 8535 3215 8565 3235
rect 8585 3215 8615 3235
rect 8635 3215 8715 3235
rect 8735 3215 8765 3235
rect 8785 3215 8815 3235
rect 8835 3215 8865 3235
rect 8885 3215 8915 3235
rect 8935 3215 9015 3235
rect 9035 3215 9065 3235
rect 9085 3215 9115 3235
rect 9135 3215 9165 3235
rect 9185 3215 9215 3235
rect 9235 3215 9315 3235
rect 9335 3215 9365 3235
rect 9385 3215 9415 3235
rect 9435 3215 9465 3235
rect 9485 3215 9515 3235
rect 9535 3215 9615 3235
rect 9635 3215 9665 3235
rect 9685 3215 9715 3235
rect 9735 3215 9765 3235
rect 9785 3215 9815 3235
rect 9835 3215 9915 3235
rect 9935 3215 9965 3235
rect 9985 3215 10015 3235
rect 10035 3215 10065 3235
rect 10085 3215 10115 3235
rect 10135 3215 10215 3235
rect 10235 3215 10265 3235
rect 10285 3215 10315 3235
rect 10335 3215 10365 3235
rect 10385 3215 10415 3235
rect 10435 3215 10515 3235
rect 10535 3215 10565 3235
rect 10585 3215 10615 3235
rect 10635 3215 10665 3235
rect 10685 3215 10715 3235
rect 10735 3215 10750 3235
rect 8400 3200 10750 3215
rect 10800 3235 11050 3250
rect 10800 3215 10815 3235
rect 10835 3215 10865 3235
rect 10885 3215 10915 3235
rect 10935 3215 10965 3235
rect 10985 3215 11015 3235
rect 11035 3215 11050 3235
rect 10800 3200 11050 3215
rect 11100 3235 11350 3250
rect 11100 3215 11115 3235
rect 11135 3215 11165 3235
rect 11185 3215 11215 3235
rect 11235 3215 11265 3235
rect 11285 3215 11315 3235
rect 11335 3215 11350 3235
rect 11100 3200 11350 3215
rect 11400 3235 11650 3250
rect 11400 3215 11415 3235
rect 11435 3215 11465 3235
rect 11485 3215 11515 3235
rect 11535 3215 11565 3235
rect 11585 3215 11615 3235
rect 11635 3215 11650 3235
rect 11400 3200 11650 3215
rect 11700 3235 11950 3250
rect 11700 3215 11715 3235
rect 11735 3215 11765 3235
rect 11785 3215 11815 3235
rect 11835 3215 11865 3235
rect 11885 3215 11915 3235
rect 11935 3215 11950 3235
rect 11700 3200 11950 3215
rect 12000 3235 12250 3250
rect 12000 3215 12015 3235
rect 12035 3215 12065 3235
rect 12085 3215 12115 3235
rect 12135 3215 12165 3235
rect 12185 3215 12215 3235
rect 12235 3215 12250 3235
rect 12000 3200 12250 3215
rect 12300 3235 12550 3250
rect 12300 3215 12315 3235
rect 12335 3215 12365 3235
rect 12385 3215 12415 3235
rect 12435 3215 12465 3235
rect 12485 3215 12515 3235
rect 12535 3215 12550 3235
rect 12300 3200 12550 3215
rect 12600 3235 12850 3250
rect 12600 3215 12615 3235
rect 12635 3215 12665 3235
rect 12685 3215 12715 3235
rect 12735 3215 12765 3235
rect 12785 3215 12815 3235
rect 12835 3215 12850 3235
rect 12600 3200 12850 3215
rect 12900 3235 13150 3250
rect 12900 3215 12915 3235
rect 12935 3215 12965 3235
rect 12985 3215 13015 3235
rect 13035 3215 13065 3235
rect 13085 3215 13115 3235
rect 13135 3215 13150 3235
rect 12900 3200 13150 3215
rect 13200 3235 13450 3250
rect 13200 3215 13215 3235
rect 13235 3215 13265 3235
rect 13285 3215 13315 3235
rect 13335 3215 13365 3235
rect 13385 3215 13415 3235
rect 13435 3215 13450 3235
rect 13200 3200 13450 3215
rect 13500 3235 13750 3250
rect 13500 3215 13515 3235
rect 13535 3215 13565 3235
rect 13585 3215 13615 3235
rect 13635 3215 13665 3235
rect 13685 3215 13715 3235
rect 13735 3215 13750 3235
rect 13500 3200 13750 3215
rect 13800 3235 14050 3250
rect 13800 3215 13815 3235
rect 13835 3215 13865 3235
rect 13885 3215 13915 3235
rect 13935 3215 13965 3235
rect 13985 3215 14015 3235
rect 14035 3215 14050 3235
rect 13800 3200 14050 3215
rect 14100 3235 14350 3250
rect 14100 3215 14115 3235
rect 14135 3215 14165 3235
rect 14185 3215 14215 3235
rect 14235 3215 14265 3235
rect 14285 3215 14315 3235
rect 14335 3215 14350 3235
rect 14100 3200 14350 3215
rect 14400 3235 14650 3250
rect 14400 3215 14415 3235
rect 14435 3215 14465 3235
rect 14485 3215 14515 3235
rect 14535 3215 14565 3235
rect 14585 3215 14615 3235
rect 14635 3215 14650 3235
rect 14400 3200 14650 3215
rect 14700 3235 14950 3250
rect 14700 3215 14715 3235
rect 14735 3215 14765 3235
rect 14785 3215 14815 3235
rect 14835 3215 14865 3235
rect 14885 3215 14915 3235
rect 14935 3215 14950 3235
rect 14700 3200 14950 3215
rect 15000 3235 15250 3250
rect 15000 3215 15015 3235
rect 15035 3215 15065 3235
rect 15085 3215 15115 3235
rect 15135 3215 15165 3235
rect 15185 3215 15215 3235
rect 15235 3215 15250 3235
rect 15000 3200 15250 3215
rect 15300 3235 15550 3250
rect 15300 3215 15315 3235
rect 15335 3215 15365 3235
rect 15385 3215 15415 3235
rect 15435 3215 15465 3235
rect 15485 3215 15515 3235
rect 15535 3215 15550 3235
rect 15300 3200 15550 3215
rect 15600 3235 15850 3250
rect 15600 3215 15615 3235
rect 15635 3215 15665 3235
rect 15685 3215 15715 3235
rect 15735 3215 15765 3235
rect 15785 3215 15815 3235
rect 15835 3215 15850 3235
rect 15600 3200 15850 3215
rect 15900 3235 16150 3250
rect 15900 3215 15915 3235
rect 15935 3215 15965 3235
rect 15985 3215 16015 3235
rect 16035 3215 16065 3235
rect 16085 3215 16115 3235
rect 16135 3215 16150 3235
rect 15900 3200 16150 3215
rect 16200 3235 16450 3250
rect 16200 3215 16215 3235
rect 16235 3215 16265 3235
rect 16285 3215 16315 3235
rect 16335 3215 16365 3235
rect 16385 3215 16415 3235
rect 16435 3215 16450 3235
rect 16200 3200 16450 3215
rect 16500 3235 16750 3250
rect 16500 3215 16515 3235
rect 16535 3215 16565 3235
rect 16585 3215 16615 3235
rect 16635 3215 16665 3235
rect 16685 3215 16715 3235
rect 16735 3215 16750 3235
rect 16500 3200 16750 3215
rect 16800 3235 17050 3250
rect 16800 3215 16815 3235
rect 16835 3215 16865 3235
rect 16885 3215 16915 3235
rect 16935 3215 16965 3235
rect 16985 3215 17015 3235
rect 17035 3215 17050 3235
rect 16800 3200 17050 3215
rect 17100 3235 17350 3250
rect 17100 3215 17115 3235
rect 17135 3215 17165 3235
rect 17185 3215 17215 3235
rect 17235 3215 17265 3235
rect 17285 3215 17315 3235
rect 17335 3215 17350 3235
rect 17100 3200 17350 3215
rect 17400 3235 17650 3250
rect 17400 3215 17415 3235
rect 17435 3215 17465 3235
rect 17485 3215 17515 3235
rect 17535 3215 17565 3235
rect 17585 3215 17615 3235
rect 17635 3215 17650 3235
rect 17400 3200 17650 3215
rect 17700 3235 17950 3250
rect 17700 3215 17715 3235
rect 17735 3215 17765 3235
rect 17785 3215 17815 3235
rect 17835 3215 17865 3235
rect 17885 3215 17915 3235
rect 17935 3215 17950 3235
rect 17700 3200 17950 3215
rect 18000 3235 18250 3250
rect 18000 3215 18015 3235
rect 18035 3215 18065 3235
rect 18085 3215 18115 3235
rect 18135 3215 18165 3235
rect 18185 3215 18215 3235
rect 18235 3215 18250 3235
rect 18000 3200 18250 3215
rect 18300 3235 18550 3250
rect 18300 3215 18315 3235
rect 18335 3215 18365 3235
rect 18385 3215 18415 3235
rect 18435 3215 18465 3235
rect 18485 3215 18515 3235
rect 18535 3215 18550 3235
rect 18300 3200 18550 3215
rect 18600 3235 18850 3250
rect 18600 3215 18615 3235
rect 18635 3215 18665 3235
rect 18685 3215 18715 3235
rect 18735 3215 18765 3235
rect 18785 3215 18815 3235
rect 18835 3215 18850 3235
rect 18600 3200 18850 3215
rect 18900 3235 19150 3250
rect 18900 3215 18915 3235
rect 18935 3215 18965 3235
rect 18985 3215 19015 3235
rect 19035 3215 19065 3235
rect 19085 3215 19115 3235
rect 19135 3215 19150 3235
rect 18900 3200 19150 3215
rect 19200 3235 19450 3250
rect 19200 3215 19215 3235
rect 19235 3215 19265 3235
rect 19285 3215 19315 3235
rect 19335 3215 19365 3235
rect 19385 3215 19415 3235
rect 19435 3215 19450 3235
rect 19200 3200 19450 3215
rect 19500 3235 19750 3250
rect 19500 3215 19515 3235
rect 19535 3215 19565 3235
rect 19585 3215 19615 3235
rect 19635 3215 19665 3235
rect 19685 3215 19715 3235
rect 19735 3215 19750 3235
rect 19500 3200 19750 3215
rect 19800 3235 20050 3250
rect 19800 3215 19815 3235
rect 19835 3215 19865 3235
rect 19885 3215 19915 3235
rect 19935 3215 19965 3235
rect 19985 3215 20015 3235
rect 20035 3215 20050 3235
rect 19800 3200 20050 3215
rect 20100 3235 20350 3250
rect 20100 3215 20115 3235
rect 20135 3215 20165 3235
rect 20185 3215 20215 3235
rect 20235 3215 20265 3235
rect 20285 3215 20315 3235
rect 20335 3215 20350 3235
rect 20100 3200 20350 3215
rect -650 3135 -600 3150
rect -650 3115 -635 3135
rect -615 3115 -600 3135
rect -650 3085 -600 3115
rect -650 3065 -635 3085
rect -615 3065 -600 3085
rect -650 3035 -600 3065
rect -650 3015 -635 3035
rect -615 3015 -600 3035
rect -650 2985 -600 3015
rect -650 2965 -635 2985
rect -615 2965 -600 2985
rect -650 2935 -600 2965
rect -650 2915 -635 2935
rect -615 2915 -600 2935
rect -650 2885 -600 2915
rect -650 2865 -635 2885
rect -615 2865 -600 2885
rect -650 2835 -600 2865
rect -650 2815 -635 2835
rect -615 2815 -600 2835
rect -650 2785 -600 2815
rect -650 2765 -635 2785
rect -615 2765 -600 2785
rect -650 2735 -600 2765
rect -650 2715 -635 2735
rect -615 2715 -600 2735
rect -650 2685 -600 2715
rect -650 2665 -635 2685
rect -615 2665 -600 2685
rect -650 2650 -600 2665
rect -500 3135 -450 3150
rect -500 3115 -485 3135
rect -465 3115 -450 3135
rect -500 3085 -450 3115
rect -500 3065 -485 3085
rect -465 3065 -450 3085
rect -500 3035 -450 3065
rect -500 3015 -485 3035
rect -465 3015 -450 3035
rect -500 2985 -450 3015
rect -500 2965 -485 2985
rect -465 2965 -450 2985
rect -500 2935 -450 2965
rect -500 2915 -485 2935
rect -465 2915 -450 2935
rect -500 2885 -450 2915
rect -500 2865 -485 2885
rect -465 2865 -450 2885
rect -500 2835 -450 2865
rect -500 2815 -485 2835
rect -465 2815 -450 2835
rect -500 2785 -450 2815
rect -500 2765 -485 2785
rect -465 2765 -450 2785
rect -500 2735 -450 2765
rect -500 2715 -485 2735
rect -465 2715 -450 2735
rect -500 2685 -450 2715
rect -500 2665 -485 2685
rect -465 2665 -450 2685
rect -500 2650 -450 2665
rect -350 3135 -300 3150
rect -350 3115 -335 3135
rect -315 3115 -300 3135
rect -350 3085 -300 3115
rect -350 3065 -335 3085
rect -315 3065 -300 3085
rect -350 3035 -300 3065
rect -350 3015 -335 3035
rect -315 3015 -300 3035
rect -350 2985 -300 3015
rect -350 2965 -335 2985
rect -315 2965 -300 2985
rect -350 2935 -300 2965
rect -350 2915 -335 2935
rect -315 2915 -300 2935
rect -350 2885 -300 2915
rect -350 2865 -335 2885
rect -315 2865 -300 2885
rect -350 2835 -300 2865
rect -350 2815 -335 2835
rect -315 2815 -300 2835
rect -350 2785 -300 2815
rect -350 2765 -335 2785
rect -315 2765 -300 2785
rect -350 2735 -300 2765
rect -350 2715 -335 2735
rect -315 2715 -300 2735
rect -350 2685 -300 2715
rect -350 2665 -335 2685
rect -315 2665 -300 2685
rect -350 2650 -300 2665
rect -200 3135 -150 3150
rect -200 3115 -185 3135
rect -165 3115 -150 3135
rect -200 3085 -150 3115
rect -200 3065 -185 3085
rect -165 3065 -150 3085
rect -200 3035 -150 3065
rect -200 3015 -185 3035
rect -165 3015 -150 3035
rect -200 2985 -150 3015
rect -200 2965 -185 2985
rect -165 2965 -150 2985
rect -200 2935 -150 2965
rect -200 2915 -185 2935
rect -165 2915 -150 2935
rect -200 2885 -150 2915
rect -200 2865 -185 2885
rect -165 2865 -150 2885
rect -200 2835 -150 2865
rect -200 2815 -185 2835
rect -165 2815 -150 2835
rect -200 2785 -150 2815
rect -200 2765 -185 2785
rect -165 2765 -150 2785
rect -200 2735 -150 2765
rect -200 2715 -185 2735
rect -165 2715 -150 2735
rect -200 2685 -150 2715
rect -200 2665 -185 2685
rect -165 2665 -150 2685
rect -200 2650 -150 2665
rect -50 3135 0 3150
rect -50 3115 -35 3135
rect -15 3115 0 3135
rect -50 3085 0 3115
rect -50 3065 -35 3085
rect -15 3065 0 3085
rect -50 3035 0 3065
rect -50 3015 -35 3035
rect -15 3015 0 3035
rect -50 2985 0 3015
rect -50 2965 -35 2985
rect -15 2965 0 2985
rect -50 2935 0 2965
rect -50 2915 -35 2935
rect -15 2915 0 2935
rect -50 2885 0 2915
rect -50 2865 -35 2885
rect -15 2865 0 2885
rect -50 2835 0 2865
rect -50 2815 -35 2835
rect -15 2815 0 2835
rect -50 2785 0 2815
rect -50 2765 -35 2785
rect -15 2765 0 2785
rect -50 2735 0 2765
rect -50 2715 -35 2735
rect -15 2715 0 2735
rect -50 2685 0 2715
rect -50 2665 -35 2685
rect -15 2665 0 2685
rect -50 2650 0 2665
rect 550 3135 600 3150
rect 550 3115 565 3135
rect 585 3115 600 3135
rect 550 3085 600 3115
rect 550 3065 565 3085
rect 585 3065 600 3085
rect 550 3035 600 3065
rect 550 3015 565 3035
rect 585 3015 600 3035
rect 550 2985 600 3015
rect 550 2965 565 2985
rect 585 2965 600 2985
rect 550 2935 600 2965
rect 550 2915 565 2935
rect 585 2915 600 2935
rect 550 2885 600 2915
rect 550 2865 565 2885
rect 585 2865 600 2885
rect 550 2835 600 2865
rect 550 2815 565 2835
rect 585 2815 600 2835
rect 550 2785 600 2815
rect 550 2765 565 2785
rect 585 2765 600 2785
rect 550 2735 600 2765
rect 550 2715 565 2735
rect 585 2715 600 2735
rect 550 2685 600 2715
rect 550 2665 565 2685
rect 585 2665 600 2685
rect 550 2650 600 2665
rect 700 3135 750 3150
rect 700 3115 715 3135
rect 735 3115 750 3135
rect 700 3085 750 3115
rect 700 3065 715 3085
rect 735 3065 750 3085
rect 700 3035 750 3065
rect 700 3015 715 3035
rect 735 3015 750 3035
rect 700 2985 750 3015
rect 700 2965 715 2985
rect 735 2965 750 2985
rect 700 2935 750 2965
rect 700 2915 715 2935
rect 735 2915 750 2935
rect 700 2885 750 2915
rect 700 2865 715 2885
rect 735 2865 750 2885
rect 700 2835 750 2865
rect 700 2815 715 2835
rect 735 2815 750 2835
rect 700 2785 750 2815
rect 700 2765 715 2785
rect 735 2765 750 2785
rect 700 2735 750 2765
rect 700 2715 715 2735
rect 735 2715 750 2735
rect 700 2685 750 2715
rect 700 2665 715 2685
rect 735 2665 750 2685
rect 700 2650 750 2665
rect 850 3135 900 3150
rect 850 3115 865 3135
rect 885 3115 900 3135
rect 850 3085 900 3115
rect 850 3065 865 3085
rect 885 3065 900 3085
rect 850 3035 900 3065
rect 850 3015 865 3035
rect 885 3015 900 3035
rect 850 2985 900 3015
rect 850 2965 865 2985
rect 885 2965 900 2985
rect 850 2935 900 2965
rect 850 2915 865 2935
rect 885 2915 900 2935
rect 850 2885 900 2915
rect 850 2865 865 2885
rect 885 2865 900 2885
rect 850 2835 900 2865
rect 850 2815 865 2835
rect 885 2815 900 2835
rect 850 2785 900 2815
rect 850 2765 865 2785
rect 885 2765 900 2785
rect 850 2735 900 2765
rect 850 2715 865 2735
rect 885 2715 900 2735
rect 850 2685 900 2715
rect 850 2665 865 2685
rect 885 2665 900 2685
rect 850 2650 900 2665
rect 1000 3135 1050 3150
rect 1000 3115 1015 3135
rect 1035 3115 1050 3135
rect 1000 3085 1050 3115
rect 1000 3065 1015 3085
rect 1035 3065 1050 3085
rect 1000 3035 1050 3065
rect 1000 3015 1015 3035
rect 1035 3015 1050 3035
rect 1000 2985 1050 3015
rect 1000 2965 1015 2985
rect 1035 2965 1050 2985
rect 1000 2935 1050 2965
rect 1000 2915 1015 2935
rect 1035 2915 1050 2935
rect 1000 2885 1050 2915
rect 1000 2865 1015 2885
rect 1035 2865 1050 2885
rect 1000 2835 1050 2865
rect 1000 2815 1015 2835
rect 1035 2815 1050 2835
rect 1000 2785 1050 2815
rect 1000 2765 1015 2785
rect 1035 2765 1050 2785
rect 1000 2735 1050 2765
rect 1000 2715 1015 2735
rect 1035 2715 1050 2735
rect 1000 2685 1050 2715
rect 1000 2665 1015 2685
rect 1035 2665 1050 2685
rect 1000 2650 1050 2665
rect 1150 3135 1200 3150
rect 1150 3115 1165 3135
rect 1185 3115 1200 3135
rect 1150 3085 1200 3115
rect 1150 3065 1165 3085
rect 1185 3065 1200 3085
rect 1150 3035 1200 3065
rect 1150 3015 1165 3035
rect 1185 3015 1200 3035
rect 1150 2985 1200 3015
rect 1150 2965 1165 2985
rect 1185 2965 1200 2985
rect 1150 2935 1200 2965
rect 1150 2915 1165 2935
rect 1185 2915 1200 2935
rect 1150 2885 1200 2915
rect 1150 2865 1165 2885
rect 1185 2865 1200 2885
rect 1150 2835 1200 2865
rect 1150 2815 1165 2835
rect 1185 2815 1200 2835
rect 1150 2785 1200 2815
rect 1150 2765 1165 2785
rect 1185 2765 1200 2785
rect 1150 2735 1200 2765
rect 1150 2715 1165 2735
rect 1185 2715 1200 2735
rect 1150 2685 1200 2715
rect 1150 2665 1165 2685
rect 1185 2665 1200 2685
rect 1150 2650 1200 2665
rect 1300 3135 1350 3150
rect 1300 3115 1315 3135
rect 1335 3115 1350 3135
rect 1300 3085 1350 3115
rect 1300 3065 1315 3085
rect 1335 3065 1350 3085
rect 1300 3035 1350 3065
rect 1300 3015 1315 3035
rect 1335 3015 1350 3035
rect 1300 2985 1350 3015
rect 1300 2965 1315 2985
rect 1335 2965 1350 2985
rect 1300 2935 1350 2965
rect 1300 2915 1315 2935
rect 1335 2915 1350 2935
rect 1300 2885 1350 2915
rect 1300 2865 1315 2885
rect 1335 2865 1350 2885
rect 1300 2835 1350 2865
rect 1300 2815 1315 2835
rect 1335 2815 1350 2835
rect 1300 2785 1350 2815
rect 1300 2765 1315 2785
rect 1335 2765 1350 2785
rect 1300 2735 1350 2765
rect 1300 2715 1315 2735
rect 1335 2715 1350 2735
rect 1300 2685 1350 2715
rect 1300 2665 1315 2685
rect 1335 2665 1350 2685
rect 1300 2650 1350 2665
rect 1450 3135 1500 3150
rect 1450 3115 1465 3135
rect 1485 3115 1500 3135
rect 1450 3085 1500 3115
rect 1450 3065 1465 3085
rect 1485 3065 1500 3085
rect 1450 3035 1500 3065
rect 1450 3015 1465 3035
rect 1485 3015 1500 3035
rect 1450 2985 1500 3015
rect 1450 2965 1465 2985
rect 1485 2965 1500 2985
rect 1450 2935 1500 2965
rect 1450 2915 1465 2935
rect 1485 2915 1500 2935
rect 1450 2885 1500 2915
rect 1450 2865 1465 2885
rect 1485 2865 1500 2885
rect 1450 2835 1500 2865
rect 1450 2815 1465 2835
rect 1485 2815 1500 2835
rect 1450 2785 1500 2815
rect 1450 2765 1465 2785
rect 1485 2765 1500 2785
rect 1450 2735 1500 2765
rect 1450 2715 1465 2735
rect 1485 2715 1500 2735
rect 1450 2685 1500 2715
rect 1450 2665 1465 2685
rect 1485 2665 1500 2685
rect 1450 2650 1500 2665
rect 1600 3135 1650 3150
rect 1600 3115 1615 3135
rect 1635 3115 1650 3135
rect 1600 3085 1650 3115
rect 1600 3065 1615 3085
rect 1635 3065 1650 3085
rect 1600 3035 1650 3065
rect 1600 3015 1615 3035
rect 1635 3015 1650 3035
rect 1600 2985 1650 3015
rect 1600 2965 1615 2985
rect 1635 2965 1650 2985
rect 1600 2935 1650 2965
rect 1600 2915 1615 2935
rect 1635 2915 1650 2935
rect 1600 2885 1650 2915
rect 1600 2865 1615 2885
rect 1635 2865 1650 2885
rect 1600 2835 1650 2865
rect 1600 2815 1615 2835
rect 1635 2815 1650 2835
rect 1600 2785 1650 2815
rect 1600 2765 1615 2785
rect 1635 2765 1650 2785
rect 1600 2735 1650 2765
rect 1600 2715 1615 2735
rect 1635 2715 1650 2735
rect 1600 2685 1650 2715
rect 1600 2665 1615 2685
rect 1635 2665 1650 2685
rect 1600 2650 1650 2665
rect 1750 3135 1800 3150
rect 1750 3115 1765 3135
rect 1785 3115 1800 3135
rect 1750 3085 1800 3115
rect 1750 3065 1765 3085
rect 1785 3065 1800 3085
rect 1750 3035 1800 3065
rect 1750 3015 1765 3035
rect 1785 3015 1800 3035
rect 1750 2985 1800 3015
rect 1750 2965 1765 2985
rect 1785 2965 1800 2985
rect 1750 2935 1800 2965
rect 1750 2915 1765 2935
rect 1785 2915 1800 2935
rect 1750 2885 1800 2915
rect 1750 2865 1765 2885
rect 1785 2865 1800 2885
rect 1750 2835 1800 2865
rect 1750 2815 1765 2835
rect 1785 2815 1800 2835
rect 1750 2785 1800 2815
rect 1750 2765 1765 2785
rect 1785 2765 1800 2785
rect 1750 2735 1800 2765
rect 1750 2715 1765 2735
rect 1785 2715 1800 2735
rect 1750 2685 1800 2715
rect 1750 2665 1765 2685
rect 1785 2665 1800 2685
rect 1750 2650 1800 2665
rect 1900 3135 1950 3150
rect 1900 3115 1915 3135
rect 1935 3115 1950 3135
rect 1900 3085 1950 3115
rect 1900 3065 1915 3085
rect 1935 3065 1950 3085
rect 1900 3035 1950 3065
rect 1900 3015 1915 3035
rect 1935 3015 1950 3035
rect 1900 2985 1950 3015
rect 1900 2965 1915 2985
rect 1935 2965 1950 2985
rect 1900 2935 1950 2965
rect 1900 2915 1915 2935
rect 1935 2915 1950 2935
rect 1900 2885 1950 2915
rect 1900 2865 1915 2885
rect 1935 2865 1950 2885
rect 1900 2835 1950 2865
rect 1900 2815 1915 2835
rect 1935 2815 1950 2835
rect 1900 2785 1950 2815
rect 1900 2765 1915 2785
rect 1935 2765 1950 2785
rect 1900 2735 1950 2765
rect 1900 2715 1915 2735
rect 1935 2715 1950 2735
rect 1900 2685 1950 2715
rect 1900 2665 1915 2685
rect 1935 2665 1950 2685
rect 1900 2650 1950 2665
rect 2050 3135 2100 3150
rect 2050 3115 2065 3135
rect 2085 3115 2100 3135
rect 2050 3085 2100 3115
rect 2050 3065 2065 3085
rect 2085 3065 2100 3085
rect 2050 3035 2100 3065
rect 2050 3015 2065 3035
rect 2085 3015 2100 3035
rect 2050 2985 2100 3015
rect 2050 2965 2065 2985
rect 2085 2965 2100 2985
rect 2050 2935 2100 2965
rect 2050 2915 2065 2935
rect 2085 2915 2100 2935
rect 2050 2885 2100 2915
rect 2050 2865 2065 2885
rect 2085 2865 2100 2885
rect 2050 2835 2100 2865
rect 2050 2815 2065 2835
rect 2085 2815 2100 2835
rect 2050 2785 2100 2815
rect 2050 2765 2065 2785
rect 2085 2765 2100 2785
rect 2050 2735 2100 2765
rect 2050 2715 2065 2735
rect 2085 2715 2100 2735
rect 2050 2685 2100 2715
rect 2050 2665 2065 2685
rect 2085 2665 2100 2685
rect 2050 2650 2100 2665
rect 2200 3135 2250 3150
rect 2200 3115 2215 3135
rect 2235 3115 2250 3135
rect 2200 3085 2250 3115
rect 2200 3065 2215 3085
rect 2235 3065 2250 3085
rect 2200 3035 2250 3065
rect 2200 3015 2215 3035
rect 2235 3015 2250 3035
rect 2200 2985 2250 3015
rect 2200 2965 2215 2985
rect 2235 2965 2250 2985
rect 2200 2935 2250 2965
rect 2200 2915 2215 2935
rect 2235 2915 2250 2935
rect 2200 2885 2250 2915
rect 2200 2865 2215 2885
rect 2235 2865 2250 2885
rect 2200 2835 2250 2865
rect 2200 2815 2215 2835
rect 2235 2815 2250 2835
rect 2200 2785 2250 2815
rect 2200 2765 2215 2785
rect 2235 2765 2250 2785
rect 2200 2735 2250 2765
rect 2200 2715 2215 2735
rect 2235 2715 2250 2735
rect 2200 2685 2250 2715
rect 2200 2665 2215 2685
rect 2235 2665 2250 2685
rect 2200 2650 2250 2665
rect 2350 3135 2400 3150
rect 2350 3115 2365 3135
rect 2385 3115 2400 3135
rect 2350 3085 2400 3115
rect 2350 3065 2365 3085
rect 2385 3065 2400 3085
rect 2350 3035 2400 3065
rect 2350 3015 2365 3035
rect 2385 3015 2400 3035
rect 2350 2985 2400 3015
rect 2350 2965 2365 2985
rect 2385 2965 2400 2985
rect 2350 2935 2400 2965
rect 2350 2915 2365 2935
rect 2385 2915 2400 2935
rect 2350 2885 2400 2915
rect 2350 2865 2365 2885
rect 2385 2865 2400 2885
rect 2350 2835 2400 2865
rect 2350 2815 2365 2835
rect 2385 2815 2400 2835
rect 2350 2785 2400 2815
rect 2350 2765 2365 2785
rect 2385 2765 2400 2785
rect 2350 2735 2400 2765
rect 2350 2715 2365 2735
rect 2385 2715 2400 2735
rect 2350 2685 2400 2715
rect 2350 2665 2365 2685
rect 2385 2665 2400 2685
rect 2350 2650 2400 2665
rect 2500 3135 2550 3150
rect 2500 3115 2515 3135
rect 2535 3115 2550 3135
rect 2500 3085 2550 3115
rect 2500 3065 2515 3085
rect 2535 3065 2550 3085
rect 2500 3035 2550 3065
rect 2500 3015 2515 3035
rect 2535 3015 2550 3035
rect 2500 2985 2550 3015
rect 2500 2965 2515 2985
rect 2535 2965 2550 2985
rect 2500 2935 2550 2965
rect 2500 2915 2515 2935
rect 2535 2915 2550 2935
rect 2500 2885 2550 2915
rect 2500 2865 2515 2885
rect 2535 2865 2550 2885
rect 2500 2835 2550 2865
rect 2500 2815 2515 2835
rect 2535 2815 2550 2835
rect 2500 2785 2550 2815
rect 2500 2765 2515 2785
rect 2535 2765 2550 2785
rect 2500 2735 2550 2765
rect 2500 2715 2515 2735
rect 2535 2715 2550 2735
rect 2500 2685 2550 2715
rect 2500 2665 2515 2685
rect 2535 2665 2550 2685
rect 2500 2650 2550 2665
rect 2650 3135 2700 3150
rect 2650 3115 2665 3135
rect 2685 3115 2700 3135
rect 2650 3085 2700 3115
rect 2650 3065 2665 3085
rect 2685 3065 2700 3085
rect 2650 3035 2700 3065
rect 2650 3015 2665 3035
rect 2685 3015 2700 3035
rect 2650 2985 2700 3015
rect 2650 2965 2665 2985
rect 2685 2965 2700 2985
rect 2650 2935 2700 2965
rect 2650 2915 2665 2935
rect 2685 2915 2700 2935
rect 2650 2885 2700 2915
rect 2650 2865 2665 2885
rect 2685 2865 2700 2885
rect 2650 2835 2700 2865
rect 2650 2815 2665 2835
rect 2685 2815 2700 2835
rect 2650 2785 2700 2815
rect 2650 2765 2665 2785
rect 2685 2765 2700 2785
rect 2650 2735 2700 2765
rect 2650 2715 2665 2735
rect 2685 2715 2700 2735
rect 2650 2685 2700 2715
rect 2650 2665 2665 2685
rect 2685 2665 2700 2685
rect 2650 2650 2700 2665
rect 2800 3135 2850 3150
rect 2800 3115 2815 3135
rect 2835 3115 2850 3135
rect 2800 3085 2850 3115
rect 2800 3065 2815 3085
rect 2835 3065 2850 3085
rect 2800 3035 2850 3065
rect 2800 3015 2815 3035
rect 2835 3015 2850 3035
rect 2800 2985 2850 3015
rect 2800 2965 2815 2985
rect 2835 2965 2850 2985
rect 2800 2935 2850 2965
rect 2800 2915 2815 2935
rect 2835 2915 2850 2935
rect 2800 2885 2850 2915
rect 2800 2865 2815 2885
rect 2835 2865 2850 2885
rect 2800 2835 2850 2865
rect 2800 2815 2815 2835
rect 2835 2815 2850 2835
rect 2800 2785 2850 2815
rect 2800 2765 2815 2785
rect 2835 2765 2850 2785
rect 2800 2735 2850 2765
rect 2800 2715 2815 2735
rect 2835 2715 2850 2735
rect 2800 2685 2850 2715
rect 2800 2665 2815 2685
rect 2835 2665 2850 2685
rect 2800 2650 2850 2665
rect 2950 3135 3000 3150
rect 2950 3115 2965 3135
rect 2985 3115 3000 3135
rect 2950 3085 3000 3115
rect 2950 3065 2965 3085
rect 2985 3065 3000 3085
rect 2950 3035 3000 3065
rect 2950 3015 2965 3035
rect 2985 3015 3000 3035
rect 2950 2985 3000 3015
rect 2950 2965 2965 2985
rect 2985 2965 3000 2985
rect 2950 2935 3000 2965
rect 2950 2915 2965 2935
rect 2985 2915 3000 2935
rect 2950 2885 3000 2915
rect 2950 2865 2965 2885
rect 2985 2865 3000 2885
rect 2950 2835 3000 2865
rect 2950 2815 2965 2835
rect 2985 2815 3000 2835
rect 2950 2785 3000 2815
rect 2950 2765 2965 2785
rect 2985 2765 3000 2785
rect 2950 2735 3000 2765
rect 2950 2715 2965 2735
rect 2985 2715 3000 2735
rect 2950 2685 3000 2715
rect 2950 2665 2965 2685
rect 2985 2665 3000 2685
rect 2950 2650 3000 2665
rect 3100 3135 3150 3150
rect 3100 3115 3115 3135
rect 3135 3115 3150 3135
rect 3100 3085 3150 3115
rect 3100 3065 3115 3085
rect 3135 3065 3150 3085
rect 3100 3035 3150 3065
rect 3100 3015 3115 3035
rect 3135 3015 3150 3035
rect 3100 2985 3150 3015
rect 3100 2965 3115 2985
rect 3135 2965 3150 2985
rect 3100 2935 3150 2965
rect 3100 2915 3115 2935
rect 3135 2915 3150 2935
rect 3100 2885 3150 2915
rect 3100 2865 3115 2885
rect 3135 2865 3150 2885
rect 3100 2835 3150 2865
rect 3100 2815 3115 2835
rect 3135 2815 3150 2835
rect 3100 2785 3150 2815
rect 3100 2765 3115 2785
rect 3135 2765 3150 2785
rect 3100 2735 3150 2765
rect 3100 2715 3115 2735
rect 3135 2715 3150 2735
rect 3100 2685 3150 2715
rect 3100 2665 3115 2685
rect 3135 2665 3150 2685
rect 3100 2650 3150 2665
rect 3250 3135 3300 3150
rect 3250 3115 3265 3135
rect 3285 3115 3300 3135
rect 3250 3085 3300 3115
rect 3250 3065 3265 3085
rect 3285 3065 3300 3085
rect 3250 3035 3300 3065
rect 3250 3015 3265 3035
rect 3285 3015 3300 3035
rect 3250 2985 3300 3015
rect 3250 2965 3265 2985
rect 3285 2965 3300 2985
rect 3250 2935 3300 2965
rect 3250 2915 3265 2935
rect 3285 2915 3300 2935
rect 3250 2885 3300 2915
rect 3250 2865 3265 2885
rect 3285 2865 3300 2885
rect 3250 2835 3300 2865
rect 3250 2815 3265 2835
rect 3285 2815 3300 2835
rect 3250 2785 3300 2815
rect 3250 2765 3265 2785
rect 3285 2765 3300 2785
rect 3250 2735 3300 2765
rect 3250 2715 3265 2735
rect 3285 2715 3300 2735
rect 3250 2685 3300 2715
rect 3250 2665 3265 2685
rect 3285 2665 3300 2685
rect 3250 2650 3300 2665
rect 3400 3135 3450 3150
rect 3400 3115 3415 3135
rect 3435 3115 3450 3135
rect 3400 3085 3450 3115
rect 3400 3065 3415 3085
rect 3435 3065 3450 3085
rect 3400 3035 3450 3065
rect 3400 3015 3415 3035
rect 3435 3015 3450 3035
rect 3400 2985 3450 3015
rect 3400 2965 3415 2985
rect 3435 2965 3450 2985
rect 3400 2935 3450 2965
rect 3400 2915 3415 2935
rect 3435 2915 3450 2935
rect 3400 2885 3450 2915
rect 3400 2865 3415 2885
rect 3435 2865 3450 2885
rect 3400 2835 3450 2865
rect 3400 2815 3415 2835
rect 3435 2815 3450 2835
rect 3400 2785 3450 2815
rect 3400 2765 3415 2785
rect 3435 2765 3450 2785
rect 3400 2735 3450 2765
rect 3400 2715 3415 2735
rect 3435 2715 3450 2735
rect 3400 2685 3450 2715
rect 3400 2665 3415 2685
rect 3435 2665 3450 2685
rect 3400 2650 3450 2665
rect 3550 3135 3600 3150
rect 3550 3115 3565 3135
rect 3585 3115 3600 3135
rect 3550 3085 3600 3115
rect 3550 3065 3565 3085
rect 3585 3065 3600 3085
rect 3550 3035 3600 3065
rect 3550 3015 3565 3035
rect 3585 3015 3600 3035
rect 3550 2985 3600 3015
rect 3550 2965 3565 2985
rect 3585 2965 3600 2985
rect 3550 2935 3600 2965
rect 3550 2915 3565 2935
rect 3585 2915 3600 2935
rect 3550 2885 3600 2915
rect 3550 2865 3565 2885
rect 3585 2865 3600 2885
rect 3550 2835 3600 2865
rect 3550 2815 3565 2835
rect 3585 2815 3600 2835
rect 3550 2785 3600 2815
rect 3550 2765 3565 2785
rect 3585 2765 3600 2785
rect 3550 2735 3600 2765
rect 3550 2715 3565 2735
rect 3585 2715 3600 2735
rect 3550 2685 3600 2715
rect 3550 2665 3565 2685
rect 3585 2665 3600 2685
rect 3550 2650 3600 2665
rect 4150 3135 4200 3150
rect 4150 3115 4165 3135
rect 4185 3115 4200 3135
rect 4150 3085 4200 3115
rect 4150 3065 4165 3085
rect 4185 3065 4200 3085
rect 4150 3035 4200 3065
rect 4150 3015 4165 3035
rect 4185 3015 4200 3035
rect 4150 2985 4200 3015
rect 4150 2965 4165 2985
rect 4185 2965 4200 2985
rect 4150 2935 4200 2965
rect 4150 2915 4165 2935
rect 4185 2915 4200 2935
rect 4150 2885 4200 2915
rect 4150 2865 4165 2885
rect 4185 2865 4200 2885
rect 4150 2835 4200 2865
rect 4150 2815 4165 2835
rect 4185 2815 4200 2835
rect 4150 2785 4200 2815
rect 4150 2765 4165 2785
rect 4185 2765 4200 2785
rect 4150 2735 4200 2765
rect 4150 2715 4165 2735
rect 4185 2715 4200 2735
rect 4150 2685 4200 2715
rect 4150 2665 4165 2685
rect 4185 2665 4200 2685
rect 4150 2650 4200 2665
rect 4750 3135 4800 3150
rect 4750 3115 4765 3135
rect 4785 3115 4800 3135
rect 4750 3085 4800 3115
rect 4750 3065 4765 3085
rect 4785 3065 4800 3085
rect 4750 3035 4800 3065
rect 4750 3015 4765 3035
rect 4785 3015 4800 3035
rect 4750 2985 4800 3015
rect 4750 2965 4765 2985
rect 4785 2965 4800 2985
rect 4750 2935 4800 2965
rect 4750 2915 4765 2935
rect 4785 2915 4800 2935
rect 4750 2885 4800 2915
rect 4750 2865 4765 2885
rect 4785 2865 4800 2885
rect 4750 2835 4800 2865
rect 4750 2815 4765 2835
rect 4785 2815 4800 2835
rect 4750 2785 4800 2815
rect 4750 2765 4765 2785
rect 4785 2765 4800 2785
rect 4750 2735 4800 2765
rect 4750 2715 4765 2735
rect 4785 2715 4800 2735
rect 4750 2685 4800 2715
rect 4750 2665 4765 2685
rect 4785 2665 4800 2685
rect 4750 2650 4800 2665
rect 4900 3135 4950 3150
rect 4900 3115 4915 3135
rect 4935 3115 4950 3135
rect 4900 3085 4950 3115
rect 4900 3065 4915 3085
rect 4935 3065 4950 3085
rect 4900 3035 4950 3065
rect 4900 3015 4915 3035
rect 4935 3015 4950 3035
rect 4900 2985 4950 3015
rect 4900 2965 4915 2985
rect 4935 2965 4950 2985
rect 4900 2935 4950 2965
rect 4900 2915 4915 2935
rect 4935 2915 4950 2935
rect 4900 2885 4950 2915
rect 4900 2865 4915 2885
rect 4935 2865 4950 2885
rect 4900 2835 4950 2865
rect 4900 2815 4915 2835
rect 4935 2815 4950 2835
rect 4900 2785 4950 2815
rect 4900 2765 4915 2785
rect 4935 2765 4950 2785
rect 4900 2735 4950 2765
rect 4900 2715 4915 2735
rect 4935 2715 4950 2735
rect 4900 2685 4950 2715
rect 4900 2665 4915 2685
rect 4935 2665 4950 2685
rect 4900 2650 4950 2665
rect 5050 3135 5100 3150
rect 5050 3115 5065 3135
rect 5085 3115 5100 3135
rect 5050 3085 5100 3115
rect 5050 3065 5065 3085
rect 5085 3065 5100 3085
rect 5050 3035 5100 3065
rect 5050 3015 5065 3035
rect 5085 3015 5100 3035
rect 5050 2985 5100 3015
rect 5050 2965 5065 2985
rect 5085 2965 5100 2985
rect 5050 2935 5100 2965
rect 5050 2915 5065 2935
rect 5085 2915 5100 2935
rect 5050 2885 5100 2915
rect 5050 2865 5065 2885
rect 5085 2865 5100 2885
rect 5050 2835 5100 2865
rect 5050 2815 5065 2835
rect 5085 2815 5100 2835
rect 5050 2785 5100 2815
rect 5050 2765 5065 2785
rect 5085 2765 5100 2785
rect 5050 2735 5100 2765
rect 5050 2715 5065 2735
rect 5085 2715 5100 2735
rect 5050 2685 5100 2715
rect 5050 2665 5065 2685
rect 5085 2665 5100 2685
rect 5050 2650 5100 2665
rect 5200 3135 5250 3150
rect 5200 3115 5215 3135
rect 5235 3115 5250 3135
rect 5200 3085 5250 3115
rect 5200 3065 5215 3085
rect 5235 3065 5250 3085
rect 5200 3035 5250 3065
rect 5200 3015 5215 3035
rect 5235 3015 5250 3035
rect 5200 2985 5250 3015
rect 5200 2965 5215 2985
rect 5235 2965 5250 2985
rect 5200 2935 5250 2965
rect 5200 2915 5215 2935
rect 5235 2915 5250 2935
rect 5200 2885 5250 2915
rect 5200 2865 5215 2885
rect 5235 2865 5250 2885
rect 5200 2835 5250 2865
rect 5200 2815 5215 2835
rect 5235 2815 5250 2835
rect 5200 2785 5250 2815
rect 5200 2765 5215 2785
rect 5235 2765 5250 2785
rect 5200 2735 5250 2765
rect 5200 2715 5215 2735
rect 5235 2715 5250 2735
rect 5200 2685 5250 2715
rect 5200 2665 5215 2685
rect 5235 2665 5250 2685
rect 5200 2650 5250 2665
rect 5350 3135 5400 3150
rect 5350 3115 5365 3135
rect 5385 3115 5400 3135
rect 5350 3085 5400 3115
rect 5350 3065 5365 3085
rect 5385 3065 5400 3085
rect 5350 3035 5400 3065
rect 5350 3015 5365 3035
rect 5385 3015 5400 3035
rect 5350 2985 5400 3015
rect 5350 2965 5365 2985
rect 5385 2965 5400 2985
rect 5350 2935 5400 2965
rect 5350 2915 5365 2935
rect 5385 2915 5400 2935
rect 5350 2885 5400 2915
rect 5350 2865 5365 2885
rect 5385 2865 5400 2885
rect 5350 2835 5400 2865
rect 5350 2815 5365 2835
rect 5385 2815 5400 2835
rect 5350 2785 5400 2815
rect 5350 2765 5365 2785
rect 5385 2765 5400 2785
rect 5350 2735 5400 2765
rect 5350 2715 5365 2735
rect 5385 2715 5400 2735
rect 5350 2685 5400 2715
rect 5350 2665 5365 2685
rect 5385 2665 5400 2685
rect 5350 2650 5400 2665
rect 5500 3135 5550 3150
rect 5500 3115 5515 3135
rect 5535 3115 5550 3135
rect 5500 3085 5550 3115
rect 5500 3065 5515 3085
rect 5535 3065 5550 3085
rect 5500 3035 5550 3065
rect 5500 3015 5515 3035
rect 5535 3015 5550 3035
rect 5500 2985 5550 3015
rect 5500 2965 5515 2985
rect 5535 2965 5550 2985
rect 5500 2935 5550 2965
rect 5500 2915 5515 2935
rect 5535 2915 5550 2935
rect 5500 2885 5550 2915
rect 5500 2865 5515 2885
rect 5535 2865 5550 2885
rect 5500 2835 5550 2865
rect 5500 2815 5515 2835
rect 5535 2815 5550 2835
rect 5500 2785 5550 2815
rect 5500 2765 5515 2785
rect 5535 2765 5550 2785
rect 5500 2735 5550 2765
rect 5500 2715 5515 2735
rect 5535 2715 5550 2735
rect 5500 2685 5550 2715
rect 5500 2665 5515 2685
rect 5535 2665 5550 2685
rect 5500 2650 5550 2665
rect 5650 3135 5700 3150
rect 5650 3115 5665 3135
rect 5685 3115 5700 3135
rect 5650 3085 5700 3115
rect 5650 3065 5665 3085
rect 5685 3065 5700 3085
rect 5650 3035 5700 3065
rect 5650 3015 5665 3035
rect 5685 3015 5700 3035
rect 5650 2985 5700 3015
rect 5650 2965 5665 2985
rect 5685 2965 5700 2985
rect 5650 2935 5700 2965
rect 5650 2915 5665 2935
rect 5685 2915 5700 2935
rect 5650 2885 5700 2915
rect 5650 2865 5665 2885
rect 5685 2865 5700 2885
rect 5650 2835 5700 2865
rect 5650 2815 5665 2835
rect 5685 2815 5700 2835
rect 5650 2785 5700 2815
rect 5650 2765 5665 2785
rect 5685 2765 5700 2785
rect 5650 2735 5700 2765
rect 5650 2715 5665 2735
rect 5685 2715 5700 2735
rect 5650 2685 5700 2715
rect 5650 2665 5665 2685
rect 5685 2665 5700 2685
rect 5650 2650 5700 2665
rect 5800 3135 5850 3150
rect 5800 3115 5815 3135
rect 5835 3115 5850 3135
rect 5800 3085 5850 3115
rect 5800 3065 5815 3085
rect 5835 3065 5850 3085
rect 5800 3035 5850 3065
rect 5800 3015 5815 3035
rect 5835 3015 5850 3035
rect 5800 2985 5850 3015
rect 5800 2965 5815 2985
rect 5835 2965 5850 2985
rect 5800 2935 5850 2965
rect 5800 2915 5815 2935
rect 5835 2915 5850 2935
rect 5800 2885 5850 2915
rect 5800 2865 5815 2885
rect 5835 2865 5850 2885
rect 5800 2835 5850 2865
rect 5800 2815 5815 2835
rect 5835 2815 5850 2835
rect 5800 2785 5850 2815
rect 5800 2765 5815 2785
rect 5835 2765 5850 2785
rect 5800 2735 5850 2765
rect 5800 2715 5815 2735
rect 5835 2715 5850 2735
rect 5800 2685 5850 2715
rect 5800 2665 5815 2685
rect 5835 2665 5850 2685
rect 5800 2650 5850 2665
rect 5950 3135 6000 3150
rect 5950 3115 5965 3135
rect 5985 3115 6000 3135
rect 5950 3085 6000 3115
rect 5950 3065 5965 3085
rect 5985 3065 6000 3085
rect 5950 3035 6000 3065
rect 5950 3015 5965 3035
rect 5985 3015 6000 3035
rect 5950 2985 6000 3015
rect 5950 2965 5965 2985
rect 5985 2965 6000 2985
rect 5950 2935 6000 2965
rect 5950 2915 5965 2935
rect 5985 2915 6000 2935
rect 5950 2885 6000 2915
rect 5950 2865 5965 2885
rect 5985 2865 6000 2885
rect 5950 2835 6000 2865
rect 5950 2815 5965 2835
rect 5985 2815 6000 2835
rect 5950 2785 6000 2815
rect 5950 2765 5965 2785
rect 5985 2765 6000 2785
rect 5950 2735 6000 2765
rect 5950 2715 5965 2735
rect 5985 2715 6000 2735
rect 5950 2685 6000 2715
rect 5950 2665 5965 2685
rect 5985 2665 6000 2685
rect 5950 2650 6000 2665
rect 6100 3135 6150 3150
rect 6100 3115 6115 3135
rect 6135 3115 6150 3135
rect 6100 3085 6150 3115
rect 6100 3065 6115 3085
rect 6135 3065 6150 3085
rect 6100 3035 6150 3065
rect 6100 3015 6115 3035
rect 6135 3015 6150 3035
rect 6100 2985 6150 3015
rect 6100 2965 6115 2985
rect 6135 2965 6150 2985
rect 6100 2935 6150 2965
rect 6100 2915 6115 2935
rect 6135 2915 6150 2935
rect 6100 2885 6150 2915
rect 6100 2865 6115 2885
rect 6135 2865 6150 2885
rect 6100 2835 6150 2865
rect 6100 2815 6115 2835
rect 6135 2815 6150 2835
rect 6100 2785 6150 2815
rect 6100 2765 6115 2785
rect 6135 2765 6150 2785
rect 6100 2735 6150 2765
rect 6100 2715 6115 2735
rect 6135 2715 6150 2735
rect 6100 2685 6150 2715
rect 6100 2665 6115 2685
rect 6135 2665 6150 2685
rect 6100 2650 6150 2665
rect 6250 3135 6300 3150
rect 6250 3115 6265 3135
rect 6285 3115 6300 3135
rect 6250 3085 6300 3115
rect 6250 3065 6265 3085
rect 6285 3065 6300 3085
rect 6250 3035 6300 3065
rect 6250 3015 6265 3035
rect 6285 3015 6300 3035
rect 6250 2985 6300 3015
rect 6250 2965 6265 2985
rect 6285 2965 6300 2985
rect 6250 2935 6300 2965
rect 6250 2915 6265 2935
rect 6285 2915 6300 2935
rect 6250 2885 6300 2915
rect 6250 2865 6265 2885
rect 6285 2865 6300 2885
rect 6250 2835 6300 2865
rect 6250 2815 6265 2835
rect 6285 2815 6300 2835
rect 6250 2785 6300 2815
rect 6250 2765 6265 2785
rect 6285 2765 6300 2785
rect 6250 2735 6300 2765
rect 6250 2715 6265 2735
rect 6285 2715 6300 2735
rect 6250 2685 6300 2715
rect 6250 2665 6265 2685
rect 6285 2665 6300 2685
rect 6250 2650 6300 2665
rect 6400 3135 6450 3150
rect 6400 3115 6415 3135
rect 6435 3115 6450 3135
rect 6400 3085 6450 3115
rect 6400 3065 6415 3085
rect 6435 3065 6450 3085
rect 6400 3035 6450 3065
rect 6400 3015 6415 3035
rect 6435 3015 6450 3035
rect 6400 2985 6450 3015
rect 6400 2965 6415 2985
rect 6435 2965 6450 2985
rect 6400 2935 6450 2965
rect 6400 2915 6415 2935
rect 6435 2915 6450 2935
rect 6400 2885 6450 2915
rect 6400 2865 6415 2885
rect 6435 2865 6450 2885
rect 6400 2835 6450 2865
rect 6400 2815 6415 2835
rect 6435 2815 6450 2835
rect 6400 2785 6450 2815
rect 6400 2765 6415 2785
rect 6435 2765 6450 2785
rect 6400 2735 6450 2765
rect 6400 2715 6415 2735
rect 6435 2715 6450 2735
rect 6400 2685 6450 2715
rect 6400 2665 6415 2685
rect 6435 2665 6450 2685
rect 6400 2650 6450 2665
rect 6550 3135 6600 3150
rect 6550 3115 6565 3135
rect 6585 3115 6600 3135
rect 6550 3085 6600 3115
rect 6550 3065 6565 3085
rect 6585 3065 6600 3085
rect 6550 3035 6600 3065
rect 6550 3015 6565 3035
rect 6585 3015 6600 3035
rect 6550 2985 6600 3015
rect 6550 2965 6565 2985
rect 6585 2965 6600 2985
rect 6550 2935 6600 2965
rect 6550 2915 6565 2935
rect 6585 2915 6600 2935
rect 6550 2885 6600 2915
rect 6550 2865 6565 2885
rect 6585 2865 6600 2885
rect 6550 2835 6600 2865
rect 6550 2815 6565 2835
rect 6585 2815 6600 2835
rect 6550 2785 6600 2815
rect 6550 2765 6565 2785
rect 6585 2765 6600 2785
rect 6550 2735 6600 2765
rect 6550 2715 6565 2735
rect 6585 2715 6600 2735
rect 6550 2685 6600 2715
rect 6550 2665 6565 2685
rect 6585 2665 6600 2685
rect 6550 2650 6600 2665
rect 6700 3135 6750 3150
rect 6700 3115 6715 3135
rect 6735 3115 6750 3135
rect 6700 3085 6750 3115
rect 6700 3065 6715 3085
rect 6735 3065 6750 3085
rect 6700 3035 6750 3065
rect 6700 3015 6715 3035
rect 6735 3015 6750 3035
rect 6700 2985 6750 3015
rect 6700 2965 6715 2985
rect 6735 2965 6750 2985
rect 6700 2935 6750 2965
rect 6700 2915 6715 2935
rect 6735 2915 6750 2935
rect 6700 2885 6750 2915
rect 6700 2865 6715 2885
rect 6735 2865 6750 2885
rect 6700 2835 6750 2865
rect 6700 2815 6715 2835
rect 6735 2815 6750 2835
rect 6700 2785 6750 2815
rect 6700 2765 6715 2785
rect 6735 2765 6750 2785
rect 6700 2735 6750 2765
rect 6700 2715 6715 2735
rect 6735 2715 6750 2735
rect 6700 2685 6750 2715
rect 6700 2665 6715 2685
rect 6735 2665 6750 2685
rect 6700 2650 6750 2665
rect 6850 3135 6900 3150
rect 6850 3115 6865 3135
rect 6885 3115 6900 3135
rect 6850 3085 6900 3115
rect 6850 3065 6865 3085
rect 6885 3065 6900 3085
rect 6850 3035 6900 3065
rect 6850 3015 6865 3035
rect 6885 3015 6900 3035
rect 6850 2985 6900 3015
rect 6850 2965 6865 2985
rect 6885 2965 6900 2985
rect 6850 2935 6900 2965
rect 6850 2915 6865 2935
rect 6885 2915 6900 2935
rect 6850 2885 6900 2915
rect 6850 2865 6865 2885
rect 6885 2865 6900 2885
rect 6850 2835 6900 2865
rect 6850 2815 6865 2835
rect 6885 2815 6900 2835
rect 6850 2785 6900 2815
rect 6850 2765 6865 2785
rect 6885 2765 6900 2785
rect 6850 2735 6900 2765
rect 6850 2715 6865 2735
rect 6885 2715 6900 2735
rect 6850 2685 6900 2715
rect 6850 2665 6865 2685
rect 6885 2665 6900 2685
rect 6850 2650 6900 2665
rect 7000 3135 7050 3150
rect 7000 3115 7015 3135
rect 7035 3115 7050 3135
rect 7000 3085 7050 3115
rect 7000 3065 7015 3085
rect 7035 3065 7050 3085
rect 7000 3035 7050 3065
rect 7000 3015 7015 3035
rect 7035 3015 7050 3035
rect 7000 2985 7050 3015
rect 7000 2965 7015 2985
rect 7035 2965 7050 2985
rect 7000 2935 7050 2965
rect 7000 2915 7015 2935
rect 7035 2915 7050 2935
rect 7000 2885 7050 2915
rect 7000 2865 7015 2885
rect 7035 2865 7050 2885
rect 7000 2835 7050 2865
rect 7000 2815 7015 2835
rect 7035 2815 7050 2835
rect 7000 2785 7050 2815
rect 7000 2765 7015 2785
rect 7035 2765 7050 2785
rect 7000 2735 7050 2765
rect 7000 2715 7015 2735
rect 7035 2715 7050 2735
rect 7000 2685 7050 2715
rect 7000 2665 7015 2685
rect 7035 2665 7050 2685
rect 7000 2650 7050 2665
rect 7150 3135 7200 3150
rect 7150 3115 7165 3135
rect 7185 3115 7200 3135
rect 7150 3085 7200 3115
rect 7150 3065 7165 3085
rect 7185 3065 7200 3085
rect 7150 3035 7200 3065
rect 7150 3015 7165 3035
rect 7185 3015 7200 3035
rect 7150 2985 7200 3015
rect 7150 2965 7165 2985
rect 7185 2965 7200 2985
rect 7150 2935 7200 2965
rect 7150 2915 7165 2935
rect 7185 2915 7200 2935
rect 7150 2885 7200 2915
rect 7150 2865 7165 2885
rect 7185 2865 7200 2885
rect 7150 2835 7200 2865
rect 7150 2815 7165 2835
rect 7185 2815 7200 2835
rect 7150 2785 7200 2815
rect 7150 2765 7165 2785
rect 7185 2765 7200 2785
rect 7150 2735 7200 2765
rect 7150 2715 7165 2735
rect 7185 2715 7200 2735
rect 7150 2685 7200 2715
rect 7150 2665 7165 2685
rect 7185 2665 7200 2685
rect 7150 2650 7200 2665
rect 7300 3135 7350 3150
rect 7300 3115 7315 3135
rect 7335 3115 7350 3135
rect 7300 3085 7350 3115
rect 7300 3065 7315 3085
rect 7335 3065 7350 3085
rect 7300 3035 7350 3065
rect 7300 3015 7315 3035
rect 7335 3015 7350 3035
rect 7300 2985 7350 3015
rect 7300 2965 7315 2985
rect 7335 2965 7350 2985
rect 7300 2935 7350 2965
rect 7300 2915 7315 2935
rect 7335 2915 7350 2935
rect 7300 2885 7350 2915
rect 7300 2865 7315 2885
rect 7335 2865 7350 2885
rect 7300 2835 7350 2865
rect 7300 2815 7315 2835
rect 7335 2815 7350 2835
rect 7300 2785 7350 2815
rect 7300 2765 7315 2785
rect 7335 2765 7350 2785
rect 7300 2735 7350 2765
rect 7300 2715 7315 2735
rect 7335 2715 7350 2735
rect 7300 2685 7350 2715
rect 7300 2665 7315 2685
rect 7335 2665 7350 2685
rect 7300 2650 7350 2665
rect 7450 3135 7500 3150
rect 7450 3115 7465 3135
rect 7485 3115 7500 3135
rect 7450 3085 7500 3115
rect 7450 3065 7465 3085
rect 7485 3065 7500 3085
rect 7450 3035 7500 3065
rect 7450 3015 7465 3035
rect 7485 3015 7500 3035
rect 7450 2985 7500 3015
rect 7450 2965 7465 2985
rect 7485 2965 7500 2985
rect 7450 2935 7500 2965
rect 7450 2915 7465 2935
rect 7485 2915 7500 2935
rect 7450 2885 7500 2915
rect 7450 2865 7465 2885
rect 7485 2865 7500 2885
rect 7450 2835 7500 2865
rect 7450 2815 7465 2835
rect 7485 2815 7500 2835
rect 7450 2785 7500 2815
rect 7450 2765 7465 2785
rect 7485 2765 7500 2785
rect 7450 2735 7500 2765
rect 7450 2715 7465 2735
rect 7485 2715 7500 2735
rect 7450 2685 7500 2715
rect 7450 2665 7465 2685
rect 7485 2665 7500 2685
rect 7450 2650 7500 2665
rect 7600 3135 7650 3150
rect 7600 3115 7615 3135
rect 7635 3115 7650 3135
rect 7600 3085 7650 3115
rect 7600 3065 7615 3085
rect 7635 3065 7650 3085
rect 7600 3035 7650 3065
rect 7600 3015 7615 3035
rect 7635 3015 7650 3035
rect 7600 2985 7650 3015
rect 7600 2965 7615 2985
rect 7635 2965 7650 2985
rect 7600 2935 7650 2965
rect 7600 2915 7615 2935
rect 7635 2915 7650 2935
rect 7600 2885 7650 2915
rect 7600 2865 7615 2885
rect 7635 2865 7650 2885
rect 7600 2835 7650 2865
rect 7600 2815 7615 2835
rect 7635 2815 7650 2835
rect 7600 2785 7650 2815
rect 7600 2765 7615 2785
rect 7635 2765 7650 2785
rect 7600 2735 7650 2765
rect 7600 2715 7615 2735
rect 7635 2715 7650 2735
rect 7600 2685 7650 2715
rect 7600 2665 7615 2685
rect 7635 2665 7650 2685
rect 7600 2650 7650 2665
rect 7750 3135 7800 3150
rect 7750 3115 7765 3135
rect 7785 3115 7800 3135
rect 7750 3085 7800 3115
rect 7750 3065 7765 3085
rect 7785 3065 7800 3085
rect 7750 3035 7800 3065
rect 7750 3015 7765 3035
rect 7785 3015 7800 3035
rect 7750 2985 7800 3015
rect 7750 2965 7765 2985
rect 7785 2965 7800 2985
rect 7750 2935 7800 2965
rect 7750 2915 7765 2935
rect 7785 2915 7800 2935
rect 7750 2885 7800 2915
rect 7750 2865 7765 2885
rect 7785 2865 7800 2885
rect 7750 2835 7800 2865
rect 7750 2815 7765 2835
rect 7785 2815 7800 2835
rect 7750 2785 7800 2815
rect 7750 2765 7765 2785
rect 7785 2765 7800 2785
rect 7750 2735 7800 2765
rect 7750 2715 7765 2735
rect 7785 2715 7800 2735
rect 7750 2685 7800 2715
rect 7750 2665 7765 2685
rect 7785 2665 7800 2685
rect 7750 2650 7800 2665
rect 8350 3135 8400 3150
rect 8350 3115 8365 3135
rect 8385 3115 8400 3135
rect 8350 3085 8400 3115
rect 8350 3065 8365 3085
rect 8385 3065 8400 3085
rect 8350 3035 8400 3065
rect 8350 3015 8365 3035
rect 8385 3015 8400 3035
rect 8350 2985 8400 3015
rect 8350 2965 8365 2985
rect 8385 2965 8400 2985
rect 8350 2935 8400 2965
rect 8350 2915 8365 2935
rect 8385 2915 8400 2935
rect 8350 2885 8400 2915
rect 8350 2865 8365 2885
rect 8385 2865 8400 2885
rect 8350 2835 8400 2865
rect 8350 2815 8365 2835
rect 8385 2815 8400 2835
rect 8350 2785 8400 2815
rect 8350 2765 8365 2785
rect 8385 2765 8400 2785
rect 8350 2735 8400 2765
rect 8350 2715 8365 2735
rect 8385 2715 8400 2735
rect 8350 2685 8400 2715
rect 8350 2665 8365 2685
rect 8385 2665 8400 2685
rect 8350 2650 8400 2665
rect 8500 3135 8550 3200
rect 8500 3115 8515 3135
rect 8535 3115 8550 3135
rect 8500 3085 8550 3115
rect 8500 3065 8515 3085
rect 8535 3065 8550 3085
rect 8500 3035 8550 3065
rect 8500 3015 8515 3035
rect 8535 3015 8550 3035
rect 8500 2985 8550 3015
rect 8500 2965 8515 2985
rect 8535 2965 8550 2985
rect 8500 2935 8550 2965
rect 8500 2915 8515 2935
rect 8535 2915 8550 2935
rect 8500 2885 8550 2915
rect 8500 2865 8515 2885
rect 8535 2865 8550 2885
rect 8500 2835 8550 2865
rect 8500 2815 8515 2835
rect 8535 2815 8550 2835
rect 8500 2785 8550 2815
rect 8500 2765 8515 2785
rect 8535 2765 8550 2785
rect 8500 2735 8550 2765
rect 8500 2715 8515 2735
rect 8535 2715 8550 2735
rect 8500 2685 8550 2715
rect 8500 2665 8515 2685
rect 8535 2665 8550 2685
rect 8500 2650 8550 2665
rect 8650 3135 8700 3150
rect 8650 3115 8665 3135
rect 8685 3115 8700 3135
rect 8650 3085 8700 3115
rect 8650 3065 8665 3085
rect 8685 3065 8700 3085
rect 8650 3035 8700 3065
rect 8650 3015 8665 3035
rect 8685 3015 8700 3035
rect 8650 2985 8700 3015
rect 8650 2965 8665 2985
rect 8685 2965 8700 2985
rect 8650 2935 8700 2965
rect 8650 2915 8665 2935
rect 8685 2915 8700 2935
rect 8650 2885 8700 2915
rect 8650 2865 8665 2885
rect 8685 2865 8700 2885
rect 8650 2835 8700 2865
rect 8650 2815 8665 2835
rect 8685 2815 8700 2835
rect 8650 2785 8700 2815
rect 8650 2765 8665 2785
rect 8685 2765 8700 2785
rect 8650 2735 8700 2765
rect 8650 2715 8665 2735
rect 8685 2715 8700 2735
rect 8650 2685 8700 2715
rect 8650 2665 8665 2685
rect 8685 2665 8700 2685
rect 8650 2650 8700 2665
rect 8800 3135 8850 3200
rect 8800 3115 8815 3135
rect 8835 3115 8850 3135
rect 8800 3085 8850 3115
rect 8800 3065 8815 3085
rect 8835 3065 8850 3085
rect 8800 3035 8850 3065
rect 8800 3015 8815 3035
rect 8835 3015 8850 3035
rect 8800 2985 8850 3015
rect 8800 2965 8815 2985
rect 8835 2965 8850 2985
rect 8800 2935 8850 2965
rect 8800 2915 8815 2935
rect 8835 2915 8850 2935
rect 8800 2885 8850 2915
rect 8800 2865 8815 2885
rect 8835 2865 8850 2885
rect 8800 2835 8850 2865
rect 8800 2815 8815 2835
rect 8835 2815 8850 2835
rect 8800 2785 8850 2815
rect 8800 2765 8815 2785
rect 8835 2765 8850 2785
rect 8800 2735 8850 2765
rect 8800 2715 8815 2735
rect 8835 2715 8850 2735
rect 8800 2685 8850 2715
rect 8800 2665 8815 2685
rect 8835 2665 8850 2685
rect 8800 2650 8850 2665
rect 8950 3135 9000 3150
rect 8950 3115 8965 3135
rect 8985 3115 9000 3135
rect 8950 3085 9000 3115
rect 8950 3065 8965 3085
rect 8985 3065 9000 3085
rect 8950 3035 9000 3065
rect 8950 3015 8965 3035
rect 8985 3015 9000 3035
rect 8950 2985 9000 3015
rect 8950 2965 8965 2985
rect 8985 2965 9000 2985
rect 8950 2935 9000 2965
rect 8950 2915 8965 2935
rect 8985 2915 9000 2935
rect 8950 2885 9000 2915
rect 8950 2865 8965 2885
rect 8985 2865 9000 2885
rect 8950 2835 9000 2865
rect 8950 2815 8965 2835
rect 8985 2815 9000 2835
rect 8950 2785 9000 2815
rect 8950 2765 8965 2785
rect 8985 2765 9000 2785
rect 8950 2735 9000 2765
rect 8950 2715 8965 2735
rect 8985 2715 9000 2735
rect 8950 2685 9000 2715
rect 8950 2665 8965 2685
rect 8985 2665 9000 2685
rect 8950 2650 9000 2665
rect 9100 3135 9150 3200
rect 9100 3115 9115 3135
rect 9135 3115 9150 3135
rect 9100 3085 9150 3115
rect 9100 3065 9115 3085
rect 9135 3065 9150 3085
rect 9100 3035 9150 3065
rect 9100 3015 9115 3035
rect 9135 3015 9150 3035
rect 9100 2985 9150 3015
rect 9100 2965 9115 2985
rect 9135 2965 9150 2985
rect 9100 2935 9150 2965
rect 9100 2915 9115 2935
rect 9135 2915 9150 2935
rect 9100 2885 9150 2915
rect 9100 2865 9115 2885
rect 9135 2865 9150 2885
rect 9100 2835 9150 2865
rect 9100 2815 9115 2835
rect 9135 2815 9150 2835
rect 9100 2785 9150 2815
rect 9100 2765 9115 2785
rect 9135 2765 9150 2785
rect 9100 2735 9150 2765
rect 9100 2715 9115 2735
rect 9135 2715 9150 2735
rect 9100 2685 9150 2715
rect 9100 2665 9115 2685
rect 9135 2665 9150 2685
rect 9100 2650 9150 2665
rect 9250 3135 9300 3150
rect 9250 3115 9265 3135
rect 9285 3115 9300 3135
rect 9250 3085 9300 3115
rect 9250 3065 9265 3085
rect 9285 3065 9300 3085
rect 9250 3035 9300 3065
rect 9250 3015 9265 3035
rect 9285 3015 9300 3035
rect 9250 2985 9300 3015
rect 9250 2965 9265 2985
rect 9285 2965 9300 2985
rect 9250 2935 9300 2965
rect 9250 2915 9265 2935
rect 9285 2915 9300 2935
rect 9250 2885 9300 2915
rect 9250 2865 9265 2885
rect 9285 2865 9300 2885
rect 9250 2835 9300 2865
rect 9250 2815 9265 2835
rect 9285 2815 9300 2835
rect 9250 2785 9300 2815
rect 9250 2765 9265 2785
rect 9285 2765 9300 2785
rect 9250 2735 9300 2765
rect 9250 2715 9265 2735
rect 9285 2715 9300 2735
rect 9250 2685 9300 2715
rect 9250 2665 9265 2685
rect 9285 2665 9300 2685
rect 9250 2650 9300 2665
rect 9400 3135 9450 3200
rect 9400 3115 9415 3135
rect 9435 3115 9450 3135
rect 9400 3085 9450 3115
rect 9400 3065 9415 3085
rect 9435 3065 9450 3085
rect 9400 3035 9450 3065
rect 9400 3015 9415 3035
rect 9435 3015 9450 3035
rect 9400 2985 9450 3015
rect 9400 2965 9415 2985
rect 9435 2965 9450 2985
rect 9400 2935 9450 2965
rect 9400 2915 9415 2935
rect 9435 2915 9450 2935
rect 9400 2885 9450 2915
rect 9400 2865 9415 2885
rect 9435 2865 9450 2885
rect 9400 2835 9450 2865
rect 9400 2815 9415 2835
rect 9435 2815 9450 2835
rect 9400 2785 9450 2815
rect 9400 2765 9415 2785
rect 9435 2765 9450 2785
rect 9400 2735 9450 2765
rect 9400 2715 9415 2735
rect 9435 2715 9450 2735
rect 9400 2685 9450 2715
rect 9400 2665 9415 2685
rect 9435 2665 9450 2685
rect 9400 2650 9450 2665
rect 9550 3135 9600 3150
rect 9550 3115 9565 3135
rect 9585 3115 9600 3135
rect 9550 3085 9600 3115
rect 9550 3065 9565 3085
rect 9585 3065 9600 3085
rect 9550 3035 9600 3065
rect 9550 3015 9565 3035
rect 9585 3015 9600 3035
rect 9550 2985 9600 3015
rect 9550 2965 9565 2985
rect 9585 2965 9600 2985
rect 9550 2935 9600 2965
rect 9550 2915 9565 2935
rect 9585 2915 9600 2935
rect 9550 2885 9600 2915
rect 9550 2865 9565 2885
rect 9585 2865 9600 2885
rect 9550 2835 9600 2865
rect 9550 2815 9565 2835
rect 9585 2815 9600 2835
rect 9550 2785 9600 2815
rect 9550 2765 9565 2785
rect 9585 2765 9600 2785
rect 9550 2735 9600 2765
rect 9550 2715 9565 2735
rect 9585 2715 9600 2735
rect 9550 2685 9600 2715
rect 9550 2665 9565 2685
rect 9585 2665 9600 2685
rect 9550 2650 9600 2665
rect 9700 3135 9750 3200
rect 9700 3115 9715 3135
rect 9735 3115 9750 3135
rect 9700 3085 9750 3115
rect 9700 3065 9715 3085
rect 9735 3065 9750 3085
rect 9700 3035 9750 3065
rect 9700 3015 9715 3035
rect 9735 3015 9750 3035
rect 9700 2985 9750 3015
rect 9700 2965 9715 2985
rect 9735 2965 9750 2985
rect 9700 2935 9750 2965
rect 9700 2915 9715 2935
rect 9735 2915 9750 2935
rect 9700 2885 9750 2915
rect 9700 2865 9715 2885
rect 9735 2865 9750 2885
rect 9700 2835 9750 2865
rect 9700 2815 9715 2835
rect 9735 2815 9750 2835
rect 9700 2785 9750 2815
rect 9700 2765 9715 2785
rect 9735 2765 9750 2785
rect 9700 2735 9750 2765
rect 9700 2715 9715 2735
rect 9735 2715 9750 2735
rect 9700 2685 9750 2715
rect 9700 2665 9715 2685
rect 9735 2665 9750 2685
rect 9700 2650 9750 2665
rect 9850 3135 9900 3150
rect 9850 3115 9865 3135
rect 9885 3115 9900 3135
rect 9850 3085 9900 3115
rect 9850 3065 9865 3085
rect 9885 3065 9900 3085
rect 9850 3035 9900 3065
rect 9850 3015 9865 3035
rect 9885 3015 9900 3035
rect 9850 2985 9900 3015
rect 9850 2965 9865 2985
rect 9885 2965 9900 2985
rect 9850 2935 9900 2965
rect 9850 2915 9865 2935
rect 9885 2915 9900 2935
rect 9850 2885 9900 2915
rect 9850 2865 9865 2885
rect 9885 2865 9900 2885
rect 9850 2835 9900 2865
rect 9850 2815 9865 2835
rect 9885 2815 9900 2835
rect 9850 2785 9900 2815
rect 9850 2765 9865 2785
rect 9885 2765 9900 2785
rect 9850 2735 9900 2765
rect 9850 2715 9865 2735
rect 9885 2715 9900 2735
rect 9850 2685 9900 2715
rect 9850 2665 9865 2685
rect 9885 2665 9900 2685
rect 9850 2650 9900 2665
rect 10000 3135 10050 3200
rect 10000 3115 10015 3135
rect 10035 3115 10050 3135
rect 10000 3085 10050 3115
rect 10000 3065 10015 3085
rect 10035 3065 10050 3085
rect 10000 3035 10050 3065
rect 10000 3015 10015 3035
rect 10035 3015 10050 3035
rect 10000 2985 10050 3015
rect 10000 2965 10015 2985
rect 10035 2965 10050 2985
rect 10000 2935 10050 2965
rect 10000 2915 10015 2935
rect 10035 2915 10050 2935
rect 10000 2885 10050 2915
rect 10000 2865 10015 2885
rect 10035 2865 10050 2885
rect 10000 2835 10050 2865
rect 10000 2815 10015 2835
rect 10035 2815 10050 2835
rect 10000 2785 10050 2815
rect 10000 2765 10015 2785
rect 10035 2765 10050 2785
rect 10000 2735 10050 2765
rect 10000 2715 10015 2735
rect 10035 2715 10050 2735
rect 10000 2685 10050 2715
rect 10000 2665 10015 2685
rect 10035 2665 10050 2685
rect 10000 2650 10050 2665
rect 10150 3135 10200 3150
rect 10150 3115 10165 3135
rect 10185 3115 10200 3135
rect 10150 3085 10200 3115
rect 10150 3065 10165 3085
rect 10185 3065 10200 3085
rect 10150 3035 10200 3065
rect 10150 3015 10165 3035
rect 10185 3015 10200 3035
rect 10150 2985 10200 3015
rect 10150 2965 10165 2985
rect 10185 2965 10200 2985
rect 10150 2935 10200 2965
rect 10150 2915 10165 2935
rect 10185 2915 10200 2935
rect 10150 2885 10200 2915
rect 10150 2865 10165 2885
rect 10185 2865 10200 2885
rect 10150 2835 10200 2865
rect 10150 2815 10165 2835
rect 10185 2815 10200 2835
rect 10150 2785 10200 2815
rect 10150 2765 10165 2785
rect 10185 2765 10200 2785
rect 10150 2735 10200 2765
rect 10150 2715 10165 2735
rect 10185 2715 10200 2735
rect 10150 2685 10200 2715
rect 10150 2665 10165 2685
rect 10185 2665 10200 2685
rect 10150 2650 10200 2665
rect 10300 3135 10350 3200
rect 10300 3115 10315 3135
rect 10335 3115 10350 3135
rect 10300 3085 10350 3115
rect 10300 3065 10315 3085
rect 10335 3065 10350 3085
rect 10300 3035 10350 3065
rect 10300 3015 10315 3035
rect 10335 3015 10350 3035
rect 10300 2985 10350 3015
rect 10300 2965 10315 2985
rect 10335 2965 10350 2985
rect 10300 2935 10350 2965
rect 10300 2915 10315 2935
rect 10335 2915 10350 2935
rect 10300 2885 10350 2915
rect 10300 2865 10315 2885
rect 10335 2865 10350 2885
rect 10300 2835 10350 2865
rect 10300 2815 10315 2835
rect 10335 2815 10350 2835
rect 10300 2785 10350 2815
rect 10300 2765 10315 2785
rect 10335 2765 10350 2785
rect 10300 2735 10350 2765
rect 10300 2715 10315 2735
rect 10335 2715 10350 2735
rect 10300 2685 10350 2715
rect 10300 2665 10315 2685
rect 10335 2665 10350 2685
rect 10300 2650 10350 2665
rect 10450 3135 10500 3150
rect 10450 3115 10465 3135
rect 10485 3115 10500 3135
rect 10450 3085 10500 3115
rect 10450 3065 10465 3085
rect 10485 3065 10500 3085
rect 10450 3035 10500 3065
rect 10450 3015 10465 3035
rect 10485 3015 10500 3035
rect 10450 2985 10500 3015
rect 10450 2965 10465 2985
rect 10485 2965 10500 2985
rect 10450 2935 10500 2965
rect 10450 2915 10465 2935
rect 10485 2915 10500 2935
rect 10450 2885 10500 2915
rect 10450 2865 10465 2885
rect 10485 2865 10500 2885
rect 10450 2835 10500 2865
rect 10450 2815 10465 2835
rect 10485 2815 10500 2835
rect 10450 2785 10500 2815
rect 10450 2765 10465 2785
rect 10485 2765 10500 2785
rect 10450 2735 10500 2765
rect 10450 2715 10465 2735
rect 10485 2715 10500 2735
rect 10450 2685 10500 2715
rect 10450 2665 10465 2685
rect 10485 2665 10500 2685
rect 10450 2650 10500 2665
rect 10600 3135 10650 3200
rect 10600 3115 10615 3135
rect 10635 3115 10650 3135
rect 10600 3085 10650 3115
rect 10600 3065 10615 3085
rect 10635 3065 10650 3085
rect 10600 3035 10650 3065
rect 10600 3015 10615 3035
rect 10635 3015 10650 3035
rect 10600 2985 10650 3015
rect 10600 2965 10615 2985
rect 10635 2965 10650 2985
rect 10600 2935 10650 2965
rect 10600 2915 10615 2935
rect 10635 2915 10650 2935
rect 10600 2885 10650 2915
rect 10600 2865 10615 2885
rect 10635 2865 10650 2885
rect 10600 2835 10650 2865
rect 10600 2815 10615 2835
rect 10635 2815 10650 2835
rect 10600 2785 10650 2815
rect 10600 2765 10615 2785
rect 10635 2765 10650 2785
rect 10600 2735 10650 2765
rect 10600 2715 10615 2735
rect 10635 2715 10650 2735
rect 10600 2685 10650 2715
rect 10600 2665 10615 2685
rect 10635 2665 10650 2685
rect 10600 2650 10650 2665
rect 10750 3135 10800 3150
rect 10750 3115 10765 3135
rect 10785 3115 10800 3135
rect 10750 3085 10800 3115
rect 10750 3065 10765 3085
rect 10785 3065 10800 3085
rect 10750 3035 10800 3065
rect 10750 3015 10765 3035
rect 10785 3015 10800 3035
rect 10750 2985 10800 3015
rect 10750 2965 10765 2985
rect 10785 2965 10800 2985
rect 10750 2935 10800 2965
rect 10750 2915 10765 2935
rect 10785 2915 10800 2935
rect 10750 2885 10800 2915
rect 10750 2865 10765 2885
rect 10785 2865 10800 2885
rect 10750 2835 10800 2865
rect 10750 2815 10765 2835
rect 10785 2815 10800 2835
rect 10750 2785 10800 2815
rect 10750 2765 10765 2785
rect 10785 2765 10800 2785
rect 10750 2735 10800 2765
rect 10750 2715 10765 2735
rect 10785 2715 10800 2735
rect 10750 2685 10800 2715
rect 10750 2665 10765 2685
rect 10785 2665 10800 2685
rect 10750 2650 10800 2665
rect 11350 3135 11400 3150
rect 11350 3115 11365 3135
rect 11385 3115 11400 3135
rect 11350 3085 11400 3115
rect 11350 3065 11365 3085
rect 11385 3065 11400 3085
rect 11350 3035 11400 3065
rect 11350 3015 11365 3035
rect 11385 3015 11400 3035
rect 11350 2985 11400 3015
rect 11350 2965 11365 2985
rect 11385 2965 11400 2985
rect 11350 2935 11400 2965
rect 11350 2915 11365 2935
rect 11385 2915 11400 2935
rect 11350 2885 11400 2915
rect 11350 2865 11365 2885
rect 11385 2865 11400 2885
rect 11350 2835 11400 2865
rect 11350 2815 11365 2835
rect 11385 2815 11400 2835
rect 11350 2785 11400 2815
rect 11350 2765 11365 2785
rect 11385 2765 11400 2785
rect 11350 2735 11400 2765
rect 11350 2715 11365 2735
rect 11385 2715 11400 2735
rect 11350 2685 11400 2715
rect 11350 2665 11365 2685
rect 11385 2665 11400 2685
rect 11350 2650 11400 2665
rect 11950 3135 12000 3150
rect 11950 3115 11965 3135
rect 11985 3115 12000 3135
rect 11950 3085 12000 3115
rect 11950 3065 11965 3085
rect 11985 3065 12000 3085
rect 11950 3035 12000 3065
rect 11950 3015 11965 3035
rect 11985 3015 12000 3035
rect 11950 2985 12000 3015
rect 11950 2965 11965 2985
rect 11985 2965 12000 2985
rect 11950 2935 12000 2965
rect 11950 2915 11965 2935
rect 11985 2915 12000 2935
rect 11950 2885 12000 2915
rect 11950 2865 11965 2885
rect 11985 2865 12000 2885
rect 11950 2835 12000 2865
rect 11950 2815 11965 2835
rect 11985 2815 12000 2835
rect 11950 2785 12000 2815
rect 11950 2765 11965 2785
rect 11985 2765 12000 2785
rect 11950 2735 12000 2765
rect 11950 2715 11965 2735
rect 11985 2715 12000 2735
rect 11950 2685 12000 2715
rect 11950 2665 11965 2685
rect 11985 2665 12000 2685
rect 11950 2650 12000 2665
rect 12550 3135 12600 3150
rect 12550 3115 12565 3135
rect 12585 3115 12600 3135
rect 12550 3085 12600 3115
rect 12550 3065 12565 3085
rect 12585 3065 12600 3085
rect 12550 3035 12600 3065
rect 12550 3015 12565 3035
rect 12585 3015 12600 3035
rect 12550 2985 12600 3015
rect 12550 2965 12565 2985
rect 12585 2965 12600 2985
rect 12550 2935 12600 2965
rect 12550 2915 12565 2935
rect 12585 2915 12600 2935
rect 12550 2885 12600 2915
rect 12550 2865 12565 2885
rect 12585 2865 12600 2885
rect 12550 2835 12600 2865
rect 12550 2815 12565 2835
rect 12585 2815 12600 2835
rect 12550 2785 12600 2815
rect 12550 2765 12565 2785
rect 12585 2765 12600 2785
rect 12550 2735 12600 2765
rect 12550 2715 12565 2735
rect 12585 2715 12600 2735
rect 12550 2685 12600 2715
rect 12550 2665 12565 2685
rect 12585 2665 12600 2685
rect 12550 2650 12600 2665
rect 13150 3135 13200 3150
rect 13150 3115 13165 3135
rect 13185 3115 13200 3135
rect 13150 3085 13200 3115
rect 13150 3065 13165 3085
rect 13185 3065 13200 3085
rect 13150 3035 13200 3065
rect 13150 3015 13165 3035
rect 13185 3015 13200 3035
rect 13150 2985 13200 3015
rect 13150 2965 13165 2985
rect 13185 2965 13200 2985
rect 13150 2935 13200 2965
rect 13150 2915 13165 2935
rect 13185 2915 13200 2935
rect 13150 2885 13200 2915
rect 13150 2865 13165 2885
rect 13185 2865 13200 2885
rect 13150 2835 13200 2865
rect 13150 2815 13165 2835
rect 13185 2815 13200 2835
rect 13150 2785 13200 2815
rect 13150 2765 13165 2785
rect 13185 2765 13200 2785
rect 13150 2735 13200 2765
rect 13150 2715 13165 2735
rect 13185 2715 13200 2735
rect 13150 2685 13200 2715
rect 13150 2665 13165 2685
rect 13185 2665 13200 2685
rect 13150 2650 13200 2665
rect 13750 3135 13800 3150
rect 13750 3115 13765 3135
rect 13785 3115 13800 3135
rect 13750 3085 13800 3115
rect 13750 3065 13765 3085
rect 13785 3065 13800 3085
rect 13750 3035 13800 3065
rect 13750 3015 13765 3035
rect 13785 3015 13800 3035
rect 13750 2985 13800 3015
rect 13750 2965 13765 2985
rect 13785 2965 13800 2985
rect 13750 2935 13800 2965
rect 13750 2915 13765 2935
rect 13785 2915 13800 2935
rect 13750 2885 13800 2915
rect 13750 2865 13765 2885
rect 13785 2865 13800 2885
rect 13750 2835 13800 2865
rect 13750 2815 13765 2835
rect 13785 2815 13800 2835
rect 13750 2785 13800 2815
rect 13750 2765 13765 2785
rect 13785 2765 13800 2785
rect 13750 2735 13800 2765
rect 13750 2715 13765 2735
rect 13785 2715 13800 2735
rect 13750 2685 13800 2715
rect 13750 2665 13765 2685
rect 13785 2665 13800 2685
rect 13750 2650 13800 2665
rect 14350 3135 14400 3150
rect 14350 3115 14365 3135
rect 14385 3115 14400 3135
rect 14350 3085 14400 3115
rect 14350 3065 14365 3085
rect 14385 3065 14400 3085
rect 14350 3035 14400 3065
rect 14350 3015 14365 3035
rect 14385 3015 14400 3035
rect 14350 2985 14400 3015
rect 14350 2965 14365 2985
rect 14385 2965 14400 2985
rect 14350 2935 14400 2965
rect 14350 2915 14365 2935
rect 14385 2915 14400 2935
rect 14350 2885 14400 2915
rect 14350 2865 14365 2885
rect 14385 2865 14400 2885
rect 14350 2835 14400 2865
rect 14350 2815 14365 2835
rect 14385 2815 14400 2835
rect 14350 2785 14400 2815
rect 14350 2765 14365 2785
rect 14385 2765 14400 2785
rect 14350 2735 14400 2765
rect 14350 2715 14365 2735
rect 14385 2715 14400 2735
rect 14350 2685 14400 2715
rect 14350 2665 14365 2685
rect 14385 2665 14400 2685
rect 14350 2650 14400 2665
rect 14950 3135 15000 3150
rect 14950 3115 14965 3135
rect 14985 3115 15000 3135
rect 14950 3085 15000 3115
rect 14950 3065 14965 3085
rect 14985 3065 15000 3085
rect 14950 3035 15000 3065
rect 14950 3015 14965 3035
rect 14985 3015 15000 3035
rect 14950 2985 15000 3015
rect 14950 2965 14965 2985
rect 14985 2965 15000 2985
rect 14950 2935 15000 2965
rect 14950 2915 14965 2935
rect 14985 2915 15000 2935
rect 14950 2885 15000 2915
rect 14950 2865 14965 2885
rect 14985 2865 15000 2885
rect 14950 2835 15000 2865
rect 14950 2815 14965 2835
rect 14985 2815 15000 2835
rect 14950 2785 15000 2815
rect 14950 2765 14965 2785
rect 14985 2765 15000 2785
rect 14950 2735 15000 2765
rect 14950 2715 14965 2735
rect 14985 2715 15000 2735
rect 14950 2685 15000 2715
rect 14950 2665 14965 2685
rect 14985 2665 15000 2685
rect 14950 2650 15000 2665
rect 15550 3135 15600 3150
rect 15550 3115 15565 3135
rect 15585 3115 15600 3135
rect 15550 3085 15600 3115
rect 15550 3065 15565 3085
rect 15585 3065 15600 3085
rect 15550 3035 15600 3065
rect 15550 3015 15565 3035
rect 15585 3015 15600 3035
rect 15550 2985 15600 3015
rect 15550 2965 15565 2985
rect 15585 2965 15600 2985
rect 15550 2935 15600 2965
rect 15550 2915 15565 2935
rect 15585 2915 15600 2935
rect 15550 2885 15600 2915
rect 15550 2865 15565 2885
rect 15585 2865 15600 2885
rect 15550 2835 15600 2865
rect 15550 2815 15565 2835
rect 15585 2815 15600 2835
rect 15550 2785 15600 2815
rect 15550 2765 15565 2785
rect 15585 2765 15600 2785
rect 15550 2735 15600 2765
rect 15550 2715 15565 2735
rect 15585 2715 15600 2735
rect 15550 2685 15600 2715
rect 15550 2665 15565 2685
rect 15585 2665 15600 2685
rect 15550 2650 15600 2665
rect 16150 3135 16200 3150
rect 16150 3115 16165 3135
rect 16185 3115 16200 3135
rect 16150 3085 16200 3115
rect 16150 3065 16165 3085
rect 16185 3065 16200 3085
rect 16150 3035 16200 3065
rect 16150 3015 16165 3035
rect 16185 3015 16200 3035
rect 16150 2985 16200 3015
rect 16150 2965 16165 2985
rect 16185 2965 16200 2985
rect 16150 2935 16200 2965
rect 16150 2915 16165 2935
rect 16185 2915 16200 2935
rect 16150 2885 16200 2915
rect 16150 2865 16165 2885
rect 16185 2865 16200 2885
rect 16150 2835 16200 2865
rect 16150 2815 16165 2835
rect 16185 2815 16200 2835
rect 16150 2785 16200 2815
rect 16150 2765 16165 2785
rect 16185 2765 16200 2785
rect 16150 2735 16200 2765
rect 16150 2715 16165 2735
rect 16185 2715 16200 2735
rect 16150 2685 16200 2715
rect 16150 2665 16165 2685
rect 16185 2665 16200 2685
rect 16150 2650 16200 2665
rect 16300 3135 16350 3150
rect 16300 3115 16315 3135
rect 16335 3115 16350 3135
rect 16300 3085 16350 3115
rect 16300 3065 16315 3085
rect 16335 3065 16350 3085
rect 16300 3035 16350 3065
rect 16300 3015 16315 3035
rect 16335 3015 16350 3035
rect 16300 2985 16350 3015
rect 16300 2965 16315 2985
rect 16335 2965 16350 2985
rect 16300 2935 16350 2965
rect 16300 2915 16315 2935
rect 16335 2915 16350 2935
rect 16300 2885 16350 2915
rect 16300 2865 16315 2885
rect 16335 2865 16350 2885
rect 16300 2835 16350 2865
rect 16300 2815 16315 2835
rect 16335 2815 16350 2835
rect 16300 2785 16350 2815
rect 16300 2765 16315 2785
rect 16335 2765 16350 2785
rect 16300 2735 16350 2765
rect 16300 2715 16315 2735
rect 16335 2715 16350 2735
rect 16300 2685 16350 2715
rect 16300 2665 16315 2685
rect 16335 2665 16350 2685
rect 16300 2650 16350 2665
rect 16450 3135 16500 3150
rect 16450 3115 16465 3135
rect 16485 3115 16500 3135
rect 16450 3085 16500 3115
rect 16450 3065 16465 3085
rect 16485 3065 16500 3085
rect 16450 3035 16500 3065
rect 16450 3015 16465 3035
rect 16485 3015 16500 3035
rect 16450 2985 16500 3015
rect 16450 2965 16465 2985
rect 16485 2965 16500 2985
rect 16450 2935 16500 2965
rect 16450 2915 16465 2935
rect 16485 2915 16500 2935
rect 16450 2885 16500 2915
rect 16450 2865 16465 2885
rect 16485 2865 16500 2885
rect 16450 2835 16500 2865
rect 16450 2815 16465 2835
rect 16485 2815 16500 2835
rect 16450 2785 16500 2815
rect 16450 2765 16465 2785
rect 16485 2765 16500 2785
rect 16450 2735 16500 2765
rect 16450 2715 16465 2735
rect 16485 2715 16500 2735
rect 16450 2685 16500 2715
rect 16450 2665 16465 2685
rect 16485 2665 16500 2685
rect 16450 2650 16500 2665
rect 16600 3135 16650 3150
rect 16600 3115 16615 3135
rect 16635 3115 16650 3135
rect 16600 3085 16650 3115
rect 16600 3065 16615 3085
rect 16635 3065 16650 3085
rect 16600 3035 16650 3065
rect 16600 3015 16615 3035
rect 16635 3015 16650 3035
rect 16600 2985 16650 3015
rect 16600 2965 16615 2985
rect 16635 2965 16650 2985
rect 16600 2935 16650 2965
rect 16600 2915 16615 2935
rect 16635 2915 16650 2935
rect 16600 2885 16650 2915
rect 16600 2865 16615 2885
rect 16635 2865 16650 2885
rect 16600 2835 16650 2865
rect 16600 2815 16615 2835
rect 16635 2815 16650 2835
rect 16600 2785 16650 2815
rect 16600 2765 16615 2785
rect 16635 2765 16650 2785
rect 16600 2735 16650 2765
rect 16600 2715 16615 2735
rect 16635 2715 16650 2735
rect 16600 2685 16650 2715
rect 16600 2665 16615 2685
rect 16635 2665 16650 2685
rect 16600 2650 16650 2665
rect 16750 3135 16800 3150
rect 16750 3115 16765 3135
rect 16785 3115 16800 3135
rect 16750 3085 16800 3115
rect 16750 3065 16765 3085
rect 16785 3065 16800 3085
rect 16750 3035 16800 3065
rect 16750 3015 16765 3035
rect 16785 3015 16800 3035
rect 16750 2985 16800 3015
rect 16750 2965 16765 2985
rect 16785 2965 16800 2985
rect 16750 2935 16800 2965
rect 16750 2915 16765 2935
rect 16785 2915 16800 2935
rect 16750 2885 16800 2915
rect 16750 2865 16765 2885
rect 16785 2865 16800 2885
rect 16750 2835 16800 2865
rect 16750 2815 16765 2835
rect 16785 2815 16800 2835
rect 16750 2785 16800 2815
rect 16750 2765 16765 2785
rect 16785 2765 16800 2785
rect 16750 2735 16800 2765
rect 16750 2715 16765 2735
rect 16785 2715 16800 2735
rect 16750 2685 16800 2715
rect 16750 2665 16765 2685
rect 16785 2665 16800 2685
rect 16750 2650 16800 2665
rect 16900 3135 16950 3150
rect 16900 3115 16915 3135
rect 16935 3115 16950 3135
rect 16900 3085 16950 3115
rect 16900 3065 16915 3085
rect 16935 3065 16950 3085
rect 16900 3035 16950 3065
rect 16900 3015 16915 3035
rect 16935 3015 16950 3035
rect 16900 2985 16950 3015
rect 16900 2965 16915 2985
rect 16935 2965 16950 2985
rect 16900 2935 16950 2965
rect 16900 2915 16915 2935
rect 16935 2915 16950 2935
rect 16900 2885 16950 2915
rect 16900 2865 16915 2885
rect 16935 2865 16950 2885
rect 16900 2835 16950 2865
rect 16900 2815 16915 2835
rect 16935 2815 16950 2835
rect 16900 2785 16950 2815
rect 16900 2765 16915 2785
rect 16935 2765 16950 2785
rect 16900 2735 16950 2765
rect 16900 2715 16915 2735
rect 16935 2715 16950 2735
rect 16900 2685 16950 2715
rect 16900 2665 16915 2685
rect 16935 2665 16950 2685
rect 16900 2650 16950 2665
rect 17050 3135 17100 3150
rect 17050 3115 17065 3135
rect 17085 3115 17100 3135
rect 17050 3085 17100 3115
rect 17050 3065 17065 3085
rect 17085 3065 17100 3085
rect 17050 3035 17100 3065
rect 17050 3015 17065 3035
rect 17085 3015 17100 3035
rect 17050 2985 17100 3015
rect 17050 2965 17065 2985
rect 17085 2965 17100 2985
rect 17050 2935 17100 2965
rect 17050 2915 17065 2935
rect 17085 2915 17100 2935
rect 17050 2885 17100 2915
rect 17050 2865 17065 2885
rect 17085 2865 17100 2885
rect 17050 2835 17100 2865
rect 17050 2815 17065 2835
rect 17085 2815 17100 2835
rect 17050 2785 17100 2815
rect 17050 2765 17065 2785
rect 17085 2765 17100 2785
rect 17050 2735 17100 2765
rect 17050 2715 17065 2735
rect 17085 2715 17100 2735
rect 17050 2685 17100 2715
rect 17050 2665 17065 2685
rect 17085 2665 17100 2685
rect 17050 2650 17100 2665
rect 17200 3135 17250 3150
rect 17200 3115 17215 3135
rect 17235 3115 17250 3135
rect 17200 3085 17250 3115
rect 17200 3065 17215 3085
rect 17235 3065 17250 3085
rect 17200 3035 17250 3065
rect 17200 3015 17215 3035
rect 17235 3015 17250 3035
rect 17200 2985 17250 3015
rect 17200 2965 17215 2985
rect 17235 2965 17250 2985
rect 17200 2935 17250 2965
rect 17200 2915 17215 2935
rect 17235 2915 17250 2935
rect 17200 2885 17250 2915
rect 17200 2865 17215 2885
rect 17235 2865 17250 2885
rect 17200 2835 17250 2865
rect 17200 2815 17215 2835
rect 17235 2815 17250 2835
rect 17200 2785 17250 2815
rect 17200 2765 17215 2785
rect 17235 2765 17250 2785
rect 17200 2735 17250 2765
rect 17200 2715 17215 2735
rect 17235 2715 17250 2735
rect 17200 2685 17250 2715
rect 17200 2665 17215 2685
rect 17235 2665 17250 2685
rect 17200 2650 17250 2665
rect 17350 3135 17400 3150
rect 17350 3115 17365 3135
rect 17385 3115 17400 3135
rect 17350 3085 17400 3115
rect 17350 3065 17365 3085
rect 17385 3065 17400 3085
rect 17350 3035 17400 3065
rect 17350 3015 17365 3035
rect 17385 3015 17400 3035
rect 17350 2985 17400 3015
rect 17350 2965 17365 2985
rect 17385 2965 17400 2985
rect 17350 2935 17400 2965
rect 17350 2915 17365 2935
rect 17385 2915 17400 2935
rect 17350 2885 17400 2915
rect 17350 2865 17365 2885
rect 17385 2865 17400 2885
rect 17350 2835 17400 2865
rect 17350 2815 17365 2835
rect 17385 2815 17400 2835
rect 17350 2785 17400 2815
rect 17350 2765 17365 2785
rect 17385 2765 17400 2785
rect 17350 2735 17400 2765
rect 17350 2715 17365 2735
rect 17385 2715 17400 2735
rect 17350 2685 17400 2715
rect 17350 2665 17365 2685
rect 17385 2665 17400 2685
rect 17350 2650 17400 2665
rect 17950 3135 18000 3150
rect 17950 3115 17965 3135
rect 17985 3115 18000 3135
rect 17950 3085 18000 3115
rect 17950 3065 17965 3085
rect 17985 3065 18000 3085
rect 17950 3035 18000 3065
rect 17950 3015 17965 3035
rect 17985 3015 18000 3035
rect 17950 2985 18000 3015
rect 17950 2965 17965 2985
rect 17985 2965 18000 2985
rect 17950 2935 18000 2965
rect 17950 2915 17965 2935
rect 17985 2915 18000 2935
rect 17950 2885 18000 2915
rect 17950 2865 17965 2885
rect 17985 2865 18000 2885
rect 17950 2835 18000 2865
rect 17950 2815 17965 2835
rect 17985 2815 18000 2835
rect 17950 2785 18000 2815
rect 17950 2765 17965 2785
rect 17985 2765 18000 2785
rect 17950 2735 18000 2765
rect 17950 2715 17965 2735
rect 17985 2715 18000 2735
rect 17950 2685 18000 2715
rect 17950 2665 17965 2685
rect 17985 2665 18000 2685
rect 17950 2650 18000 2665
rect 18550 3135 18600 3150
rect 18550 3115 18565 3135
rect 18585 3115 18600 3135
rect 18550 3085 18600 3115
rect 18550 3065 18565 3085
rect 18585 3065 18600 3085
rect 18550 3035 18600 3065
rect 18550 3015 18565 3035
rect 18585 3015 18600 3035
rect 18550 2985 18600 3015
rect 18550 2965 18565 2985
rect 18585 2965 18600 2985
rect 18550 2935 18600 2965
rect 18550 2915 18565 2935
rect 18585 2915 18600 2935
rect 18550 2885 18600 2915
rect 18550 2865 18565 2885
rect 18585 2865 18600 2885
rect 18550 2835 18600 2865
rect 18550 2815 18565 2835
rect 18585 2815 18600 2835
rect 18550 2785 18600 2815
rect 18550 2765 18565 2785
rect 18585 2765 18600 2785
rect 18550 2735 18600 2765
rect 18550 2715 18565 2735
rect 18585 2715 18600 2735
rect 18550 2685 18600 2715
rect 18550 2665 18565 2685
rect 18585 2665 18600 2685
rect 18550 2650 18600 2665
rect 18700 3135 18750 3150
rect 18700 3115 18715 3135
rect 18735 3115 18750 3135
rect 18700 3085 18750 3115
rect 18700 3065 18715 3085
rect 18735 3065 18750 3085
rect 18700 3035 18750 3065
rect 18700 3015 18715 3035
rect 18735 3015 18750 3035
rect 18700 2985 18750 3015
rect 18700 2965 18715 2985
rect 18735 2965 18750 2985
rect 18700 2935 18750 2965
rect 18700 2915 18715 2935
rect 18735 2915 18750 2935
rect 18700 2885 18750 2915
rect 18700 2865 18715 2885
rect 18735 2865 18750 2885
rect 18700 2835 18750 2865
rect 18700 2815 18715 2835
rect 18735 2815 18750 2835
rect 18700 2785 18750 2815
rect 18700 2765 18715 2785
rect 18735 2765 18750 2785
rect 18700 2735 18750 2765
rect 18700 2715 18715 2735
rect 18735 2715 18750 2735
rect 18700 2685 18750 2715
rect 18700 2665 18715 2685
rect 18735 2665 18750 2685
rect 18700 2650 18750 2665
rect 18850 3135 18900 3150
rect 18850 3115 18865 3135
rect 18885 3115 18900 3135
rect 18850 3085 18900 3115
rect 18850 3065 18865 3085
rect 18885 3065 18900 3085
rect 18850 3035 18900 3065
rect 18850 3015 18865 3035
rect 18885 3015 18900 3035
rect 18850 2985 18900 3015
rect 18850 2965 18865 2985
rect 18885 2965 18900 2985
rect 18850 2935 18900 2965
rect 18850 2915 18865 2935
rect 18885 2915 18900 2935
rect 18850 2885 18900 2915
rect 18850 2865 18865 2885
rect 18885 2865 18900 2885
rect 18850 2835 18900 2865
rect 18850 2815 18865 2835
rect 18885 2815 18900 2835
rect 18850 2785 18900 2815
rect 18850 2765 18865 2785
rect 18885 2765 18900 2785
rect 18850 2735 18900 2765
rect 18850 2715 18865 2735
rect 18885 2715 18900 2735
rect 18850 2685 18900 2715
rect 18850 2665 18865 2685
rect 18885 2665 18900 2685
rect 18850 2650 18900 2665
rect 19000 3135 19050 3150
rect 19000 3115 19015 3135
rect 19035 3115 19050 3135
rect 19000 3085 19050 3115
rect 19000 3065 19015 3085
rect 19035 3065 19050 3085
rect 19000 3035 19050 3065
rect 19000 3015 19015 3035
rect 19035 3015 19050 3035
rect 19000 2985 19050 3015
rect 19000 2965 19015 2985
rect 19035 2965 19050 2985
rect 19000 2935 19050 2965
rect 19000 2915 19015 2935
rect 19035 2915 19050 2935
rect 19000 2885 19050 2915
rect 19000 2865 19015 2885
rect 19035 2865 19050 2885
rect 19000 2835 19050 2865
rect 19000 2815 19015 2835
rect 19035 2815 19050 2835
rect 19000 2785 19050 2815
rect 19000 2765 19015 2785
rect 19035 2765 19050 2785
rect 19000 2735 19050 2765
rect 19000 2715 19015 2735
rect 19035 2715 19050 2735
rect 19000 2685 19050 2715
rect 19000 2665 19015 2685
rect 19035 2665 19050 2685
rect 19000 2650 19050 2665
rect 19150 3135 19200 3150
rect 19150 3115 19165 3135
rect 19185 3115 19200 3135
rect 19150 3085 19200 3115
rect 19150 3065 19165 3085
rect 19185 3065 19200 3085
rect 19150 3035 19200 3065
rect 19150 3015 19165 3035
rect 19185 3015 19200 3035
rect 19150 2985 19200 3015
rect 19150 2965 19165 2985
rect 19185 2965 19200 2985
rect 19150 2935 19200 2965
rect 19150 2915 19165 2935
rect 19185 2915 19200 2935
rect 19150 2885 19200 2915
rect 19150 2865 19165 2885
rect 19185 2865 19200 2885
rect 19150 2835 19200 2865
rect 19150 2815 19165 2835
rect 19185 2815 19200 2835
rect 19150 2785 19200 2815
rect 19150 2765 19165 2785
rect 19185 2765 19200 2785
rect 19150 2735 19200 2765
rect 19150 2715 19165 2735
rect 19185 2715 19200 2735
rect 19150 2685 19200 2715
rect 19150 2665 19165 2685
rect 19185 2665 19200 2685
rect 19150 2650 19200 2665
rect 19300 3135 19350 3150
rect 19300 3115 19315 3135
rect 19335 3115 19350 3135
rect 19300 3085 19350 3115
rect 19300 3065 19315 3085
rect 19335 3065 19350 3085
rect 19300 3035 19350 3065
rect 19300 3015 19315 3035
rect 19335 3015 19350 3035
rect 19300 2985 19350 3015
rect 19300 2965 19315 2985
rect 19335 2965 19350 2985
rect 19300 2935 19350 2965
rect 19300 2915 19315 2935
rect 19335 2915 19350 2935
rect 19300 2885 19350 2915
rect 19300 2865 19315 2885
rect 19335 2865 19350 2885
rect 19300 2835 19350 2865
rect 19300 2815 19315 2835
rect 19335 2815 19350 2835
rect 19300 2785 19350 2815
rect 19300 2765 19315 2785
rect 19335 2765 19350 2785
rect 19300 2735 19350 2765
rect 19300 2715 19315 2735
rect 19335 2715 19350 2735
rect 19300 2685 19350 2715
rect 19300 2665 19315 2685
rect 19335 2665 19350 2685
rect 19300 2650 19350 2665
rect 19450 3135 19500 3150
rect 19450 3115 19465 3135
rect 19485 3115 19500 3135
rect 19450 3085 19500 3115
rect 19450 3065 19465 3085
rect 19485 3065 19500 3085
rect 19450 3035 19500 3065
rect 19450 3015 19465 3035
rect 19485 3015 19500 3035
rect 19450 2985 19500 3015
rect 19450 2965 19465 2985
rect 19485 2965 19500 2985
rect 19450 2935 19500 2965
rect 19450 2915 19465 2935
rect 19485 2915 19500 2935
rect 19450 2885 19500 2915
rect 19450 2865 19465 2885
rect 19485 2865 19500 2885
rect 19450 2835 19500 2865
rect 19450 2815 19465 2835
rect 19485 2815 19500 2835
rect 19450 2785 19500 2815
rect 19450 2765 19465 2785
rect 19485 2765 19500 2785
rect 19450 2735 19500 2765
rect 19450 2715 19465 2735
rect 19485 2715 19500 2735
rect 19450 2685 19500 2715
rect 19450 2665 19465 2685
rect 19485 2665 19500 2685
rect 19450 2650 19500 2665
rect 19600 3135 19650 3150
rect 19600 3115 19615 3135
rect 19635 3115 19650 3135
rect 19600 3085 19650 3115
rect 19600 3065 19615 3085
rect 19635 3065 19650 3085
rect 19600 3035 19650 3065
rect 19600 3015 19615 3035
rect 19635 3015 19650 3035
rect 19600 2985 19650 3015
rect 19600 2965 19615 2985
rect 19635 2965 19650 2985
rect 19600 2935 19650 2965
rect 19600 2915 19615 2935
rect 19635 2915 19650 2935
rect 19600 2885 19650 2915
rect 19600 2865 19615 2885
rect 19635 2865 19650 2885
rect 19600 2835 19650 2865
rect 19600 2815 19615 2835
rect 19635 2815 19650 2835
rect 19600 2785 19650 2815
rect 19600 2765 19615 2785
rect 19635 2765 19650 2785
rect 19600 2735 19650 2765
rect 19600 2715 19615 2735
rect 19635 2715 19650 2735
rect 19600 2685 19650 2715
rect 19600 2665 19615 2685
rect 19635 2665 19650 2685
rect 19600 2650 19650 2665
rect 19750 3135 19800 3150
rect 19750 3115 19765 3135
rect 19785 3115 19800 3135
rect 19750 3085 19800 3115
rect 19750 3065 19765 3085
rect 19785 3065 19800 3085
rect 19750 3035 19800 3065
rect 19750 3015 19765 3035
rect 19785 3015 19800 3035
rect 19750 2985 19800 3015
rect 19750 2965 19765 2985
rect 19785 2965 19800 2985
rect 19750 2935 19800 2965
rect 19750 2915 19765 2935
rect 19785 2915 19800 2935
rect 19750 2885 19800 2915
rect 19750 2865 19765 2885
rect 19785 2865 19800 2885
rect 19750 2835 19800 2865
rect 19750 2815 19765 2835
rect 19785 2815 19800 2835
rect 19750 2785 19800 2815
rect 19750 2765 19765 2785
rect 19785 2765 19800 2785
rect 19750 2735 19800 2765
rect 19750 2715 19765 2735
rect 19785 2715 19800 2735
rect 19750 2685 19800 2715
rect 19750 2665 19765 2685
rect 19785 2665 19800 2685
rect 19750 2650 19800 2665
rect 20350 3135 20400 3150
rect 20350 3115 20365 3135
rect 20385 3115 20400 3135
rect 20350 3085 20400 3115
rect 20350 3065 20365 3085
rect 20385 3065 20400 3085
rect 20350 3035 20400 3065
rect 20350 3015 20365 3035
rect 20385 3015 20400 3035
rect 20350 2985 20400 3015
rect 20350 2965 20365 2985
rect 20385 2965 20400 2985
rect 20350 2935 20400 2965
rect 20350 2915 20365 2935
rect 20385 2915 20400 2935
rect 20350 2885 20400 2915
rect 20350 2865 20365 2885
rect 20385 2865 20400 2885
rect 20350 2835 20400 2865
rect 20350 2815 20365 2835
rect 20385 2815 20400 2835
rect 20350 2785 20400 2815
rect 20350 2765 20365 2785
rect 20385 2765 20400 2785
rect 20350 2735 20400 2765
rect 20350 2715 20365 2735
rect 20385 2715 20400 2735
rect 20350 2685 20400 2715
rect 20350 2665 20365 2685
rect 20385 2665 20400 2685
rect 20350 2650 20400 2665
rect -650 2585 20400 2600
rect -650 2565 -635 2585
rect -615 2565 -585 2585
rect -565 2565 -535 2585
rect -515 2565 -485 2585
rect -465 2565 -435 2585
rect -415 2565 -385 2585
rect -365 2565 -335 2585
rect -315 2565 -285 2585
rect -265 2565 -235 2585
rect -215 2565 -185 2585
rect -165 2565 -135 2585
rect -115 2565 -85 2585
rect -65 2565 -35 2585
rect -15 2565 15 2585
rect 35 2565 65 2585
rect 85 2565 115 2585
rect 135 2565 165 2585
rect 185 2565 215 2585
rect 235 2565 265 2585
rect 285 2565 315 2585
rect 335 2565 365 2585
rect 385 2565 415 2585
rect 435 2565 465 2585
rect 485 2565 515 2585
rect 535 2565 565 2585
rect 585 2565 615 2585
rect 635 2565 665 2585
rect 685 2565 715 2585
rect 735 2565 765 2585
rect 785 2565 815 2585
rect 835 2565 865 2585
rect 885 2565 915 2585
rect 935 2565 965 2585
rect 985 2565 1015 2585
rect 1035 2565 1065 2585
rect 1085 2565 1115 2585
rect 1135 2565 1165 2585
rect 1185 2565 1215 2585
rect 1235 2565 1265 2585
rect 1285 2565 1315 2585
rect 1335 2565 1365 2585
rect 1385 2565 1415 2585
rect 1435 2565 1465 2585
rect 1485 2565 1515 2585
rect 1535 2565 1565 2585
rect 1585 2565 1615 2585
rect 1635 2565 1665 2585
rect 1685 2565 1715 2585
rect 1735 2565 1765 2585
rect 1785 2565 1815 2585
rect 1835 2565 1865 2585
rect 1885 2565 1915 2585
rect 1935 2565 1965 2585
rect 1985 2565 2015 2585
rect 2035 2565 2065 2585
rect 2085 2565 2115 2585
rect 2135 2565 2165 2585
rect 2185 2565 2215 2585
rect 2235 2565 2265 2585
rect 2285 2565 2315 2585
rect 2335 2565 2365 2585
rect 2385 2565 2415 2585
rect 2435 2565 2465 2585
rect 2485 2565 2515 2585
rect 2535 2565 2565 2585
rect 2585 2565 2615 2585
rect 2635 2565 2665 2585
rect 2685 2565 2715 2585
rect 2735 2565 2765 2585
rect 2785 2565 2815 2585
rect 2835 2565 2865 2585
rect 2885 2565 2915 2585
rect 2935 2565 2965 2585
rect 2985 2565 3015 2585
rect 3035 2565 3065 2585
rect 3085 2565 3115 2585
rect 3135 2565 3165 2585
rect 3185 2565 3215 2585
rect 3235 2565 3265 2585
rect 3285 2565 3315 2585
rect 3335 2565 3365 2585
rect 3385 2565 3415 2585
rect 3435 2565 3465 2585
rect 3485 2565 3515 2585
rect 3535 2565 3565 2585
rect 3585 2565 3615 2585
rect 3635 2565 3665 2585
rect 3685 2565 3715 2585
rect 3735 2565 3765 2585
rect 3785 2565 3815 2585
rect 3835 2565 3865 2585
rect 3885 2565 3915 2585
rect 3935 2565 3965 2585
rect 3985 2565 4015 2585
rect 4035 2565 4065 2585
rect 4085 2565 4115 2585
rect 4135 2565 4165 2585
rect 4185 2565 4215 2585
rect 4235 2565 4265 2585
rect 4285 2565 4315 2585
rect 4335 2565 4365 2585
rect 4385 2565 4415 2585
rect 4435 2565 4465 2585
rect 4485 2565 4515 2585
rect 4535 2565 4565 2585
rect 4585 2565 4615 2585
rect 4635 2565 4665 2585
rect 4685 2565 4715 2585
rect 4735 2565 4765 2585
rect 4785 2565 4815 2585
rect 4835 2565 4865 2585
rect 4885 2565 4915 2585
rect 4935 2565 4965 2585
rect 4985 2565 5015 2585
rect 5035 2565 5065 2585
rect 5085 2565 5115 2585
rect 5135 2565 5165 2585
rect 5185 2565 5215 2585
rect 5235 2565 5265 2585
rect 5285 2565 5315 2585
rect 5335 2565 5365 2585
rect 5385 2565 5415 2585
rect 5435 2565 5465 2585
rect 5485 2565 5515 2585
rect 5535 2565 5565 2585
rect 5585 2565 5615 2585
rect 5635 2565 5665 2585
rect 5685 2565 5715 2585
rect 5735 2565 5765 2585
rect 5785 2565 5815 2585
rect 5835 2565 5865 2585
rect 5885 2565 5915 2585
rect 5935 2565 5965 2585
rect 5985 2565 6015 2585
rect 6035 2565 6065 2585
rect 6085 2565 6115 2585
rect 6135 2565 6165 2585
rect 6185 2565 6215 2585
rect 6235 2565 6265 2585
rect 6285 2565 6315 2585
rect 6335 2565 6365 2585
rect 6385 2565 6415 2585
rect 6435 2565 6465 2585
rect 6485 2565 6515 2585
rect 6535 2565 6565 2585
rect 6585 2565 6615 2585
rect 6635 2565 6665 2585
rect 6685 2565 6715 2585
rect 6735 2565 6765 2585
rect 6785 2565 6815 2585
rect 6835 2565 6865 2585
rect 6885 2565 6915 2585
rect 6935 2565 6965 2585
rect 6985 2565 7015 2585
rect 7035 2565 7065 2585
rect 7085 2565 7115 2585
rect 7135 2565 7165 2585
rect 7185 2565 7215 2585
rect 7235 2565 7265 2585
rect 7285 2565 7315 2585
rect 7335 2565 7365 2585
rect 7385 2565 7415 2585
rect 7435 2565 7465 2585
rect 7485 2565 7515 2585
rect 7535 2565 7565 2585
rect 7585 2565 7615 2585
rect 7635 2565 7665 2585
rect 7685 2565 7715 2585
rect 7735 2565 7765 2585
rect 7785 2565 7815 2585
rect 7835 2565 7865 2585
rect 7885 2565 7915 2585
rect 7935 2565 7965 2585
rect 7985 2565 8015 2585
rect 8035 2565 8065 2585
rect 8085 2565 8115 2585
rect 8135 2565 8165 2585
rect 8185 2565 8215 2585
rect 8235 2565 8265 2585
rect 8285 2565 8315 2585
rect 8335 2565 8365 2585
rect 8385 2565 8415 2585
rect 8435 2565 8465 2585
rect 8485 2565 8515 2585
rect 8535 2565 8565 2585
rect 8585 2565 8615 2585
rect 8635 2565 8665 2585
rect 8685 2565 8715 2585
rect 8735 2565 8765 2585
rect 8785 2565 8815 2585
rect 8835 2565 8865 2585
rect 8885 2565 8915 2585
rect 8935 2565 8965 2585
rect 8985 2565 9015 2585
rect 9035 2565 9065 2585
rect 9085 2565 9115 2585
rect 9135 2565 9165 2585
rect 9185 2565 9215 2585
rect 9235 2565 9265 2585
rect 9285 2565 9315 2585
rect 9335 2565 9365 2585
rect 9385 2565 9415 2585
rect 9435 2565 9465 2585
rect 9485 2565 9515 2585
rect 9535 2565 9565 2585
rect 9585 2565 9615 2585
rect 9635 2565 9665 2585
rect 9685 2565 9715 2585
rect 9735 2565 9765 2585
rect 9785 2565 9815 2585
rect 9835 2565 9865 2585
rect 9885 2565 9915 2585
rect 9935 2565 9965 2585
rect 9985 2565 10015 2585
rect 10035 2565 10065 2585
rect 10085 2565 10115 2585
rect 10135 2565 10165 2585
rect 10185 2565 10215 2585
rect 10235 2565 10265 2585
rect 10285 2565 10315 2585
rect 10335 2565 10365 2585
rect 10385 2565 10415 2585
rect 10435 2565 10465 2585
rect 10485 2565 10515 2585
rect 10535 2565 10565 2585
rect 10585 2565 10615 2585
rect 10635 2565 10665 2585
rect 10685 2565 10715 2585
rect 10735 2565 10765 2585
rect 10785 2565 10815 2585
rect 10835 2565 10865 2585
rect 10885 2565 10915 2585
rect 10935 2565 10965 2585
rect 10985 2565 11015 2585
rect 11035 2565 11065 2585
rect 11085 2565 11115 2585
rect 11135 2565 11165 2585
rect 11185 2565 11215 2585
rect 11235 2565 11265 2585
rect 11285 2565 11315 2585
rect 11335 2565 11365 2585
rect 11385 2565 11415 2585
rect 11435 2565 11465 2585
rect 11485 2565 11515 2585
rect 11535 2565 11565 2585
rect 11585 2565 11615 2585
rect 11635 2565 11665 2585
rect 11685 2565 11715 2585
rect 11735 2565 11765 2585
rect 11785 2565 11815 2585
rect 11835 2565 11865 2585
rect 11885 2565 11915 2585
rect 11935 2565 11965 2585
rect 11985 2565 12015 2585
rect 12035 2565 12065 2585
rect 12085 2565 12115 2585
rect 12135 2565 12165 2585
rect 12185 2565 12215 2585
rect 12235 2565 12265 2585
rect 12285 2565 12315 2585
rect 12335 2565 12365 2585
rect 12385 2565 12415 2585
rect 12435 2565 12465 2585
rect 12485 2565 12515 2585
rect 12535 2565 12565 2585
rect 12585 2565 12615 2585
rect 12635 2565 12665 2585
rect 12685 2565 12715 2585
rect 12735 2565 12765 2585
rect 12785 2565 12815 2585
rect 12835 2565 12865 2585
rect 12885 2565 12915 2585
rect 12935 2565 12965 2585
rect 12985 2565 13015 2585
rect 13035 2565 13065 2585
rect 13085 2565 13115 2585
rect 13135 2565 13165 2585
rect 13185 2565 13215 2585
rect 13235 2565 13265 2585
rect 13285 2565 13315 2585
rect 13335 2565 13365 2585
rect 13385 2565 13415 2585
rect 13435 2565 13465 2585
rect 13485 2565 13515 2585
rect 13535 2565 13565 2585
rect 13585 2565 13615 2585
rect 13635 2565 13665 2585
rect 13685 2565 13715 2585
rect 13735 2565 13765 2585
rect 13785 2565 13815 2585
rect 13835 2565 13865 2585
rect 13885 2565 13915 2585
rect 13935 2565 13965 2585
rect 13985 2565 14015 2585
rect 14035 2565 14065 2585
rect 14085 2565 14115 2585
rect 14135 2565 14165 2585
rect 14185 2565 14215 2585
rect 14235 2565 14265 2585
rect 14285 2565 14315 2585
rect 14335 2565 14365 2585
rect 14385 2565 14415 2585
rect 14435 2565 14465 2585
rect 14485 2565 14515 2585
rect 14535 2565 14565 2585
rect 14585 2565 14615 2585
rect 14635 2565 14665 2585
rect 14685 2565 14715 2585
rect 14735 2565 14765 2585
rect 14785 2565 14815 2585
rect 14835 2565 14865 2585
rect 14885 2565 14915 2585
rect 14935 2565 14965 2585
rect 14985 2565 15015 2585
rect 15035 2565 15065 2585
rect 15085 2565 15115 2585
rect 15135 2565 15165 2585
rect 15185 2565 15215 2585
rect 15235 2565 15265 2585
rect 15285 2565 15315 2585
rect 15335 2565 15365 2585
rect 15385 2565 15415 2585
rect 15435 2565 15465 2585
rect 15485 2565 15515 2585
rect 15535 2565 15565 2585
rect 15585 2565 15615 2585
rect 15635 2565 15665 2585
rect 15685 2565 15715 2585
rect 15735 2565 15765 2585
rect 15785 2565 15815 2585
rect 15835 2565 15865 2585
rect 15885 2565 15915 2585
rect 15935 2565 15965 2585
rect 15985 2565 16015 2585
rect 16035 2565 16065 2585
rect 16085 2565 16115 2585
rect 16135 2565 16165 2585
rect 16185 2565 16215 2585
rect 16235 2565 16265 2585
rect 16285 2565 16315 2585
rect 16335 2565 16365 2585
rect 16385 2565 16415 2585
rect 16435 2565 16465 2585
rect 16485 2565 16515 2585
rect 16535 2565 16565 2585
rect 16585 2565 16615 2585
rect 16635 2565 16665 2585
rect 16685 2565 16715 2585
rect 16735 2565 16765 2585
rect 16785 2565 16815 2585
rect 16835 2565 16865 2585
rect 16885 2565 16915 2585
rect 16935 2565 16965 2585
rect 16985 2565 17015 2585
rect 17035 2565 17065 2585
rect 17085 2565 17115 2585
rect 17135 2565 17165 2585
rect 17185 2565 17215 2585
rect 17235 2565 17265 2585
rect 17285 2565 17315 2585
rect 17335 2565 17365 2585
rect 17385 2565 17415 2585
rect 17435 2565 17465 2585
rect 17485 2565 17515 2585
rect 17535 2565 17565 2585
rect 17585 2565 17615 2585
rect 17635 2565 17665 2585
rect 17685 2565 17715 2585
rect 17735 2565 17765 2585
rect 17785 2565 17815 2585
rect 17835 2565 17865 2585
rect 17885 2565 17915 2585
rect 17935 2565 17965 2585
rect 17985 2565 18015 2585
rect 18035 2565 18065 2585
rect 18085 2565 18115 2585
rect 18135 2565 18165 2585
rect 18185 2565 18215 2585
rect 18235 2565 18265 2585
rect 18285 2565 18315 2585
rect 18335 2565 18365 2585
rect 18385 2565 18415 2585
rect 18435 2565 18465 2585
rect 18485 2565 18515 2585
rect 18535 2565 18565 2585
rect 18585 2565 18615 2585
rect 18635 2565 18665 2585
rect 18685 2565 18715 2585
rect 18735 2565 18765 2585
rect 18785 2565 18815 2585
rect 18835 2565 18865 2585
rect 18885 2565 18915 2585
rect 18935 2565 18965 2585
rect 18985 2565 19015 2585
rect 19035 2565 19065 2585
rect 19085 2565 19115 2585
rect 19135 2565 19165 2585
rect 19185 2565 19215 2585
rect 19235 2565 19265 2585
rect 19285 2565 19315 2585
rect 19335 2565 19365 2585
rect 19385 2565 19415 2585
rect 19435 2565 19465 2585
rect 19485 2565 19515 2585
rect 19535 2565 19565 2585
rect 19585 2565 19615 2585
rect 19635 2565 19665 2585
rect 19685 2565 19715 2585
rect 19735 2565 19765 2585
rect 19785 2565 19815 2585
rect 19835 2565 19865 2585
rect 19885 2565 19915 2585
rect 19935 2565 19965 2585
rect 19985 2565 20015 2585
rect 20035 2565 20065 2585
rect 20085 2565 20115 2585
rect 20135 2565 20165 2585
rect 20185 2565 20215 2585
rect 20235 2565 20265 2585
rect 20285 2565 20315 2585
rect 20335 2565 20365 2585
rect 20385 2565 20400 2585
rect -650 2550 20400 2565
rect -900 2435 20400 2450
rect -900 2415 -885 2435
rect -865 2415 -835 2435
rect -815 2415 -785 2435
rect -765 2415 -735 2435
rect -715 2415 -685 2435
rect -665 2415 -635 2435
rect -615 2415 -585 2435
rect -565 2415 -535 2435
rect -515 2415 -485 2435
rect -465 2415 -435 2435
rect -415 2415 -385 2435
rect -365 2415 -335 2435
rect -315 2415 -285 2435
rect -265 2415 -235 2435
rect -215 2415 -185 2435
rect -165 2415 -135 2435
rect -115 2415 -85 2435
rect -65 2415 -35 2435
rect -15 2415 15 2435
rect 35 2415 65 2435
rect 85 2415 115 2435
rect 135 2415 165 2435
rect 185 2415 215 2435
rect 235 2415 265 2435
rect 285 2415 315 2435
rect 335 2415 365 2435
rect 385 2415 415 2435
rect 435 2415 465 2435
rect 485 2415 515 2435
rect 535 2415 565 2435
rect 585 2415 615 2435
rect 635 2415 665 2435
rect 685 2415 715 2435
rect 735 2415 765 2435
rect 785 2415 815 2435
rect 835 2415 865 2435
rect 885 2415 915 2435
rect 935 2415 965 2435
rect 985 2415 1015 2435
rect 1035 2415 1065 2435
rect 1085 2415 1115 2435
rect 1135 2415 1165 2435
rect 1185 2415 1215 2435
rect 1235 2415 1265 2435
rect 1285 2415 1315 2435
rect 1335 2415 1365 2435
rect 1385 2415 1415 2435
rect 1435 2415 1465 2435
rect 1485 2415 1515 2435
rect 1535 2415 1565 2435
rect 1585 2415 1615 2435
rect 1635 2415 1665 2435
rect 1685 2415 1715 2435
rect 1735 2415 1765 2435
rect 1785 2415 1815 2435
rect 1835 2415 1865 2435
rect 1885 2415 1915 2435
rect 1935 2415 1965 2435
rect 1985 2415 2015 2435
rect 2035 2415 2065 2435
rect 2085 2415 2115 2435
rect 2135 2415 2165 2435
rect 2185 2415 2215 2435
rect 2235 2415 2265 2435
rect 2285 2415 2315 2435
rect 2335 2415 2365 2435
rect 2385 2415 2415 2435
rect 2435 2415 2465 2435
rect 2485 2415 2515 2435
rect 2535 2415 2565 2435
rect 2585 2415 2615 2435
rect 2635 2415 2665 2435
rect 2685 2415 2715 2435
rect 2735 2415 2765 2435
rect 2785 2415 2815 2435
rect 2835 2415 2865 2435
rect 2885 2415 2915 2435
rect 2935 2415 2965 2435
rect 2985 2415 3015 2435
rect 3035 2415 3065 2435
rect 3085 2415 3115 2435
rect 3135 2415 3165 2435
rect 3185 2415 3215 2435
rect 3235 2415 3265 2435
rect 3285 2415 3315 2435
rect 3335 2415 3365 2435
rect 3385 2415 3415 2435
rect 3435 2415 3465 2435
rect 3485 2415 3515 2435
rect 3535 2415 3565 2435
rect 3585 2415 3615 2435
rect 3635 2415 3665 2435
rect 3685 2415 3715 2435
rect 3735 2415 3765 2435
rect 3785 2415 3815 2435
rect 3835 2415 3865 2435
rect 3885 2415 3915 2435
rect 3935 2415 3965 2435
rect 3985 2415 4015 2435
rect 4035 2415 4065 2435
rect 4085 2415 4115 2435
rect 4135 2415 4165 2435
rect 4185 2415 4215 2435
rect 4235 2415 4265 2435
rect 4285 2415 4315 2435
rect 4335 2415 4365 2435
rect 4385 2415 4415 2435
rect 4435 2415 4465 2435
rect 4485 2415 4515 2435
rect 4535 2415 4565 2435
rect 4585 2415 4615 2435
rect 4635 2415 4665 2435
rect 4685 2415 4715 2435
rect 4735 2415 4765 2435
rect 4785 2415 4815 2435
rect 4835 2415 4865 2435
rect 4885 2415 4915 2435
rect 4935 2415 4965 2435
rect 4985 2415 5015 2435
rect 5035 2415 5065 2435
rect 5085 2415 5115 2435
rect 5135 2415 5165 2435
rect 5185 2415 5215 2435
rect 5235 2415 5265 2435
rect 5285 2415 5315 2435
rect 5335 2415 5365 2435
rect 5385 2415 5415 2435
rect 5435 2415 5465 2435
rect 5485 2415 5515 2435
rect 5535 2415 5565 2435
rect 5585 2415 5615 2435
rect 5635 2415 5665 2435
rect 5685 2415 5715 2435
rect 5735 2415 5765 2435
rect 5785 2415 5815 2435
rect 5835 2415 5865 2435
rect 5885 2415 5915 2435
rect 5935 2415 5965 2435
rect 5985 2415 6015 2435
rect 6035 2415 6065 2435
rect 6085 2415 6115 2435
rect 6135 2415 6165 2435
rect 6185 2415 6215 2435
rect 6235 2415 6265 2435
rect 6285 2415 6315 2435
rect 6335 2415 6365 2435
rect 6385 2415 6415 2435
rect 6435 2415 6465 2435
rect 6485 2415 6515 2435
rect 6535 2415 6565 2435
rect 6585 2415 6615 2435
rect 6635 2415 6665 2435
rect 6685 2415 6715 2435
rect 6735 2415 6765 2435
rect 6785 2415 6815 2435
rect 6835 2415 6865 2435
rect 6885 2415 6915 2435
rect 6935 2415 6965 2435
rect 6985 2415 7015 2435
rect 7035 2415 7065 2435
rect 7085 2415 7115 2435
rect 7135 2415 7165 2435
rect 7185 2415 7215 2435
rect 7235 2415 7265 2435
rect 7285 2415 7315 2435
rect 7335 2415 7365 2435
rect 7385 2415 7415 2435
rect 7435 2415 7465 2435
rect 7485 2415 7515 2435
rect 7535 2415 7565 2435
rect 7585 2415 7615 2435
rect 7635 2415 7665 2435
rect 7685 2415 7715 2435
rect 7735 2415 7765 2435
rect 7785 2415 7815 2435
rect 7835 2415 7865 2435
rect 7885 2415 7915 2435
rect 7935 2415 7965 2435
rect 7985 2415 8015 2435
rect 8035 2415 8065 2435
rect 8085 2415 8115 2435
rect 8135 2415 8165 2435
rect 8185 2415 8215 2435
rect 8235 2415 8265 2435
rect 8285 2415 8315 2435
rect 8335 2415 8365 2435
rect 8385 2415 8415 2435
rect 8435 2415 8465 2435
rect 8485 2415 8515 2435
rect 8535 2415 8565 2435
rect 8585 2415 8615 2435
rect 8635 2415 8665 2435
rect 8685 2415 8715 2435
rect 8735 2415 8765 2435
rect 8785 2415 8815 2435
rect 8835 2415 8865 2435
rect 8885 2415 8915 2435
rect 8935 2415 8965 2435
rect 8985 2415 9015 2435
rect 9035 2415 9065 2435
rect 9085 2415 9115 2435
rect 9135 2415 9165 2435
rect 9185 2415 9215 2435
rect 9235 2415 9265 2435
rect 9285 2415 9315 2435
rect 9335 2415 9365 2435
rect 9385 2415 9415 2435
rect 9435 2415 9465 2435
rect 9485 2415 9515 2435
rect 9535 2415 9565 2435
rect 9585 2415 9615 2435
rect 9635 2415 9665 2435
rect 9685 2415 9715 2435
rect 9735 2415 9765 2435
rect 9785 2415 9815 2435
rect 9835 2415 9865 2435
rect 9885 2415 9915 2435
rect 9935 2415 9965 2435
rect 9985 2415 10015 2435
rect 10035 2415 10065 2435
rect 10085 2415 10115 2435
rect 10135 2415 10165 2435
rect 10185 2415 10215 2435
rect 10235 2415 10265 2435
rect 10285 2415 10315 2435
rect 10335 2415 10365 2435
rect 10385 2415 10415 2435
rect 10435 2415 10465 2435
rect 10485 2415 10515 2435
rect 10535 2415 10565 2435
rect 10585 2415 10615 2435
rect 10635 2415 10665 2435
rect 10685 2415 10715 2435
rect 10735 2415 10765 2435
rect 10785 2415 10815 2435
rect 10835 2415 10865 2435
rect 10885 2415 10915 2435
rect 10935 2415 10965 2435
rect 10985 2415 11015 2435
rect 11035 2415 11065 2435
rect 11085 2415 11115 2435
rect 11135 2415 11165 2435
rect 11185 2415 11215 2435
rect 11235 2415 11265 2435
rect 11285 2415 11315 2435
rect 11335 2415 11365 2435
rect 11385 2415 11415 2435
rect 11435 2415 11465 2435
rect 11485 2415 11515 2435
rect 11535 2415 11565 2435
rect 11585 2415 11615 2435
rect 11635 2415 11665 2435
rect 11685 2415 11715 2435
rect 11735 2415 11765 2435
rect 11785 2415 11815 2435
rect 11835 2415 11865 2435
rect 11885 2415 11915 2435
rect 11935 2415 11965 2435
rect 11985 2415 12015 2435
rect 12035 2415 12065 2435
rect 12085 2415 12115 2435
rect 12135 2415 12165 2435
rect 12185 2415 12215 2435
rect 12235 2415 12265 2435
rect 12285 2415 12315 2435
rect 12335 2415 12365 2435
rect 12385 2415 12415 2435
rect 12435 2415 12465 2435
rect 12485 2415 12515 2435
rect 12535 2415 12565 2435
rect 12585 2415 12615 2435
rect 12635 2415 12665 2435
rect 12685 2415 12715 2435
rect 12735 2415 12765 2435
rect 12785 2415 12815 2435
rect 12835 2415 12865 2435
rect 12885 2415 12915 2435
rect 12935 2415 12965 2435
rect 12985 2415 13015 2435
rect 13035 2415 13065 2435
rect 13085 2415 13115 2435
rect 13135 2415 13165 2435
rect 13185 2415 13215 2435
rect 13235 2415 13265 2435
rect 13285 2415 13315 2435
rect 13335 2415 13365 2435
rect 13385 2415 13415 2435
rect 13435 2415 13465 2435
rect 13485 2415 13515 2435
rect 13535 2415 13565 2435
rect 13585 2415 13615 2435
rect 13635 2415 13665 2435
rect 13685 2415 13715 2435
rect 13735 2415 13765 2435
rect 13785 2415 13815 2435
rect 13835 2415 13865 2435
rect 13885 2415 13915 2435
rect 13935 2415 13965 2435
rect 13985 2415 14015 2435
rect 14035 2415 14065 2435
rect 14085 2415 14115 2435
rect 14135 2415 14165 2435
rect 14185 2415 14215 2435
rect 14235 2415 14265 2435
rect 14285 2415 14315 2435
rect 14335 2415 14365 2435
rect 14385 2415 14415 2435
rect 14435 2415 14465 2435
rect 14485 2415 14515 2435
rect 14535 2415 14565 2435
rect 14585 2415 14615 2435
rect 14635 2415 14665 2435
rect 14685 2415 14715 2435
rect 14735 2415 14765 2435
rect 14785 2415 14815 2435
rect 14835 2415 14865 2435
rect 14885 2415 14915 2435
rect 14935 2415 14965 2435
rect 14985 2415 15015 2435
rect 15035 2415 15065 2435
rect 15085 2415 15115 2435
rect 15135 2415 15165 2435
rect 15185 2415 15215 2435
rect 15235 2415 15265 2435
rect 15285 2415 15315 2435
rect 15335 2415 15365 2435
rect 15385 2415 15415 2435
rect 15435 2415 15465 2435
rect 15485 2415 15515 2435
rect 15535 2415 15565 2435
rect 15585 2415 15615 2435
rect 15635 2415 15665 2435
rect 15685 2415 15715 2435
rect 15735 2415 15765 2435
rect 15785 2415 15815 2435
rect 15835 2415 15865 2435
rect 15885 2415 15915 2435
rect 15935 2415 15965 2435
rect 15985 2415 16015 2435
rect 16035 2415 16065 2435
rect 16085 2415 16115 2435
rect 16135 2415 16165 2435
rect 16185 2415 16215 2435
rect 16235 2415 16265 2435
rect 16285 2415 16315 2435
rect 16335 2415 16365 2435
rect 16385 2415 16415 2435
rect 16435 2415 16465 2435
rect 16485 2415 16515 2435
rect 16535 2415 16565 2435
rect 16585 2415 16615 2435
rect 16635 2415 16665 2435
rect 16685 2415 16715 2435
rect 16735 2415 16765 2435
rect 16785 2415 16815 2435
rect 16835 2415 16865 2435
rect 16885 2415 16915 2435
rect 16935 2415 16965 2435
rect 16985 2415 17015 2435
rect 17035 2415 17065 2435
rect 17085 2415 17115 2435
rect 17135 2415 17165 2435
rect 17185 2415 17215 2435
rect 17235 2415 17265 2435
rect 17285 2415 17315 2435
rect 17335 2415 17365 2435
rect 17385 2415 17415 2435
rect 17435 2415 17465 2435
rect 17485 2415 17515 2435
rect 17535 2415 17565 2435
rect 17585 2415 17615 2435
rect 17635 2415 17665 2435
rect 17685 2415 17715 2435
rect 17735 2415 17765 2435
rect 17785 2415 17815 2435
rect 17835 2415 17865 2435
rect 17885 2415 17915 2435
rect 17935 2415 17965 2435
rect 17985 2415 18015 2435
rect 18035 2415 18065 2435
rect 18085 2415 18115 2435
rect 18135 2415 18165 2435
rect 18185 2415 18215 2435
rect 18235 2415 18265 2435
rect 18285 2415 18315 2435
rect 18335 2415 18365 2435
rect 18385 2415 18415 2435
rect 18435 2415 18465 2435
rect 18485 2415 18515 2435
rect 18535 2415 18565 2435
rect 18585 2415 18615 2435
rect 18635 2415 18665 2435
rect 18685 2415 18715 2435
rect 18735 2415 18765 2435
rect 18785 2415 18815 2435
rect 18835 2415 18865 2435
rect 18885 2415 18915 2435
rect 18935 2415 18965 2435
rect 18985 2415 19015 2435
rect 19035 2415 19065 2435
rect 19085 2415 19115 2435
rect 19135 2415 19165 2435
rect 19185 2415 19215 2435
rect 19235 2415 19265 2435
rect 19285 2415 19315 2435
rect 19335 2415 19365 2435
rect 19385 2415 19415 2435
rect 19435 2415 19465 2435
rect 19485 2415 19515 2435
rect 19535 2415 19565 2435
rect 19585 2415 19615 2435
rect 19635 2415 19665 2435
rect 19685 2415 19715 2435
rect 19735 2415 19765 2435
rect 19785 2415 19815 2435
rect 19835 2415 19865 2435
rect 19885 2415 19915 2435
rect 19935 2415 19965 2435
rect 19985 2415 20015 2435
rect 20035 2415 20065 2435
rect 20085 2415 20115 2435
rect 20135 2415 20165 2435
rect 20185 2415 20215 2435
rect 20235 2415 20265 2435
rect 20285 2415 20315 2435
rect 20335 2415 20365 2435
rect 20385 2415 20400 2435
rect -900 2400 20400 2415
rect -900 2035 20400 2050
rect -900 2015 -885 2035
rect -865 2015 -835 2035
rect -815 2015 -785 2035
rect -765 2015 -735 2035
rect -715 2015 -685 2035
rect -665 2015 -635 2035
rect -615 2015 -585 2035
rect -565 2015 -535 2035
rect -515 2015 -485 2035
rect -465 2015 -435 2035
rect -415 2015 -385 2035
rect -365 2015 -335 2035
rect -315 2015 -285 2035
rect -265 2015 -235 2035
rect -215 2015 -185 2035
rect -165 2015 -135 2035
rect -115 2015 -85 2035
rect -65 2015 -35 2035
rect -15 2015 15 2035
rect 35 2015 65 2035
rect 85 2015 115 2035
rect 135 2015 165 2035
rect 185 2015 215 2035
rect 235 2015 265 2035
rect 285 2015 315 2035
rect 335 2015 365 2035
rect 385 2015 415 2035
rect 435 2015 465 2035
rect 485 2015 515 2035
rect 535 2015 565 2035
rect 585 2015 615 2035
rect 635 2015 665 2035
rect 685 2015 715 2035
rect 735 2015 765 2035
rect 785 2015 815 2035
rect 835 2015 865 2035
rect 885 2015 915 2035
rect 935 2015 965 2035
rect 985 2015 1015 2035
rect 1035 2015 1065 2035
rect 1085 2015 1115 2035
rect 1135 2015 1165 2035
rect 1185 2015 1215 2035
rect 1235 2015 1265 2035
rect 1285 2015 1315 2035
rect 1335 2015 1365 2035
rect 1385 2015 1415 2035
rect 1435 2015 1465 2035
rect 1485 2015 1515 2035
rect 1535 2015 1565 2035
rect 1585 2015 1615 2035
rect 1635 2015 1665 2035
rect 1685 2015 1715 2035
rect 1735 2015 1765 2035
rect 1785 2015 1815 2035
rect 1835 2015 1865 2035
rect 1885 2015 1915 2035
rect 1935 2015 1965 2035
rect 1985 2015 2015 2035
rect 2035 2015 2065 2035
rect 2085 2015 2115 2035
rect 2135 2015 2165 2035
rect 2185 2015 2215 2035
rect 2235 2015 2265 2035
rect 2285 2015 2315 2035
rect 2335 2015 2365 2035
rect 2385 2015 2415 2035
rect 2435 2015 2465 2035
rect 2485 2015 2515 2035
rect 2535 2015 2565 2035
rect 2585 2015 2615 2035
rect 2635 2015 2665 2035
rect 2685 2015 2715 2035
rect 2735 2015 2765 2035
rect 2785 2015 2815 2035
rect 2835 2015 2865 2035
rect 2885 2015 2915 2035
rect 2935 2015 2965 2035
rect 2985 2015 3015 2035
rect 3035 2015 3065 2035
rect 3085 2015 3115 2035
rect 3135 2015 3165 2035
rect 3185 2015 3215 2035
rect 3235 2015 3265 2035
rect 3285 2015 3315 2035
rect 3335 2015 3365 2035
rect 3385 2015 3415 2035
rect 3435 2015 3465 2035
rect 3485 2015 3515 2035
rect 3535 2015 3565 2035
rect 3585 2015 3615 2035
rect 3635 2015 3665 2035
rect 3685 2015 3715 2035
rect 3735 2015 3765 2035
rect 3785 2015 3815 2035
rect 3835 2015 3865 2035
rect 3885 2015 3915 2035
rect 3935 2015 3965 2035
rect 3985 2015 4015 2035
rect 4035 2015 4065 2035
rect 4085 2015 4115 2035
rect 4135 2015 4165 2035
rect 4185 2015 4215 2035
rect 4235 2015 4265 2035
rect 4285 2015 4315 2035
rect 4335 2015 4365 2035
rect 4385 2015 4415 2035
rect 4435 2015 4465 2035
rect 4485 2015 4515 2035
rect 4535 2015 4565 2035
rect 4585 2015 4615 2035
rect 4635 2015 4665 2035
rect 4685 2015 4715 2035
rect 4735 2015 4765 2035
rect 4785 2015 4815 2035
rect 4835 2015 4865 2035
rect 4885 2015 4915 2035
rect 4935 2015 4965 2035
rect 4985 2015 5015 2035
rect 5035 2015 5065 2035
rect 5085 2015 5115 2035
rect 5135 2015 5165 2035
rect 5185 2015 5215 2035
rect 5235 2015 5265 2035
rect 5285 2015 5315 2035
rect 5335 2015 5365 2035
rect 5385 2015 5415 2035
rect 5435 2015 5465 2035
rect 5485 2015 5515 2035
rect 5535 2015 5565 2035
rect 5585 2015 5615 2035
rect 5635 2015 5665 2035
rect 5685 2015 5715 2035
rect 5735 2015 5765 2035
rect 5785 2015 5815 2035
rect 5835 2015 5865 2035
rect 5885 2015 5915 2035
rect 5935 2015 5965 2035
rect 5985 2015 6015 2035
rect 6035 2015 6065 2035
rect 6085 2015 6115 2035
rect 6135 2015 6165 2035
rect 6185 2015 6215 2035
rect 6235 2015 6265 2035
rect 6285 2015 6315 2035
rect 6335 2015 6365 2035
rect 6385 2015 6415 2035
rect 6435 2015 6465 2035
rect 6485 2015 6515 2035
rect 6535 2015 6565 2035
rect 6585 2015 6615 2035
rect 6635 2015 6665 2035
rect 6685 2015 6715 2035
rect 6735 2015 6765 2035
rect 6785 2015 6815 2035
rect 6835 2015 6865 2035
rect 6885 2015 6915 2035
rect 6935 2015 6965 2035
rect 6985 2015 7015 2035
rect 7035 2015 7065 2035
rect 7085 2015 7115 2035
rect 7135 2015 7165 2035
rect 7185 2015 7215 2035
rect 7235 2015 7265 2035
rect 7285 2015 7315 2035
rect 7335 2015 7365 2035
rect 7385 2015 7415 2035
rect 7435 2015 7465 2035
rect 7485 2015 7515 2035
rect 7535 2015 7565 2035
rect 7585 2015 7615 2035
rect 7635 2015 7665 2035
rect 7685 2015 7715 2035
rect 7735 2015 7765 2035
rect 7785 2015 7815 2035
rect 7835 2015 7865 2035
rect 7885 2015 7915 2035
rect 7935 2015 7965 2035
rect 7985 2015 8015 2035
rect 8035 2015 8065 2035
rect 8085 2015 8115 2035
rect 8135 2015 8165 2035
rect 8185 2015 8215 2035
rect 8235 2015 8265 2035
rect 8285 2015 8315 2035
rect 8335 2015 8365 2035
rect 8385 2015 8415 2035
rect 8435 2015 8465 2035
rect 8485 2015 8515 2035
rect 8535 2015 8565 2035
rect 8585 2015 8615 2035
rect 8635 2015 8665 2035
rect 8685 2015 8715 2035
rect 8735 2015 8765 2035
rect 8785 2015 8815 2035
rect 8835 2015 8865 2035
rect 8885 2015 8915 2035
rect 8935 2015 8965 2035
rect 8985 2015 9015 2035
rect 9035 2015 9065 2035
rect 9085 2015 9115 2035
rect 9135 2015 9165 2035
rect 9185 2015 9215 2035
rect 9235 2015 9265 2035
rect 9285 2015 9315 2035
rect 9335 2015 9365 2035
rect 9385 2015 9415 2035
rect 9435 2015 9465 2035
rect 9485 2015 9515 2035
rect 9535 2015 9565 2035
rect 9585 2015 9615 2035
rect 9635 2015 9665 2035
rect 9685 2015 9715 2035
rect 9735 2015 9765 2035
rect 9785 2015 9815 2035
rect 9835 2015 9865 2035
rect 9885 2015 9915 2035
rect 9935 2015 9965 2035
rect 9985 2015 10015 2035
rect 10035 2015 10065 2035
rect 10085 2015 10115 2035
rect 10135 2015 10165 2035
rect 10185 2015 10215 2035
rect 10235 2015 10265 2035
rect 10285 2015 10315 2035
rect 10335 2015 10365 2035
rect 10385 2015 10415 2035
rect 10435 2015 10465 2035
rect 10485 2015 10515 2035
rect 10535 2015 10565 2035
rect 10585 2015 10615 2035
rect 10635 2015 10665 2035
rect 10685 2015 10715 2035
rect 10735 2015 10765 2035
rect 10785 2015 10815 2035
rect 10835 2015 10865 2035
rect 10885 2015 10915 2035
rect 10935 2015 10965 2035
rect 10985 2015 11015 2035
rect 11035 2015 11065 2035
rect 11085 2015 11115 2035
rect 11135 2015 11165 2035
rect 11185 2015 11215 2035
rect 11235 2015 11265 2035
rect 11285 2015 11315 2035
rect 11335 2015 11365 2035
rect 11385 2015 11415 2035
rect 11435 2015 11465 2035
rect 11485 2015 11515 2035
rect 11535 2015 11565 2035
rect 11585 2015 11615 2035
rect 11635 2015 11665 2035
rect 11685 2015 11715 2035
rect 11735 2015 11765 2035
rect 11785 2015 11815 2035
rect 11835 2015 11865 2035
rect 11885 2015 11915 2035
rect 11935 2015 11965 2035
rect 11985 2015 12015 2035
rect 12035 2015 12065 2035
rect 12085 2015 12115 2035
rect 12135 2015 12165 2035
rect 12185 2015 12215 2035
rect 12235 2015 12265 2035
rect 12285 2015 12315 2035
rect 12335 2015 12365 2035
rect 12385 2015 12415 2035
rect 12435 2015 12465 2035
rect 12485 2015 12515 2035
rect 12535 2015 12565 2035
rect 12585 2015 12615 2035
rect 12635 2015 12665 2035
rect 12685 2015 12715 2035
rect 12735 2015 12765 2035
rect 12785 2015 12815 2035
rect 12835 2015 12865 2035
rect 12885 2015 12915 2035
rect 12935 2015 12965 2035
rect 12985 2015 13015 2035
rect 13035 2015 13065 2035
rect 13085 2015 13115 2035
rect 13135 2015 13165 2035
rect 13185 2015 13215 2035
rect 13235 2015 13265 2035
rect 13285 2015 13315 2035
rect 13335 2015 13365 2035
rect 13385 2015 13415 2035
rect 13435 2015 13465 2035
rect 13485 2015 13515 2035
rect 13535 2015 13565 2035
rect 13585 2015 13615 2035
rect 13635 2015 13665 2035
rect 13685 2015 13715 2035
rect 13735 2015 13765 2035
rect 13785 2015 13815 2035
rect 13835 2015 13865 2035
rect 13885 2015 13915 2035
rect 13935 2015 13965 2035
rect 13985 2015 14015 2035
rect 14035 2015 14065 2035
rect 14085 2015 14115 2035
rect 14135 2015 14165 2035
rect 14185 2015 14215 2035
rect 14235 2015 14265 2035
rect 14285 2015 14315 2035
rect 14335 2015 14365 2035
rect 14385 2015 14415 2035
rect 14435 2015 14465 2035
rect 14485 2015 14515 2035
rect 14535 2015 14565 2035
rect 14585 2015 14615 2035
rect 14635 2015 14665 2035
rect 14685 2015 14715 2035
rect 14735 2015 14765 2035
rect 14785 2015 14815 2035
rect 14835 2015 14865 2035
rect 14885 2015 14915 2035
rect 14935 2015 14965 2035
rect 14985 2015 15015 2035
rect 15035 2015 15065 2035
rect 15085 2015 15115 2035
rect 15135 2015 15165 2035
rect 15185 2015 15215 2035
rect 15235 2015 15265 2035
rect 15285 2015 15315 2035
rect 15335 2015 15365 2035
rect 15385 2015 15415 2035
rect 15435 2015 15465 2035
rect 15485 2015 15515 2035
rect 15535 2015 15565 2035
rect 15585 2015 15615 2035
rect 15635 2015 15665 2035
rect 15685 2015 15715 2035
rect 15735 2015 15765 2035
rect 15785 2015 15815 2035
rect 15835 2015 15865 2035
rect 15885 2015 15915 2035
rect 15935 2015 15965 2035
rect 15985 2015 16015 2035
rect 16035 2015 16065 2035
rect 16085 2015 16115 2035
rect 16135 2015 16165 2035
rect 16185 2015 16215 2035
rect 16235 2015 16265 2035
rect 16285 2015 16315 2035
rect 16335 2015 16365 2035
rect 16385 2015 16415 2035
rect 16435 2015 16465 2035
rect 16485 2015 16515 2035
rect 16535 2015 16565 2035
rect 16585 2015 16615 2035
rect 16635 2015 16665 2035
rect 16685 2015 16715 2035
rect 16735 2015 16765 2035
rect 16785 2015 16815 2035
rect 16835 2015 16865 2035
rect 16885 2015 16915 2035
rect 16935 2015 16965 2035
rect 16985 2015 17015 2035
rect 17035 2015 17065 2035
rect 17085 2015 17115 2035
rect 17135 2015 17165 2035
rect 17185 2015 17215 2035
rect 17235 2015 17265 2035
rect 17285 2015 17315 2035
rect 17335 2015 17365 2035
rect 17385 2015 17415 2035
rect 17435 2015 17465 2035
rect 17485 2015 17515 2035
rect 17535 2015 17565 2035
rect 17585 2015 17615 2035
rect 17635 2015 17665 2035
rect 17685 2015 17715 2035
rect 17735 2015 17765 2035
rect 17785 2015 17815 2035
rect 17835 2015 17865 2035
rect 17885 2015 17915 2035
rect 17935 2015 17965 2035
rect 17985 2015 18015 2035
rect 18035 2015 18065 2035
rect 18085 2015 18115 2035
rect 18135 2015 18165 2035
rect 18185 2015 18215 2035
rect 18235 2015 18265 2035
rect 18285 2015 18315 2035
rect 18335 2015 18365 2035
rect 18385 2015 18415 2035
rect 18435 2015 18465 2035
rect 18485 2015 18515 2035
rect 18535 2015 18565 2035
rect 18585 2015 18615 2035
rect 18635 2015 18665 2035
rect 18685 2015 18715 2035
rect 18735 2015 18765 2035
rect 18785 2015 18815 2035
rect 18835 2015 18865 2035
rect 18885 2015 18915 2035
rect 18935 2015 18965 2035
rect 18985 2015 19015 2035
rect 19035 2015 19065 2035
rect 19085 2015 19115 2035
rect 19135 2015 19165 2035
rect 19185 2015 19215 2035
rect 19235 2015 19265 2035
rect 19285 2015 19315 2035
rect 19335 2015 19365 2035
rect 19385 2015 19415 2035
rect 19435 2015 19465 2035
rect 19485 2015 19515 2035
rect 19535 2015 19565 2035
rect 19585 2015 19615 2035
rect 19635 2015 19665 2035
rect 19685 2015 19715 2035
rect 19735 2015 19765 2035
rect 19785 2015 19815 2035
rect 19835 2015 19865 2035
rect 19885 2015 19915 2035
rect 19935 2015 19965 2035
rect 19985 2015 20015 2035
rect 20035 2015 20065 2035
rect 20085 2015 20115 2035
rect 20135 2015 20165 2035
rect 20185 2015 20215 2035
rect 20235 2015 20265 2035
rect 20285 2015 20315 2035
rect 20335 2015 20365 2035
rect 20385 2015 20400 2035
rect -900 2000 20400 2015
rect -650 1835 20400 1850
rect -650 1815 -635 1835
rect -615 1815 -585 1835
rect -565 1815 -535 1835
rect -515 1815 -485 1835
rect -465 1815 -435 1835
rect -415 1815 -385 1835
rect -365 1815 -335 1835
rect -315 1815 -285 1835
rect -265 1815 -235 1835
rect -215 1815 -185 1835
rect -165 1815 -135 1835
rect -115 1815 -85 1835
rect -65 1815 -35 1835
rect -15 1815 15 1835
rect 35 1815 65 1835
rect 85 1815 115 1835
rect 135 1815 165 1835
rect 185 1815 215 1835
rect 235 1815 265 1835
rect 285 1815 315 1835
rect 335 1815 365 1835
rect 385 1815 415 1835
rect 435 1815 465 1835
rect 485 1815 515 1835
rect 535 1815 565 1835
rect 585 1815 615 1835
rect 635 1815 665 1835
rect 685 1815 715 1835
rect 735 1815 765 1835
rect 785 1815 815 1835
rect 835 1815 865 1835
rect 885 1815 915 1835
rect 935 1815 965 1835
rect 985 1815 1015 1835
rect 1035 1815 1065 1835
rect 1085 1815 1115 1835
rect 1135 1815 1165 1835
rect 1185 1815 1215 1835
rect 1235 1815 1265 1835
rect 1285 1815 1315 1835
rect 1335 1815 1365 1835
rect 1385 1815 1415 1835
rect 1435 1815 1465 1835
rect 1485 1815 1515 1835
rect 1535 1815 1565 1835
rect 1585 1815 1615 1835
rect 1635 1815 1665 1835
rect 1685 1815 1715 1835
rect 1735 1815 1765 1835
rect 1785 1815 1815 1835
rect 1835 1815 1865 1835
rect 1885 1815 1915 1835
rect 1935 1815 1965 1835
rect 1985 1815 2015 1835
rect 2035 1815 2065 1835
rect 2085 1815 2115 1835
rect 2135 1815 2165 1835
rect 2185 1815 2215 1835
rect 2235 1815 2265 1835
rect 2285 1815 2315 1835
rect 2335 1815 2365 1835
rect 2385 1815 2415 1835
rect 2435 1815 2465 1835
rect 2485 1815 2515 1835
rect 2535 1815 2565 1835
rect 2585 1815 2615 1835
rect 2635 1815 2665 1835
rect 2685 1815 2715 1835
rect 2735 1815 2765 1835
rect 2785 1815 2815 1835
rect 2835 1815 2865 1835
rect 2885 1815 2915 1835
rect 2935 1815 2965 1835
rect 2985 1815 3015 1835
rect 3035 1815 3065 1835
rect 3085 1815 3115 1835
rect 3135 1815 3165 1835
rect 3185 1815 3215 1835
rect 3235 1815 3265 1835
rect 3285 1815 3315 1835
rect 3335 1815 3365 1835
rect 3385 1815 3415 1835
rect 3435 1815 3465 1835
rect 3485 1815 3515 1835
rect 3535 1815 3565 1835
rect 3585 1815 3615 1835
rect 3635 1815 3665 1835
rect 3685 1815 3715 1835
rect 3735 1815 3765 1835
rect 3785 1815 3815 1835
rect 3835 1815 3865 1835
rect 3885 1815 3915 1835
rect 3935 1815 3965 1835
rect 3985 1815 4015 1835
rect 4035 1815 4065 1835
rect 4085 1815 4115 1835
rect 4135 1815 4165 1835
rect 4185 1815 4215 1835
rect 4235 1815 4265 1835
rect 4285 1815 4315 1835
rect 4335 1815 4365 1835
rect 4385 1815 4415 1835
rect 4435 1815 4465 1835
rect 4485 1815 4515 1835
rect 4535 1815 4565 1835
rect 4585 1815 4615 1835
rect 4635 1815 4665 1835
rect 4685 1815 4715 1835
rect 4735 1815 4765 1835
rect 4785 1815 4815 1835
rect 4835 1815 4865 1835
rect 4885 1815 4915 1835
rect 4935 1815 4965 1835
rect 4985 1815 5015 1835
rect 5035 1815 5065 1835
rect 5085 1815 5115 1835
rect 5135 1815 5165 1835
rect 5185 1815 5215 1835
rect 5235 1815 5265 1835
rect 5285 1815 5315 1835
rect 5335 1815 5365 1835
rect 5385 1815 5415 1835
rect 5435 1815 5465 1835
rect 5485 1815 5515 1835
rect 5535 1815 5565 1835
rect 5585 1815 5615 1835
rect 5635 1815 5665 1835
rect 5685 1815 5715 1835
rect 5735 1815 5765 1835
rect 5785 1815 5815 1835
rect 5835 1815 5865 1835
rect 5885 1815 5915 1835
rect 5935 1815 5965 1835
rect 5985 1815 6015 1835
rect 6035 1815 6065 1835
rect 6085 1815 6115 1835
rect 6135 1815 6165 1835
rect 6185 1815 6215 1835
rect 6235 1815 6265 1835
rect 6285 1815 6315 1835
rect 6335 1815 6365 1835
rect 6385 1815 6415 1835
rect 6435 1815 6465 1835
rect 6485 1815 6515 1835
rect 6535 1815 6565 1835
rect 6585 1815 6615 1835
rect 6635 1815 6665 1835
rect 6685 1815 6715 1835
rect 6735 1815 6765 1835
rect 6785 1815 6815 1835
rect 6835 1815 6865 1835
rect 6885 1815 6915 1835
rect 6935 1815 6965 1835
rect 6985 1815 7015 1835
rect 7035 1815 7065 1835
rect 7085 1815 7115 1835
rect 7135 1815 7165 1835
rect 7185 1815 7215 1835
rect 7235 1815 7265 1835
rect 7285 1815 7315 1835
rect 7335 1815 7365 1835
rect 7385 1815 7415 1835
rect 7435 1815 7465 1835
rect 7485 1815 7515 1835
rect 7535 1815 7565 1835
rect 7585 1815 7615 1835
rect 7635 1815 7665 1835
rect 7685 1815 7715 1835
rect 7735 1815 7765 1835
rect 7785 1815 7815 1835
rect 7835 1815 7865 1835
rect 7885 1815 7915 1835
rect 7935 1815 7965 1835
rect 7985 1815 8015 1835
rect 8035 1815 8065 1835
rect 8085 1815 8115 1835
rect 8135 1815 8165 1835
rect 8185 1815 8215 1835
rect 8235 1815 8265 1835
rect 8285 1815 8315 1835
rect 8335 1815 8365 1835
rect 8385 1815 8415 1835
rect 8435 1815 8465 1835
rect 8485 1815 8515 1835
rect 8535 1815 8565 1835
rect 8585 1815 8615 1835
rect 8635 1815 8665 1835
rect 8685 1815 8715 1835
rect 8735 1815 8765 1835
rect 8785 1815 8815 1835
rect 8835 1815 8865 1835
rect 8885 1815 8915 1835
rect 8935 1815 8965 1835
rect 8985 1815 9015 1835
rect 9035 1815 9065 1835
rect 9085 1815 9115 1835
rect 9135 1815 9165 1835
rect 9185 1815 9215 1835
rect 9235 1815 9265 1835
rect 9285 1815 9315 1835
rect 9335 1815 9365 1835
rect 9385 1815 9415 1835
rect 9435 1815 9465 1835
rect 9485 1815 9515 1835
rect 9535 1815 9565 1835
rect 9585 1815 9615 1835
rect 9635 1815 9665 1835
rect 9685 1815 9715 1835
rect 9735 1815 9765 1835
rect 9785 1815 9815 1835
rect 9835 1815 9865 1835
rect 9885 1815 9915 1835
rect 9935 1815 9965 1835
rect 9985 1815 10015 1835
rect 10035 1815 10065 1835
rect 10085 1815 10115 1835
rect 10135 1815 10165 1835
rect 10185 1815 10215 1835
rect 10235 1815 10265 1835
rect 10285 1815 10315 1835
rect 10335 1815 10365 1835
rect 10385 1815 10415 1835
rect 10435 1815 10465 1835
rect 10485 1815 10515 1835
rect 10535 1815 10565 1835
rect 10585 1815 10615 1835
rect 10635 1815 10665 1835
rect 10685 1815 10715 1835
rect 10735 1815 10765 1835
rect 10785 1815 10815 1835
rect 10835 1815 10865 1835
rect 10885 1815 10915 1835
rect 10935 1815 10965 1835
rect 10985 1815 11015 1835
rect 11035 1815 11065 1835
rect 11085 1815 11115 1835
rect 11135 1815 11165 1835
rect 11185 1815 11215 1835
rect 11235 1815 11265 1835
rect 11285 1815 11315 1835
rect 11335 1815 11365 1835
rect 11385 1815 11415 1835
rect 11435 1815 11465 1835
rect 11485 1815 11515 1835
rect 11535 1815 11565 1835
rect 11585 1815 11615 1835
rect 11635 1815 11665 1835
rect 11685 1815 11715 1835
rect 11735 1815 11765 1835
rect 11785 1815 11815 1835
rect 11835 1815 11865 1835
rect 11885 1815 11915 1835
rect 11935 1815 11965 1835
rect 11985 1815 12015 1835
rect 12035 1815 12065 1835
rect 12085 1815 12115 1835
rect 12135 1815 12165 1835
rect 12185 1815 12215 1835
rect 12235 1815 12265 1835
rect 12285 1815 12315 1835
rect 12335 1815 12365 1835
rect 12385 1815 12415 1835
rect 12435 1815 12465 1835
rect 12485 1815 12515 1835
rect 12535 1815 12565 1835
rect 12585 1815 12615 1835
rect 12635 1815 12665 1835
rect 12685 1815 12715 1835
rect 12735 1815 12765 1835
rect 12785 1815 12815 1835
rect 12835 1815 12865 1835
rect 12885 1815 12915 1835
rect 12935 1815 12965 1835
rect 12985 1815 13015 1835
rect 13035 1815 13065 1835
rect 13085 1815 13115 1835
rect 13135 1815 13165 1835
rect 13185 1815 13215 1835
rect 13235 1815 13265 1835
rect 13285 1815 13315 1835
rect 13335 1815 13365 1835
rect 13385 1815 13415 1835
rect 13435 1815 13465 1835
rect 13485 1815 13515 1835
rect 13535 1815 13565 1835
rect 13585 1815 13615 1835
rect 13635 1815 13665 1835
rect 13685 1815 13715 1835
rect 13735 1815 13765 1835
rect 13785 1815 13815 1835
rect 13835 1815 13865 1835
rect 13885 1815 13915 1835
rect 13935 1815 13965 1835
rect 13985 1815 14015 1835
rect 14035 1815 14065 1835
rect 14085 1815 14115 1835
rect 14135 1815 14165 1835
rect 14185 1815 14215 1835
rect 14235 1815 14265 1835
rect 14285 1815 14315 1835
rect 14335 1815 14365 1835
rect 14385 1815 14415 1835
rect 14435 1815 14465 1835
rect 14485 1815 14515 1835
rect 14535 1815 14565 1835
rect 14585 1815 14615 1835
rect 14635 1815 14665 1835
rect 14685 1815 14715 1835
rect 14735 1815 14765 1835
rect 14785 1815 14815 1835
rect 14835 1815 14865 1835
rect 14885 1815 14915 1835
rect 14935 1815 14965 1835
rect 14985 1815 15015 1835
rect 15035 1815 15065 1835
rect 15085 1815 15115 1835
rect 15135 1815 15165 1835
rect 15185 1815 15215 1835
rect 15235 1815 15265 1835
rect 15285 1815 15315 1835
rect 15335 1815 15365 1835
rect 15385 1815 15415 1835
rect 15435 1815 15465 1835
rect 15485 1815 15515 1835
rect 15535 1815 15565 1835
rect 15585 1815 15615 1835
rect 15635 1815 15665 1835
rect 15685 1815 15715 1835
rect 15735 1815 15765 1835
rect 15785 1815 15815 1835
rect 15835 1815 15865 1835
rect 15885 1815 15915 1835
rect 15935 1815 15965 1835
rect 15985 1815 16015 1835
rect 16035 1815 16065 1835
rect 16085 1815 16115 1835
rect 16135 1815 16165 1835
rect 16185 1815 16215 1835
rect 16235 1815 16265 1835
rect 16285 1815 16315 1835
rect 16335 1815 16365 1835
rect 16385 1815 16415 1835
rect 16435 1815 16465 1835
rect 16485 1815 16515 1835
rect 16535 1815 16565 1835
rect 16585 1815 16615 1835
rect 16635 1815 16665 1835
rect 16685 1815 16715 1835
rect 16735 1815 16765 1835
rect 16785 1815 16815 1835
rect 16835 1815 16865 1835
rect 16885 1815 16915 1835
rect 16935 1815 16965 1835
rect 16985 1815 17015 1835
rect 17035 1815 17065 1835
rect 17085 1815 17115 1835
rect 17135 1815 17165 1835
rect 17185 1815 17215 1835
rect 17235 1815 17265 1835
rect 17285 1815 17315 1835
rect 17335 1815 17365 1835
rect 17385 1815 17415 1835
rect 17435 1815 17465 1835
rect 17485 1815 17515 1835
rect 17535 1815 17565 1835
rect 17585 1815 17615 1835
rect 17635 1815 17665 1835
rect 17685 1815 17715 1835
rect 17735 1815 17765 1835
rect 17785 1815 17815 1835
rect 17835 1815 17865 1835
rect 17885 1815 17915 1835
rect 17935 1815 17965 1835
rect 17985 1815 18015 1835
rect 18035 1815 18065 1835
rect 18085 1815 18115 1835
rect 18135 1815 18165 1835
rect 18185 1815 18215 1835
rect 18235 1815 18265 1835
rect 18285 1815 18315 1835
rect 18335 1815 18365 1835
rect 18385 1815 18415 1835
rect 18435 1815 18465 1835
rect 18485 1815 18515 1835
rect 18535 1815 18565 1835
rect 18585 1815 18615 1835
rect 18635 1815 18665 1835
rect 18685 1815 18715 1835
rect 18735 1815 18765 1835
rect 18785 1815 18815 1835
rect 18835 1815 18865 1835
rect 18885 1815 18915 1835
rect 18935 1815 18965 1835
rect 18985 1815 19015 1835
rect 19035 1815 19065 1835
rect 19085 1815 19115 1835
rect 19135 1815 19165 1835
rect 19185 1815 19215 1835
rect 19235 1815 19265 1835
rect 19285 1815 19315 1835
rect 19335 1815 19365 1835
rect 19385 1815 19415 1835
rect 19435 1815 19465 1835
rect 19485 1815 19515 1835
rect 19535 1815 19565 1835
rect 19585 1815 19615 1835
rect 19635 1815 19665 1835
rect 19685 1815 19715 1835
rect 19735 1815 19765 1835
rect 19785 1815 19815 1835
rect 19835 1815 19865 1835
rect 19885 1815 19915 1835
rect 19935 1815 19965 1835
rect 19985 1815 20015 1835
rect 20035 1815 20065 1835
rect 20085 1815 20115 1835
rect 20135 1815 20165 1835
rect 20185 1815 20215 1835
rect 20235 1815 20265 1835
rect 20285 1815 20315 1835
rect 20335 1815 20365 1835
rect 20385 1815 20400 1835
rect -650 1800 20400 1815
rect -650 1685 20400 1700
rect -650 1665 -635 1685
rect -615 1665 -585 1685
rect -565 1665 -535 1685
rect -515 1665 -485 1685
rect -465 1665 -435 1685
rect -415 1665 -385 1685
rect -365 1665 -335 1685
rect -315 1665 -285 1685
rect -265 1665 -235 1685
rect -215 1665 -185 1685
rect -165 1665 -135 1685
rect -115 1665 -85 1685
rect -65 1665 -35 1685
rect -15 1665 15 1685
rect 35 1665 65 1685
rect 85 1665 115 1685
rect 135 1665 165 1685
rect 185 1665 215 1685
rect 235 1665 265 1685
rect 285 1665 315 1685
rect 335 1665 365 1685
rect 385 1665 415 1685
rect 435 1665 465 1685
rect 485 1665 515 1685
rect 535 1665 565 1685
rect 585 1665 615 1685
rect 635 1665 665 1685
rect 685 1665 715 1685
rect 735 1665 765 1685
rect 785 1665 815 1685
rect 835 1665 865 1685
rect 885 1665 915 1685
rect 935 1665 965 1685
rect 985 1665 1015 1685
rect 1035 1665 1065 1685
rect 1085 1665 1115 1685
rect 1135 1665 1165 1685
rect 1185 1665 1215 1685
rect 1235 1665 1265 1685
rect 1285 1665 1315 1685
rect 1335 1665 1365 1685
rect 1385 1665 1415 1685
rect 1435 1665 1465 1685
rect 1485 1665 1515 1685
rect 1535 1665 1565 1685
rect 1585 1665 1615 1685
rect 1635 1665 1665 1685
rect 1685 1665 1715 1685
rect 1735 1665 1765 1685
rect 1785 1665 1815 1685
rect 1835 1665 1865 1685
rect 1885 1665 1915 1685
rect 1935 1665 1965 1685
rect 1985 1665 2015 1685
rect 2035 1665 2065 1685
rect 2085 1665 2115 1685
rect 2135 1665 2165 1685
rect 2185 1665 2215 1685
rect 2235 1665 2265 1685
rect 2285 1665 2315 1685
rect 2335 1665 2365 1685
rect 2385 1665 2415 1685
rect 2435 1665 2465 1685
rect 2485 1665 2515 1685
rect 2535 1665 2565 1685
rect 2585 1665 2615 1685
rect 2635 1665 2665 1685
rect 2685 1665 2715 1685
rect 2735 1665 2765 1685
rect 2785 1665 2815 1685
rect 2835 1665 2865 1685
rect 2885 1665 2915 1685
rect 2935 1665 2965 1685
rect 2985 1665 3015 1685
rect 3035 1665 3065 1685
rect 3085 1665 3115 1685
rect 3135 1665 3165 1685
rect 3185 1665 3215 1685
rect 3235 1665 3265 1685
rect 3285 1665 3315 1685
rect 3335 1665 3365 1685
rect 3385 1665 3415 1685
rect 3435 1665 3465 1685
rect 3485 1665 3515 1685
rect 3535 1665 3565 1685
rect 3585 1665 3615 1685
rect 3635 1665 3665 1685
rect 3685 1665 3715 1685
rect 3735 1665 3765 1685
rect 3785 1665 3815 1685
rect 3835 1665 3865 1685
rect 3885 1665 3915 1685
rect 3935 1665 3965 1685
rect 3985 1665 4015 1685
rect 4035 1665 4065 1685
rect 4085 1665 4115 1685
rect 4135 1665 4165 1685
rect 4185 1665 4215 1685
rect 4235 1665 4265 1685
rect 4285 1665 4315 1685
rect 4335 1665 4365 1685
rect 4385 1665 4415 1685
rect 4435 1665 4465 1685
rect 4485 1665 4515 1685
rect 4535 1665 4565 1685
rect 4585 1665 4615 1685
rect 4635 1665 4665 1685
rect 4685 1665 4715 1685
rect 4735 1665 4765 1685
rect 4785 1665 4815 1685
rect 4835 1665 4865 1685
rect 4885 1665 4915 1685
rect 4935 1665 4965 1685
rect 4985 1665 5015 1685
rect 5035 1665 5065 1685
rect 5085 1665 5115 1685
rect 5135 1665 5165 1685
rect 5185 1665 5215 1685
rect 5235 1665 5265 1685
rect 5285 1665 5315 1685
rect 5335 1665 5365 1685
rect 5385 1665 5415 1685
rect 5435 1665 5465 1685
rect 5485 1665 5515 1685
rect 5535 1665 5565 1685
rect 5585 1665 5615 1685
rect 5635 1665 5665 1685
rect 5685 1665 5715 1685
rect 5735 1665 5765 1685
rect 5785 1665 5815 1685
rect 5835 1665 5865 1685
rect 5885 1665 5915 1685
rect 5935 1665 5965 1685
rect 5985 1665 6015 1685
rect 6035 1665 6065 1685
rect 6085 1665 6115 1685
rect 6135 1665 6165 1685
rect 6185 1665 6215 1685
rect 6235 1665 6265 1685
rect 6285 1665 6315 1685
rect 6335 1665 6365 1685
rect 6385 1665 6415 1685
rect 6435 1665 6465 1685
rect 6485 1665 6515 1685
rect 6535 1665 6565 1685
rect 6585 1665 6615 1685
rect 6635 1665 6665 1685
rect 6685 1665 6715 1685
rect 6735 1665 6765 1685
rect 6785 1665 6815 1685
rect 6835 1665 6865 1685
rect 6885 1665 6915 1685
rect 6935 1665 6965 1685
rect 6985 1665 7015 1685
rect 7035 1665 7065 1685
rect 7085 1665 7115 1685
rect 7135 1665 7165 1685
rect 7185 1665 7215 1685
rect 7235 1665 7265 1685
rect 7285 1665 7315 1685
rect 7335 1665 7365 1685
rect 7385 1665 7415 1685
rect 7435 1665 7465 1685
rect 7485 1665 7515 1685
rect 7535 1665 7565 1685
rect 7585 1665 7615 1685
rect 7635 1665 7665 1685
rect 7685 1665 7715 1685
rect 7735 1665 7765 1685
rect 7785 1665 7815 1685
rect 7835 1665 7865 1685
rect 7885 1665 7915 1685
rect 7935 1665 7965 1685
rect 7985 1665 8015 1685
rect 8035 1665 8065 1685
rect 8085 1665 8115 1685
rect 8135 1665 8165 1685
rect 8185 1665 8215 1685
rect 8235 1665 8265 1685
rect 8285 1665 8315 1685
rect 8335 1665 8365 1685
rect 8385 1665 8415 1685
rect 8435 1665 8465 1685
rect 8485 1665 8515 1685
rect 8535 1665 8565 1685
rect 8585 1665 8615 1685
rect 8635 1665 8665 1685
rect 8685 1665 8715 1685
rect 8735 1665 8765 1685
rect 8785 1665 8815 1685
rect 8835 1665 8865 1685
rect 8885 1665 8915 1685
rect 8935 1665 8965 1685
rect 8985 1665 9015 1685
rect 9035 1665 9065 1685
rect 9085 1665 9115 1685
rect 9135 1665 9165 1685
rect 9185 1665 9215 1685
rect 9235 1665 9265 1685
rect 9285 1665 9315 1685
rect 9335 1665 9365 1685
rect 9385 1665 9415 1685
rect 9435 1665 9465 1685
rect 9485 1665 9515 1685
rect 9535 1665 9565 1685
rect 9585 1665 9615 1685
rect 9635 1665 9665 1685
rect 9685 1665 9715 1685
rect 9735 1665 9765 1685
rect 9785 1665 9815 1685
rect 9835 1665 9865 1685
rect 9885 1665 9915 1685
rect 9935 1665 9965 1685
rect 9985 1665 10015 1685
rect 10035 1665 10065 1685
rect 10085 1665 10115 1685
rect 10135 1665 10165 1685
rect 10185 1665 10215 1685
rect 10235 1665 10265 1685
rect 10285 1665 10315 1685
rect 10335 1665 10365 1685
rect 10385 1665 10415 1685
rect 10435 1665 10465 1685
rect 10485 1665 10515 1685
rect 10535 1665 10565 1685
rect 10585 1665 10615 1685
rect 10635 1665 10665 1685
rect 10685 1665 10715 1685
rect 10735 1665 10765 1685
rect 10785 1665 10815 1685
rect 10835 1665 10865 1685
rect 10885 1665 10915 1685
rect 10935 1665 10965 1685
rect 10985 1665 11015 1685
rect 11035 1665 11065 1685
rect 11085 1665 11115 1685
rect 11135 1665 11165 1685
rect 11185 1665 11215 1685
rect 11235 1665 11265 1685
rect 11285 1665 11315 1685
rect 11335 1665 11365 1685
rect 11385 1665 11415 1685
rect 11435 1665 11465 1685
rect 11485 1665 11515 1685
rect 11535 1665 11565 1685
rect 11585 1665 11615 1685
rect 11635 1665 11665 1685
rect 11685 1665 11715 1685
rect 11735 1665 11765 1685
rect 11785 1665 11815 1685
rect 11835 1665 11865 1685
rect 11885 1665 11915 1685
rect 11935 1665 11965 1685
rect 11985 1665 12015 1685
rect 12035 1665 12065 1685
rect 12085 1665 12115 1685
rect 12135 1665 12165 1685
rect 12185 1665 12215 1685
rect 12235 1665 12265 1685
rect 12285 1665 12315 1685
rect 12335 1665 12365 1685
rect 12385 1665 12415 1685
rect 12435 1665 12465 1685
rect 12485 1665 12515 1685
rect 12535 1665 12565 1685
rect 12585 1665 12615 1685
rect 12635 1665 12665 1685
rect 12685 1665 12715 1685
rect 12735 1665 12765 1685
rect 12785 1665 12815 1685
rect 12835 1665 12865 1685
rect 12885 1665 12915 1685
rect 12935 1665 12965 1685
rect 12985 1665 13015 1685
rect 13035 1665 13065 1685
rect 13085 1665 13115 1685
rect 13135 1665 13165 1685
rect 13185 1665 13215 1685
rect 13235 1665 13265 1685
rect 13285 1665 13315 1685
rect 13335 1665 13365 1685
rect 13385 1665 13415 1685
rect 13435 1665 13465 1685
rect 13485 1665 13515 1685
rect 13535 1665 13565 1685
rect 13585 1665 13615 1685
rect 13635 1665 13665 1685
rect 13685 1665 13715 1685
rect 13735 1665 13765 1685
rect 13785 1665 13815 1685
rect 13835 1665 13865 1685
rect 13885 1665 13915 1685
rect 13935 1665 13965 1685
rect 13985 1665 14015 1685
rect 14035 1665 14065 1685
rect 14085 1665 14115 1685
rect 14135 1665 14165 1685
rect 14185 1665 14215 1685
rect 14235 1665 14265 1685
rect 14285 1665 14315 1685
rect 14335 1665 14365 1685
rect 14385 1665 14415 1685
rect 14435 1665 14465 1685
rect 14485 1665 14515 1685
rect 14535 1665 14565 1685
rect 14585 1665 14615 1685
rect 14635 1665 14665 1685
rect 14685 1665 14715 1685
rect 14735 1665 14765 1685
rect 14785 1665 14815 1685
rect 14835 1665 14865 1685
rect 14885 1665 14915 1685
rect 14935 1665 14965 1685
rect 14985 1665 15015 1685
rect 15035 1665 15065 1685
rect 15085 1665 15115 1685
rect 15135 1665 15165 1685
rect 15185 1665 15215 1685
rect 15235 1665 15265 1685
rect 15285 1665 15315 1685
rect 15335 1665 15365 1685
rect 15385 1665 15415 1685
rect 15435 1665 15465 1685
rect 15485 1665 15515 1685
rect 15535 1665 15565 1685
rect 15585 1665 15615 1685
rect 15635 1665 15665 1685
rect 15685 1665 15715 1685
rect 15735 1665 15765 1685
rect 15785 1665 15815 1685
rect 15835 1665 15865 1685
rect 15885 1665 15915 1685
rect 15935 1665 15965 1685
rect 15985 1665 16015 1685
rect 16035 1665 16065 1685
rect 16085 1665 16115 1685
rect 16135 1665 16165 1685
rect 16185 1665 16215 1685
rect 16235 1665 16265 1685
rect 16285 1665 16315 1685
rect 16335 1665 16365 1685
rect 16385 1665 16415 1685
rect 16435 1665 16465 1685
rect 16485 1665 16515 1685
rect 16535 1665 16565 1685
rect 16585 1665 16615 1685
rect 16635 1665 16665 1685
rect 16685 1665 16715 1685
rect 16735 1665 16765 1685
rect 16785 1665 16815 1685
rect 16835 1665 16865 1685
rect 16885 1665 16915 1685
rect 16935 1665 16965 1685
rect 16985 1665 17015 1685
rect 17035 1665 17065 1685
rect 17085 1665 17115 1685
rect 17135 1665 17165 1685
rect 17185 1665 17215 1685
rect 17235 1665 17265 1685
rect 17285 1665 17315 1685
rect 17335 1665 17365 1685
rect 17385 1665 17415 1685
rect 17435 1665 17465 1685
rect 17485 1665 17515 1685
rect 17535 1665 17565 1685
rect 17585 1665 17615 1685
rect 17635 1665 17665 1685
rect 17685 1665 17715 1685
rect 17735 1665 17765 1685
rect 17785 1665 17815 1685
rect 17835 1665 17865 1685
rect 17885 1665 17915 1685
rect 17935 1665 17965 1685
rect 17985 1665 18015 1685
rect 18035 1665 18065 1685
rect 18085 1665 18115 1685
rect 18135 1665 18165 1685
rect 18185 1665 18215 1685
rect 18235 1665 18265 1685
rect 18285 1665 18315 1685
rect 18335 1665 18365 1685
rect 18385 1665 18415 1685
rect 18435 1665 18465 1685
rect 18485 1665 18515 1685
rect 18535 1665 18565 1685
rect 18585 1665 18615 1685
rect 18635 1665 18665 1685
rect 18685 1665 18715 1685
rect 18735 1665 18765 1685
rect 18785 1665 18815 1685
rect 18835 1665 18865 1685
rect 18885 1665 18915 1685
rect 18935 1665 18965 1685
rect 18985 1665 19015 1685
rect 19035 1665 19065 1685
rect 19085 1665 19115 1685
rect 19135 1665 19165 1685
rect 19185 1665 19215 1685
rect 19235 1665 19265 1685
rect 19285 1665 19315 1685
rect 19335 1665 19365 1685
rect 19385 1665 19415 1685
rect 19435 1665 19465 1685
rect 19485 1665 19515 1685
rect 19535 1665 19565 1685
rect 19585 1665 19615 1685
rect 19635 1665 19665 1685
rect 19685 1665 19715 1685
rect 19735 1665 19765 1685
rect 19785 1665 19815 1685
rect 19835 1665 19865 1685
rect 19885 1665 19915 1685
rect 19935 1665 19965 1685
rect 19985 1665 20015 1685
rect 20035 1665 20065 1685
rect 20085 1665 20115 1685
rect 20135 1665 20165 1685
rect 20185 1665 20215 1685
rect 20235 1665 20265 1685
rect 20285 1665 20315 1685
rect 20335 1665 20365 1685
rect 20385 1665 20400 1685
rect -650 1650 20400 1665
rect -650 1585 -600 1600
rect -650 1565 -635 1585
rect -615 1565 -600 1585
rect -650 1535 -600 1565
rect -650 1515 -635 1535
rect -615 1515 -600 1535
rect -650 1485 -600 1515
rect -650 1465 -635 1485
rect -615 1465 -600 1485
rect -650 1435 -600 1465
rect -650 1415 -635 1435
rect -615 1415 -600 1435
rect -650 1385 -600 1415
rect -650 1365 -635 1385
rect -615 1365 -600 1385
rect -650 1335 -600 1365
rect -650 1315 -635 1335
rect -615 1315 -600 1335
rect -650 1285 -600 1315
rect -650 1265 -635 1285
rect -615 1265 -600 1285
rect -650 1235 -600 1265
rect -650 1215 -635 1235
rect -615 1215 -600 1235
rect -650 1185 -600 1215
rect -650 1165 -635 1185
rect -615 1165 -600 1185
rect -650 1135 -600 1165
rect -650 1115 -635 1135
rect -615 1115 -600 1135
rect -650 1085 -600 1115
rect -650 1065 -635 1085
rect -615 1065 -600 1085
rect -650 1035 -600 1065
rect -650 1015 -635 1035
rect -615 1015 -600 1035
rect -650 985 -600 1015
rect -650 965 -635 985
rect -615 965 -600 985
rect -650 935 -600 965
rect -650 915 -635 935
rect -615 915 -600 935
rect -650 900 -600 915
rect -500 1585 -450 1600
rect -500 1565 -485 1585
rect -465 1565 -450 1585
rect -500 1535 -450 1565
rect -500 1515 -485 1535
rect -465 1515 -450 1535
rect -500 1485 -450 1515
rect -500 1465 -485 1485
rect -465 1465 -450 1485
rect -500 1435 -450 1465
rect -500 1415 -485 1435
rect -465 1415 -450 1435
rect -500 1385 -450 1415
rect -500 1365 -485 1385
rect -465 1365 -450 1385
rect -500 1335 -450 1365
rect -500 1315 -485 1335
rect -465 1315 -450 1335
rect -500 1285 -450 1315
rect -500 1265 -485 1285
rect -465 1265 -450 1285
rect -500 1235 -450 1265
rect -500 1215 -485 1235
rect -465 1215 -450 1235
rect -500 1185 -450 1215
rect -500 1165 -485 1185
rect -465 1165 -450 1185
rect -500 1135 -450 1165
rect -500 1115 -485 1135
rect -465 1115 -450 1135
rect -500 1085 -450 1115
rect -500 1065 -485 1085
rect -465 1065 -450 1085
rect -500 1035 -450 1065
rect -500 1015 -485 1035
rect -465 1015 -450 1035
rect -500 985 -450 1015
rect -500 965 -485 985
rect -465 965 -450 985
rect -500 935 -450 965
rect -500 915 -485 935
rect -465 915 -450 935
rect -500 900 -450 915
rect -350 1585 -300 1600
rect -350 1565 -335 1585
rect -315 1565 -300 1585
rect -350 1535 -300 1565
rect -350 1515 -335 1535
rect -315 1515 -300 1535
rect -350 1485 -300 1515
rect -350 1465 -335 1485
rect -315 1465 -300 1485
rect -350 1435 -300 1465
rect -350 1415 -335 1435
rect -315 1415 -300 1435
rect -350 1385 -300 1415
rect -350 1365 -335 1385
rect -315 1365 -300 1385
rect -350 1335 -300 1365
rect -350 1315 -335 1335
rect -315 1315 -300 1335
rect -350 1285 -300 1315
rect -350 1265 -335 1285
rect -315 1265 -300 1285
rect -350 1235 -300 1265
rect -350 1215 -335 1235
rect -315 1215 -300 1235
rect -350 1185 -300 1215
rect -350 1165 -335 1185
rect -315 1165 -300 1185
rect -350 1135 -300 1165
rect -350 1115 -335 1135
rect -315 1115 -300 1135
rect -350 1085 -300 1115
rect -350 1065 -335 1085
rect -315 1065 -300 1085
rect -350 1035 -300 1065
rect -350 1015 -335 1035
rect -315 1015 -300 1035
rect -350 985 -300 1015
rect -350 965 -335 985
rect -315 965 -300 985
rect -350 935 -300 965
rect -350 915 -335 935
rect -315 915 -300 935
rect -350 900 -300 915
rect -200 1585 -150 1600
rect -200 1565 -185 1585
rect -165 1565 -150 1585
rect -200 1535 -150 1565
rect -200 1515 -185 1535
rect -165 1515 -150 1535
rect -200 1485 -150 1515
rect -200 1465 -185 1485
rect -165 1465 -150 1485
rect -200 1435 -150 1465
rect -200 1415 -185 1435
rect -165 1415 -150 1435
rect -200 1385 -150 1415
rect -200 1365 -185 1385
rect -165 1365 -150 1385
rect -200 1335 -150 1365
rect -200 1315 -185 1335
rect -165 1315 -150 1335
rect -200 1285 -150 1315
rect -200 1265 -185 1285
rect -165 1265 -150 1285
rect -200 1235 -150 1265
rect -200 1215 -185 1235
rect -165 1215 -150 1235
rect -200 1185 -150 1215
rect -200 1165 -185 1185
rect -165 1165 -150 1185
rect -200 1135 -150 1165
rect -200 1115 -185 1135
rect -165 1115 -150 1135
rect -200 1085 -150 1115
rect -200 1065 -185 1085
rect -165 1065 -150 1085
rect -200 1035 -150 1065
rect -200 1015 -185 1035
rect -165 1015 -150 1035
rect -200 985 -150 1015
rect -200 965 -185 985
rect -165 965 -150 985
rect -200 935 -150 965
rect -200 915 -185 935
rect -165 915 -150 935
rect -200 900 -150 915
rect -50 1585 0 1600
rect -50 1565 -35 1585
rect -15 1565 0 1585
rect -50 1535 0 1565
rect -50 1515 -35 1535
rect -15 1515 0 1535
rect -50 1485 0 1515
rect -50 1465 -35 1485
rect -15 1465 0 1485
rect -50 1435 0 1465
rect -50 1415 -35 1435
rect -15 1415 0 1435
rect -50 1385 0 1415
rect -50 1365 -35 1385
rect -15 1365 0 1385
rect -50 1335 0 1365
rect -50 1315 -35 1335
rect -15 1315 0 1335
rect -50 1285 0 1315
rect -50 1265 -35 1285
rect -15 1265 0 1285
rect -50 1235 0 1265
rect -50 1215 -35 1235
rect -15 1215 0 1235
rect -50 1185 0 1215
rect -50 1165 -35 1185
rect -15 1165 0 1185
rect -50 1135 0 1165
rect -50 1115 -35 1135
rect -15 1115 0 1135
rect -50 1085 0 1115
rect -50 1065 -35 1085
rect -15 1065 0 1085
rect -50 1035 0 1065
rect -50 1015 -35 1035
rect -15 1015 0 1035
rect -50 985 0 1015
rect -50 965 -35 985
rect -15 965 0 985
rect -50 935 0 965
rect -50 915 -35 935
rect -15 915 0 935
rect -50 900 0 915
rect 1150 1585 1200 1600
rect 1150 1565 1165 1585
rect 1185 1565 1200 1585
rect 1150 1535 1200 1565
rect 1150 1515 1165 1535
rect 1185 1515 1200 1535
rect 1150 1485 1200 1515
rect 1150 1465 1165 1485
rect 1185 1465 1200 1485
rect 1150 1435 1200 1465
rect 1150 1415 1165 1435
rect 1185 1415 1200 1435
rect 1150 1385 1200 1415
rect 1150 1365 1165 1385
rect 1185 1365 1200 1385
rect 1150 1335 1200 1365
rect 1150 1315 1165 1335
rect 1185 1315 1200 1335
rect 1150 1285 1200 1315
rect 1150 1265 1165 1285
rect 1185 1265 1200 1285
rect 1150 1235 1200 1265
rect 1150 1215 1165 1235
rect 1185 1215 1200 1235
rect 1150 1185 1200 1215
rect 1150 1165 1165 1185
rect 1185 1165 1200 1185
rect 1150 1135 1200 1165
rect 1150 1115 1165 1135
rect 1185 1115 1200 1135
rect 1150 1085 1200 1115
rect 1150 1065 1165 1085
rect 1185 1065 1200 1085
rect 1150 1035 1200 1065
rect 1150 1015 1165 1035
rect 1185 1015 1200 1035
rect 1150 985 1200 1015
rect 1150 965 1165 985
rect 1185 965 1200 985
rect 1150 935 1200 965
rect 1150 915 1165 935
rect 1185 915 1200 935
rect 1150 900 1200 915
rect 1450 1585 1500 1600
rect 1450 1565 1465 1585
rect 1485 1565 1500 1585
rect 1450 1535 1500 1565
rect 1450 1515 1465 1535
rect 1485 1515 1500 1535
rect 1450 1485 1500 1515
rect 1450 1465 1465 1485
rect 1485 1465 1500 1485
rect 1450 1435 1500 1465
rect 1450 1415 1465 1435
rect 1485 1415 1500 1435
rect 1450 1385 1500 1415
rect 1450 1365 1465 1385
rect 1485 1365 1500 1385
rect 1450 1335 1500 1365
rect 1450 1315 1465 1335
rect 1485 1315 1500 1335
rect 1450 1285 1500 1315
rect 1450 1265 1465 1285
rect 1485 1265 1500 1285
rect 1450 1235 1500 1265
rect 1450 1215 1465 1235
rect 1485 1215 1500 1235
rect 1450 1185 1500 1215
rect 1450 1165 1465 1185
rect 1485 1165 1500 1185
rect 1450 1135 1500 1165
rect 1450 1115 1465 1135
rect 1485 1115 1500 1135
rect 1450 1085 1500 1115
rect 1450 1065 1465 1085
rect 1485 1065 1500 1085
rect 1450 1035 1500 1065
rect 1450 1015 1465 1035
rect 1485 1015 1500 1035
rect 1450 985 1500 1015
rect 1450 965 1465 985
rect 1485 965 1500 985
rect 1450 935 1500 965
rect 1450 915 1465 935
rect 1485 915 1500 935
rect 1450 900 1500 915
rect 1750 1585 1800 1600
rect 1750 1565 1765 1585
rect 1785 1565 1800 1585
rect 1750 1535 1800 1565
rect 1750 1515 1765 1535
rect 1785 1515 1800 1535
rect 1750 1485 1800 1515
rect 1750 1465 1765 1485
rect 1785 1465 1800 1485
rect 1750 1435 1800 1465
rect 1750 1415 1765 1435
rect 1785 1415 1800 1435
rect 1750 1385 1800 1415
rect 1750 1365 1765 1385
rect 1785 1365 1800 1385
rect 1750 1335 1800 1365
rect 1750 1315 1765 1335
rect 1785 1315 1800 1335
rect 1750 1285 1800 1315
rect 1750 1265 1765 1285
rect 1785 1265 1800 1285
rect 1750 1235 1800 1265
rect 1750 1215 1765 1235
rect 1785 1215 1800 1235
rect 1750 1185 1800 1215
rect 1750 1165 1765 1185
rect 1785 1165 1800 1185
rect 1750 1135 1800 1165
rect 1750 1115 1765 1135
rect 1785 1115 1800 1135
rect 1750 1085 1800 1115
rect 1750 1065 1765 1085
rect 1785 1065 1800 1085
rect 1750 1035 1800 1065
rect 1750 1015 1765 1035
rect 1785 1015 1800 1035
rect 1750 985 1800 1015
rect 1750 965 1765 985
rect 1785 965 1800 985
rect 1750 935 1800 965
rect 1750 915 1765 935
rect 1785 915 1800 935
rect 1750 900 1800 915
rect 2050 1585 2100 1600
rect 2050 1565 2065 1585
rect 2085 1565 2100 1585
rect 2050 1535 2100 1565
rect 2050 1515 2065 1535
rect 2085 1515 2100 1535
rect 2050 1485 2100 1515
rect 2050 1465 2065 1485
rect 2085 1465 2100 1485
rect 2050 1435 2100 1465
rect 2050 1415 2065 1435
rect 2085 1415 2100 1435
rect 2050 1385 2100 1415
rect 2050 1365 2065 1385
rect 2085 1365 2100 1385
rect 2050 1335 2100 1365
rect 2050 1315 2065 1335
rect 2085 1315 2100 1335
rect 2050 1285 2100 1315
rect 2050 1265 2065 1285
rect 2085 1265 2100 1285
rect 2050 1235 2100 1265
rect 2050 1215 2065 1235
rect 2085 1215 2100 1235
rect 2050 1185 2100 1215
rect 2050 1165 2065 1185
rect 2085 1165 2100 1185
rect 2050 1135 2100 1165
rect 2050 1115 2065 1135
rect 2085 1115 2100 1135
rect 2050 1085 2100 1115
rect 2050 1065 2065 1085
rect 2085 1065 2100 1085
rect 2050 1035 2100 1065
rect 2050 1015 2065 1035
rect 2085 1015 2100 1035
rect 2050 985 2100 1015
rect 2050 965 2065 985
rect 2085 965 2100 985
rect 2050 935 2100 965
rect 2050 915 2065 935
rect 2085 915 2100 935
rect 2050 900 2100 915
rect 2350 1585 2400 1600
rect 2350 1565 2365 1585
rect 2385 1565 2400 1585
rect 2350 1535 2400 1565
rect 2350 1515 2365 1535
rect 2385 1515 2400 1535
rect 2350 1485 2400 1515
rect 2350 1465 2365 1485
rect 2385 1465 2400 1485
rect 2350 1435 2400 1465
rect 2350 1415 2365 1435
rect 2385 1415 2400 1435
rect 2350 1385 2400 1415
rect 2350 1365 2365 1385
rect 2385 1365 2400 1385
rect 2350 1335 2400 1365
rect 2350 1315 2365 1335
rect 2385 1315 2400 1335
rect 2350 1285 2400 1315
rect 2350 1265 2365 1285
rect 2385 1265 2400 1285
rect 2350 1235 2400 1265
rect 2350 1215 2365 1235
rect 2385 1215 2400 1235
rect 2350 1185 2400 1215
rect 2350 1165 2365 1185
rect 2385 1165 2400 1185
rect 2350 1135 2400 1165
rect 2350 1115 2365 1135
rect 2385 1115 2400 1135
rect 2350 1085 2400 1115
rect 2350 1065 2365 1085
rect 2385 1065 2400 1085
rect 2350 1035 2400 1065
rect 2350 1015 2365 1035
rect 2385 1015 2400 1035
rect 2350 985 2400 1015
rect 2350 965 2365 985
rect 2385 965 2400 985
rect 2350 935 2400 965
rect 2350 915 2365 935
rect 2385 915 2400 935
rect 2350 900 2400 915
rect 2650 1585 2700 1600
rect 2650 1565 2665 1585
rect 2685 1565 2700 1585
rect 2650 1535 2700 1565
rect 2650 1515 2665 1535
rect 2685 1515 2700 1535
rect 2650 1485 2700 1515
rect 2650 1465 2665 1485
rect 2685 1465 2700 1485
rect 2650 1435 2700 1465
rect 2650 1415 2665 1435
rect 2685 1415 2700 1435
rect 2650 1385 2700 1415
rect 2650 1365 2665 1385
rect 2685 1365 2700 1385
rect 2650 1335 2700 1365
rect 2650 1315 2665 1335
rect 2685 1315 2700 1335
rect 2650 1285 2700 1315
rect 2650 1265 2665 1285
rect 2685 1265 2700 1285
rect 2650 1235 2700 1265
rect 2650 1215 2665 1235
rect 2685 1215 2700 1235
rect 2650 1185 2700 1215
rect 2650 1165 2665 1185
rect 2685 1165 2700 1185
rect 2650 1135 2700 1165
rect 2650 1115 2665 1135
rect 2685 1115 2700 1135
rect 2650 1085 2700 1115
rect 2650 1065 2665 1085
rect 2685 1065 2700 1085
rect 2650 1035 2700 1065
rect 2650 1015 2665 1035
rect 2685 1015 2700 1035
rect 2650 985 2700 1015
rect 2650 965 2665 985
rect 2685 965 2700 985
rect 2650 935 2700 965
rect 2650 915 2665 935
rect 2685 915 2700 935
rect 2650 900 2700 915
rect 2950 1585 3000 1600
rect 2950 1565 2965 1585
rect 2985 1565 3000 1585
rect 2950 1535 3000 1565
rect 2950 1515 2965 1535
rect 2985 1515 3000 1535
rect 2950 1485 3000 1515
rect 2950 1465 2965 1485
rect 2985 1465 3000 1485
rect 2950 1435 3000 1465
rect 2950 1415 2965 1435
rect 2985 1415 3000 1435
rect 2950 1385 3000 1415
rect 2950 1365 2965 1385
rect 2985 1365 3000 1385
rect 2950 1335 3000 1365
rect 2950 1315 2965 1335
rect 2985 1315 3000 1335
rect 2950 1285 3000 1315
rect 2950 1265 2965 1285
rect 2985 1265 3000 1285
rect 2950 1235 3000 1265
rect 2950 1215 2965 1235
rect 2985 1215 3000 1235
rect 2950 1185 3000 1215
rect 2950 1165 2965 1185
rect 2985 1165 3000 1185
rect 2950 1135 3000 1165
rect 2950 1115 2965 1135
rect 2985 1115 3000 1135
rect 2950 1085 3000 1115
rect 2950 1065 2965 1085
rect 2985 1065 3000 1085
rect 2950 1035 3000 1065
rect 2950 1015 2965 1035
rect 2985 1015 3000 1035
rect 2950 985 3000 1015
rect 2950 965 2965 985
rect 2985 965 3000 985
rect 2950 935 3000 965
rect 2950 915 2965 935
rect 2985 915 3000 935
rect 2950 900 3000 915
rect 3250 1585 3300 1600
rect 3250 1565 3265 1585
rect 3285 1565 3300 1585
rect 3250 1535 3300 1565
rect 3250 1515 3265 1535
rect 3285 1515 3300 1535
rect 3250 1485 3300 1515
rect 3250 1465 3265 1485
rect 3285 1465 3300 1485
rect 3250 1435 3300 1465
rect 3250 1415 3265 1435
rect 3285 1415 3300 1435
rect 3250 1385 3300 1415
rect 3250 1365 3265 1385
rect 3285 1365 3300 1385
rect 3250 1335 3300 1365
rect 3250 1315 3265 1335
rect 3285 1315 3300 1335
rect 3250 1285 3300 1315
rect 3250 1265 3265 1285
rect 3285 1265 3300 1285
rect 3250 1235 3300 1265
rect 3250 1215 3265 1235
rect 3285 1215 3300 1235
rect 3250 1185 3300 1215
rect 3250 1165 3265 1185
rect 3285 1165 3300 1185
rect 3250 1135 3300 1165
rect 3250 1115 3265 1135
rect 3285 1115 3300 1135
rect 3250 1085 3300 1115
rect 3250 1065 3265 1085
rect 3285 1065 3300 1085
rect 3250 1035 3300 1065
rect 3250 1015 3265 1035
rect 3285 1015 3300 1035
rect 3250 985 3300 1015
rect 3250 965 3265 985
rect 3285 965 3300 985
rect 3250 935 3300 965
rect 3250 915 3265 935
rect 3285 915 3300 935
rect 3250 900 3300 915
rect 3550 1585 3600 1600
rect 3550 1565 3565 1585
rect 3585 1565 3600 1585
rect 3550 1535 3600 1565
rect 3550 1515 3565 1535
rect 3585 1515 3600 1535
rect 3550 1485 3600 1515
rect 3550 1465 3565 1485
rect 3585 1465 3600 1485
rect 3550 1435 3600 1465
rect 3550 1415 3565 1435
rect 3585 1415 3600 1435
rect 3550 1385 3600 1415
rect 3550 1365 3565 1385
rect 3585 1365 3600 1385
rect 3550 1335 3600 1365
rect 3550 1315 3565 1335
rect 3585 1315 3600 1335
rect 3550 1285 3600 1315
rect 3550 1265 3565 1285
rect 3585 1265 3600 1285
rect 3550 1235 3600 1265
rect 3550 1215 3565 1235
rect 3585 1215 3600 1235
rect 3550 1185 3600 1215
rect 3550 1165 3565 1185
rect 3585 1165 3600 1185
rect 3550 1135 3600 1165
rect 3550 1115 3565 1135
rect 3585 1115 3600 1135
rect 3550 1085 3600 1115
rect 3550 1065 3565 1085
rect 3585 1065 3600 1085
rect 3550 1035 3600 1065
rect 3550 1015 3565 1035
rect 3585 1015 3600 1035
rect 3550 985 3600 1015
rect 3550 965 3565 985
rect 3585 965 3600 985
rect 3550 935 3600 965
rect 3550 915 3565 935
rect 3585 915 3600 935
rect 3550 900 3600 915
rect 3700 1585 3750 1600
rect 3700 1565 3715 1585
rect 3735 1565 3750 1585
rect 3700 1535 3750 1565
rect 3700 1515 3715 1535
rect 3735 1515 3750 1535
rect 3700 1485 3750 1515
rect 3700 1465 3715 1485
rect 3735 1465 3750 1485
rect 3700 1435 3750 1465
rect 3700 1415 3715 1435
rect 3735 1415 3750 1435
rect 3700 1385 3750 1415
rect 3700 1365 3715 1385
rect 3735 1365 3750 1385
rect 3700 1335 3750 1365
rect 3700 1315 3715 1335
rect 3735 1315 3750 1335
rect 3700 1285 3750 1315
rect 3700 1265 3715 1285
rect 3735 1265 3750 1285
rect 3700 1235 3750 1265
rect 3700 1215 3715 1235
rect 3735 1215 3750 1235
rect 3700 1185 3750 1215
rect 3700 1165 3715 1185
rect 3735 1165 3750 1185
rect 3700 1135 3750 1165
rect 3700 1115 3715 1135
rect 3735 1115 3750 1135
rect 3700 1085 3750 1115
rect 3700 1065 3715 1085
rect 3735 1065 3750 1085
rect 3700 1035 3750 1065
rect 3700 1015 3715 1035
rect 3735 1015 3750 1035
rect 3700 985 3750 1015
rect 3700 965 3715 985
rect 3735 965 3750 985
rect 3700 935 3750 965
rect 3700 915 3715 935
rect 3735 915 3750 935
rect 3700 900 3750 915
rect 3850 1585 3900 1600
rect 3850 1565 3865 1585
rect 3885 1565 3900 1585
rect 3850 1535 3900 1565
rect 3850 1515 3865 1535
rect 3885 1515 3900 1535
rect 3850 1485 3900 1515
rect 3850 1465 3865 1485
rect 3885 1465 3900 1485
rect 3850 1435 3900 1465
rect 3850 1415 3865 1435
rect 3885 1415 3900 1435
rect 3850 1385 3900 1415
rect 3850 1365 3865 1385
rect 3885 1365 3900 1385
rect 3850 1335 3900 1365
rect 3850 1315 3865 1335
rect 3885 1315 3900 1335
rect 3850 1285 3900 1315
rect 3850 1265 3865 1285
rect 3885 1265 3900 1285
rect 3850 1235 3900 1265
rect 3850 1215 3865 1235
rect 3885 1215 3900 1235
rect 3850 1185 3900 1215
rect 3850 1165 3865 1185
rect 3885 1165 3900 1185
rect 3850 1135 3900 1165
rect 3850 1115 3865 1135
rect 3885 1115 3900 1135
rect 3850 1085 3900 1115
rect 3850 1065 3865 1085
rect 3885 1065 3900 1085
rect 3850 1035 3900 1065
rect 3850 1015 3865 1035
rect 3885 1015 3900 1035
rect 3850 985 3900 1015
rect 3850 965 3865 985
rect 3885 965 3900 985
rect 3850 935 3900 965
rect 3850 915 3865 935
rect 3885 915 3900 935
rect 3850 900 3900 915
rect 4000 1585 4050 1600
rect 4000 1565 4015 1585
rect 4035 1565 4050 1585
rect 4000 1535 4050 1565
rect 4000 1515 4015 1535
rect 4035 1515 4050 1535
rect 4000 1485 4050 1515
rect 4000 1465 4015 1485
rect 4035 1465 4050 1485
rect 4000 1435 4050 1465
rect 4000 1415 4015 1435
rect 4035 1415 4050 1435
rect 4000 1385 4050 1415
rect 4000 1365 4015 1385
rect 4035 1365 4050 1385
rect 4000 1335 4050 1365
rect 4000 1315 4015 1335
rect 4035 1315 4050 1335
rect 4000 1285 4050 1315
rect 4000 1265 4015 1285
rect 4035 1265 4050 1285
rect 4000 1235 4050 1265
rect 4000 1215 4015 1235
rect 4035 1215 4050 1235
rect 4000 1185 4050 1215
rect 4000 1165 4015 1185
rect 4035 1165 4050 1185
rect 4000 1135 4050 1165
rect 4000 1115 4015 1135
rect 4035 1115 4050 1135
rect 4000 1085 4050 1115
rect 4000 1065 4015 1085
rect 4035 1065 4050 1085
rect 4000 1035 4050 1065
rect 4000 1015 4015 1035
rect 4035 1015 4050 1035
rect 4000 985 4050 1015
rect 4000 965 4015 985
rect 4035 965 4050 985
rect 4000 935 4050 965
rect 4000 915 4015 935
rect 4035 915 4050 935
rect 4000 900 4050 915
rect 4150 1585 4200 1600
rect 4150 1565 4165 1585
rect 4185 1565 4200 1585
rect 4150 1535 4200 1565
rect 4150 1515 4165 1535
rect 4185 1515 4200 1535
rect 4150 1485 4200 1515
rect 4150 1465 4165 1485
rect 4185 1465 4200 1485
rect 4150 1435 4200 1465
rect 4150 1415 4165 1435
rect 4185 1415 4200 1435
rect 4150 1385 4200 1415
rect 4150 1365 4165 1385
rect 4185 1365 4200 1385
rect 4150 1335 4200 1365
rect 4150 1315 4165 1335
rect 4185 1315 4200 1335
rect 4150 1285 4200 1315
rect 4150 1265 4165 1285
rect 4185 1265 4200 1285
rect 4150 1235 4200 1265
rect 4150 1215 4165 1235
rect 4185 1215 4200 1235
rect 4150 1185 4200 1215
rect 4150 1165 4165 1185
rect 4185 1165 4200 1185
rect 4150 1135 4200 1165
rect 4150 1115 4165 1135
rect 4185 1115 4200 1135
rect 4150 1085 4200 1115
rect 4150 1065 4165 1085
rect 4185 1065 4200 1085
rect 4150 1035 4200 1065
rect 4150 1015 4165 1035
rect 4185 1015 4200 1035
rect 4150 985 4200 1015
rect 4150 965 4165 985
rect 4185 965 4200 985
rect 4150 935 4200 965
rect 4150 915 4165 935
rect 4185 915 4200 935
rect 4150 900 4200 915
rect 4300 1585 4350 1600
rect 4300 1565 4315 1585
rect 4335 1565 4350 1585
rect 4300 1535 4350 1565
rect 4300 1515 4315 1535
rect 4335 1515 4350 1535
rect 4300 1485 4350 1515
rect 4300 1465 4315 1485
rect 4335 1465 4350 1485
rect 4300 1435 4350 1465
rect 4300 1415 4315 1435
rect 4335 1415 4350 1435
rect 4300 1385 4350 1415
rect 4300 1365 4315 1385
rect 4335 1365 4350 1385
rect 4300 1335 4350 1365
rect 4300 1315 4315 1335
rect 4335 1315 4350 1335
rect 4300 1285 4350 1315
rect 4300 1265 4315 1285
rect 4335 1265 4350 1285
rect 4300 1235 4350 1265
rect 4300 1215 4315 1235
rect 4335 1215 4350 1235
rect 4300 1185 4350 1215
rect 4300 1165 4315 1185
rect 4335 1165 4350 1185
rect 4300 1135 4350 1165
rect 4300 1115 4315 1135
rect 4335 1115 4350 1135
rect 4300 1085 4350 1115
rect 4300 1065 4315 1085
rect 4335 1065 4350 1085
rect 4300 1035 4350 1065
rect 4300 1015 4315 1035
rect 4335 1015 4350 1035
rect 4300 985 4350 1015
rect 4300 965 4315 985
rect 4335 965 4350 985
rect 4300 935 4350 965
rect 4300 915 4315 935
rect 4335 915 4350 935
rect 4300 900 4350 915
rect 4450 1585 4500 1600
rect 4450 1565 4465 1585
rect 4485 1565 4500 1585
rect 4450 1535 4500 1565
rect 4450 1515 4465 1535
rect 4485 1515 4500 1535
rect 4450 1485 4500 1515
rect 4450 1465 4465 1485
rect 4485 1465 4500 1485
rect 4450 1435 4500 1465
rect 4450 1415 4465 1435
rect 4485 1415 4500 1435
rect 4450 1385 4500 1415
rect 4450 1365 4465 1385
rect 4485 1365 4500 1385
rect 4450 1335 4500 1365
rect 4450 1315 4465 1335
rect 4485 1315 4500 1335
rect 4450 1285 4500 1315
rect 4450 1265 4465 1285
rect 4485 1265 4500 1285
rect 4450 1235 4500 1265
rect 4450 1215 4465 1235
rect 4485 1215 4500 1235
rect 4450 1185 4500 1215
rect 4450 1165 4465 1185
rect 4485 1165 4500 1185
rect 4450 1135 4500 1165
rect 4450 1115 4465 1135
rect 4485 1115 4500 1135
rect 4450 1085 4500 1115
rect 4450 1065 4465 1085
rect 4485 1065 4500 1085
rect 4450 1035 4500 1065
rect 4450 1015 4465 1035
rect 4485 1015 4500 1035
rect 4450 985 4500 1015
rect 4450 965 4465 985
rect 4485 965 4500 985
rect 4450 935 4500 965
rect 4450 915 4465 935
rect 4485 915 4500 935
rect 4450 900 4500 915
rect 4600 1585 4650 1600
rect 4600 1565 4615 1585
rect 4635 1565 4650 1585
rect 4600 1535 4650 1565
rect 4600 1515 4615 1535
rect 4635 1515 4650 1535
rect 4600 1485 4650 1515
rect 4600 1465 4615 1485
rect 4635 1465 4650 1485
rect 4600 1435 4650 1465
rect 4600 1415 4615 1435
rect 4635 1415 4650 1435
rect 4600 1385 4650 1415
rect 4600 1365 4615 1385
rect 4635 1365 4650 1385
rect 4600 1335 4650 1365
rect 4600 1315 4615 1335
rect 4635 1315 4650 1335
rect 4600 1285 4650 1315
rect 4600 1265 4615 1285
rect 4635 1265 4650 1285
rect 4600 1235 4650 1265
rect 4600 1215 4615 1235
rect 4635 1215 4650 1235
rect 4600 1185 4650 1215
rect 4600 1165 4615 1185
rect 4635 1165 4650 1185
rect 4600 1135 4650 1165
rect 4600 1115 4615 1135
rect 4635 1115 4650 1135
rect 4600 1085 4650 1115
rect 4600 1065 4615 1085
rect 4635 1065 4650 1085
rect 4600 1035 4650 1065
rect 4600 1015 4615 1035
rect 4635 1015 4650 1035
rect 4600 985 4650 1015
rect 4600 965 4615 985
rect 4635 965 4650 985
rect 4600 935 4650 965
rect 4600 915 4615 935
rect 4635 915 4650 935
rect 4600 900 4650 915
rect 4750 1585 4800 1600
rect 4750 1565 4765 1585
rect 4785 1565 4800 1585
rect 4750 1535 4800 1565
rect 4750 1515 4765 1535
rect 4785 1515 4800 1535
rect 4750 1485 4800 1515
rect 4750 1465 4765 1485
rect 4785 1465 4800 1485
rect 4750 1435 4800 1465
rect 4750 1415 4765 1435
rect 4785 1415 4800 1435
rect 4750 1385 4800 1415
rect 4750 1365 4765 1385
rect 4785 1365 4800 1385
rect 4750 1335 4800 1365
rect 4750 1315 4765 1335
rect 4785 1315 4800 1335
rect 4750 1285 4800 1315
rect 4750 1265 4765 1285
rect 4785 1265 4800 1285
rect 4750 1235 4800 1265
rect 4750 1215 4765 1235
rect 4785 1215 4800 1235
rect 4750 1185 4800 1215
rect 4750 1165 4765 1185
rect 4785 1165 4800 1185
rect 4750 1135 4800 1165
rect 4750 1115 4765 1135
rect 4785 1115 4800 1135
rect 4750 1085 4800 1115
rect 4750 1065 4765 1085
rect 4785 1065 4800 1085
rect 4750 1035 4800 1065
rect 4750 1015 4765 1035
rect 4785 1015 4800 1035
rect 4750 985 4800 1015
rect 4750 965 4765 985
rect 4785 965 4800 985
rect 4750 935 4800 965
rect 4750 915 4765 935
rect 4785 915 4800 935
rect 4750 900 4800 915
rect 5050 1585 5100 1600
rect 5050 1565 5065 1585
rect 5085 1565 5100 1585
rect 5050 1535 5100 1565
rect 5050 1515 5065 1535
rect 5085 1515 5100 1535
rect 5050 1485 5100 1515
rect 5050 1465 5065 1485
rect 5085 1465 5100 1485
rect 5050 1435 5100 1465
rect 5050 1415 5065 1435
rect 5085 1415 5100 1435
rect 5050 1385 5100 1415
rect 5050 1365 5065 1385
rect 5085 1365 5100 1385
rect 5050 1335 5100 1365
rect 5050 1315 5065 1335
rect 5085 1315 5100 1335
rect 5050 1285 5100 1315
rect 5050 1265 5065 1285
rect 5085 1265 5100 1285
rect 5050 1235 5100 1265
rect 5050 1215 5065 1235
rect 5085 1215 5100 1235
rect 5050 1185 5100 1215
rect 5050 1165 5065 1185
rect 5085 1165 5100 1185
rect 5050 1135 5100 1165
rect 5050 1115 5065 1135
rect 5085 1115 5100 1135
rect 5050 1085 5100 1115
rect 5050 1065 5065 1085
rect 5085 1065 5100 1085
rect 5050 1035 5100 1065
rect 5050 1015 5065 1035
rect 5085 1015 5100 1035
rect 5050 985 5100 1015
rect 5050 965 5065 985
rect 5085 965 5100 985
rect 5050 935 5100 965
rect 5050 915 5065 935
rect 5085 915 5100 935
rect 5050 900 5100 915
rect 5350 1585 5400 1600
rect 5350 1565 5365 1585
rect 5385 1565 5400 1585
rect 5350 1535 5400 1565
rect 5350 1515 5365 1535
rect 5385 1515 5400 1535
rect 5350 1485 5400 1515
rect 5350 1465 5365 1485
rect 5385 1465 5400 1485
rect 5350 1435 5400 1465
rect 5350 1415 5365 1435
rect 5385 1415 5400 1435
rect 5350 1385 5400 1415
rect 5350 1365 5365 1385
rect 5385 1365 5400 1385
rect 5350 1335 5400 1365
rect 5350 1315 5365 1335
rect 5385 1315 5400 1335
rect 5350 1285 5400 1315
rect 5350 1265 5365 1285
rect 5385 1265 5400 1285
rect 5350 1235 5400 1265
rect 5350 1215 5365 1235
rect 5385 1215 5400 1235
rect 5350 1185 5400 1215
rect 5350 1165 5365 1185
rect 5385 1165 5400 1185
rect 5350 1135 5400 1165
rect 5350 1115 5365 1135
rect 5385 1115 5400 1135
rect 5350 1085 5400 1115
rect 5350 1065 5365 1085
rect 5385 1065 5400 1085
rect 5350 1035 5400 1065
rect 5350 1015 5365 1035
rect 5385 1015 5400 1035
rect 5350 985 5400 1015
rect 5350 965 5365 985
rect 5385 965 5400 985
rect 5350 935 5400 965
rect 5350 915 5365 935
rect 5385 915 5400 935
rect 5350 900 5400 915
rect 5650 1585 5700 1600
rect 5650 1565 5665 1585
rect 5685 1565 5700 1585
rect 5650 1535 5700 1565
rect 5650 1515 5665 1535
rect 5685 1515 5700 1535
rect 5650 1485 5700 1515
rect 5650 1465 5665 1485
rect 5685 1465 5700 1485
rect 5650 1435 5700 1465
rect 5650 1415 5665 1435
rect 5685 1415 5700 1435
rect 5650 1385 5700 1415
rect 5650 1365 5665 1385
rect 5685 1365 5700 1385
rect 5650 1335 5700 1365
rect 5650 1315 5665 1335
rect 5685 1315 5700 1335
rect 5650 1285 5700 1315
rect 5650 1265 5665 1285
rect 5685 1265 5700 1285
rect 5650 1235 5700 1265
rect 5650 1215 5665 1235
rect 5685 1215 5700 1235
rect 5650 1185 5700 1215
rect 5650 1165 5665 1185
rect 5685 1165 5700 1185
rect 5650 1135 5700 1165
rect 5650 1115 5665 1135
rect 5685 1115 5700 1135
rect 5650 1085 5700 1115
rect 5650 1065 5665 1085
rect 5685 1065 5700 1085
rect 5650 1035 5700 1065
rect 5650 1015 5665 1035
rect 5685 1015 5700 1035
rect 5650 985 5700 1015
rect 5650 965 5665 985
rect 5685 965 5700 985
rect 5650 935 5700 965
rect 5650 915 5665 935
rect 5685 915 5700 935
rect 5650 900 5700 915
rect 5950 1585 6000 1600
rect 5950 1565 5965 1585
rect 5985 1565 6000 1585
rect 5950 1535 6000 1565
rect 5950 1515 5965 1535
rect 5985 1515 6000 1535
rect 5950 1485 6000 1515
rect 5950 1465 5965 1485
rect 5985 1465 6000 1485
rect 5950 1435 6000 1465
rect 5950 1415 5965 1435
rect 5985 1415 6000 1435
rect 5950 1385 6000 1415
rect 5950 1365 5965 1385
rect 5985 1365 6000 1385
rect 5950 1335 6000 1365
rect 5950 1315 5965 1335
rect 5985 1315 6000 1335
rect 5950 1285 6000 1315
rect 5950 1265 5965 1285
rect 5985 1265 6000 1285
rect 5950 1235 6000 1265
rect 5950 1215 5965 1235
rect 5985 1215 6000 1235
rect 5950 1185 6000 1215
rect 5950 1165 5965 1185
rect 5985 1165 6000 1185
rect 5950 1135 6000 1165
rect 5950 1115 5965 1135
rect 5985 1115 6000 1135
rect 5950 1085 6000 1115
rect 5950 1065 5965 1085
rect 5985 1065 6000 1085
rect 5950 1035 6000 1065
rect 5950 1015 5965 1035
rect 5985 1015 6000 1035
rect 5950 985 6000 1015
rect 5950 965 5965 985
rect 5985 965 6000 985
rect 5950 935 6000 965
rect 5950 915 5965 935
rect 5985 915 6000 935
rect 5950 900 6000 915
rect 6250 1585 6300 1600
rect 6250 1565 6265 1585
rect 6285 1565 6300 1585
rect 6250 1535 6300 1565
rect 6250 1515 6265 1535
rect 6285 1515 6300 1535
rect 6250 1485 6300 1515
rect 6250 1465 6265 1485
rect 6285 1465 6300 1485
rect 6250 1435 6300 1465
rect 6250 1415 6265 1435
rect 6285 1415 6300 1435
rect 6250 1385 6300 1415
rect 6250 1365 6265 1385
rect 6285 1365 6300 1385
rect 6250 1335 6300 1365
rect 6250 1315 6265 1335
rect 6285 1315 6300 1335
rect 6250 1285 6300 1315
rect 6250 1265 6265 1285
rect 6285 1265 6300 1285
rect 6250 1235 6300 1265
rect 6250 1215 6265 1235
rect 6285 1215 6300 1235
rect 6250 1185 6300 1215
rect 6250 1165 6265 1185
rect 6285 1165 6300 1185
rect 6250 1135 6300 1165
rect 6250 1115 6265 1135
rect 6285 1115 6300 1135
rect 6250 1085 6300 1115
rect 6250 1065 6265 1085
rect 6285 1065 6300 1085
rect 6250 1035 6300 1065
rect 6250 1015 6265 1035
rect 6285 1015 6300 1035
rect 6250 985 6300 1015
rect 6250 965 6265 985
rect 6285 965 6300 985
rect 6250 935 6300 965
rect 6250 915 6265 935
rect 6285 915 6300 935
rect 6250 900 6300 915
rect 6550 1585 6600 1600
rect 6550 1565 6565 1585
rect 6585 1565 6600 1585
rect 6550 1535 6600 1565
rect 6550 1515 6565 1535
rect 6585 1515 6600 1535
rect 6550 1485 6600 1515
rect 6550 1465 6565 1485
rect 6585 1465 6600 1485
rect 6550 1435 6600 1465
rect 6550 1415 6565 1435
rect 6585 1415 6600 1435
rect 6550 1385 6600 1415
rect 6550 1365 6565 1385
rect 6585 1365 6600 1385
rect 6550 1335 6600 1365
rect 6550 1315 6565 1335
rect 6585 1315 6600 1335
rect 6550 1285 6600 1315
rect 6550 1265 6565 1285
rect 6585 1265 6600 1285
rect 6550 1235 6600 1265
rect 6550 1215 6565 1235
rect 6585 1215 6600 1235
rect 6550 1185 6600 1215
rect 6550 1165 6565 1185
rect 6585 1165 6600 1185
rect 6550 1135 6600 1165
rect 6550 1115 6565 1135
rect 6585 1115 6600 1135
rect 6550 1085 6600 1115
rect 6550 1065 6565 1085
rect 6585 1065 6600 1085
rect 6550 1035 6600 1065
rect 6550 1015 6565 1035
rect 6585 1015 6600 1035
rect 6550 985 6600 1015
rect 6550 965 6565 985
rect 6585 965 6600 985
rect 6550 935 6600 965
rect 6550 915 6565 935
rect 6585 915 6600 935
rect 6550 900 6600 915
rect 6850 1585 6900 1600
rect 6850 1565 6865 1585
rect 6885 1565 6900 1585
rect 6850 1535 6900 1565
rect 6850 1515 6865 1535
rect 6885 1515 6900 1535
rect 6850 1485 6900 1515
rect 6850 1465 6865 1485
rect 6885 1465 6900 1485
rect 6850 1435 6900 1465
rect 6850 1415 6865 1435
rect 6885 1415 6900 1435
rect 6850 1385 6900 1415
rect 6850 1365 6865 1385
rect 6885 1365 6900 1385
rect 6850 1335 6900 1365
rect 6850 1315 6865 1335
rect 6885 1315 6900 1335
rect 6850 1285 6900 1315
rect 6850 1265 6865 1285
rect 6885 1265 6900 1285
rect 6850 1235 6900 1265
rect 6850 1215 6865 1235
rect 6885 1215 6900 1235
rect 6850 1185 6900 1215
rect 6850 1165 6865 1185
rect 6885 1165 6900 1185
rect 6850 1135 6900 1165
rect 6850 1115 6865 1135
rect 6885 1115 6900 1135
rect 6850 1085 6900 1115
rect 6850 1065 6865 1085
rect 6885 1065 6900 1085
rect 6850 1035 6900 1065
rect 6850 1015 6865 1035
rect 6885 1015 6900 1035
rect 6850 985 6900 1015
rect 6850 965 6865 985
rect 6885 965 6900 985
rect 6850 935 6900 965
rect 6850 915 6865 935
rect 6885 915 6900 935
rect 6850 900 6900 915
rect 7150 1585 7200 1600
rect 7150 1565 7165 1585
rect 7185 1565 7200 1585
rect 7150 1535 7200 1565
rect 7150 1515 7165 1535
rect 7185 1515 7200 1535
rect 7150 1485 7200 1515
rect 7150 1465 7165 1485
rect 7185 1465 7200 1485
rect 7150 1435 7200 1465
rect 7150 1415 7165 1435
rect 7185 1415 7200 1435
rect 7150 1385 7200 1415
rect 7150 1365 7165 1385
rect 7185 1365 7200 1385
rect 7150 1335 7200 1365
rect 7150 1315 7165 1335
rect 7185 1315 7200 1335
rect 7150 1285 7200 1315
rect 7150 1265 7165 1285
rect 7185 1265 7200 1285
rect 7150 1235 7200 1265
rect 7150 1215 7165 1235
rect 7185 1215 7200 1235
rect 7150 1185 7200 1215
rect 7150 1165 7165 1185
rect 7185 1165 7200 1185
rect 7150 1135 7200 1165
rect 7150 1115 7165 1135
rect 7185 1115 7200 1135
rect 7150 1085 7200 1115
rect 7150 1065 7165 1085
rect 7185 1065 7200 1085
rect 7150 1035 7200 1065
rect 7150 1015 7165 1035
rect 7185 1015 7200 1035
rect 7150 985 7200 1015
rect 7150 965 7165 985
rect 7185 965 7200 985
rect 7150 935 7200 965
rect 7150 915 7165 935
rect 7185 915 7200 935
rect 7150 900 7200 915
rect 8350 1585 8400 1600
rect 8350 1565 8365 1585
rect 8385 1565 8400 1585
rect 8350 1535 8400 1565
rect 8350 1515 8365 1535
rect 8385 1515 8400 1535
rect 8350 1485 8400 1515
rect 8350 1465 8365 1485
rect 8385 1465 8400 1485
rect 8350 1435 8400 1465
rect 8350 1415 8365 1435
rect 8385 1415 8400 1435
rect 8350 1385 8400 1415
rect 8350 1365 8365 1385
rect 8385 1365 8400 1385
rect 8350 1335 8400 1365
rect 8350 1315 8365 1335
rect 8385 1315 8400 1335
rect 8350 1285 8400 1315
rect 8350 1265 8365 1285
rect 8385 1265 8400 1285
rect 8350 1235 8400 1265
rect 8350 1215 8365 1235
rect 8385 1215 8400 1235
rect 8350 1185 8400 1215
rect 8350 1165 8365 1185
rect 8385 1165 8400 1185
rect 8350 1135 8400 1165
rect 8350 1115 8365 1135
rect 8385 1115 8400 1135
rect 8350 1085 8400 1115
rect 8350 1065 8365 1085
rect 8385 1065 8400 1085
rect 8350 1035 8400 1065
rect 8350 1015 8365 1035
rect 8385 1015 8400 1035
rect 8350 985 8400 1015
rect 8350 965 8365 985
rect 8385 965 8400 985
rect 8350 935 8400 965
rect 8350 915 8365 935
rect 8385 915 8400 935
rect 8350 900 8400 915
rect 9550 1585 9600 1600
rect 9550 1565 9565 1585
rect 9585 1565 9600 1585
rect 9550 1535 9600 1565
rect 9550 1515 9565 1535
rect 9585 1515 9600 1535
rect 9550 1485 9600 1515
rect 9550 1465 9565 1485
rect 9585 1465 9600 1485
rect 9550 1435 9600 1465
rect 9550 1415 9565 1435
rect 9585 1415 9600 1435
rect 9550 1385 9600 1415
rect 9550 1365 9565 1385
rect 9585 1365 9600 1385
rect 9550 1335 9600 1365
rect 9550 1315 9565 1335
rect 9585 1315 9600 1335
rect 9550 1285 9600 1315
rect 9550 1265 9565 1285
rect 9585 1265 9600 1285
rect 9550 1235 9600 1265
rect 9550 1215 9565 1235
rect 9585 1215 9600 1235
rect 9550 1185 9600 1215
rect 9550 1165 9565 1185
rect 9585 1165 9600 1185
rect 9550 1135 9600 1165
rect 9550 1115 9565 1135
rect 9585 1115 9600 1135
rect 9550 1085 9600 1115
rect 9550 1065 9565 1085
rect 9585 1065 9600 1085
rect 9550 1035 9600 1065
rect 9550 1015 9565 1035
rect 9585 1015 9600 1035
rect 9550 985 9600 1015
rect 9550 965 9565 985
rect 9585 965 9600 985
rect 9550 935 9600 965
rect 9550 915 9565 935
rect 9585 915 9600 935
rect 9550 900 9600 915
rect 10750 1585 10800 1600
rect 10750 1565 10765 1585
rect 10785 1565 10800 1585
rect 10750 1535 10800 1565
rect 10750 1515 10765 1535
rect 10785 1515 10800 1535
rect 10750 1485 10800 1515
rect 10750 1465 10765 1485
rect 10785 1465 10800 1485
rect 10750 1435 10800 1465
rect 10750 1415 10765 1435
rect 10785 1415 10800 1435
rect 10750 1385 10800 1415
rect 10750 1365 10765 1385
rect 10785 1365 10800 1385
rect 10750 1335 10800 1365
rect 10750 1315 10765 1335
rect 10785 1315 10800 1335
rect 10750 1285 10800 1315
rect 10750 1265 10765 1285
rect 10785 1265 10800 1285
rect 10750 1235 10800 1265
rect 10750 1215 10765 1235
rect 10785 1215 10800 1235
rect 10750 1185 10800 1215
rect 10750 1165 10765 1185
rect 10785 1165 10800 1185
rect 10750 1135 10800 1165
rect 10750 1115 10765 1135
rect 10785 1115 10800 1135
rect 10750 1085 10800 1115
rect 10750 1065 10765 1085
rect 10785 1065 10800 1085
rect 10750 1035 10800 1065
rect 10750 1015 10765 1035
rect 10785 1015 10800 1035
rect 10750 985 10800 1015
rect 10750 965 10765 985
rect 10785 965 10800 985
rect 10750 935 10800 965
rect 10750 915 10765 935
rect 10785 915 10800 935
rect 10750 900 10800 915
rect 11950 1585 12000 1600
rect 11950 1565 11965 1585
rect 11985 1565 12000 1585
rect 11950 1535 12000 1565
rect 11950 1515 11965 1535
rect 11985 1515 12000 1535
rect 11950 1485 12000 1515
rect 11950 1465 11965 1485
rect 11985 1465 12000 1485
rect 11950 1435 12000 1465
rect 11950 1415 11965 1435
rect 11985 1415 12000 1435
rect 11950 1385 12000 1415
rect 11950 1365 11965 1385
rect 11985 1365 12000 1385
rect 11950 1335 12000 1365
rect 11950 1315 11965 1335
rect 11985 1315 12000 1335
rect 11950 1285 12000 1315
rect 11950 1265 11965 1285
rect 11985 1265 12000 1285
rect 11950 1235 12000 1265
rect 11950 1215 11965 1235
rect 11985 1215 12000 1235
rect 11950 1185 12000 1215
rect 11950 1165 11965 1185
rect 11985 1165 12000 1185
rect 11950 1135 12000 1165
rect 11950 1115 11965 1135
rect 11985 1115 12000 1135
rect 11950 1085 12000 1115
rect 11950 1065 11965 1085
rect 11985 1065 12000 1085
rect 11950 1035 12000 1065
rect 11950 1015 11965 1035
rect 11985 1015 12000 1035
rect 11950 985 12000 1015
rect 11950 965 11965 985
rect 11985 965 12000 985
rect 11950 935 12000 965
rect 11950 915 11965 935
rect 11985 915 12000 935
rect 11950 900 12000 915
rect 12250 1585 12300 1600
rect 12250 1565 12265 1585
rect 12285 1565 12300 1585
rect 12250 1535 12300 1565
rect 12250 1515 12265 1535
rect 12285 1515 12300 1535
rect 12250 1485 12300 1515
rect 12250 1465 12265 1485
rect 12285 1465 12300 1485
rect 12250 1435 12300 1465
rect 12250 1415 12265 1435
rect 12285 1415 12300 1435
rect 12250 1385 12300 1415
rect 12250 1365 12265 1385
rect 12285 1365 12300 1385
rect 12250 1335 12300 1365
rect 12250 1315 12265 1335
rect 12285 1315 12300 1335
rect 12250 1285 12300 1315
rect 12250 1265 12265 1285
rect 12285 1265 12300 1285
rect 12250 1235 12300 1265
rect 12250 1215 12265 1235
rect 12285 1215 12300 1235
rect 12250 1185 12300 1215
rect 12250 1165 12265 1185
rect 12285 1165 12300 1185
rect 12250 1135 12300 1165
rect 12250 1115 12265 1135
rect 12285 1115 12300 1135
rect 12250 1085 12300 1115
rect 12250 1065 12265 1085
rect 12285 1065 12300 1085
rect 12250 1035 12300 1065
rect 12250 1015 12265 1035
rect 12285 1015 12300 1035
rect 12250 985 12300 1015
rect 12250 965 12265 985
rect 12285 965 12300 985
rect 12250 935 12300 965
rect 12250 915 12265 935
rect 12285 915 12300 935
rect 12250 900 12300 915
rect 12550 1585 12600 1600
rect 12550 1565 12565 1585
rect 12585 1565 12600 1585
rect 12550 1535 12600 1565
rect 12550 1515 12565 1535
rect 12585 1515 12600 1535
rect 12550 1485 12600 1515
rect 12550 1465 12565 1485
rect 12585 1465 12600 1485
rect 12550 1435 12600 1465
rect 12550 1415 12565 1435
rect 12585 1415 12600 1435
rect 12550 1385 12600 1415
rect 12550 1365 12565 1385
rect 12585 1365 12600 1385
rect 12550 1335 12600 1365
rect 12550 1315 12565 1335
rect 12585 1315 12600 1335
rect 12550 1285 12600 1315
rect 12550 1265 12565 1285
rect 12585 1265 12600 1285
rect 12550 1235 12600 1265
rect 12550 1215 12565 1235
rect 12585 1215 12600 1235
rect 12550 1185 12600 1215
rect 12550 1165 12565 1185
rect 12585 1165 12600 1185
rect 12550 1135 12600 1165
rect 12550 1115 12565 1135
rect 12585 1115 12600 1135
rect 12550 1085 12600 1115
rect 12550 1065 12565 1085
rect 12585 1065 12600 1085
rect 12550 1035 12600 1065
rect 12550 1015 12565 1035
rect 12585 1015 12600 1035
rect 12550 985 12600 1015
rect 12550 965 12565 985
rect 12585 965 12600 985
rect 12550 935 12600 965
rect 12550 915 12565 935
rect 12585 915 12600 935
rect 12550 900 12600 915
rect 12850 1585 12900 1600
rect 12850 1565 12865 1585
rect 12885 1565 12900 1585
rect 12850 1535 12900 1565
rect 12850 1515 12865 1535
rect 12885 1515 12900 1535
rect 12850 1485 12900 1515
rect 12850 1465 12865 1485
rect 12885 1465 12900 1485
rect 12850 1435 12900 1465
rect 12850 1415 12865 1435
rect 12885 1415 12900 1435
rect 12850 1385 12900 1415
rect 12850 1365 12865 1385
rect 12885 1365 12900 1385
rect 12850 1335 12900 1365
rect 12850 1315 12865 1335
rect 12885 1315 12900 1335
rect 12850 1285 12900 1315
rect 12850 1265 12865 1285
rect 12885 1265 12900 1285
rect 12850 1235 12900 1265
rect 12850 1215 12865 1235
rect 12885 1215 12900 1235
rect 12850 1185 12900 1215
rect 12850 1165 12865 1185
rect 12885 1165 12900 1185
rect 12850 1135 12900 1165
rect 12850 1115 12865 1135
rect 12885 1115 12900 1135
rect 12850 1085 12900 1115
rect 12850 1065 12865 1085
rect 12885 1065 12900 1085
rect 12850 1035 12900 1065
rect 12850 1015 12865 1035
rect 12885 1015 12900 1035
rect 12850 985 12900 1015
rect 12850 965 12865 985
rect 12885 965 12900 985
rect 12850 935 12900 965
rect 12850 915 12865 935
rect 12885 915 12900 935
rect 12850 900 12900 915
rect 13150 1585 13200 1600
rect 13150 1565 13165 1585
rect 13185 1565 13200 1585
rect 13150 1535 13200 1565
rect 13150 1515 13165 1535
rect 13185 1515 13200 1535
rect 13150 1485 13200 1515
rect 13150 1465 13165 1485
rect 13185 1465 13200 1485
rect 13150 1435 13200 1465
rect 13150 1415 13165 1435
rect 13185 1415 13200 1435
rect 13150 1385 13200 1415
rect 13150 1365 13165 1385
rect 13185 1365 13200 1385
rect 13150 1335 13200 1365
rect 13150 1315 13165 1335
rect 13185 1315 13200 1335
rect 13150 1285 13200 1315
rect 13150 1265 13165 1285
rect 13185 1265 13200 1285
rect 13150 1235 13200 1265
rect 13150 1215 13165 1235
rect 13185 1215 13200 1235
rect 13150 1185 13200 1215
rect 13150 1165 13165 1185
rect 13185 1165 13200 1185
rect 13150 1135 13200 1165
rect 13150 1115 13165 1135
rect 13185 1115 13200 1135
rect 13150 1085 13200 1115
rect 13150 1065 13165 1085
rect 13185 1065 13200 1085
rect 13150 1035 13200 1065
rect 13150 1015 13165 1035
rect 13185 1015 13200 1035
rect 13150 985 13200 1015
rect 13150 965 13165 985
rect 13185 965 13200 985
rect 13150 935 13200 965
rect 13150 915 13165 935
rect 13185 915 13200 935
rect 13150 900 13200 915
rect 13450 1585 13500 1600
rect 13450 1565 13465 1585
rect 13485 1565 13500 1585
rect 13450 1535 13500 1565
rect 13450 1515 13465 1535
rect 13485 1515 13500 1535
rect 13450 1485 13500 1515
rect 13450 1465 13465 1485
rect 13485 1465 13500 1485
rect 13450 1435 13500 1465
rect 13450 1415 13465 1435
rect 13485 1415 13500 1435
rect 13450 1385 13500 1415
rect 13450 1365 13465 1385
rect 13485 1365 13500 1385
rect 13450 1335 13500 1365
rect 13450 1315 13465 1335
rect 13485 1315 13500 1335
rect 13450 1285 13500 1315
rect 13450 1265 13465 1285
rect 13485 1265 13500 1285
rect 13450 1235 13500 1265
rect 13450 1215 13465 1235
rect 13485 1215 13500 1235
rect 13450 1185 13500 1215
rect 13450 1165 13465 1185
rect 13485 1165 13500 1185
rect 13450 1135 13500 1165
rect 13450 1115 13465 1135
rect 13485 1115 13500 1135
rect 13450 1085 13500 1115
rect 13450 1065 13465 1085
rect 13485 1065 13500 1085
rect 13450 1035 13500 1065
rect 13450 1015 13465 1035
rect 13485 1015 13500 1035
rect 13450 985 13500 1015
rect 13450 965 13465 985
rect 13485 965 13500 985
rect 13450 935 13500 965
rect 13450 915 13465 935
rect 13485 915 13500 935
rect 13450 900 13500 915
rect 13750 1585 13800 1600
rect 13750 1565 13765 1585
rect 13785 1565 13800 1585
rect 13750 1535 13800 1565
rect 13750 1515 13765 1535
rect 13785 1515 13800 1535
rect 13750 1485 13800 1515
rect 13750 1465 13765 1485
rect 13785 1465 13800 1485
rect 13750 1435 13800 1465
rect 13750 1415 13765 1435
rect 13785 1415 13800 1435
rect 13750 1385 13800 1415
rect 13750 1365 13765 1385
rect 13785 1365 13800 1385
rect 13750 1335 13800 1365
rect 13750 1315 13765 1335
rect 13785 1315 13800 1335
rect 13750 1285 13800 1315
rect 13750 1265 13765 1285
rect 13785 1265 13800 1285
rect 13750 1235 13800 1265
rect 13750 1215 13765 1235
rect 13785 1215 13800 1235
rect 13750 1185 13800 1215
rect 13750 1165 13765 1185
rect 13785 1165 13800 1185
rect 13750 1135 13800 1165
rect 13750 1115 13765 1135
rect 13785 1115 13800 1135
rect 13750 1085 13800 1115
rect 13750 1065 13765 1085
rect 13785 1065 13800 1085
rect 13750 1035 13800 1065
rect 13750 1015 13765 1035
rect 13785 1015 13800 1035
rect 13750 985 13800 1015
rect 13750 965 13765 985
rect 13785 965 13800 985
rect 13750 935 13800 965
rect 13750 915 13765 935
rect 13785 915 13800 935
rect 13750 900 13800 915
rect 14050 1585 14100 1600
rect 14050 1565 14065 1585
rect 14085 1565 14100 1585
rect 14050 1535 14100 1565
rect 14050 1515 14065 1535
rect 14085 1515 14100 1535
rect 14050 1485 14100 1515
rect 14050 1465 14065 1485
rect 14085 1465 14100 1485
rect 14050 1435 14100 1465
rect 14050 1415 14065 1435
rect 14085 1415 14100 1435
rect 14050 1385 14100 1415
rect 14050 1365 14065 1385
rect 14085 1365 14100 1385
rect 14050 1335 14100 1365
rect 14050 1315 14065 1335
rect 14085 1315 14100 1335
rect 14050 1285 14100 1315
rect 14050 1265 14065 1285
rect 14085 1265 14100 1285
rect 14050 1235 14100 1265
rect 14050 1215 14065 1235
rect 14085 1215 14100 1235
rect 14050 1185 14100 1215
rect 14050 1165 14065 1185
rect 14085 1165 14100 1185
rect 14050 1135 14100 1165
rect 14050 1115 14065 1135
rect 14085 1115 14100 1135
rect 14050 1085 14100 1115
rect 14050 1065 14065 1085
rect 14085 1065 14100 1085
rect 14050 1035 14100 1065
rect 14050 1015 14065 1035
rect 14085 1015 14100 1035
rect 14050 985 14100 1015
rect 14050 965 14065 985
rect 14085 965 14100 985
rect 14050 935 14100 965
rect 14050 915 14065 935
rect 14085 915 14100 935
rect 14050 900 14100 915
rect 14350 1585 14400 1600
rect 14350 1565 14365 1585
rect 14385 1565 14400 1585
rect 14350 1535 14400 1565
rect 14350 1515 14365 1535
rect 14385 1515 14400 1535
rect 14350 1485 14400 1515
rect 14350 1465 14365 1485
rect 14385 1465 14400 1485
rect 14350 1435 14400 1465
rect 14350 1415 14365 1435
rect 14385 1415 14400 1435
rect 14350 1385 14400 1415
rect 14350 1365 14365 1385
rect 14385 1365 14400 1385
rect 14350 1335 14400 1365
rect 14350 1315 14365 1335
rect 14385 1315 14400 1335
rect 14350 1285 14400 1315
rect 14350 1265 14365 1285
rect 14385 1265 14400 1285
rect 14350 1235 14400 1265
rect 14350 1215 14365 1235
rect 14385 1215 14400 1235
rect 14350 1185 14400 1215
rect 14350 1165 14365 1185
rect 14385 1165 14400 1185
rect 14350 1135 14400 1165
rect 14350 1115 14365 1135
rect 14385 1115 14400 1135
rect 14350 1085 14400 1115
rect 14350 1065 14365 1085
rect 14385 1065 14400 1085
rect 14350 1035 14400 1065
rect 14350 1015 14365 1035
rect 14385 1015 14400 1035
rect 14350 985 14400 1015
rect 14350 965 14365 985
rect 14385 965 14400 985
rect 14350 935 14400 965
rect 14350 915 14365 935
rect 14385 915 14400 935
rect 14350 900 14400 915
rect 15550 1585 15600 1600
rect 15550 1565 15565 1585
rect 15585 1565 15600 1585
rect 15550 1535 15600 1565
rect 15550 1515 15565 1535
rect 15585 1515 15600 1535
rect 15550 1485 15600 1515
rect 15550 1465 15565 1485
rect 15585 1465 15600 1485
rect 15550 1435 15600 1465
rect 15550 1415 15565 1435
rect 15585 1415 15600 1435
rect 15550 1385 15600 1415
rect 15550 1365 15565 1385
rect 15585 1365 15600 1385
rect 15550 1335 15600 1365
rect 15550 1315 15565 1335
rect 15585 1315 15600 1335
rect 15550 1285 15600 1315
rect 15550 1265 15565 1285
rect 15585 1265 15600 1285
rect 15550 1235 15600 1265
rect 15550 1215 15565 1235
rect 15585 1215 15600 1235
rect 15550 1185 15600 1215
rect 15550 1165 15565 1185
rect 15585 1165 15600 1185
rect 15550 1135 15600 1165
rect 15550 1115 15565 1135
rect 15585 1115 15600 1135
rect 15550 1085 15600 1115
rect 15550 1065 15565 1085
rect 15585 1065 15600 1085
rect 15550 1035 15600 1065
rect 15550 1015 15565 1035
rect 15585 1015 15600 1035
rect 15550 985 15600 1015
rect 15550 965 15565 985
rect 15585 965 15600 985
rect 15550 935 15600 965
rect 15550 915 15565 935
rect 15585 915 15600 935
rect 15550 900 15600 915
rect 16750 1585 16800 1600
rect 16750 1565 16765 1585
rect 16785 1565 16800 1585
rect 16750 1535 16800 1565
rect 16750 1515 16765 1535
rect 16785 1515 16800 1535
rect 16750 1485 16800 1515
rect 16750 1465 16765 1485
rect 16785 1465 16800 1485
rect 16750 1435 16800 1465
rect 16750 1415 16765 1435
rect 16785 1415 16800 1435
rect 16750 1385 16800 1415
rect 16750 1365 16765 1385
rect 16785 1365 16800 1385
rect 16750 1335 16800 1365
rect 16750 1315 16765 1335
rect 16785 1315 16800 1335
rect 16750 1285 16800 1315
rect 16750 1265 16765 1285
rect 16785 1265 16800 1285
rect 16750 1235 16800 1265
rect 16750 1215 16765 1235
rect 16785 1215 16800 1235
rect 16750 1185 16800 1215
rect 16750 1165 16765 1185
rect 16785 1165 16800 1185
rect 16750 1135 16800 1165
rect 16750 1115 16765 1135
rect 16785 1115 16800 1135
rect 16750 1085 16800 1115
rect 16750 1065 16765 1085
rect 16785 1065 16800 1085
rect 16750 1035 16800 1065
rect 16750 1015 16765 1035
rect 16785 1015 16800 1035
rect 16750 985 16800 1015
rect 16750 965 16765 985
rect 16785 965 16800 985
rect 16750 935 16800 965
rect 16750 915 16765 935
rect 16785 915 16800 935
rect 16750 900 16800 915
rect 17950 1585 18000 1600
rect 17950 1565 17965 1585
rect 17985 1565 18000 1585
rect 17950 1535 18000 1565
rect 17950 1515 17965 1535
rect 17985 1515 18000 1535
rect 17950 1485 18000 1515
rect 17950 1465 17965 1485
rect 17985 1465 18000 1485
rect 17950 1435 18000 1465
rect 17950 1415 17965 1435
rect 17985 1415 18000 1435
rect 17950 1385 18000 1415
rect 17950 1365 17965 1385
rect 17985 1365 18000 1385
rect 17950 1335 18000 1365
rect 17950 1315 17965 1335
rect 17985 1315 18000 1335
rect 17950 1285 18000 1315
rect 17950 1265 17965 1285
rect 17985 1265 18000 1285
rect 17950 1235 18000 1265
rect 17950 1215 17965 1235
rect 17985 1215 18000 1235
rect 17950 1185 18000 1215
rect 17950 1165 17965 1185
rect 17985 1165 18000 1185
rect 17950 1135 18000 1165
rect 17950 1115 17965 1135
rect 17985 1115 18000 1135
rect 17950 1085 18000 1115
rect 17950 1065 17965 1085
rect 17985 1065 18000 1085
rect 17950 1035 18000 1065
rect 17950 1015 17965 1035
rect 17985 1015 18000 1035
rect 17950 985 18000 1015
rect 17950 965 17965 985
rect 17985 965 18000 985
rect 17950 935 18000 965
rect 17950 915 17965 935
rect 17985 915 18000 935
rect 17950 900 18000 915
rect 19150 1585 19200 1600
rect 19150 1565 19165 1585
rect 19185 1565 19200 1585
rect 19150 1535 19200 1565
rect 19150 1515 19165 1535
rect 19185 1515 19200 1535
rect 19150 1485 19200 1515
rect 19150 1465 19165 1485
rect 19185 1465 19200 1485
rect 19150 1435 19200 1465
rect 19150 1415 19165 1435
rect 19185 1415 19200 1435
rect 19150 1385 19200 1415
rect 19150 1365 19165 1385
rect 19185 1365 19200 1385
rect 19150 1335 19200 1365
rect 19150 1315 19165 1335
rect 19185 1315 19200 1335
rect 19150 1285 19200 1315
rect 19150 1265 19165 1285
rect 19185 1265 19200 1285
rect 19150 1235 19200 1265
rect 19150 1215 19165 1235
rect 19185 1215 19200 1235
rect 19150 1185 19200 1215
rect 19150 1165 19165 1185
rect 19185 1165 19200 1185
rect 19150 1135 19200 1165
rect 19150 1115 19165 1135
rect 19185 1115 19200 1135
rect 19150 1085 19200 1115
rect 19150 1065 19165 1085
rect 19185 1065 19200 1085
rect 19150 1035 19200 1065
rect 19150 1015 19165 1035
rect 19185 1015 19200 1035
rect 19150 985 19200 1015
rect 19150 965 19165 985
rect 19185 965 19200 985
rect 19150 935 19200 965
rect 19150 915 19165 935
rect 19185 915 19200 935
rect 19150 900 19200 915
rect 20350 1585 20400 1600
rect 20350 1565 20365 1585
rect 20385 1565 20400 1585
rect 20350 1535 20400 1565
rect 20350 1515 20365 1535
rect 20385 1515 20400 1535
rect 20350 1485 20400 1515
rect 20350 1465 20365 1485
rect 20385 1465 20400 1485
rect 20350 1435 20400 1465
rect 20350 1415 20365 1435
rect 20385 1415 20400 1435
rect 20350 1385 20400 1415
rect 20350 1365 20365 1385
rect 20385 1365 20400 1385
rect 20350 1335 20400 1365
rect 20350 1315 20365 1335
rect 20385 1315 20400 1335
rect 20350 1285 20400 1315
rect 20350 1265 20365 1285
rect 20385 1265 20400 1285
rect 20350 1235 20400 1265
rect 20350 1215 20365 1235
rect 20385 1215 20400 1235
rect 20350 1185 20400 1215
rect 20350 1165 20365 1185
rect 20385 1165 20400 1185
rect 20350 1135 20400 1165
rect 20350 1115 20365 1135
rect 20385 1115 20400 1135
rect 20350 1085 20400 1115
rect 20350 1065 20365 1085
rect 20385 1065 20400 1085
rect 20350 1035 20400 1065
rect 20350 1015 20365 1035
rect 20385 1015 20400 1035
rect 20350 985 20400 1015
rect 20350 965 20365 985
rect 20385 965 20400 985
rect 20350 935 20400 965
rect 20350 915 20365 935
rect 20385 915 20400 935
rect 20350 900 20400 915
rect -600 835 -350 850
rect -600 815 -585 835
rect -565 815 -535 835
rect -515 815 -485 835
rect -465 815 -435 835
rect -415 815 -385 835
rect -365 815 -350 835
rect -600 800 -350 815
rect -300 835 -50 850
rect -300 815 -285 835
rect -265 815 -235 835
rect -215 815 -185 835
rect -165 815 -135 835
rect -115 815 -85 835
rect -65 815 -50 835
rect -300 800 -50 815
rect 0 835 250 850
rect 0 815 15 835
rect 35 815 65 835
rect 85 815 115 835
rect 135 815 165 835
rect 185 815 215 835
rect 235 815 250 835
rect 0 800 250 815
rect 300 835 550 850
rect 300 815 315 835
rect 335 815 365 835
rect 385 815 415 835
rect 435 815 465 835
rect 485 815 515 835
rect 535 815 550 835
rect 300 800 550 815
rect 600 835 850 850
rect 600 815 615 835
rect 635 815 665 835
rect 685 815 715 835
rect 735 815 765 835
rect 785 815 815 835
rect 835 815 850 835
rect 600 800 850 815
rect 900 835 1150 850
rect 900 815 915 835
rect 935 815 965 835
rect 985 815 1015 835
rect 1035 815 1065 835
rect 1085 815 1115 835
rect 1135 815 1150 835
rect 900 800 1150 815
rect 1200 835 1450 850
rect 1200 815 1215 835
rect 1235 815 1265 835
rect 1285 815 1315 835
rect 1335 815 1365 835
rect 1385 815 1415 835
rect 1435 815 1450 835
rect 1200 800 1450 815
rect 1500 835 1750 850
rect 1500 815 1515 835
rect 1535 815 1565 835
rect 1585 815 1615 835
rect 1635 815 1665 835
rect 1685 815 1715 835
rect 1735 815 1750 835
rect 1500 800 1750 815
rect 1800 835 2050 850
rect 1800 815 1815 835
rect 1835 815 1865 835
rect 1885 815 1915 835
rect 1935 815 1965 835
rect 1985 815 2015 835
rect 2035 815 2050 835
rect 1800 800 2050 815
rect 2100 835 2350 850
rect 2100 815 2115 835
rect 2135 815 2165 835
rect 2185 815 2215 835
rect 2235 815 2265 835
rect 2285 815 2315 835
rect 2335 815 2350 835
rect 2100 800 2350 815
rect 2400 835 2650 850
rect 2400 815 2415 835
rect 2435 815 2465 835
rect 2485 815 2515 835
rect 2535 815 2565 835
rect 2585 815 2615 835
rect 2635 815 2650 835
rect 2400 800 2650 815
rect 2700 835 2950 850
rect 2700 815 2715 835
rect 2735 815 2765 835
rect 2785 815 2815 835
rect 2835 815 2865 835
rect 2885 815 2915 835
rect 2935 815 2950 835
rect 2700 800 2950 815
rect 3000 835 3250 850
rect 3000 815 3015 835
rect 3035 815 3065 835
rect 3085 815 3115 835
rect 3135 815 3165 835
rect 3185 815 3215 835
rect 3235 815 3250 835
rect 3000 800 3250 815
rect 3300 835 3550 850
rect 3300 815 3315 835
rect 3335 815 3365 835
rect 3385 815 3415 835
rect 3435 815 3465 835
rect 3485 815 3515 835
rect 3535 815 3550 835
rect 3300 800 3550 815
rect 3600 835 3850 850
rect 3600 815 3615 835
rect 3635 815 3665 835
rect 3685 815 3715 835
rect 3735 815 3765 835
rect 3785 815 3815 835
rect 3835 815 3850 835
rect 3600 800 3850 815
rect 3900 835 4150 850
rect 3900 815 3915 835
rect 3935 815 3965 835
rect 3985 815 4015 835
rect 4035 815 4065 835
rect 4085 815 4115 835
rect 4135 815 4150 835
rect 3900 800 4150 815
rect 4200 835 4450 850
rect 4200 815 4215 835
rect 4235 815 4265 835
rect 4285 815 4315 835
rect 4335 815 4365 835
rect 4385 815 4415 835
rect 4435 815 4450 835
rect 4200 800 4450 815
rect 4500 835 4750 850
rect 4500 815 4515 835
rect 4535 815 4565 835
rect 4585 815 4615 835
rect 4635 815 4665 835
rect 4685 815 4715 835
rect 4735 815 4750 835
rect 4500 800 4750 815
rect 4800 835 5050 850
rect 4800 815 4815 835
rect 4835 815 4865 835
rect 4885 815 4915 835
rect 4935 815 4965 835
rect 4985 815 5015 835
rect 5035 815 5050 835
rect 4800 800 5050 815
rect 5100 835 5350 850
rect 5100 815 5115 835
rect 5135 815 5165 835
rect 5185 815 5215 835
rect 5235 815 5265 835
rect 5285 815 5315 835
rect 5335 815 5350 835
rect 5100 800 5350 815
rect 5400 835 5650 850
rect 5400 815 5415 835
rect 5435 815 5465 835
rect 5485 815 5515 835
rect 5535 815 5565 835
rect 5585 815 5615 835
rect 5635 815 5650 835
rect 5400 800 5650 815
rect 5700 835 5950 850
rect 5700 815 5715 835
rect 5735 815 5765 835
rect 5785 815 5815 835
rect 5835 815 5865 835
rect 5885 815 5915 835
rect 5935 815 5950 835
rect 5700 800 5950 815
rect 6000 835 6250 850
rect 6000 815 6015 835
rect 6035 815 6065 835
rect 6085 815 6115 835
rect 6135 815 6165 835
rect 6185 815 6215 835
rect 6235 815 6250 835
rect 6000 800 6250 815
rect 6300 835 6550 850
rect 6300 815 6315 835
rect 6335 815 6365 835
rect 6385 815 6415 835
rect 6435 815 6465 835
rect 6485 815 6515 835
rect 6535 815 6550 835
rect 6300 800 6550 815
rect 6600 835 6850 850
rect 6600 815 6615 835
rect 6635 815 6665 835
rect 6685 815 6715 835
rect 6735 815 6765 835
rect 6785 815 6815 835
rect 6835 815 6850 835
rect 6600 800 6850 815
rect 6900 835 7150 850
rect 6900 815 6915 835
rect 6935 815 6965 835
rect 6985 815 7015 835
rect 7035 815 7065 835
rect 7085 815 7115 835
rect 7135 815 7150 835
rect 6900 800 7150 815
rect 7200 835 7450 850
rect 7200 815 7215 835
rect 7235 815 7265 835
rect 7285 815 7315 835
rect 7335 815 7365 835
rect 7385 815 7415 835
rect 7435 815 7450 835
rect 7200 800 7450 815
rect 7500 835 7750 850
rect 7500 815 7515 835
rect 7535 815 7565 835
rect 7585 815 7615 835
rect 7635 815 7665 835
rect 7685 815 7715 835
rect 7735 815 7750 835
rect 7500 800 7750 815
rect 7800 835 8050 850
rect 7800 815 7815 835
rect 7835 815 7865 835
rect 7885 815 7915 835
rect 7935 815 7965 835
rect 7985 815 8015 835
rect 8035 815 8050 835
rect 7800 800 8050 815
rect 8100 835 8350 850
rect 8100 815 8115 835
rect 8135 815 8165 835
rect 8185 815 8215 835
rect 8235 815 8265 835
rect 8285 815 8315 835
rect 8335 815 8350 835
rect 8100 800 8350 815
rect 8400 835 8650 850
rect 8400 815 8415 835
rect 8435 815 8465 835
rect 8485 815 8515 835
rect 8535 815 8565 835
rect 8585 815 8615 835
rect 8635 815 8650 835
rect 8400 800 8650 815
rect 8700 835 8950 850
rect 8700 815 8715 835
rect 8735 815 8765 835
rect 8785 815 8815 835
rect 8835 815 8865 835
rect 8885 815 8915 835
rect 8935 815 8950 835
rect 8700 800 8950 815
rect 9000 835 9250 850
rect 9000 815 9015 835
rect 9035 815 9065 835
rect 9085 815 9115 835
rect 9135 815 9165 835
rect 9185 815 9215 835
rect 9235 815 9250 835
rect 9000 800 9250 815
rect 9300 835 9550 850
rect 9300 815 9315 835
rect 9335 815 9365 835
rect 9385 815 9415 835
rect 9435 815 9465 835
rect 9485 815 9515 835
rect 9535 815 9550 835
rect 9300 800 9550 815
rect 9600 835 9850 850
rect 9600 815 9615 835
rect 9635 815 9665 835
rect 9685 815 9715 835
rect 9735 815 9765 835
rect 9785 815 9815 835
rect 9835 815 9850 835
rect 9600 800 9850 815
rect 9900 835 10150 850
rect 9900 815 9915 835
rect 9935 815 9965 835
rect 9985 815 10015 835
rect 10035 815 10065 835
rect 10085 815 10115 835
rect 10135 815 10150 835
rect 9900 800 10150 815
rect 10200 835 10450 850
rect 10200 815 10215 835
rect 10235 815 10265 835
rect 10285 815 10315 835
rect 10335 815 10365 835
rect 10385 815 10415 835
rect 10435 815 10450 835
rect 10200 800 10450 815
rect 10500 835 10750 850
rect 10500 815 10515 835
rect 10535 815 10565 835
rect 10585 815 10615 835
rect 10635 815 10665 835
rect 10685 815 10715 835
rect 10735 815 10750 835
rect 10500 800 10750 815
rect 10800 835 11050 850
rect 10800 815 10815 835
rect 10835 815 10865 835
rect 10885 815 10915 835
rect 10935 815 10965 835
rect 10985 815 11015 835
rect 11035 815 11050 835
rect 10800 800 11050 815
rect 11100 835 11350 850
rect 11100 815 11115 835
rect 11135 815 11165 835
rect 11185 815 11215 835
rect 11235 815 11265 835
rect 11285 815 11315 835
rect 11335 815 11350 835
rect 11100 800 11350 815
rect 11400 835 11650 850
rect 11400 815 11415 835
rect 11435 815 11465 835
rect 11485 815 11515 835
rect 11535 815 11565 835
rect 11585 815 11615 835
rect 11635 815 11650 835
rect 11400 800 11650 815
rect 11700 835 11950 850
rect 11700 815 11715 835
rect 11735 815 11765 835
rect 11785 815 11815 835
rect 11835 815 11865 835
rect 11885 815 11915 835
rect 11935 815 11950 835
rect 11700 800 11950 815
rect 12000 835 12250 850
rect 12000 815 12015 835
rect 12035 815 12065 835
rect 12085 815 12115 835
rect 12135 815 12165 835
rect 12185 815 12215 835
rect 12235 815 12250 835
rect 12000 800 12250 815
rect 12300 835 12550 850
rect 12300 815 12315 835
rect 12335 815 12365 835
rect 12385 815 12415 835
rect 12435 815 12465 835
rect 12485 815 12515 835
rect 12535 815 12550 835
rect 12300 800 12550 815
rect 12600 835 12850 850
rect 12600 815 12615 835
rect 12635 815 12665 835
rect 12685 815 12715 835
rect 12735 815 12765 835
rect 12785 815 12815 835
rect 12835 815 12850 835
rect 12600 800 12850 815
rect 12900 835 13150 850
rect 12900 815 12915 835
rect 12935 815 12965 835
rect 12985 815 13015 835
rect 13035 815 13065 835
rect 13085 815 13115 835
rect 13135 815 13150 835
rect 12900 800 13150 815
rect 13200 835 13450 850
rect 13200 815 13215 835
rect 13235 815 13265 835
rect 13285 815 13315 835
rect 13335 815 13365 835
rect 13385 815 13415 835
rect 13435 815 13450 835
rect 13200 800 13450 815
rect 13500 835 13750 850
rect 13500 815 13515 835
rect 13535 815 13565 835
rect 13585 815 13615 835
rect 13635 815 13665 835
rect 13685 815 13715 835
rect 13735 815 13750 835
rect 13500 800 13750 815
rect 13800 835 14050 850
rect 13800 815 13815 835
rect 13835 815 13865 835
rect 13885 815 13915 835
rect 13935 815 13965 835
rect 13985 815 14015 835
rect 14035 815 14050 835
rect 13800 800 14050 815
rect 14100 835 14350 850
rect 14100 815 14115 835
rect 14135 815 14165 835
rect 14185 815 14215 835
rect 14235 815 14265 835
rect 14285 815 14315 835
rect 14335 815 14350 835
rect 14100 800 14350 815
rect 14400 835 14650 850
rect 14400 815 14415 835
rect 14435 815 14465 835
rect 14485 815 14515 835
rect 14535 815 14565 835
rect 14585 815 14615 835
rect 14635 815 14650 835
rect 14400 800 14650 815
rect 14700 835 14950 850
rect 14700 815 14715 835
rect 14735 815 14765 835
rect 14785 815 14815 835
rect 14835 815 14865 835
rect 14885 815 14915 835
rect 14935 815 14950 835
rect 14700 800 14950 815
rect 15000 835 15250 850
rect 15000 815 15015 835
rect 15035 815 15065 835
rect 15085 815 15115 835
rect 15135 815 15165 835
rect 15185 815 15215 835
rect 15235 815 15250 835
rect 15000 800 15250 815
rect 15300 835 15550 850
rect 15300 815 15315 835
rect 15335 815 15365 835
rect 15385 815 15415 835
rect 15435 815 15465 835
rect 15485 815 15515 835
rect 15535 815 15550 835
rect 15300 800 15550 815
rect 15600 835 15850 850
rect 15600 815 15615 835
rect 15635 815 15665 835
rect 15685 815 15715 835
rect 15735 815 15765 835
rect 15785 815 15815 835
rect 15835 815 15850 835
rect 15600 800 15850 815
rect 15900 835 16150 850
rect 15900 815 15915 835
rect 15935 815 15965 835
rect 15985 815 16015 835
rect 16035 815 16065 835
rect 16085 815 16115 835
rect 16135 815 16150 835
rect 15900 800 16150 815
rect 16200 835 16450 850
rect 16200 815 16215 835
rect 16235 815 16265 835
rect 16285 815 16315 835
rect 16335 815 16365 835
rect 16385 815 16415 835
rect 16435 815 16450 835
rect 16200 800 16450 815
rect 16500 835 16750 850
rect 16500 815 16515 835
rect 16535 815 16565 835
rect 16585 815 16615 835
rect 16635 815 16665 835
rect 16685 815 16715 835
rect 16735 815 16750 835
rect 16500 800 16750 815
rect 16800 835 17050 850
rect 16800 815 16815 835
rect 16835 815 16865 835
rect 16885 815 16915 835
rect 16935 815 16965 835
rect 16985 815 17015 835
rect 17035 815 17050 835
rect 16800 800 17050 815
rect 17100 835 17350 850
rect 17100 815 17115 835
rect 17135 815 17165 835
rect 17185 815 17215 835
rect 17235 815 17265 835
rect 17285 815 17315 835
rect 17335 815 17350 835
rect 17100 800 17350 815
rect 17400 835 17650 850
rect 17400 815 17415 835
rect 17435 815 17465 835
rect 17485 815 17515 835
rect 17535 815 17565 835
rect 17585 815 17615 835
rect 17635 815 17650 835
rect 17400 800 17650 815
rect 17700 835 17950 850
rect 17700 815 17715 835
rect 17735 815 17765 835
rect 17785 815 17815 835
rect 17835 815 17865 835
rect 17885 815 17915 835
rect 17935 815 17950 835
rect 17700 800 17950 815
rect 18000 835 18250 850
rect 18000 815 18015 835
rect 18035 815 18065 835
rect 18085 815 18115 835
rect 18135 815 18165 835
rect 18185 815 18215 835
rect 18235 815 18250 835
rect 18000 800 18250 815
rect 18300 835 18550 850
rect 18300 815 18315 835
rect 18335 815 18365 835
rect 18385 815 18415 835
rect 18435 815 18465 835
rect 18485 815 18515 835
rect 18535 815 18550 835
rect 18300 800 18550 815
rect 18600 835 18850 850
rect 18600 815 18615 835
rect 18635 815 18665 835
rect 18685 815 18715 835
rect 18735 815 18765 835
rect 18785 815 18815 835
rect 18835 815 18850 835
rect 18600 800 18850 815
rect 18900 835 19150 850
rect 18900 815 18915 835
rect 18935 815 18965 835
rect 18985 815 19015 835
rect 19035 815 19065 835
rect 19085 815 19115 835
rect 19135 815 19150 835
rect 18900 800 19150 815
rect 19200 835 19450 850
rect 19200 815 19215 835
rect 19235 815 19265 835
rect 19285 815 19315 835
rect 19335 815 19365 835
rect 19385 815 19415 835
rect 19435 815 19450 835
rect 19200 800 19450 815
rect 19500 835 19750 850
rect 19500 815 19515 835
rect 19535 815 19565 835
rect 19585 815 19615 835
rect 19635 815 19665 835
rect 19685 815 19715 835
rect 19735 815 19750 835
rect 19500 800 19750 815
rect 19800 835 20050 850
rect 19800 815 19815 835
rect 19835 815 19865 835
rect 19885 815 19915 835
rect 19935 815 19965 835
rect 19985 815 20015 835
rect 20035 815 20050 835
rect 19800 800 20050 815
rect 20100 835 20350 850
rect 20100 815 20115 835
rect 20135 815 20165 835
rect 20185 815 20215 835
rect 20235 815 20265 835
rect 20285 815 20315 835
rect 20335 815 20350 835
rect 20100 800 20350 815
rect -650 735 -600 750
rect -650 715 -635 735
rect -615 715 -600 735
rect -650 685 -600 715
rect -650 665 -635 685
rect -615 665 -600 685
rect -650 635 -600 665
rect -650 615 -635 635
rect -615 615 -600 635
rect -650 585 -600 615
rect -650 565 -635 585
rect -615 565 -600 585
rect -650 535 -600 565
rect -650 515 -635 535
rect -615 515 -600 535
rect -650 485 -600 515
rect -650 465 -635 485
rect -615 465 -600 485
rect -650 435 -600 465
rect -650 415 -635 435
rect -615 415 -600 435
rect -650 385 -600 415
rect -650 365 -635 385
rect -615 365 -600 385
rect -650 335 -600 365
rect -650 315 -635 335
rect -615 315 -600 335
rect -650 285 -600 315
rect -650 265 -635 285
rect -615 265 -600 285
rect -650 235 -600 265
rect -650 215 -635 235
rect -615 215 -600 235
rect -650 185 -600 215
rect -650 165 -635 185
rect -615 165 -600 185
rect -650 135 -600 165
rect -650 115 -635 135
rect -615 115 -600 135
rect -650 85 -600 115
rect -650 65 -635 85
rect -615 65 -600 85
rect -650 50 -600 65
rect -500 735 -450 750
rect -500 715 -485 735
rect -465 715 -450 735
rect -500 685 -450 715
rect -500 665 -485 685
rect -465 665 -450 685
rect -500 635 -450 665
rect -500 615 -485 635
rect -465 615 -450 635
rect -500 585 -450 615
rect -500 565 -485 585
rect -465 565 -450 585
rect -500 535 -450 565
rect -500 515 -485 535
rect -465 515 -450 535
rect -500 485 -450 515
rect -500 465 -485 485
rect -465 465 -450 485
rect -500 435 -450 465
rect -500 415 -485 435
rect -465 415 -450 435
rect -500 385 -450 415
rect -500 365 -485 385
rect -465 365 -450 385
rect -500 335 -450 365
rect -500 315 -485 335
rect -465 315 -450 335
rect -500 285 -450 315
rect -500 265 -485 285
rect -465 265 -450 285
rect -500 235 -450 265
rect -500 215 -485 235
rect -465 215 -450 235
rect -500 185 -450 215
rect -500 165 -485 185
rect -465 165 -450 185
rect -500 135 -450 165
rect -500 115 -485 135
rect -465 115 -450 135
rect -500 85 -450 115
rect -500 65 -485 85
rect -465 65 -450 85
rect -500 50 -450 65
rect -350 735 -300 750
rect -350 715 -335 735
rect -315 715 -300 735
rect -350 685 -300 715
rect -350 665 -335 685
rect -315 665 -300 685
rect -350 635 -300 665
rect -350 615 -335 635
rect -315 615 -300 635
rect -350 585 -300 615
rect -350 565 -335 585
rect -315 565 -300 585
rect -350 535 -300 565
rect -350 515 -335 535
rect -315 515 -300 535
rect -350 485 -300 515
rect -350 465 -335 485
rect -315 465 -300 485
rect -350 435 -300 465
rect -350 415 -335 435
rect -315 415 -300 435
rect -350 385 -300 415
rect -350 365 -335 385
rect -315 365 -300 385
rect -350 335 -300 365
rect -350 315 -335 335
rect -315 315 -300 335
rect -350 285 -300 315
rect -350 265 -335 285
rect -315 265 -300 285
rect -350 235 -300 265
rect -350 215 -335 235
rect -315 215 -300 235
rect -350 185 -300 215
rect -350 165 -335 185
rect -315 165 -300 185
rect -350 135 -300 165
rect -350 115 -335 135
rect -315 115 -300 135
rect -350 85 -300 115
rect -350 65 -335 85
rect -315 65 -300 85
rect -350 50 -300 65
rect -200 735 -150 750
rect -200 715 -185 735
rect -165 715 -150 735
rect -200 685 -150 715
rect -200 665 -185 685
rect -165 665 -150 685
rect -200 635 -150 665
rect -200 615 -185 635
rect -165 615 -150 635
rect -200 585 -150 615
rect -200 565 -185 585
rect -165 565 -150 585
rect -200 535 -150 565
rect -200 515 -185 535
rect -165 515 -150 535
rect -200 485 -150 515
rect -200 465 -185 485
rect -165 465 -150 485
rect -200 435 -150 465
rect -200 415 -185 435
rect -165 415 -150 435
rect -200 385 -150 415
rect -200 365 -185 385
rect -165 365 -150 385
rect -200 335 -150 365
rect -200 315 -185 335
rect -165 315 -150 335
rect -200 285 -150 315
rect -200 265 -185 285
rect -165 265 -150 285
rect -200 235 -150 265
rect -200 215 -185 235
rect -165 215 -150 235
rect -200 185 -150 215
rect -200 165 -185 185
rect -165 165 -150 185
rect -200 135 -150 165
rect -200 115 -185 135
rect -165 115 -150 135
rect -200 85 -150 115
rect -200 65 -185 85
rect -165 65 -150 85
rect -200 50 -150 65
rect -50 735 0 750
rect -50 715 -35 735
rect -15 715 0 735
rect -50 685 0 715
rect -50 665 -35 685
rect -15 665 0 685
rect -50 635 0 665
rect -50 615 -35 635
rect -15 615 0 635
rect -50 585 0 615
rect -50 565 -35 585
rect -15 565 0 585
rect -50 535 0 565
rect -50 515 -35 535
rect -15 515 0 535
rect -50 485 0 515
rect -50 465 -35 485
rect -15 465 0 485
rect -50 435 0 465
rect -50 415 -35 435
rect -15 415 0 435
rect -50 385 0 415
rect -50 365 -35 385
rect -15 365 0 385
rect -50 335 0 365
rect -50 315 -35 335
rect -15 315 0 335
rect -50 285 0 315
rect -50 265 -35 285
rect -15 265 0 285
rect -50 235 0 265
rect -50 215 -35 235
rect -15 215 0 235
rect -50 185 0 215
rect -50 165 -35 185
rect -15 165 0 185
rect -50 135 0 165
rect -50 115 -35 135
rect -15 115 0 135
rect -50 85 0 115
rect -50 65 -35 85
rect -15 65 0 85
rect -50 50 0 65
rect 1150 735 1200 750
rect 1150 715 1165 735
rect 1185 715 1200 735
rect 1150 685 1200 715
rect 1150 665 1165 685
rect 1185 665 1200 685
rect 1150 635 1200 665
rect 1150 615 1165 635
rect 1185 615 1200 635
rect 1150 585 1200 615
rect 1150 565 1165 585
rect 1185 565 1200 585
rect 1150 535 1200 565
rect 1150 515 1165 535
rect 1185 515 1200 535
rect 1150 485 1200 515
rect 1150 465 1165 485
rect 1185 465 1200 485
rect 1150 435 1200 465
rect 1150 415 1165 435
rect 1185 415 1200 435
rect 1150 385 1200 415
rect 1150 365 1165 385
rect 1185 365 1200 385
rect 1150 335 1200 365
rect 1150 315 1165 335
rect 1185 315 1200 335
rect 1150 285 1200 315
rect 1150 265 1165 285
rect 1185 265 1200 285
rect 1150 235 1200 265
rect 1150 215 1165 235
rect 1185 215 1200 235
rect 1150 185 1200 215
rect 1150 165 1165 185
rect 1185 165 1200 185
rect 1150 135 1200 165
rect 1150 115 1165 135
rect 1185 115 1200 135
rect 1150 85 1200 115
rect 1150 65 1165 85
rect 1185 65 1200 85
rect 1150 50 1200 65
rect 1450 735 1500 750
rect 1450 715 1465 735
rect 1485 715 1500 735
rect 1450 685 1500 715
rect 1450 665 1465 685
rect 1485 665 1500 685
rect 1450 635 1500 665
rect 1450 615 1465 635
rect 1485 615 1500 635
rect 1450 585 1500 615
rect 1450 565 1465 585
rect 1485 565 1500 585
rect 1450 535 1500 565
rect 1450 515 1465 535
rect 1485 515 1500 535
rect 1450 485 1500 515
rect 1450 465 1465 485
rect 1485 465 1500 485
rect 1450 435 1500 465
rect 1450 415 1465 435
rect 1485 415 1500 435
rect 1450 385 1500 415
rect 1450 365 1465 385
rect 1485 365 1500 385
rect 1450 335 1500 365
rect 1450 315 1465 335
rect 1485 315 1500 335
rect 1450 285 1500 315
rect 1450 265 1465 285
rect 1485 265 1500 285
rect 1450 235 1500 265
rect 1450 215 1465 235
rect 1485 215 1500 235
rect 1450 185 1500 215
rect 1450 165 1465 185
rect 1485 165 1500 185
rect 1450 135 1500 165
rect 1450 115 1465 135
rect 1485 115 1500 135
rect 1450 85 1500 115
rect 1450 65 1465 85
rect 1485 65 1500 85
rect 1450 50 1500 65
rect 1750 735 1800 750
rect 1750 715 1765 735
rect 1785 715 1800 735
rect 1750 685 1800 715
rect 1750 665 1765 685
rect 1785 665 1800 685
rect 1750 635 1800 665
rect 1750 615 1765 635
rect 1785 615 1800 635
rect 1750 585 1800 615
rect 1750 565 1765 585
rect 1785 565 1800 585
rect 1750 535 1800 565
rect 1750 515 1765 535
rect 1785 515 1800 535
rect 1750 485 1800 515
rect 1750 465 1765 485
rect 1785 465 1800 485
rect 1750 435 1800 465
rect 1750 415 1765 435
rect 1785 415 1800 435
rect 1750 385 1800 415
rect 1750 365 1765 385
rect 1785 365 1800 385
rect 1750 335 1800 365
rect 1750 315 1765 335
rect 1785 315 1800 335
rect 1750 285 1800 315
rect 1750 265 1765 285
rect 1785 265 1800 285
rect 1750 235 1800 265
rect 1750 215 1765 235
rect 1785 215 1800 235
rect 1750 185 1800 215
rect 1750 165 1765 185
rect 1785 165 1800 185
rect 1750 135 1800 165
rect 1750 115 1765 135
rect 1785 115 1800 135
rect 1750 85 1800 115
rect 1750 65 1765 85
rect 1785 65 1800 85
rect 1750 50 1800 65
rect 2050 735 2100 750
rect 2050 715 2065 735
rect 2085 715 2100 735
rect 2050 685 2100 715
rect 2050 665 2065 685
rect 2085 665 2100 685
rect 2050 635 2100 665
rect 2050 615 2065 635
rect 2085 615 2100 635
rect 2050 585 2100 615
rect 2050 565 2065 585
rect 2085 565 2100 585
rect 2050 535 2100 565
rect 2050 515 2065 535
rect 2085 515 2100 535
rect 2050 485 2100 515
rect 2050 465 2065 485
rect 2085 465 2100 485
rect 2050 435 2100 465
rect 2050 415 2065 435
rect 2085 415 2100 435
rect 2050 385 2100 415
rect 2050 365 2065 385
rect 2085 365 2100 385
rect 2050 335 2100 365
rect 2050 315 2065 335
rect 2085 315 2100 335
rect 2050 285 2100 315
rect 2050 265 2065 285
rect 2085 265 2100 285
rect 2050 235 2100 265
rect 2050 215 2065 235
rect 2085 215 2100 235
rect 2050 185 2100 215
rect 2050 165 2065 185
rect 2085 165 2100 185
rect 2050 135 2100 165
rect 2050 115 2065 135
rect 2085 115 2100 135
rect 2050 85 2100 115
rect 2050 65 2065 85
rect 2085 65 2100 85
rect 2050 50 2100 65
rect 2350 735 2400 750
rect 2350 715 2365 735
rect 2385 715 2400 735
rect 2350 685 2400 715
rect 2350 665 2365 685
rect 2385 665 2400 685
rect 2350 635 2400 665
rect 2350 615 2365 635
rect 2385 615 2400 635
rect 2350 585 2400 615
rect 2350 565 2365 585
rect 2385 565 2400 585
rect 2350 535 2400 565
rect 2350 515 2365 535
rect 2385 515 2400 535
rect 2350 485 2400 515
rect 2350 465 2365 485
rect 2385 465 2400 485
rect 2350 435 2400 465
rect 2350 415 2365 435
rect 2385 415 2400 435
rect 2350 385 2400 415
rect 2350 365 2365 385
rect 2385 365 2400 385
rect 2350 335 2400 365
rect 2350 315 2365 335
rect 2385 315 2400 335
rect 2350 285 2400 315
rect 2350 265 2365 285
rect 2385 265 2400 285
rect 2350 235 2400 265
rect 2350 215 2365 235
rect 2385 215 2400 235
rect 2350 185 2400 215
rect 2350 165 2365 185
rect 2385 165 2400 185
rect 2350 135 2400 165
rect 2350 115 2365 135
rect 2385 115 2400 135
rect 2350 85 2400 115
rect 2350 65 2365 85
rect 2385 65 2400 85
rect 2350 50 2400 65
rect 2650 735 2700 750
rect 2650 715 2665 735
rect 2685 715 2700 735
rect 2650 685 2700 715
rect 2650 665 2665 685
rect 2685 665 2700 685
rect 2650 635 2700 665
rect 2650 615 2665 635
rect 2685 615 2700 635
rect 2650 585 2700 615
rect 2650 565 2665 585
rect 2685 565 2700 585
rect 2650 535 2700 565
rect 2650 515 2665 535
rect 2685 515 2700 535
rect 2650 485 2700 515
rect 2650 465 2665 485
rect 2685 465 2700 485
rect 2650 435 2700 465
rect 2650 415 2665 435
rect 2685 415 2700 435
rect 2650 385 2700 415
rect 2650 365 2665 385
rect 2685 365 2700 385
rect 2650 335 2700 365
rect 2650 315 2665 335
rect 2685 315 2700 335
rect 2650 285 2700 315
rect 2650 265 2665 285
rect 2685 265 2700 285
rect 2650 235 2700 265
rect 2650 215 2665 235
rect 2685 215 2700 235
rect 2650 185 2700 215
rect 2650 165 2665 185
rect 2685 165 2700 185
rect 2650 135 2700 165
rect 2650 115 2665 135
rect 2685 115 2700 135
rect 2650 85 2700 115
rect 2650 65 2665 85
rect 2685 65 2700 85
rect 2650 50 2700 65
rect 2950 735 3000 750
rect 2950 715 2965 735
rect 2985 715 3000 735
rect 2950 685 3000 715
rect 2950 665 2965 685
rect 2985 665 3000 685
rect 2950 635 3000 665
rect 2950 615 2965 635
rect 2985 615 3000 635
rect 2950 585 3000 615
rect 2950 565 2965 585
rect 2985 565 3000 585
rect 2950 535 3000 565
rect 2950 515 2965 535
rect 2985 515 3000 535
rect 2950 485 3000 515
rect 2950 465 2965 485
rect 2985 465 3000 485
rect 2950 435 3000 465
rect 2950 415 2965 435
rect 2985 415 3000 435
rect 2950 385 3000 415
rect 2950 365 2965 385
rect 2985 365 3000 385
rect 2950 335 3000 365
rect 2950 315 2965 335
rect 2985 315 3000 335
rect 2950 285 3000 315
rect 2950 265 2965 285
rect 2985 265 3000 285
rect 2950 235 3000 265
rect 2950 215 2965 235
rect 2985 215 3000 235
rect 2950 185 3000 215
rect 2950 165 2965 185
rect 2985 165 3000 185
rect 2950 135 3000 165
rect 2950 115 2965 135
rect 2985 115 3000 135
rect 2950 85 3000 115
rect 2950 65 2965 85
rect 2985 65 3000 85
rect 2950 50 3000 65
rect 3250 735 3300 750
rect 3250 715 3265 735
rect 3285 715 3300 735
rect 3250 685 3300 715
rect 3250 665 3265 685
rect 3285 665 3300 685
rect 3250 635 3300 665
rect 3250 615 3265 635
rect 3285 615 3300 635
rect 3250 585 3300 615
rect 3250 565 3265 585
rect 3285 565 3300 585
rect 3250 535 3300 565
rect 3250 515 3265 535
rect 3285 515 3300 535
rect 3250 485 3300 515
rect 3250 465 3265 485
rect 3285 465 3300 485
rect 3250 435 3300 465
rect 3250 415 3265 435
rect 3285 415 3300 435
rect 3250 385 3300 415
rect 3250 365 3265 385
rect 3285 365 3300 385
rect 3250 335 3300 365
rect 3250 315 3265 335
rect 3285 315 3300 335
rect 3250 285 3300 315
rect 3250 265 3265 285
rect 3285 265 3300 285
rect 3250 235 3300 265
rect 3250 215 3265 235
rect 3285 215 3300 235
rect 3250 185 3300 215
rect 3250 165 3265 185
rect 3285 165 3300 185
rect 3250 135 3300 165
rect 3250 115 3265 135
rect 3285 115 3300 135
rect 3250 85 3300 115
rect 3250 65 3265 85
rect 3285 65 3300 85
rect 3250 50 3300 65
rect 3550 735 3600 750
rect 3550 715 3565 735
rect 3585 715 3600 735
rect 3550 685 3600 715
rect 3550 665 3565 685
rect 3585 665 3600 685
rect 3550 635 3600 665
rect 3550 615 3565 635
rect 3585 615 3600 635
rect 3550 585 3600 615
rect 3550 565 3565 585
rect 3585 565 3600 585
rect 3550 535 3600 565
rect 3550 515 3565 535
rect 3585 515 3600 535
rect 3550 485 3600 515
rect 3550 465 3565 485
rect 3585 465 3600 485
rect 3550 435 3600 465
rect 3550 415 3565 435
rect 3585 415 3600 435
rect 3550 385 3600 415
rect 3550 365 3565 385
rect 3585 365 3600 385
rect 3550 335 3600 365
rect 3550 315 3565 335
rect 3585 315 3600 335
rect 3550 285 3600 315
rect 3550 265 3565 285
rect 3585 265 3600 285
rect 3550 235 3600 265
rect 3550 215 3565 235
rect 3585 215 3600 235
rect 3550 185 3600 215
rect 3550 165 3565 185
rect 3585 165 3600 185
rect 3550 135 3600 165
rect 3550 115 3565 135
rect 3585 115 3600 135
rect 3550 85 3600 115
rect 3550 65 3565 85
rect 3585 65 3600 85
rect 3550 50 3600 65
rect 3700 735 3750 750
rect 3700 715 3715 735
rect 3735 715 3750 735
rect 3700 685 3750 715
rect 3700 665 3715 685
rect 3735 665 3750 685
rect 3700 635 3750 665
rect 3700 615 3715 635
rect 3735 615 3750 635
rect 3700 585 3750 615
rect 3700 565 3715 585
rect 3735 565 3750 585
rect 3700 535 3750 565
rect 3700 515 3715 535
rect 3735 515 3750 535
rect 3700 485 3750 515
rect 3700 465 3715 485
rect 3735 465 3750 485
rect 3700 435 3750 465
rect 3700 415 3715 435
rect 3735 415 3750 435
rect 3700 385 3750 415
rect 3700 365 3715 385
rect 3735 365 3750 385
rect 3700 335 3750 365
rect 3700 315 3715 335
rect 3735 315 3750 335
rect 3700 285 3750 315
rect 3700 265 3715 285
rect 3735 265 3750 285
rect 3700 235 3750 265
rect 3700 215 3715 235
rect 3735 215 3750 235
rect 3700 185 3750 215
rect 3700 165 3715 185
rect 3735 165 3750 185
rect 3700 135 3750 165
rect 3700 115 3715 135
rect 3735 115 3750 135
rect 3700 85 3750 115
rect 3700 65 3715 85
rect 3735 65 3750 85
rect 3700 50 3750 65
rect 3850 735 3900 750
rect 3850 715 3865 735
rect 3885 715 3900 735
rect 3850 685 3900 715
rect 3850 665 3865 685
rect 3885 665 3900 685
rect 3850 635 3900 665
rect 3850 615 3865 635
rect 3885 615 3900 635
rect 3850 585 3900 615
rect 3850 565 3865 585
rect 3885 565 3900 585
rect 3850 535 3900 565
rect 3850 515 3865 535
rect 3885 515 3900 535
rect 3850 485 3900 515
rect 3850 465 3865 485
rect 3885 465 3900 485
rect 3850 435 3900 465
rect 3850 415 3865 435
rect 3885 415 3900 435
rect 3850 385 3900 415
rect 3850 365 3865 385
rect 3885 365 3900 385
rect 3850 335 3900 365
rect 3850 315 3865 335
rect 3885 315 3900 335
rect 3850 285 3900 315
rect 3850 265 3865 285
rect 3885 265 3900 285
rect 3850 235 3900 265
rect 3850 215 3865 235
rect 3885 215 3900 235
rect 3850 185 3900 215
rect 3850 165 3865 185
rect 3885 165 3900 185
rect 3850 135 3900 165
rect 3850 115 3865 135
rect 3885 115 3900 135
rect 3850 85 3900 115
rect 3850 65 3865 85
rect 3885 65 3900 85
rect 3850 50 3900 65
rect 4000 735 4050 750
rect 4000 715 4015 735
rect 4035 715 4050 735
rect 4000 685 4050 715
rect 4000 665 4015 685
rect 4035 665 4050 685
rect 4000 635 4050 665
rect 4000 615 4015 635
rect 4035 615 4050 635
rect 4000 585 4050 615
rect 4000 565 4015 585
rect 4035 565 4050 585
rect 4000 535 4050 565
rect 4000 515 4015 535
rect 4035 515 4050 535
rect 4000 485 4050 515
rect 4000 465 4015 485
rect 4035 465 4050 485
rect 4000 435 4050 465
rect 4000 415 4015 435
rect 4035 415 4050 435
rect 4000 385 4050 415
rect 4000 365 4015 385
rect 4035 365 4050 385
rect 4000 335 4050 365
rect 4000 315 4015 335
rect 4035 315 4050 335
rect 4000 285 4050 315
rect 4000 265 4015 285
rect 4035 265 4050 285
rect 4000 235 4050 265
rect 4000 215 4015 235
rect 4035 215 4050 235
rect 4000 185 4050 215
rect 4000 165 4015 185
rect 4035 165 4050 185
rect 4000 135 4050 165
rect 4000 115 4015 135
rect 4035 115 4050 135
rect 4000 85 4050 115
rect 4000 65 4015 85
rect 4035 65 4050 85
rect 4000 50 4050 65
rect 4150 735 4200 750
rect 4150 715 4165 735
rect 4185 715 4200 735
rect 4150 685 4200 715
rect 4150 665 4165 685
rect 4185 665 4200 685
rect 4150 635 4200 665
rect 4150 615 4165 635
rect 4185 615 4200 635
rect 4150 585 4200 615
rect 4150 565 4165 585
rect 4185 565 4200 585
rect 4150 535 4200 565
rect 4150 515 4165 535
rect 4185 515 4200 535
rect 4150 485 4200 515
rect 4150 465 4165 485
rect 4185 465 4200 485
rect 4150 435 4200 465
rect 4150 415 4165 435
rect 4185 415 4200 435
rect 4150 385 4200 415
rect 4150 365 4165 385
rect 4185 365 4200 385
rect 4150 335 4200 365
rect 4150 315 4165 335
rect 4185 315 4200 335
rect 4150 285 4200 315
rect 4150 265 4165 285
rect 4185 265 4200 285
rect 4150 235 4200 265
rect 4150 215 4165 235
rect 4185 215 4200 235
rect 4150 185 4200 215
rect 4150 165 4165 185
rect 4185 165 4200 185
rect 4150 135 4200 165
rect 4150 115 4165 135
rect 4185 115 4200 135
rect 4150 85 4200 115
rect 4150 65 4165 85
rect 4185 65 4200 85
rect 4150 50 4200 65
rect 4300 735 4350 750
rect 4300 715 4315 735
rect 4335 715 4350 735
rect 4300 685 4350 715
rect 4300 665 4315 685
rect 4335 665 4350 685
rect 4300 635 4350 665
rect 4300 615 4315 635
rect 4335 615 4350 635
rect 4300 585 4350 615
rect 4300 565 4315 585
rect 4335 565 4350 585
rect 4300 535 4350 565
rect 4300 515 4315 535
rect 4335 515 4350 535
rect 4300 485 4350 515
rect 4300 465 4315 485
rect 4335 465 4350 485
rect 4300 435 4350 465
rect 4300 415 4315 435
rect 4335 415 4350 435
rect 4300 385 4350 415
rect 4300 365 4315 385
rect 4335 365 4350 385
rect 4300 335 4350 365
rect 4300 315 4315 335
rect 4335 315 4350 335
rect 4300 285 4350 315
rect 4300 265 4315 285
rect 4335 265 4350 285
rect 4300 235 4350 265
rect 4300 215 4315 235
rect 4335 215 4350 235
rect 4300 185 4350 215
rect 4300 165 4315 185
rect 4335 165 4350 185
rect 4300 135 4350 165
rect 4300 115 4315 135
rect 4335 115 4350 135
rect 4300 85 4350 115
rect 4300 65 4315 85
rect 4335 65 4350 85
rect 4300 50 4350 65
rect 4450 735 4500 750
rect 4450 715 4465 735
rect 4485 715 4500 735
rect 4450 685 4500 715
rect 4450 665 4465 685
rect 4485 665 4500 685
rect 4450 635 4500 665
rect 4450 615 4465 635
rect 4485 615 4500 635
rect 4450 585 4500 615
rect 4450 565 4465 585
rect 4485 565 4500 585
rect 4450 535 4500 565
rect 4450 515 4465 535
rect 4485 515 4500 535
rect 4450 485 4500 515
rect 4450 465 4465 485
rect 4485 465 4500 485
rect 4450 435 4500 465
rect 4450 415 4465 435
rect 4485 415 4500 435
rect 4450 385 4500 415
rect 4450 365 4465 385
rect 4485 365 4500 385
rect 4450 335 4500 365
rect 4450 315 4465 335
rect 4485 315 4500 335
rect 4450 285 4500 315
rect 4450 265 4465 285
rect 4485 265 4500 285
rect 4450 235 4500 265
rect 4450 215 4465 235
rect 4485 215 4500 235
rect 4450 185 4500 215
rect 4450 165 4465 185
rect 4485 165 4500 185
rect 4450 135 4500 165
rect 4450 115 4465 135
rect 4485 115 4500 135
rect 4450 85 4500 115
rect 4450 65 4465 85
rect 4485 65 4500 85
rect 4450 50 4500 65
rect 4600 735 4650 750
rect 4600 715 4615 735
rect 4635 715 4650 735
rect 4600 685 4650 715
rect 4600 665 4615 685
rect 4635 665 4650 685
rect 4600 635 4650 665
rect 4600 615 4615 635
rect 4635 615 4650 635
rect 4600 585 4650 615
rect 4600 565 4615 585
rect 4635 565 4650 585
rect 4600 535 4650 565
rect 4600 515 4615 535
rect 4635 515 4650 535
rect 4600 485 4650 515
rect 4600 465 4615 485
rect 4635 465 4650 485
rect 4600 435 4650 465
rect 4600 415 4615 435
rect 4635 415 4650 435
rect 4600 385 4650 415
rect 4600 365 4615 385
rect 4635 365 4650 385
rect 4600 335 4650 365
rect 4600 315 4615 335
rect 4635 315 4650 335
rect 4600 285 4650 315
rect 4600 265 4615 285
rect 4635 265 4650 285
rect 4600 235 4650 265
rect 4600 215 4615 235
rect 4635 215 4650 235
rect 4600 185 4650 215
rect 4600 165 4615 185
rect 4635 165 4650 185
rect 4600 135 4650 165
rect 4600 115 4615 135
rect 4635 115 4650 135
rect 4600 85 4650 115
rect 4600 65 4615 85
rect 4635 65 4650 85
rect 4600 50 4650 65
rect 4750 735 4800 750
rect 4750 715 4765 735
rect 4785 715 4800 735
rect 4750 685 4800 715
rect 4750 665 4765 685
rect 4785 665 4800 685
rect 4750 635 4800 665
rect 4750 615 4765 635
rect 4785 615 4800 635
rect 4750 585 4800 615
rect 4750 565 4765 585
rect 4785 565 4800 585
rect 4750 535 4800 565
rect 4750 515 4765 535
rect 4785 515 4800 535
rect 4750 485 4800 515
rect 4750 465 4765 485
rect 4785 465 4800 485
rect 4750 435 4800 465
rect 4750 415 4765 435
rect 4785 415 4800 435
rect 4750 385 4800 415
rect 4750 365 4765 385
rect 4785 365 4800 385
rect 4750 335 4800 365
rect 4750 315 4765 335
rect 4785 315 4800 335
rect 4750 285 4800 315
rect 4750 265 4765 285
rect 4785 265 4800 285
rect 4750 235 4800 265
rect 4750 215 4765 235
rect 4785 215 4800 235
rect 4750 185 4800 215
rect 4750 165 4765 185
rect 4785 165 4800 185
rect 4750 135 4800 165
rect 4750 115 4765 135
rect 4785 115 4800 135
rect 4750 85 4800 115
rect 4750 65 4765 85
rect 4785 65 4800 85
rect 4750 50 4800 65
rect 5050 735 5100 750
rect 5050 715 5065 735
rect 5085 715 5100 735
rect 5050 685 5100 715
rect 5050 665 5065 685
rect 5085 665 5100 685
rect 5050 635 5100 665
rect 5050 615 5065 635
rect 5085 615 5100 635
rect 5050 585 5100 615
rect 5050 565 5065 585
rect 5085 565 5100 585
rect 5050 535 5100 565
rect 5050 515 5065 535
rect 5085 515 5100 535
rect 5050 485 5100 515
rect 5050 465 5065 485
rect 5085 465 5100 485
rect 5050 435 5100 465
rect 5050 415 5065 435
rect 5085 415 5100 435
rect 5050 385 5100 415
rect 5050 365 5065 385
rect 5085 365 5100 385
rect 5050 335 5100 365
rect 5050 315 5065 335
rect 5085 315 5100 335
rect 5050 285 5100 315
rect 5050 265 5065 285
rect 5085 265 5100 285
rect 5050 235 5100 265
rect 5050 215 5065 235
rect 5085 215 5100 235
rect 5050 185 5100 215
rect 5050 165 5065 185
rect 5085 165 5100 185
rect 5050 135 5100 165
rect 5050 115 5065 135
rect 5085 115 5100 135
rect 5050 85 5100 115
rect 5050 65 5065 85
rect 5085 65 5100 85
rect 5050 50 5100 65
rect 5350 735 5400 750
rect 5350 715 5365 735
rect 5385 715 5400 735
rect 5350 685 5400 715
rect 5350 665 5365 685
rect 5385 665 5400 685
rect 5350 635 5400 665
rect 5350 615 5365 635
rect 5385 615 5400 635
rect 5350 585 5400 615
rect 5350 565 5365 585
rect 5385 565 5400 585
rect 5350 535 5400 565
rect 5350 515 5365 535
rect 5385 515 5400 535
rect 5350 485 5400 515
rect 5350 465 5365 485
rect 5385 465 5400 485
rect 5350 435 5400 465
rect 5350 415 5365 435
rect 5385 415 5400 435
rect 5350 385 5400 415
rect 5350 365 5365 385
rect 5385 365 5400 385
rect 5350 335 5400 365
rect 5350 315 5365 335
rect 5385 315 5400 335
rect 5350 285 5400 315
rect 5350 265 5365 285
rect 5385 265 5400 285
rect 5350 235 5400 265
rect 5350 215 5365 235
rect 5385 215 5400 235
rect 5350 185 5400 215
rect 5350 165 5365 185
rect 5385 165 5400 185
rect 5350 135 5400 165
rect 5350 115 5365 135
rect 5385 115 5400 135
rect 5350 85 5400 115
rect 5350 65 5365 85
rect 5385 65 5400 85
rect 5350 50 5400 65
rect 5650 735 5700 750
rect 5650 715 5665 735
rect 5685 715 5700 735
rect 5650 685 5700 715
rect 5650 665 5665 685
rect 5685 665 5700 685
rect 5650 635 5700 665
rect 5650 615 5665 635
rect 5685 615 5700 635
rect 5650 585 5700 615
rect 5650 565 5665 585
rect 5685 565 5700 585
rect 5650 535 5700 565
rect 5650 515 5665 535
rect 5685 515 5700 535
rect 5650 485 5700 515
rect 5650 465 5665 485
rect 5685 465 5700 485
rect 5650 435 5700 465
rect 5650 415 5665 435
rect 5685 415 5700 435
rect 5650 385 5700 415
rect 5650 365 5665 385
rect 5685 365 5700 385
rect 5650 335 5700 365
rect 5650 315 5665 335
rect 5685 315 5700 335
rect 5650 285 5700 315
rect 5650 265 5665 285
rect 5685 265 5700 285
rect 5650 235 5700 265
rect 5650 215 5665 235
rect 5685 215 5700 235
rect 5650 185 5700 215
rect 5650 165 5665 185
rect 5685 165 5700 185
rect 5650 135 5700 165
rect 5650 115 5665 135
rect 5685 115 5700 135
rect 5650 85 5700 115
rect 5650 65 5665 85
rect 5685 65 5700 85
rect 5650 50 5700 65
rect 5950 735 6000 750
rect 5950 715 5965 735
rect 5985 715 6000 735
rect 5950 685 6000 715
rect 5950 665 5965 685
rect 5985 665 6000 685
rect 5950 635 6000 665
rect 5950 615 5965 635
rect 5985 615 6000 635
rect 5950 585 6000 615
rect 5950 565 5965 585
rect 5985 565 6000 585
rect 5950 535 6000 565
rect 5950 515 5965 535
rect 5985 515 6000 535
rect 5950 485 6000 515
rect 5950 465 5965 485
rect 5985 465 6000 485
rect 5950 435 6000 465
rect 5950 415 5965 435
rect 5985 415 6000 435
rect 5950 385 6000 415
rect 5950 365 5965 385
rect 5985 365 6000 385
rect 5950 335 6000 365
rect 5950 315 5965 335
rect 5985 315 6000 335
rect 5950 285 6000 315
rect 5950 265 5965 285
rect 5985 265 6000 285
rect 5950 235 6000 265
rect 5950 215 5965 235
rect 5985 215 6000 235
rect 5950 185 6000 215
rect 5950 165 5965 185
rect 5985 165 6000 185
rect 5950 135 6000 165
rect 5950 115 5965 135
rect 5985 115 6000 135
rect 5950 85 6000 115
rect 5950 65 5965 85
rect 5985 65 6000 85
rect 5950 50 6000 65
rect 6250 735 6300 750
rect 6250 715 6265 735
rect 6285 715 6300 735
rect 6250 685 6300 715
rect 6250 665 6265 685
rect 6285 665 6300 685
rect 6250 635 6300 665
rect 6250 615 6265 635
rect 6285 615 6300 635
rect 6250 585 6300 615
rect 6250 565 6265 585
rect 6285 565 6300 585
rect 6250 535 6300 565
rect 6250 515 6265 535
rect 6285 515 6300 535
rect 6250 485 6300 515
rect 6250 465 6265 485
rect 6285 465 6300 485
rect 6250 435 6300 465
rect 6250 415 6265 435
rect 6285 415 6300 435
rect 6250 385 6300 415
rect 6250 365 6265 385
rect 6285 365 6300 385
rect 6250 335 6300 365
rect 6250 315 6265 335
rect 6285 315 6300 335
rect 6250 285 6300 315
rect 6250 265 6265 285
rect 6285 265 6300 285
rect 6250 235 6300 265
rect 6250 215 6265 235
rect 6285 215 6300 235
rect 6250 185 6300 215
rect 6250 165 6265 185
rect 6285 165 6300 185
rect 6250 135 6300 165
rect 6250 115 6265 135
rect 6285 115 6300 135
rect 6250 85 6300 115
rect 6250 65 6265 85
rect 6285 65 6300 85
rect 6250 50 6300 65
rect 6550 735 6600 750
rect 6550 715 6565 735
rect 6585 715 6600 735
rect 6550 685 6600 715
rect 6550 665 6565 685
rect 6585 665 6600 685
rect 6550 635 6600 665
rect 6550 615 6565 635
rect 6585 615 6600 635
rect 6550 585 6600 615
rect 6550 565 6565 585
rect 6585 565 6600 585
rect 6550 535 6600 565
rect 6550 515 6565 535
rect 6585 515 6600 535
rect 6550 485 6600 515
rect 6550 465 6565 485
rect 6585 465 6600 485
rect 6550 435 6600 465
rect 6550 415 6565 435
rect 6585 415 6600 435
rect 6550 385 6600 415
rect 6550 365 6565 385
rect 6585 365 6600 385
rect 6550 335 6600 365
rect 6550 315 6565 335
rect 6585 315 6600 335
rect 6550 285 6600 315
rect 6550 265 6565 285
rect 6585 265 6600 285
rect 6550 235 6600 265
rect 6550 215 6565 235
rect 6585 215 6600 235
rect 6550 185 6600 215
rect 6550 165 6565 185
rect 6585 165 6600 185
rect 6550 135 6600 165
rect 6550 115 6565 135
rect 6585 115 6600 135
rect 6550 85 6600 115
rect 6550 65 6565 85
rect 6585 65 6600 85
rect 6550 50 6600 65
rect 6850 735 6900 750
rect 6850 715 6865 735
rect 6885 715 6900 735
rect 6850 685 6900 715
rect 6850 665 6865 685
rect 6885 665 6900 685
rect 6850 635 6900 665
rect 6850 615 6865 635
rect 6885 615 6900 635
rect 6850 585 6900 615
rect 6850 565 6865 585
rect 6885 565 6900 585
rect 6850 535 6900 565
rect 6850 515 6865 535
rect 6885 515 6900 535
rect 6850 485 6900 515
rect 6850 465 6865 485
rect 6885 465 6900 485
rect 6850 435 6900 465
rect 6850 415 6865 435
rect 6885 415 6900 435
rect 6850 385 6900 415
rect 6850 365 6865 385
rect 6885 365 6900 385
rect 6850 335 6900 365
rect 6850 315 6865 335
rect 6885 315 6900 335
rect 6850 285 6900 315
rect 6850 265 6865 285
rect 6885 265 6900 285
rect 6850 235 6900 265
rect 6850 215 6865 235
rect 6885 215 6900 235
rect 6850 185 6900 215
rect 6850 165 6865 185
rect 6885 165 6900 185
rect 6850 135 6900 165
rect 6850 115 6865 135
rect 6885 115 6900 135
rect 6850 85 6900 115
rect 6850 65 6865 85
rect 6885 65 6900 85
rect 6850 50 6900 65
rect 7150 735 7200 750
rect 7150 715 7165 735
rect 7185 715 7200 735
rect 7150 685 7200 715
rect 7150 665 7165 685
rect 7185 665 7200 685
rect 7150 635 7200 665
rect 7150 615 7165 635
rect 7185 615 7200 635
rect 7150 585 7200 615
rect 7150 565 7165 585
rect 7185 565 7200 585
rect 7150 535 7200 565
rect 7150 515 7165 535
rect 7185 515 7200 535
rect 7150 485 7200 515
rect 7150 465 7165 485
rect 7185 465 7200 485
rect 7150 435 7200 465
rect 7150 415 7165 435
rect 7185 415 7200 435
rect 7150 385 7200 415
rect 7150 365 7165 385
rect 7185 365 7200 385
rect 7150 335 7200 365
rect 7150 315 7165 335
rect 7185 315 7200 335
rect 7150 285 7200 315
rect 7150 265 7165 285
rect 7185 265 7200 285
rect 7150 235 7200 265
rect 7150 215 7165 235
rect 7185 215 7200 235
rect 7150 185 7200 215
rect 7150 165 7165 185
rect 7185 165 7200 185
rect 7150 135 7200 165
rect 7150 115 7165 135
rect 7185 115 7200 135
rect 7150 85 7200 115
rect 7150 65 7165 85
rect 7185 65 7200 85
rect 7150 50 7200 65
rect 8350 735 8400 750
rect 8350 715 8365 735
rect 8385 715 8400 735
rect 8350 685 8400 715
rect 8350 665 8365 685
rect 8385 665 8400 685
rect 8350 635 8400 665
rect 8350 615 8365 635
rect 8385 615 8400 635
rect 8350 585 8400 615
rect 8350 565 8365 585
rect 8385 565 8400 585
rect 8350 535 8400 565
rect 8350 515 8365 535
rect 8385 515 8400 535
rect 8350 485 8400 515
rect 8350 465 8365 485
rect 8385 465 8400 485
rect 8350 435 8400 465
rect 8350 415 8365 435
rect 8385 415 8400 435
rect 8350 385 8400 415
rect 8350 365 8365 385
rect 8385 365 8400 385
rect 8350 335 8400 365
rect 8350 315 8365 335
rect 8385 315 8400 335
rect 8350 285 8400 315
rect 8350 265 8365 285
rect 8385 265 8400 285
rect 8350 235 8400 265
rect 8350 215 8365 235
rect 8385 215 8400 235
rect 8350 185 8400 215
rect 8350 165 8365 185
rect 8385 165 8400 185
rect 8350 135 8400 165
rect 8350 115 8365 135
rect 8385 115 8400 135
rect 8350 85 8400 115
rect 8350 65 8365 85
rect 8385 65 8400 85
rect 8350 50 8400 65
rect 9550 735 9600 750
rect 9550 715 9565 735
rect 9585 715 9600 735
rect 9550 685 9600 715
rect 9550 665 9565 685
rect 9585 665 9600 685
rect 9550 635 9600 665
rect 9550 615 9565 635
rect 9585 615 9600 635
rect 9550 585 9600 615
rect 9550 565 9565 585
rect 9585 565 9600 585
rect 9550 535 9600 565
rect 9550 515 9565 535
rect 9585 515 9600 535
rect 9550 485 9600 515
rect 9550 465 9565 485
rect 9585 465 9600 485
rect 9550 435 9600 465
rect 9550 415 9565 435
rect 9585 415 9600 435
rect 9550 385 9600 415
rect 9550 365 9565 385
rect 9585 365 9600 385
rect 9550 335 9600 365
rect 9550 315 9565 335
rect 9585 315 9600 335
rect 9550 285 9600 315
rect 9550 265 9565 285
rect 9585 265 9600 285
rect 9550 235 9600 265
rect 9550 215 9565 235
rect 9585 215 9600 235
rect 9550 185 9600 215
rect 9550 165 9565 185
rect 9585 165 9600 185
rect 9550 135 9600 165
rect 9550 115 9565 135
rect 9585 115 9600 135
rect 9550 85 9600 115
rect 9550 65 9565 85
rect 9585 65 9600 85
rect 9550 50 9600 65
rect 10750 735 10800 750
rect 10750 715 10765 735
rect 10785 715 10800 735
rect 10750 685 10800 715
rect 10750 665 10765 685
rect 10785 665 10800 685
rect 10750 635 10800 665
rect 10750 615 10765 635
rect 10785 615 10800 635
rect 10750 585 10800 615
rect 10750 565 10765 585
rect 10785 565 10800 585
rect 10750 535 10800 565
rect 10750 515 10765 535
rect 10785 515 10800 535
rect 10750 485 10800 515
rect 10750 465 10765 485
rect 10785 465 10800 485
rect 10750 435 10800 465
rect 10750 415 10765 435
rect 10785 415 10800 435
rect 10750 385 10800 415
rect 10750 365 10765 385
rect 10785 365 10800 385
rect 10750 335 10800 365
rect 10750 315 10765 335
rect 10785 315 10800 335
rect 10750 285 10800 315
rect 10750 265 10765 285
rect 10785 265 10800 285
rect 10750 235 10800 265
rect 10750 215 10765 235
rect 10785 215 10800 235
rect 10750 185 10800 215
rect 10750 165 10765 185
rect 10785 165 10800 185
rect 10750 135 10800 165
rect 10750 115 10765 135
rect 10785 115 10800 135
rect 10750 85 10800 115
rect 10750 65 10765 85
rect 10785 65 10800 85
rect 10750 50 10800 65
rect 11950 735 12000 750
rect 11950 715 11965 735
rect 11985 715 12000 735
rect 11950 685 12000 715
rect 11950 665 11965 685
rect 11985 665 12000 685
rect 11950 635 12000 665
rect 11950 615 11965 635
rect 11985 615 12000 635
rect 11950 585 12000 615
rect 11950 565 11965 585
rect 11985 565 12000 585
rect 11950 535 12000 565
rect 11950 515 11965 535
rect 11985 515 12000 535
rect 11950 485 12000 515
rect 11950 465 11965 485
rect 11985 465 12000 485
rect 11950 435 12000 465
rect 11950 415 11965 435
rect 11985 415 12000 435
rect 11950 385 12000 415
rect 11950 365 11965 385
rect 11985 365 12000 385
rect 11950 335 12000 365
rect 11950 315 11965 335
rect 11985 315 12000 335
rect 11950 285 12000 315
rect 11950 265 11965 285
rect 11985 265 12000 285
rect 11950 235 12000 265
rect 11950 215 11965 235
rect 11985 215 12000 235
rect 11950 185 12000 215
rect 11950 165 11965 185
rect 11985 165 12000 185
rect 11950 135 12000 165
rect 11950 115 11965 135
rect 11985 115 12000 135
rect 11950 85 12000 115
rect 11950 65 11965 85
rect 11985 65 12000 85
rect 11950 50 12000 65
rect 12250 735 12300 750
rect 12250 715 12265 735
rect 12285 715 12300 735
rect 12250 685 12300 715
rect 12250 665 12265 685
rect 12285 665 12300 685
rect 12250 635 12300 665
rect 12250 615 12265 635
rect 12285 615 12300 635
rect 12250 585 12300 615
rect 12250 565 12265 585
rect 12285 565 12300 585
rect 12250 535 12300 565
rect 12250 515 12265 535
rect 12285 515 12300 535
rect 12250 485 12300 515
rect 12250 465 12265 485
rect 12285 465 12300 485
rect 12250 435 12300 465
rect 12250 415 12265 435
rect 12285 415 12300 435
rect 12250 385 12300 415
rect 12250 365 12265 385
rect 12285 365 12300 385
rect 12250 335 12300 365
rect 12250 315 12265 335
rect 12285 315 12300 335
rect 12250 285 12300 315
rect 12250 265 12265 285
rect 12285 265 12300 285
rect 12250 235 12300 265
rect 12250 215 12265 235
rect 12285 215 12300 235
rect 12250 185 12300 215
rect 12250 165 12265 185
rect 12285 165 12300 185
rect 12250 135 12300 165
rect 12250 115 12265 135
rect 12285 115 12300 135
rect 12250 85 12300 115
rect 12250 65 12265 85
rect 12285 65 12300 85
rect 12250 50 12300 65
rect 12550 735 12600 750
rect 12550 715 12565 735
rect 12585 715 12600 735
rect 12550 685 12600 715
rect 12550 665 12565 685
rect 12585 665 12600 685
rect 12550 635 12600 665
rect 12550 615 12565 635
rect 12585 615 12600 635
rect 12550 585 12600 615
rect 12550 565 12565 585
rect 12585 565 12600 585
rect 12550 535 12600 565
rect 12550 515 12565 535
rect 12585 515 12600 535
rect 12550 485 12600 515
rect 12550 465 12565 485
rect 12585 465 12600 485
rect 12550 435 12600 465
rect 12550 415 12565 435
rect 12585 415 12600 435
rect 12550 385 12600 415
rect 12550 365 12565 385
rect 12585 365 12600 385
rect 12550 335 12600 365
rect 12550 315 12565 335
rect 12585 315 12600 335
rect 12550 285 12600 315
rect 12550 265 12565 285
rect 12585 265 12600 285
rect 12550 235 12600 265
rect 12550 215 12565 235
rect 12585 215 12600 235
rect 12550 185 12600 215
rect 12550 165 12565 185
rect 12585 165 12600 185
rect 12550 135 12600 165
rect 12550 115 12565 135
rect 12585 115 12600 135
rect 12550 85 12600 115
rect 12550 65 12565 85
rect 12585 65 12600 85
rect 12550 50 12600 65
rect 12850 735 12900 750
rect 12850 715 12865 735
rect 12885 715 12900 735
rect 12850 685 12900 715
rect 12850 665 12865 685
rect 12885 665 12900 685
rect 12850 635 12900 665
rect 12850 615 12865 635
rect 12885 615 12900 635
rect 12850 585 12900 615
rect 12850 565 12865 585
rect 12885 565 12900 585
rect 12850 535 12900 565
rect 12850 515 12865 535
rect 12885 515 12900 535
rect 12850 485 12900 515
rect 12850 465 12865 485
rect 12885 465 12900 485
rect 12850 435 12900 465
rect 12850 415 12865 435
rect 12885 415 12900 435
rect 12850 385 12900 415
rect 12850 365 12865 385
rect 12885 365 12900 385
rect 12850 335 12900 365
rect 12850 315 12865 335
rect 12885 315 12900 335
rect 12850 285 12900 315
rect 12850 265 12865 285
rect 12885 265 12900 285
rect 12850 235 12900 265
rect 12850 215 12865 235
rect 12885 215 12900 235
rect 12850 185 12900 215
rect 12850 165 12865 185
rect 12885 165 12900 185
rect 12850 135 12900 165
rect 12850 115 12865 135
rect 12885 115 12900 135
rect 12850 85 12900 115
rect 12850 65 12865 85
rect 12885 65 12900 85
rect 12850 50 12900 65
rect 13150 735 13200 750
rect 13150 715 13165 735
rect 13185 715 13200 735
rect 13150 685 13200 715
rect 13150 665 13165 685
rect 13185 665 13200 685
rect 13150 635 13200 665
rect 13150 615 13165 635
rect 13185 615 13200 635
rect 13150 585 13200 615
rect 13150 565 13165 585
rect 13185 565 13200 585
rect 13150 535 13200 565
rect 13150 515 13165 535
rect 13185 515 13200 535
rect 13150 485 13200 515
rect 13150 465 13165 485
rect 13185 465 13200 485
rect 13150 435 13200 465
rect 13150 415 13165 435
rect 13185 415 13200 435
rect 13150 385 13200 415
rect 13150 365 13165 385
rect 13185 365 13200 385
rect 13150 335 13200 365
rect 13150 315 13165 335
rect 13185 315 13200 335
rect 13150 285 13200 315
rect 13150 265 13165 285
rect 13185 265 13200 285
rect 13150 235 13200 265
rect 13150 215 13165 235
rect 13185 215 13200 235
rect 13150 185 13200 215
rect 13150 165 13165 185
rect 13185 165 13200 185
rect 13150 135 13200 165
rect 13150 115 13165 135
rect 13185 115 13200 135
rect 13150 85 13200 115
rect 13150 65 13165 85
rect 13185 65 13200 85
rect 13150 50 13200 65
rect 13450 735 13500 750
rect 13450 715 13465 735
rect 13485 715 13500 735
rect 13450 685 13500 715
rect 13450 665 13465 685
rect 13485 665 13500 685
rect 13450 635 13500 665
rect 13450 615 13465 635
rect 13485 615 13500 635
rect 13450 585 13500 615
rect 13450 565 13465 585
rect 13485 565 13500 585
rect 13450 535 13500 565
rect 13450 515 13465 535
rect 13485 515 13500 535
rect 13450 485 13500 515
rect 13450 465 13465 485
rect 13485 465 13500 485
rect 13450 435 13500 465
rect 13450 415 13465 435
rect 13485 415 13500 435
rect 13450 385 13500 415
rect 13450 365 13465 385
rect 13485 365 13500 385
rect 13450 335 13500 365
rect 13450 315 13465 335
rect 13485 315 13500 335
rect 13450 285 13500 315
rect 13450 265 13465 285
rect 13485 265 13500 285
rect 13450 235 13500 265
rect 13450 215 13465 235
rect 13485 215 13500 235
rect 13450 185 13500 215
rect 13450 165 13465 185
rect 13485 165 13500 185
rect 13450 135 13500 165
rect 13450 115 13465 135
rect 13485 115 13500 135
rect 13450 85 13500 115
rect 13450 65 13465 85
rect 13485 65 13500 85
rect 13450 50 13500 65
rect 13750 735 13800 750
rect 13750 715 13765 735
rect 13785 715 13800 735
rect 13750 685 13800 715
rect 13750 665 13765 685
rect 13785 665 13800 685
rect 13750 635 13800 665
rect 13750 615 13765 635
rect 13785 615 13800 635
rect 13750 585 13800 615
rect 13750 565 13765 585
rect 13785 565 13800 585
rect 13750 535 13800 565
rect 13750 515 13765 535
rect 13785 515 13800 535
rect 13750 485 13800 515
rect 13750 465 13765 485
rect 13785 465 13800 485
rect 13750 435 13800 465
rect 13750 415 13765 435
rect 13785 415 13800 435
rect 13750 385 13800 415
rect 13750 365 13765 385
rect 13785 365 13800 385
rect 13750 335 13800 365
rect 13750 315 13765 335
rect 13785 315 13800 335
rect 13750 285 13800 315
rect 13750 265 13765 285
rect 13785 265 13800 285
rect 13750 235 13800 265
rect 13750 215 13765 235
rect 13785 215 13800 235
rect 13750 185 13800 215
rect 13750 165 13765 185
rect 13785 165 13800 185
rect 13750 135 13800 165
rect 13750 115 13765 135
rect 13785 115 13800 135
rect 13750 85 13800 115
rect 13750 65 13765 85
rect 13785 65 13800 85
rect 13750 50 13800 65
rect 14050 735 14100 750
rect 14050 715 14065 735
rect 14085 715 14100 735
rect 14050 685 14100 715
rect 14050 665 14065 685
rect 14085 665 14100 685
rect 14050 635 14100 665
rect 14050 615 14065 635
rect 14085 615 14100 635
rect 14050 585 14100 615
rect 14050 565 14065 585
rect 14085 565 14100 585
rect 14050 535 14100 565
rect 14050 515 14065 535
rect 14085 515 14100 535
rect 14050 485 14100 515
rect 14050 465 14065 485
rect 14085 465 14100 485
rect 14050 435 14100 465
rect 14050 415 14065 435
rect 14085 415 14100 435
rect 14050 385 14100 415
rect 14050 365 14065 385
rect 14085 365 14100 385
rect 14050 335 14100 365
rect 14050 315 14065 335
rect 14085 315 14100 335
rect 14050 285 14100 315
rect 14050 265 14065 285
rect 14085 265 14100 285
rect 14050 235 14100 265
rect 14050 215 14065 235
rect 14085 215 14100 235
rect 14050 185 14100 215
rect 14050 165 14065 185
rect 14085 165 14100 185
rect 14050 135 14100 165
rect 14050 115 14065 135
rect 14085 115 14100 135
rect 14050 85 14100 115
rect 14050 65 14065 85
rect 14085 65 14100 85
rect 14050 50 14100 65
rect 14350 735 14400 750
rect 14350 715 14365 735
rect 14385 715 14400 735
rect 14350 685 14400 715
rect 14350 665 14365 685
rect 14385 665 14400 685
rect 14350 635 14400 665
rect 14350 615 14365 635
rect 14385 615 14400 635
rect 14350 585 14400 615
rect 14350 565 14365 585
rect 14385 565 14400 585
rect 14350 535 14400 565
rect 14350 515 14365 535
rect 14385 515 14400 535
rect 14350 485 14400 515
rect 14350 465 14365 485
rect 14385 465 14400 485
rect 14350 435 14400 465
rect 14350 415 14365 435
rect 14385 415 14400 435
rect 14350 385 14400 415
rect 14350 365 14365 385
rect 14385 365 14400 385
rect 14350 335 14400 365
rect 14350 315 14365 335
rect 14385 315 14400 335
rect 14350 285 14400 315
rect 14350 265 14365 285
rect 14385 265 14400 285
rect 14350 235 14400 265
rect 14350 215 14365 235
rect 14385 215 14400 235
rect 14350 185 14400 215
rect 14350 165 14365 185
rect 14385 165 14400 185
rect 14350 135 14400 165
rect 14350 115 14365 135
rect 14385 115 14400 135
rect 14350 85 14400 115
rect 14350 65 14365 85
rect 14385 65 14400 85
rect 14350 50 14400 65
rect 15550 735 15600 750
rect 15550 715 15565 735
rect 15585 715 15600 735
rect 15550 685 15600 715
rect 15550 665 15565 685
rect 15585 665 15600 685
rect 15550 635 15600 665
rect 15550 615 15565 635
rect 15585 615 15600 635
rect 15550 585 15600 615
rect 15550 565 15565 585
rect 15585 565 15600 585
rect 15550 535 15600 565
rect 15550 515 15565 535
rect 15585 515 15600 535
rect 15550 485 15600 515
rect 15550 465 15565 485
rect 15585 465 15600 485
rect 15550 435 15600 465
rect 15550 415 15565 435
rect 15585 415 15600 435
rect 15550 385 15600 415
rect 15550 365 15565 385
rect 15585 365 15600 385
rect 15550 335 15600 365
rect 15550 315 15565 335
rect 15585 315 15600 335
rect 15550 285 15600 315
rect 15550 265 15565 285
rect 15585 265 15600 285
rect 15550 235 15600 265
rect 15550 215 15565 235
rect 15585 215 15600 235
rect 15550 185 15600 215
rect 15550 165 15565 185
rect 15585 165 15600 185
rect 15550 135 15600 165
rect 15550 115 15565 135
rect 15585 115 15600 135
rect 15550 85 15600 115
rect 15550 65 15565 85
rect 15585 65 15600 85
rect 15550 50 15600 65
rect 16750 735 16800 750
rect 16750 715 16765 735
rect 16785 715 16800 735
rect 16750 685 16800 715
rect 16750 665 16765 685
rect 16785 665 16800 685
rect 16750 635 16800 665
rect 16750 615 16765 635
rect 16785 615 16800 635
rect 16750 585 16800 615
rect 16750 565 16765 585
rect 16785 565 16800 585
rect 16750 535 16800 565
rect 16750 515 16765 535
rect 16785 515 16800 535
rect 16750 485 16800 515
rect 16750 465 16765 485
rect 16785 465 16800 485
rect 16750 435 16800 465
rect 16750 415 16765 435
rect 16785 415 16800 435
rect 16750 385 16800 415
rect 16750 365 16765 385
rect 16785 365 16800 385
rect 16750 335 16800 365
rect 16750 315 16765 335
rect 16785 315 16800 335
rect 16750 285 16800 315
rect 16750 265 16765 285
rect 16785 265 16800 285
rect 16750 235 16800 265
rect 16750 215 16765 235
rect 16785 215 16800 235
rect 16750 185 16800 215
rect 16750 165 16765 185
rect 16785 165 16800 185
rect 16750 135 16800 165
rect 16750 115 16765 135
rect 16785 115 16800 135
rect 16750 85 16800 115
rect 16750 65 16765 85
rect 16785 65 16800 85
rect 16750 50 16800 65
rect 17950 735 18000 750
rect 17950 715 17965 735
rect 17985 715 18000 735
rect 17950 685 18000 715
rect 17950 665 17965 685
rect 17985 665 18000 685
rect 17950 635 18000 665
rect 17950 615 17965 635
rect 17985 615 18000 635
rect 17950 585 18000 615
rect 17950 565 17965 585
rect 17985 565 18000 585
rect 17950 535 18000 565
rect 17950 515 17965 535
rect 17985 515 18000 535
rect 17950 485 18000 515
rect 17950 465 17965 485
rect 17985 465 18000 485
rect 17950 435 18000 465
rect 17950 415 17965 435
rect 17985 415 18000 435
rect 17950 385 18000 415
rect 17950 365 17965 385
rect 17985 365 18000 385
rect 17950 335 18000 365
rect 17950 315 17965 335
rect 17985 315 18000 335
rect 17950 285 18000 315
rect 17950 265 17965 285
rect 17985 265 18000 285
rect 17950 235 18000 265
rect 17950 215 17965 235
rect 17985 215 18000 235
rect 17950 185 18000 215
rect 17950 165 17965 185
rect 17985 165 18000 185
rect 17950 135 18000 165
rect 17950 115 17965 135
rect 17985 115 18000 135
rect 17950 85 18000 115
rect 17950 65 17965 85
rect 17985 65 18000 85
rect 17950 50 18000 65
rect 19150 735 19200 750
rect 19150 715 19165 735
rect 19185 715 19200 735
rect 19150 685 19200 715
rect 19150 665 19165 685
rect 19185 665 19200 685
rect 19150 635 19200 665
rect 19150 615 19165 635
rect 19185 615 19200 635
rect 19150 585 19200 615
rect 19150 565 19165 585
rect 19185 565 19200 585
rect 19150 535 19200 565
rect 19150 515 19165 535
rect 19185 515 19200 535
rect 19150 485 19200 515
rect 19150 465 19165 485
rect 19185 465 19200 485
rect 19150 435 19200 465
rect 19150 415 19165 435
rect 19185 415 19200 435
rect 19150 385 19200 415
rect 19150 365 19165 385
rect 19185 365 19200 385
rect 19150 335 19200 365
rect 19150 315 19165 335
rect 19185 315 19200 335
rect 19150 285 19200 315
rect 19150 265 19165 285
rect 19185 265 19200 285
rect 19150 235 19200 265
rect 19150 215 19165 235
rect 19185 215 19200 235
rect 19150 185 19200 215
rect 19150 165 19165 185
rect 19185 165 19200 185
rect 19150 135 19200 165
rect 19150 115 19165 135
rect 19185 115 19200 135
rect 19150 85 19200 115
rect 19150 65 19165 85
rect 19185 65 19200 85
rect 19150 50 19200 65
rect 20350 735 20400 750
rect 20350 715 20365 735
rect 20385 715 20400 735
rect 20350 685 20400 715
rect 20350 665 20365 685
rect 20385 665 20400 685
rect 20350 635 20400 665
rect 20350 615 20365 635
rect 20385 615 20400 635
rect 20350 585 20400 615
rect 20350 565 20365 585
rect 20385 565 20400 585
rect 20350 535 20400 565
rect 20350 515 20365 535
rect 20385 515 20400 535
rect 20350 485 20400 515
rect 20350 465 20365 485
rect 20385 465 20400 485
rect 20350 435 20400 465
rect 20350 415 20365 435
rect 20385 415 20400 435
rect 20350 385 20400 415
rect 20350 365 20365 385
rect 20385 365 20400 385
rect 20350 335 20400 365
rect 20350 315 20365 335
rect 20385 315 20400 335
rect 20350 285 20400 315
rect 20350 265 20365 285
rect 20385 265 20400 285
rect 20350 235 20400 265
rect 20350 215 20365 235
rect 20385 215 20400 235
rect 20350 185 20400 215
rect 20350 165 20365 185
rect 20385 165 20400 185
rect 20350 135 20400 165
rect 20350 115 20365 135
rect 20385 115 20400 135
rect 20350 85 20400 115
rect 20350 65 20365 85
rect 20385 65 20400 85
rect 20350 50 20400 65
rect -650 -15 20400 0
rect -650 -35 -635 -15
rect -615 -35 -585 -15
rect -565 -35 -535 -15
rect -515 -35 -485 -15
rect -465 -35 -435 -15
rect -415 -35 -385 -15
rect -365 -35 -335 -15
rect -315 -35 -285 -15
rect -265 -35 -235 -15
rect -215 -35 -185 -15
rect -165 -35 -135 -15
rect -115 -35 -85 -15
rect -65 -35 -35 -15
rect -15 -35 15 -15
rect 35 -35 65 -15
rect 85 -35 115 -15
rect 135 -35 165 -15
rect 185 -35 215 -15
rect 235 -35 265 -15
rect 285 -35 315 -15
rect 335 -35 365 -15
rect 385 -35 415 -15
rect 435 -35 465 -15
rect 485 -35 515 -15
rect 535 -35 565 -15
rect 585 -35 615 -15
rect 635 -35 665 -15
rect 685 -35 715 -15
rect 735 -35 765 -15
rect 785 -35 815 -15
rect 835 -35 865 -15
rect 885 -35 915 -15
rect 935 -35 965 -15
rect 985 -35 1015 -15
rect 1035 -35 1065 -15
rect 1085 -35 1115 -15
rect 1135 -35 1165 -15
rect 1185 -35 1215 -15
rect 1235 -35 1265 -15
rect 1285 -35 1315 -15
rect 1335 -35 1365 -15
rect 1385 -35 1415 -15
rect 1435 -35 1465 -15
rect 1485 -35 1515 -15
rect 1535 -35 1565 -15
rect 1585 -35 1615 -15
rect 1635 -35 1665 -15
rect 1685 -35 1715 -15
rect 1735 -35 1765 -15
rect 1785 -35 1815 -15
rect 1835 -35 1865 -15
rect 1885 -35 1915 -15
rect 1935 -35 1965 -15
rect 1985 -35 2015 -15
rect 2035 -35 2065 -15
rect 2085 -35 2115 -15
rect 2135 -35 2165 -15
rect 2185 -35 2215 -15
rect 2235 -35 2265 -15
rect 2285 -35 2315 -15
rect 2335 -35 2365 -15
rect 2385 -35 2415 -15
rect 2435 -35 2465 -15
rect 2485 -35 2515 -15
rect 2535 -35 2565 -15
rect 2585 -35 2615 -15
rect 2635 -35 2665 -15
rect 2685 -35 2715 -15
rect 2735 -35 2765 -15
rect 2785 -35 2815 -15
rect 2835 -35 2865 -15
rect 2885 -35 2915 -15
rect 2935 -35 2965 -15
rect 2985 -35 3015 -15
rect 3035 -35 3065 -15
rect 3085 -35 3115 -15
rect 3135 -35 3165 -15
rect 3185 -35 3215 -15
rect 3235 -35 3265 -15
rect 3285 -35 3315 -15
rect 3335 -35 3365 -15
rect 3385 -35 3415 -15
rect 3435 -35 3465 -15
rect 3485 -35 3515 -15
rect 3535 -35 3565 -15
rect 3585 -35 3615 -15
rect 3635 -35 3665 -15
rect 3685 -35 3715 -15
rect 3735 -35 3765 -15
rect 3785 -35 3815 -15
rect 3835 -35 3865 -15
rect 3885 -35 3915 -15
rect 3935 -35 3965 -15
rect 3985 -35 4015 -15
rect 4035 -35 4065 -15
rect 4085 -35 4115 -15
rect 4135 -35 4165 -15
rect 4185 -35 4215 -15
rect 4235 -35 4265 -15
rect 4285 -35 4315 -15
rect 4335 -35 4365 -15
rect 4385 -35 4415 -15
rect 4435 -35 4465 -15
rect 4485 -35 4515 -15
rect 4535 -35 4565 -15
rect 4585 -35 4615 -15
rect 4635 -35 4665 -15
rect 4685 -35 4715 -15
rect 4735 -35 4765 -15
rect 4785 -35 4815 -15
rect 4835 -35 4865 -15
rect 4885 -35 4915 -15
rect 4935 -35 4965 -15
rect 4985 -35 5015 -15
rect 5035 -35 5065 -15
rect 5085 -35 5115 -15
rect 5135 -35 5165 -15
rect 5185 -35 5215 -15
rect 5235 -35 5265 -15
rect 5285 -35 5315 -15
rect 5335 -35 5365 -15
rect 5385 -35 5415 -15
rect 5435 -35 5465 -15
rect 5485 -35 5515 -15
rect 5535 -35 5565 -15
rect 5585 -35 5615 -15
rect 5635 -35 5665 -15
rect 5685 -35 5715 -15
rect 5735 -35 5765 -15
rect 5785 -35 5815 -15
rect 5835 -35 5865 -15
rect 5885 -35 5915 -15
rect 5935 -35 5965 -15
rect 5985 -35 6015 -15
rect 6035 -35 6065 -15
rect 6085 -35 6115 -15
rect 6135 -35 6165 -15
rect 6185 -35 6215 -15
rect 6235 -35 6265 -15
rect 6285 -35 6315 -15
rect 6335 -35 6365 -15
rect 6385 -35 6415 -15
rect 6435 -35 6465 -15
rect 6485 -35 6515 -15
rect 6535 -35 6565 -15
rect 6585 -35 6615 -15
rect 6635 -35 6665 -15
rect 6685 -35 6715 -15
rect 6735 -35 6765 -15
rect 6785 -35 6815 -15
rect 6835 -35 6865 -15
rect 6885 -35 6915 -15
rect 6935 -35 6965 -15
rect 6985 -35 7015 -15
rect 7035 -35 7065 -15
rect 7085 -35 7115 -15
rect 7135 -35 7165 -15
rect 7185 -35 7215 -15
rect 7235 -35 7265 -15
rect 7285 -35 7315 -15
rect 7335 -35 7365 -15
rect 7385 -35 7415 -15
rect 7435 -35 7465 -15
rect 7485 -35 7515 -15
rect 7535 -35 7565 -15
rect 7585 -35 7615 -15
rect 7635 -35 7665 -15
rect 7685 -35 7715 -15
rect 7735 -35 7765 -15
rect 7785 -35 7815 -15
rect 7835 -35 7865 -15
rect 7885 -35 7915 -15
rect 7935 -35 7965 -15
rect 7985 -35 8015 -15
rect 8035 -35 8065 -15
rect 8085 -35 8115 -15
rect 8135 -35 8165 -15
rect 8185 -35 8215 -15
rect 8235 -35 8265 -15
rect 8285 -35 8315 -15
rect 8335 -35 8365 -15
rect 8385 -35 8415 -15
rect 8435 -35 8465 -15
rect 8485 -35 8515 -15
rect 8535 -35 8565 -15
rect 8585 -35 8615 -15
rect 8635 -35 8665 -15
rect 8685 -35 8715 -15
rect 8735 -35 8765 -15
rect 8785 -35 8815 -15
rect 8835 -35 8865 -15
rect 8885 -35 8915 -15
rect 8935 -35 8965 -15
rect 8985 -35 9015 -15
rect 9035 -35 9065 -15
rect 9085 -35 9115 -15
rect 9135 -35 9165 -15
rect 9185 -35 9215 -15
rect 9235 -35 9265 -15
rect 9285 -35 9315 -15
rect 9335 -35 9365 -15
rect 9385 -35 9415 -15
rect 9435 -35 9465 -15
rect 9485 -35 9515 -15
rect 9535 -35 9565 -15
rect 9585 -35 9615 -15
rect 9635 -35 9665 -15
rect 9685 -35 9715 -15
rect 9735 -35 9765 -15
rect 9785 -35 9815 -15
rect 9835 -35 9865 -15
rect 9885 -35 9915 -15
rect 9935 -35 9965 -15
rect 9985 -35 10015 -15
rect 10035 -35 10065 -15
rect 10085 -35 10115 -15
rect 10135 -35 10165 -15
rect 10185 -35 10215 -15
rect 10235 -35 10265 -15
rect 10285 -35 10315 -15
rect 10335 -35 10365 -15
rect 10385 -35 10415 -15
rect 10435 -35 10465 -15
rect 10485 -35 10515 -15
rect 10535 -35 10565 -15
rect 10585 -35 10615 -15
rect 10635 -35 10665 -15
rect 10685 -35 10715 -15
rect 10735 -35 10765 -15
rect 10785 -35 10815 -15
rect 10835 -35 10865 -15
rect 10885 -35 10915 -15
rect 10935 -35 10965 -15
rect 10985 -35 11015 -15
rect 11035 -35 11065 -15
rect 11085 -35 11115 -15
rect 11135 -35 11165 -15
rect 11185 -35 11215 -15
rect 11235 -35 11265 -15
rect 11285 -35 11315 -15
rect 11335 -35 11365 -15
rect 11385 -35 11415 -15
rect 11435 -35 11465 -15
rect 11485 -35 11515 -15
rect 11535 -35 11565 -15
rect 11585 -35 11615 -15
rect 11635 -35 11665 -15
rect 11685 -35 11715 -15
rect 11735 -35 11765 -15
rect 11785 -35 11815 -15
rect 11835 -35 11865 -15
rect 11885 -35 11915 -15
rect 11935 -35 11965 -15
rect 11985 -35 12015 -15
rect 12035 -35 12065 -15
rect 12085 -35 12115 -15
rect 12135 -35 12165 -15
rect 12185 -35 12215 -15
rect 12235 -35 12265 -15
rect 12285 -35 12315 -15
rect 12335 -35 12365 -15
rect 12385 -35 12415 -15
rect 12435 -35 12465 -15
rect 12485 -35 12515 -15
rect 12535 -35 12565 -15
rect 12585 -35 12615 -15
rect 12635 -35 12665 -15
rect 12685 -35 12715 -15
rect 12735 -35 12765 -15
rect 12785 -35 12815 -15
rect 12835 -35 12865 -15
rect 12885 -35 12915 -15
rect 12935 -35 12965 -15
rect 12985 -35 13015 -15
rect 13035 -35 13065 -15
rect 13085 -35 13115 -15
rect 13135 -35 13165 -15
rect 13185 -35 13215 -15
rect 13235 -35 13265 -15
rect 13285 -35 13315 -15
rect 13335 -35 13365 -15
rect 13385 -35 13415 -15
rect 13435 -35 13465 -15
rect 13485 -35 13515 -15
rect 13535 -35 13565 -15
rect 13585 -35 13615 -15
rect 13635 -35 13665 -15
rect 13685 -35 13715 -15
rect 13735 -35 13765 -15
rect 13785 -35 13815 -15
rect 13835 -35 13865 -15
rect 13885 -35 13915 -15
rect 13935 -35 13965 -15
rect 13985 -35 14015 -15
rect 14035 -35 14065 -15
rect 14085 -35 14115 -15
rect 14135 -35 14165 -15
rect 14185 -35 14215 -15
rect 14235 -35 14265 -15
rect 14285 -35 14315 -15
rect 14335 -35 14365 -15
rect 14385 -35 14415 -15
rect 14435 -35 14465 -15
rect 14485 -35 14515 -15
rect 14535 -35 14565 -15
rect 14585 -35 14615 -15
rect 14635 -35 14665 -15
rect 14685 -35 14715 -15
rect 14735 -35 14765 -15
rect 14785 -35 14815 -15
rect 14835 -35 14865 -15
rect 14885 -35 14915 -15
rect 14935 -35 14965 -15
rect 14985 -35 15015 -15
rect 15035 -35 15065 -15
rect 15085 -35 15115 -15
rect 15135 -35 15165 -15
rect 15185 -35 15215 -15
rect 15235 -35 15265 -15
rect 15285 -35 15315 -15
rect 15335 -35 15365 -15
rect 15385 -35 15415 -15
rect 15435 -35 15465 -15
rect 15485 -35 15515 -15
rect 15535 -35 15565 -15
rect 15585 -35 15615 -15
rect 15635 -35 15665 -15
rect 15685 -35 15715 -15
rect 15735 -35 15765 -15
rect 15785 -35 15815 -15
rect 15835 -35 15865 -15
rect 15885 -35 15915 -15
rect 15935 -35 15965 -15
rect 15985 -35 16015 -15
rect 16035 -35 16065 -15
rect 16085 -35 16115 -15
rect 16135 -35 16165 -15
rect 16185 -35 16215 -15
rect 16235 -35 16265 -15
rect 16285 -35 16315 -15
rect 16335 -35 16365 -15
rect 16385 -35 16415 -15
rect 16435 -35 16465 -15
rect 16485 -35 16515 -15
rect 16535 -35 16565 -15
rect 16585 -35 16615 -15
rect 16635 -35 16665 -15
rect 16685 -35 16715 -15
rect 16735 -35 16765 -15
rect 16785 -35 16815 -15
rect 16835 -35 16865 -15
rect 16885 -35 16915 -15
rect 16935 -35 16965 -15
rect 16985 -35 17015 -15
rect 17035 -35 17065 -15
rect 17085 -35 17115 -15
rect 17135 -35 17165 -15
rect 17185 -35 17215 -15
rect 17235 -35 17265 -15
rect 17285 -35 17315 -15
rect 17335 -35 17365 -15
rect 17385 -35 17415 -15
rect 17435 -35 17465 -15
rect 17485 -35 17515 -15
rect 17535 -35 17565 -15
rect 17585 -35 17615 -15
rect 17635 -35 17665 -15
rect 17685 -35 17715 -15
rect 17735 -35 17765 -15
rect 17785 -35 17815 -15
rect 17835 -35 17865 -15
rect 17885 -35 17915 -15
rect 17935 -35 17965 -15
rect 17985 -35 18015 -15
rect 18035 -35 18065 -15
rect 18085 -35 18115 -15
rect 18135 -35 18165 -15
rect 18185 -35 18215 -15
rect 18235 -35 18265 -15
rect 18285 -35 18315 -15
rect 18335 -35 18365 -15
rect 18385 -35 18415 -15
rect 18435 -35 18465 -15
rect 18485 -35 18515 -15
rect 18535 -35 18565 -15
rect 18585 -35 18615 -15
rect 18635 -35 18665 -15
rect 18685 -35 18715 -15
rect 18735 -35 18765 -15
rect 18785 -35 18815 -15
rect 18835 -35 18865 -15
rect 18885 -35 18915 -15
rect 18935 -35 18965 -15
rect 18985 -35 19015 -15
rect 19035 -35 19065 -15
rect 19085 -35 19115 -15
rect 19135 -35 19165 -15
rect 19185 -35 19215 -15
rect 19235 -35 19265 -15
rect 19285 -35 19315 -15
rect 19335 -35 19365 -15
rect 19385 -35 19415 -15
rect 19435 -35 19465 -15
rect 19485 -35 19515 -15
rect 19535 -35 19565 -15
rect 19585 -35 19615 -15
rect 19635 -35 19665 -15
rect 19685 -35 19715 -15
rect 19735 -35 19765 -15
rect 19785 -35 19815 -15
rect 19835 -35 19865 -15
rect 19885 -35 19915 -15
rect 19935 -35 19965 -15
rect 19985 -35 20015 -15
rect 20035 -35 20065 -15
rect 20085 -35 20115 -15
rect 20135 -35 20165 -15
rect 20185 -35 20215 -15
rect 20235 -35 20265 -15
rect 20285 -35 20315 -15
rect 20335 -35 20365 -15
rect 20385 -35 20400 -15
rect -650 -50 20400 -35
rect -650 -115 -600 -100
rect -650 -135 -635 -115
rect -615 -135 -600 -115
rect -650 -165 -600 -135
rect -650 -185 -635 -165
rect -615 -185 -600 -165
rect -650 -215 -600 -185
rect -650 -235 -635 -215
rect -615 -235 -600 -215
rect -650 -265 -600 -235
rect -650 -285 -635 -265
rect -615 -285 -600 -265
rect -650 -315 -600 -285
rect -650 -335 -635 -315
rect -615 -335 -600 -315
rect -650 -365 -600 -335
rect -650 -385 -635 -365
rect -615 -385 -600 -365
rect -650 -415 -600 -385
rect -650 -435 -635 -415
rect -615 -435 -600 -415
rect -650 -465 -600 -435
rect -650 -485 -635 -465
rect -615 -485 -600 -465
rect -650 -515 -600 -485
rect -650 -535 -635 -515
rect -615 -535 -600 -515
rect -650 -565 -600 -535
rect -650 -585 -635 -565
rect -615 -585 -600 -565
rect -650 -615 -600 -585
rect -650 -635 -635 -615
rect -615 -635 -600 -615
rect -650 -665 -600 -635
rect -650 -685 -635 -665
rect -615 -685 -600 -665
rect -650 -715 -600 -685
rect -650 -735 -635 -715
rect -615 -735 -600 -715
rect -650 -765 -600 -735
rect -650 -785 -635 -765
rect -615 -785 -600 -765
rect -650 -800 -600 -785
rect -500 -115 -450 -100
rect -500 -135 -485 -115
rect -465 -135 -450 -115
rect -500 -165 -450 -135
rect -500 -185 -485 -165
rect -465 -185 -450 -165
rect -500 -215 -450 -185
rect -500 -235 -485 -215
rect -465 -235 -450 -215
rect -500 -265 -450 -235
rect -500 -285 -485 -265
rect -465 -285 -450 -265
rect -500 -315 -450 -285
rect -500 -335 -485 -315
rect -465 -335 -450 -315
rect -500 -365 -450 -335
rect -500 -385 -485 -365
rect -465 -385 -450 -365
rect -500 -415 -450 -385
rect -500 -435 -485 -415
rect -465 -435 -450 -415
rect -500 -465 -450 -435
rect -500 -485 -485 -465
rect -465 -485 -450 -465
rect -500 -515 -450 -485
rect -500 -535 -485 -515
rect -465 -535 -450 -515
rect -500 -565 -450 -535
rect -500 -585 -485 -565
rect -465 -585 -450 -565
rect -500 -615 -450 -585
rect -500 -635 -485 -615
rect -465 -635 -450 -615
rect -500 -665 -450 -635
rect -500 -685 -485 -665
rect -465 -685 -450 -665
rect -500 -715 -450 -685
rect -500 -735 -485 -715
rect -465 -735 -450 -715
rect -500 -765 -450 -735
rect -500 -785 -485 -765
rect -465 -785 -450 -765
rect -500 -800 -450 -785
rect -350 -115 -300 -100
rect -350 -135 -335 -115
rect -315 -135 -300 -115
rect -350 -165 -300 -135
rect -350 -185 -335 -165
rect -315 -185 -300 -165
rect -350 -215 -300 -185
rect -350 -235 -335 -215
rect -315 -235 -300 -215
rect -350 -265 -300 -235
rect -350 -285 -335 -265
rect -315 -285 -300 -265
rect -350 -315 -300 -285
rect -350 -335 -335 -315
rect -315 -335 -300 -315
rect -350 -365 -300 -335
rect -350 -385 -335 -365
rect -315 -385 -300 -365
rect -350 -415 -300 -385
rect -350 -435 -335 -415
rect -315 -435 -300 -415
rect -350 -465 -300 -435
rect -350 -485 -335 -465
rect -315 -485 -300 -465
rect -350 -515 -300 -485
rect -350 -535 -335 -515
rect -315 -535 -300 -515
rect -350 -565 -300 -535
rect -350 -585 -335 -565
rect -315 -585 -300 -565
rect -350 -615 -300 -585
rect -350 -635 -335 -615
rect -315 -635 -300 -615
rect -350 -665 -300 -635
rect -350 -685 -335 -665
rect -315 -685 -300 -665
rect -350 -715 -300 -685
rect -350 -735 -335 -715
rect -315 -735 -300 -715
rect -350 -765 -300 -735
rect -350 -785 -335 -765
rect -315 -785 -300 -765
rect -350 -800 -300 -785
rect -200 -115 -150 -100
rect -200 -135 -185 -115
rect -165 -135 -150 -115
rect -200 -165 -150 -135
rect -200 -185 -185 -165
rect -165 -185 -150 -165
rect -200 -215 -150 -185
rect -200 -235 -185 -215
rect -165 -235 -150 -215
rect -200 -265 -150 -235
rect -200 -285 -185 -265
rect -165 -285 -150 -265
rect -200 -315 -150 -285
rect -200 -335 -185 -315
rect -165 -335 -150 -315
rect -200 -365 -150 -335
rect -200 -385 -185 -365
rect -165 -385 -150 -365
rect -200 -415 -150 -385
rect -200 -435 -185 -415
rect -165 -435 -150 -415
rect -200 -465 -150 -435
rect -200 -485 -185 -465
rect -165 -485 -150 -465
rect -200 -515 -150 -485
rect -200 -535 -185 -515
rect -165 -535 -150 -515
rect -200 -565 -150 -535
rect -200 -585 -185 -565
rect -165 -585 -150 -565
rect -200 -615 -150 -585
rect -200 -635 -185 -615
rect -165 -635 -150 -615
rect -200 -665 -150 -635
rect -200 -685 -185 -665
rect -165 -685 -150 -665
rect -200 -715 -150 -685
rect -200 -735 -185 -715
rect -165 -735 -150 -715
rect -200 -765 -150 -735
rect -200 -785 -185 -765
rect -165 -785 -150 -765
rect -200 -800 -150 -785
rect -50 -115 0 -100
rect -50 -135 -35 -115
rect -15 -135 0 -115
rect -50 -165 0 -135
rect -50 -185 -35 -165
rect -15 -185 0 -165
rect -50 -215 0 -185
rect -50 -235 -35 -215
rect -15 -235 0 -215
rect -50 -265 0 -235
rect -50 -285 -35 -265
rect -15 -285 0 -265
rect -50 -315 0 -285
rect -50 -335 -35 -315
rect -15 -335 0 -315
rect -50 -365 0 -335
rect -50 -385 -35 -365
rect -15 -385 0 -365
rect -50 -415 0 -385
rect -50 -435 -35 -415
rect -15 -435 0 -415
rect -50 -465 0 -435
rect -50 -485 -35 -465
rect -15 -485 0 -465
rect -50 -515 0 -485
rect -50 -535 -35 -515
rect -15 -535 0 -515
rect -50 -565 0 -535
rect -50 -585 -35 -565
rect -15 -585 0 -565
rect -50 -615 0 -585
rect -50 -635 -35 -615
rect -15 -635 0 -615
rect -50 -665 0 -635
rect -50 -685 -35 -665
rect -15 -685 0 -665
rect -50 -715 0 -685
rect -50 -735 -35 -715
rect -15 -735 0 -715
rect -50 -765 0 -735
rect -50 -785 -35 -765
rect -15 -785 0 -765
rect -50 -800 0 -785
rect 1150 -115 1200 -100
rect 1150 -135 1165 -115
rect 1185 -135 1200 -115
rect 1150 -165 1200 -135
rect 1150 -185 1165 -165
rect 1185 -185 1200 -165
rect 1150 -215 1200 -185
rect 1150 -235 1165 -215
rect 1185 -235 1200 -215
rect 1150 -265 1200 -235
rect 1150 -285 1165 -265
rect 1185 -285 1200 -265
rect 1150 -315 1200 -285
rect 1150 -335 1165 -315
rect 1185 -335 1200 -315
rect 1150 -365 1200 -335
rect 1150 -385 1165 -365
rect 1185 -385 1200 -365
rect 1150 -415 1200 -385
rect 1150 -435 1165 -415
rect 1185 -435 1200 -415
rect 1150 -465 1200 -435
rect 1150 -485 1165 -465
rect 1185 -485 1200 -465
rect 1150 -515 1200 -485
rect 1150 -535 1165 -515
rect 1185 -535 1200 -515
rect 1150 -565 1200 -535
rect 1150 -585 1165 -565
rect 1185 -585 1200 -565
rect 1150 -615 1200 -585
rect 1150 -635 1165 -615
rect 1185 -635 1200 -615
rect 1150 -665 1200 -635
rect 1150 -685 1165 -665
rect 1185 -685 1200 -665
rect 1150 -715 1200 -685
rect 1150 -735 1165 -715
rect 1185 -735 1200 -715
rect 1150 -765 1200 -735
rect 1150 -785 1165 -765
rect 1185 -785 1200 -765
rect 1150 -800 1200 -785
rect 1450 -115 1500 -100
rect 1450 -135 1465 -115
rect 1485 -135 1500 -115
rect 1450 -165 1500 -135
rect 1450 -185 1465 -165
rect 1485 -185 1500 -165
rect 1450 -215 1500 -185
rect 1450 -235 1465 -215
rect 1485 -235 1500 -215
rect 1450 -265 1500 -235
rect 1450 -285 1465 -265
rect 1485 -285 1500 -265
rect 1450 -315 1500 -285
rect 1450 -335 1465 -315
rect 1485 -335 1500 -315
rect 1450 -365 1500 -335
rect 1450 -385 1465 -365
rect 1485 -385 1500 -365
rect 1450 -415 1500 -385
rect 1450 -435 1465 -415
rect 1485 -435 1500 -415
rect 1450 -465 1500 -435
rect 1450 -485 1465 -465
rect 1485 -485 1500 -465
rect 1450 -515 1500 -485
rect 1450 -535 1465 -515
rect 1485 -535 1500 -515
rect 1450 -565 1500 -535
rect 1450 -585 1465 -565
rect 1485 -585 1500 -565
rect 1450 -615 1500 -585
rect 1450 -635 1465 -615
rect 1485 -635 1500 -615
rect 1450 -665 1500 -635
rect 1450 -685 1465 -665
rect 1485 -685 1500 -665
rect 1450 -715 1500 -685
rect 1450 -735 1465 -715
rect 1485 -735 1500 -715
rect 1450 -765 1500 -735
rect 1450 -785 1465 -765
rect 1485 -785 1500 -765
rect 1450 -800 1500 -785
rect 1750 -115 1800 -100
rect 1750 -135 1765 -115
rect 1785 -135 1800 -115
rect 1750 -165 1800 -135
rect 1750 -185 1765 -165
rect 1785 -185 1800 -165
rect 1750 -215 1800 -185
rect 1750 -235 1765 -215
rect 1785 -235 1800 -215
rect 1750 -265 1800 -235
rect 1750 -285 1765 -265
rect 1785 -285 1800 -265
rect 1750 -315 1800 -285
rect 1750 -335 1765 -315
rect 1785 -335 1800 -315
rect 1750 -365 1800 -335
rect 1750 -385 1765 -365
rect 1785 -385 1800 -365
rect 1750 -415 1800 -385
rect 1750 -435 1765 -415
rect 1785 -435 1800 -415
rect 1750 -465 1800 -435
rect 1750 -485 1765 -465
rect 1785 -485 1800 -465
rect 1750 -515 1800 -485
rect 1750 -535 1765 -515
rect 1785 -535 1800 -515
rect 1750 -565 1800 -535
rect 1750 -585 1765 -565
rect 1785 -585 1800 -565
rect 1750 -615 1800 -585
rect 1750 -635 1765 -615
rect 1785 -635 1800 -615
rect 1750 -665 1800 -635
rect 1750 -685 1765 -665
rect 1785 -685 1800 -665
rect 1750 -715 1800 -685
rect 1750 -735 1765 -715
rect 1785 -735 1800 -715
rect 1750 -765 1800 -735
rect 1750 -785 1765 -765
rect 1785 -785 1800 -765
rect 1750 -800 1800 -785
rect 2050 -115 2100 -100
rect 2050 -135 2065 -115
rect 2085 -135 2100 -115
rect 2050 -165 2100 -135
rect 2050 -185 2065 -165
rect 2085 -185 2100 -165
rect 2050 -215 2100 -185
rect 2050 -235 2065 -215
rect 2085 -235 2100 -215
rect 2050 -265 2100 -235
rect 2050 -285 2065 -265
rect 2085 -285 2100 -265
rect 2050 -315 2100 -285
rect 2050 -335 2065 -315
rect 2085 -335 2100 -315
rect 2050 -365 2100 -335
rect 2050 -385 2065 -365
rect 2085 -385 2100 -365
rect 2050 -415 2100 -385
rect 2050 -435 2065 -415
rect 2085 -435 2100 -415
rect 2050 -465 2100 -435
rect 2050 -485 2065 -465
rect 2085 -485 2100 -465
rect 2050 -515 2100 -485
rect 2050 -535 2065 -515
rect 2085 -535 2100 -515
rect 2050 -565 2100 -535
rect 2050 -585 2065 -565
rect 2085 -585 2100 -565
rect 2050 -615 2100 -585
rect 2050 -635 2065 -615
rect 2085 -635 2100 -615
rect 2050 -665 2100 -635
rect 2050 -685 2065 -665
rect 2085 -685 2100 -665
rect 2050 -715 2100 -685
rect 2050 -735 2065 -715
rect 2085 -735 2100 -715
rect 2050 -765 2100 -735
rect 2050 -785 2065 -765
rect 2085 -785 2100 -765
rect 2050 -800 2100 -785
rect 2350 -115 2400 -100
rect 2350 -135 2365 -115
rect 2385 -135 2400 -115
rect 2350 -165 2400 -135
rect 2350 -185 2365 -165
rect 2385 -185 2400 -165
rect 2350 -215 2400 -185
rect 2350 -235 2365 -215
rect 2385 -235 2400 -215
rect 2350 -265 2400 -235
rect 2350 -285 2365 -265
rect 2385 -285 2400 -265
rect 2350 -315 2400 -285
rect 2350 -335 2365 -315
rect 2385 -335 2400 -315
rect 2350 -365 2400 -335
rect 2350 -385 2365 -365
rect 2385 -385 2400 -365
rect 2350 -415 2400 -385
rect 2350 -435 2365 -415
rect 2385 -435 2400 -415
rect 2350 -465 2400 -435
rect 2350 -485 2365 -465
rect 2385 -485 2400 -465
rect 2350 -515 2400 -485
rect 2350 -535 2365 -515
rect 2385 -535 2400 -515
rect 2350 -565 2400 -535
rect 2350 -585 2365 -565
rect 2385 -585 2400 -565
rect 2350 -615 2400 -585
rect 2350 -635 2365 -615
rect 2385 -635 2400 -615
rect 2350 -665 2400 -635
rect 2350 -685 2365 -665
rect 2385 -685 2400 -665
rect 2350 -715 2400 -685
rect 2350 -735 2365 -715
rect 2385 -735 2400 -715
rect 2350 -765 2400 -735
rect 2350 -785 2365 -765
rect 2385 -785 2400 -765
rect 2350 -800 2400 -785
rect 2650 -115 2700 -100
rect 2650 -135 2665 -115
rect 2685 -135 2700 -115
rect 2650 -165 2700 -135
rect 2650 -185 2665 -165
rect 2685 -185 2700 -165
rect 2650 -215 2700 -185
rect 2650 -235 2665 -215
rect 2685 -235 2700 -215
rect 2650 -265 2700 -235
rect 2650 -285 2665 -265
rect 2685 -285 2700 -265
rect 2650 -315 2700 -285
rect 2650 -335 2665 -315
rect 2685 -335 2700 -315
rect 2650 -365 2700 -335
rect 2650 -385 2665 -365
rect 2685 -385 2700 -365
rect 2650 -415 2700 -385
rect 2650 -435 2665 -415
rect 2685 -435 2700 -415
rect 2650 -465 2700 -435
rect 2650 -485 2665 -465
rect 2685 -485 2700 -465
rect 2650 -515 2700 -485
rect 2650 -535 2665 -515
rect 2685 -535 2700 -515
rect 2650 -565 2700 -535
rect 2650 -585 2665 -565
rect 2685 -585 2700 -565
rect 2650 -615 2700 -585
rect 2650 -635 2665 -615
rect 2685 -635 2700 -615
rect 2650 -665 2700 -635
rect 2650 -685 2665 -665
rect 2685 -685 2700 -665
rect 2650 -715 2700 -685
rect 2650 -735 2665 -715
rect 2685 -735 2700 -715
rect 2650 -765 2700 -735
rect 2650 -785 2665 -765
rect 2685 -785 2700 -765
rect 2650 -800 2700 -785
rect 2950 -115 3000 -100
rect 2950 -135 2965 -115
rect 2985 -135 3000 -115
rect 2950 -165 3000 -135
rect 2950 -185 2965 -165
rect 2985 -185 3000 -165
rect 2950 -215 3000 -185
rect 2950 -235 2965 -215
rect 2985 -235 3000 -215
rect 2950 -265 3000 -235
rect 2950 -285 2965 -265
rect 2985 -285 3000 -265
rect 2950 -315 3000 -285
rect 2950 -335 2965 -315
rect 2985 -335 3000 -315
rect 2950 -365 3000 -335
rect 2950 -385 2965 -365
rect 2985 -385 3000 -365
rect 2950 -415 3000 -385
rect 2950 -435 2965 -415
rect 2985 -435 3000 -415
rect 2950 -465 3000 -435
rect 2950 -485 2965 -465
rect 2985 -485 3000 -465
rect 2950 -515 3000 -485
rect 2950 -535 2965 -515
rect 2985 -535 3000 -515
rect 2950 -565 3000 -535
rect 2950 -585 2965 -565
rect 2985 -585 3000 -565
rect 2950 -615 3000 -585
rect 2950 -635 2965 -615
rect 2985 -635 3000 -615
rect 2950 -665 3000 -635
rect 2950 -685 2965 -665
rect 2985 -685 3000 -665
rect 2950 -715 3000 -685
rect 2950 -735 2965 -715
rect 2985 -735 3000 -715
rect 2950 -765 3000 -735
rect 2950 -785 2965 -765
rect 2985 -785 3000 -765
rect 2950 -800 3000 -785
rect 3250 -115 3300 -100
rect 3250 -135 3265 -115
rect 3285 -135 3300 -115
rect 3250 -165 3300 -135
rect 3250 -185 3265 -165
rect 3285 -185 3300 -165
rect 3250 -215 3300 -185
rect 3250 -235 3265 -215
rect 3285 -235 3300 -215
rect 3250 -265 3300 -235
rect 3250 -285 3265 -265
rect 3285 -285 3300 -265
rect 3250 -315 3300 -285
rect 3250 -335 3265 -315
rect 3285 -335 3300 -315
rect 3250 -365 3300 -335
rect 3250 -385 3265 -365
rect 3285 -385 3300 -365
rect 3250 -415 3300 -385
rect 3250 -435 3265 -415
rect 3285 -435 3300 -415
rect 3250 -465 3300 -435
rect 3250 -485 3265 -465
rect 3285 -485 3300 -465
rect 3250 -515 3300 -485
rect 3250 -535 3265 -515
rect 3285 -535 3300 -515
rect 3250 -565 3300 -535
rect 3250 -585 3265 -565
rect 3285 -585 3300 -565
rect 3250 -615 3300 -585
rect 3250 -635 3265 -615
rect 3285 -635 3300 -615
rect 3250 -665 3300 -635
rect 3250 -685 3265 -665
rect 3285 -685 3300 -665
rect 3250 -715 3300 -685
rect 3250 -735 3265 -715
rect 3285 -735 3300 -715
rect 3250 -765 3300 -735
rect 3250 -785 3265 -765
rect 3285 -785 3300 -765
rect 3250 -800 3300 -785
rect 3550 -115 3600 -100
rect 3550 -135 3565 -115
rect 3585 -135 3600 -115
rect 3550 -165 3600 -135
rect 3550 -185 3565 -165
rect 3585 -185 3600 -165
rect 3550 -215 3600 -185
rect 3550 -235 3565 -215
rect 3585 -235 3600 -215
rect 3550 -265 3600 -235
rect 3550 -285 3565 -265
rect 3585 -285 3600 -265
rect 3550 -315 3600 -285
rect 3550 -335 3565 -315
rect 3585 -335 3600 -315
rect 3550 -365 3600 -335
rect 3550 -385 3565 -365
rect 3585 -385 3600 -365
rect 3550 -415 3600 -385
rect 3550 -435 3565 -415
rect 3585 -435 3600 -415
rect 3550 -465 3600 -435
rect 3550 -485 3565 -465
rect 3585 -485 3600 -465
rect 3550 -515 3600 -485
rect 3550 -535 3565 -515
rect 3585 -535 3600 -515
rect 3550 -565 3600 -535
rect 3550 -585 3565 -565
rect 3585 -585 3600 -565
rect 3550 -615 3600 -585
rect 3550 -635 3565 -615
rect 3585 -635 3600 -615
rect 3550 -665 3600 -635
rect 3550 -685 3565 -665
rect 3585 -685 3600 -665
rect 3550 -715 3600 -685
rect 3550 -735 3565 -715
rect 3585 -735 3600 -715
rect 3550 -765 3600 -735
rect 3550 -785 3565 -765
rect 3585 -785 3600 -765
rect 3550 -800 3600 -785
rect 3700 -115 3750 -100
rect 3700 -135 3715 -115
rect 3735 -135 3750 -115
rect 3700 -165 3750 -135
rect 3700 -185 3715 -165
rect 3735 -185 3750 -165
rect 3700 -215 3750 -185
rect 3700 -235 3715 -215
rect 3735 -235 3750 -215
rect 3700 -265 3750 -235
rect 3700 -285 3715 -265
rect 3735 -285 3750 -265
rect 3700 -315 3750 -285
rect 3700 -335 3715 -315
rect 3735 -335 3750 -315
rect 3700 -365 3750 -335
rect 3700 -385 3715 -365
rect 3735 -385 3750 -365
rect 3700 -415 3750 -385
rect 3700 -435 3715 -415
rect 3735 -435 3750 -415
rect 3700 -465 3750 -435
rect 3700 -485 3715 -465
rect 3735 -485 3750 -465
rect 3700 -515 3750 -485
rect 3700 -535 3715 -515
rect 3735 -535 3750 -515
rect 3700 -565 3750 -535
rect 3700 -585 3715 -565
rect 3735 -585 3750 -565
rect 3700 -615 3750 -585
rect 3700 -635 3715 -615
rect 3735 -635 3750 -615
rect 3700 -665 3750 -635
rect 3700 -685 3715 -665
rect 3735 -685 3750 -665
rect 3700 -715 3750 -685
rect 3700 -735 3715 -715
rect 3735 -735 3750 -715
rect 3700 -765 3750 -735
rect 3700 -785 3715 -765
rect 3735 -785 3750 -765
rect 3700 -800 3750 -785
rect 3850 -115 3900 -100
rect 3850 -135 3865 -115
rect 3885 -135 3900 -115
rect 3850 -165 3900 -135
rect 3850 -185 3865 -165
rect 3885 -185 3900 -165
rect 3850 -215 3900 -185
rect 3850 -235 3865 -215
rect 3885 -235 3900 -215
rect 3850 -265 3900 -235
rect 3850 -285 3865 -265
rect 3885 -285 3900 -265
rect 3850 -315 3900 -285
rect 3850 -335 3865 -315
rect 3885 -335 3900 -315
rect 3850 -365 3900 -335
rect 3850 -385 3865 -365
rect 3885 -385 3900 -365
rect 3850 -415 3900 -385
rect 3850 -435 3865 -415
rect 3885 -435 3900 -415
rect 3850 -465 3900 -435
rect 3850 -485 3865 -465
rect 3885 -485 3900 -465
rect 3850 -515 3900 -485
rect 3850 -535 3865 -515
rect 3885 -535 3900 -515
rect 3850 -565 3900 -535
rect 3850 -585 3865 -565
rect 3885 -585 3900 -565
rect 3850 -615 3900 -585
rect 3850 -635 3865 -615
rect 3885 -635 3900 -615
rect 3850 -665 3900 -635
rect 3850 -685 3865 -665
rect 3885 -685 3900 -665
rect 3850 -715 3900 -685
rect 3850 -735 3865 -715
rect 3885 -735 3900 -715
rect 3850 -765 3900 -735
rect 3850 -785 3865 -765
rect 3885 -785 3900 -765
rect 3850 -800 3900 -785
rect 4000 -115 4050 -100
rect 4000 -135 4015 -115
rect 4035 -135 4050 -115
rect 4000 -165 4050 -135
rect 4000 -185 4015 -165
rect 4035 -185 4050 -165
rect 4000 -215 4050 -185
rect 4000 -235 4015 -215
rect 4035 -235 4050 -215
rect 4000 -265 4050 -235
rect 4000 -285 4015 -265
rect 4035 -285 4050 -265
rect 4000 -315 4050 -285
rect 4000 -335 4015 -315
rect 4035 -335 4050 -315
rect 4000 -365 4050 -335
rect 4000 -385 4015 -365
rect 4035 -385 4050 -365
rect 4000 -415 4050 -385
rect 4000 -435 4015 -415
rect 4035 -435 4050 -415
rect 4000 -465 4050 -435
rect 4000 -485 4015 -465
rect 4035 -485 4050 -465
rect 4000 -515 4050 -485
rect 4000 -535 4015 -515
rect 4035 -535 4050 -515
rect 4000 -565 4050 -535
rect 4000 -585 4015 -565
rect 4035 -585 4050 -565
rect 4000 -615 4050 -585
rect 4000 -635 4015 -615
rect 4035 -635 4050 -615
rect 4000 -665 4050 -635
rect 4000 -685 4015 -665
rect 4035 -685 4050 -665
rect 4000 -715 4050 -685
rect 4000 -735 4015 -715
rect 4035 -735 4050 -715
rect 4000 -765 4050 -735
rect 4000 -785 4015 -765
rect 4035 -785 4050 -765
rect 4000 -800 4050 -785
rect 4150 -115 4200 -100
rect 4150 -135 4165 -115
rect 4185 -135 4200 -115
rect 4150 -165 4200 -135
rect 4150 -185 4165 -165
rect 4185 -185 4200 -165
rect 4150 -215 4200 -185
rect 4150 -235 4165 -215
rect 4185 -235 4200 -215
rect 4150 -265 4200 -235
rect 4150 -285 4165 -265
rect 4185 -285 4200 -265
rect 4150 -315 4200 -285
rect 4150 -335 4165 -315
rect 4185 -335 4200 -315
rect 4150 -365 4200 -335
rect 4150 -385 4165 -365
rect 4185 -385 4200 -365
rect 4150 -415 4200 -385
rect 4150 -435 4165 -415
rect 4185 -435 4200 -415
rect 4150 -465 4200 -435
rect 4150 -485 4165 -465
rect 4185 -485 4200 -465
rect 4150 -515 4200 -485
rect 4150 -535 4165 -515
rect 4185 -535 4200 -515
rect 4150 -565 4200 -535
rect 4150 -585 4165 -565
rect 4185 -585 4200 -565
rect 4150 -615 4200 -585
rect 4150 -635 4165 -615
rect 4185 -635 4200 -615
rect 4150 -665 4200 -635
rect 4150 -685 4165 -665
rect 4185 -685 4200 -665
rect 4150 -715 4200 -685
rect 4150 -735 4165 -715
rect 4185 -735 4200 -715
rect 4150 -765 4200 -735
rect 4150 -785 4165 -765
rect 4185 -785 4200 -765
rect 4150 -800 4200 -785
rect 4300 -115 4350 -100
rect 4300 -135 4315 -115
rect 4335 -135 4350 -115
rect 4300 -165 4350 -135
rect 4300 -185 4315 -165
rect 4335 -185 4350 -165
rect 4300 -215 4350 -185
rect 4300 -235 4315 -215
rect 4335 -235 4350 -215
rect 4300 -265 4350 -235
rect 4300 -285 4315 -265
rect 4335 -285 4350 -265
rect 4300 -315 4350 -285
rect 4300 -335 4315 -315
rect 4335 -335 4350 -315
rect 4300 -365 4350 -335
rect 4300 -385 4315 -365
rect 4335 -385 4350 -365
rect 4300 -415 4350 -385
rect 4300 -435 4315 -415
rect 4335 -435 4350 -415
rect 4300 -465 4350 -435
rect 4300 -485 4315 -465
rect 4335 -485 4350 -465
rect 4300 -515 4350 -485
rect 4300 -535 4315 -515
rect 4335 -535 4350 -515
rect 4300 -565 4350 -535
rect 4300 -585 4315 -565
rect 4335 -585 4350 -565
rect 4300 -615 4350 -585
rect 4300 -635 4315 -615
rect 4335 -635 4350 -615
rect 4300 -665 4350 -635
rect 4300 -685 4315 -665
rect 4335 -685 4350 -665
rect 4300 -715 4350 -685
rect 4300 -735 4315 -715
rect 4335 -735 4350 -715
rect 4300 -765 4350 -735
rect 4300 -785 4315 -765
rect 4335 -785 4350 -765
rect 4300 -800 4350 -785
rect 4450 -115 4500 -100
rect 4450 -135 4465 -115
rect 4485 -135 4500 -115
rect 4450 -165 4500 -135
rect 4450 -185 4465 -165
rect 4485 -185 4500 -165
rect 4450 -215 4500 -185
rect 4450 -235 4465 -215
rect 4485 -235 4500 -215
rect 4450 -265 4500 -235
rect 4450 -285 4465 -265
rect 4485 -285 4500 -265
rect 4450 -315 4500 -285
rect 4450 -335 4465 -315
rect 4485 -335 4500 -315
rect 4450 -365 4500 -335
rect 4450 -385 4465 -365
rect 4485 -385 4500 -365
rect 4450 -415 4500 -385
rect 4450 -435 4465 -415
rect 4485 -435 4500 -415
rect 4450 -465 4500 -435
rect 4450 -485 4465 -465
rect 4485 -485 4500 -465
rect 4450 -515 4500 -485
rect 4450 -535 4465 -515
rect 4485 -535 4500 -515
rect 4450 -565 4500 -535
rect 4450 -585 4465 -565
rect 4485 -585 4500 -565
rect 4450 -615 4500 -585
rect 4450 -635 4465 -615
rect 4485 -635 4500 -615
rect 4450 -665 4500 -635
rect 4450 -685 4465 -665
rect 4485 -685 4500 -665
rect 4450 -715 4500 -685
rect 4450 -735 4465 -715
rect 4485 -735 4500 -715
rect 4450 -765 4500 -735
rect 4450 -785 4465 -765
rect 4485 -785 4500 -765
rect 4450 -800 4500 -785
rect 4600 -115 4650 -100
rect 4600 -135 4615 -115
rect 4635 -135 4650 -115
rect 4600 -165 4650 -135
rect 4600 -185 4615 -165
rect 4635 -185 4650 -165
rect 4600 -215 4650 -185
rect 4600 -235 4615 -215
rect 4635 -235 4650 -215
rect 4600 -265 4650 -235
rect 4600 -285 4615 -265
rect 4635 -285 4650 -265
rect 4600 -315 4650 -285
rect 4600 -335 4615 -315
rect 4635 -335 4650 -315
rect 4600 -365 4650 -335
rect 4600 -385 4615 -365
rect 4635 -385 4650 -365
rect 4600 -415 4650 -385
rect 4600 -435 4615 -415
rect 4635 -435 4650 -415
rect 4600 -465 4650 -435
rect 4600 -485 4615 -465
rect 4635 -485 4650 -465
rect 4600 -515 4650 -485
rect 4600 -535 4615 -515
rect 4635 -535 4650 -515
rect 4600 -565 4650 -535
rect 4600 -585 4615 -565
rect 4635 -585 4650 -565
rect 4600 -615 4650 -585
rect 4600 -635 4615 -615
rect 4635 -635 4650 -615
rect 4600 -665 4650 -635
rect 4600 -685 4615 -665
rect 4635 -685 4650 -665
rect 4600 -715 4650 -685
rect 4600 -735 4615 -715
rect 4635 -735 4650 -715
rect 4600 -765 4650 -735
rect 4600 -785 4615 -765
rect 4635 -785 4650 -765
rect 4600 -800 4650 -785
rect 4750 -115 4800 -100
rect 4750 -135 4765 -115
rect 4785 -135 4800 -115
rect 4750 -165 4800 -135
rect 4750 -185 4765 -165
rect 4785 -185 4800 -165
rect 4750 -215 4800 -185
rect 4750 -235 4765 -215
rect 4785 -235 4800 -215
rect 4750 -265 4800 -235
rect 4750 -285 4765 -265
rect 4785 -285 4800 -265
rect 4750 -315 4800 -285
rect 4750 -335 4765 -315
rect 4785 -335 4800 -315
rect 4750 -365 4800 -335
rect 4750 -385 4765 -365
rect 4785 -385 4800 -365
rect 4750 -415 4800 -385
rect 4750 -435 4765 -415
rect 4785 -435 4800 -415
rect 4750 -465 4800 -435
rect 4750 -485 4765 -465
rect 4785 -485 4800 -465
rect 4750 -515 4800 -485
rect 4750 -535 4765 -515
rect 4785 -535 4800 -515
rect 4750 -565 4800 -535
rect 4750 -585 4765 -565
rect 4785 -585 4800 -565
rect 4750 -615 4800 -585
rect 4750 -635 4765 -615
rect 4785 -635 4800 -615
rect 4750 -665 4800 -635
rect 4750 -685 4765 -665
rect 4785 -685 4800 -665
rect 4750 -715 4800 -685
rect 4750 -735 4765 -715
rect 4785 -735 4800 -715
rect 4750 -765 4800 -735
rect 4750 -785 4765 -765
rect 4785 -785 4800 -765
rect 4750 -800 4800 -785
rect 5050 -115 5100 -100
rect 5050 -135 5065 -115
rect 5085 -135 5100 -115
rect 5050 -165 5100 -135
rect 5050 -185 5065 -165
rect 5085 -185 5100 -165
rect 5050 -215 5100 -185
rect 5050 -235 5065 -215
rect 5085 -235 5100 -215
rect 5050 -265 5100 -235
rect 5050 -285 5065 -265
rect 5085 -285 5100 -265
rect 5050 -315 5100 -285
rect 5050 -335 5065 -315
rect 5085 -335 5100 -315
rect 5050 -365 5100 -335
rect 5050 -385 5065 -365
rect 5085 -385 5100 -365
rect 5050 -415 5100 -385
rect 5050 -435 5065 -415
rect 5085 -435 5100 -415
rect 5050 -465 5100 -435
rect 5050 -485 5065 -465
rect 5085 -485 5100 -465
rect 5050 -515 5100 -485
rect 5050 -535 5065 -515
rect 5085 -535 5100 -515
rect 5050 -565 5100 -535
rect 5050 -585 5065 -565
rect 5085 -585 5100 -565
rect 5050 -615 5100 -585
rect 5050 -635 5065 -615
rect 5085 -635 5100 -615
rect 5050 -665 5100 -635
rect 5050 -685 5065 -665
rect 5085 -685 5100 -665
rect 5050 -715 5100 -685
rect 5050 -735 5065 -715
rect 5085 -735 5100 -715
rect 5050 -765 5100 -735
rect 5050 -785 5065 -765
rect 5085 -785 5100 -765
rect 5050 -800 5100 -785
rect 5350 -115 5400 -100
rect 5350 -135 5365 -115
rect 5385 -135 5400 -115
rect 5350 -165 5400 -135
rect 5350 -185 5365 -165
rect 5385 -185 5400 -165
rect 5350 -215 5400 -185
rect 5350 -235 5365 -215
rect 5385 -235 5400 -215
rect 5350 -265 5400 -235
rect 5350 -285 5365 -265
rect 5385 -285 5400 -265
rect 5350 -315 5400 -285
rect 5350 -335 5365 -315
rect 5385 -335 5400 -315
rect 5350 -365 5400 -335
rect 5350 -385 5365 -365
rect 5385 -385 5400 -365
rect 5350 -415 5400 -385
rect 5350 -435 5365 -415
rect 5385 -435 5400 -415
rect 5350 -465 5400 -435
rect 5350 -485 5365 -465
rect 5385 -485 5400 -465
rect 5350 -515 5400 -485
rect 5350 -535 5365 -515
rect 5385 -535 5400 -515
rect 5350 -565 5400 -535
rect 5350 -585 5365 -565
rect 5385 -585 5400 -565
rect 5350 -615 5400 -585
rect 5350 -635 5365 -615
rect 5385 -635 5400 -615
rect 5350 -665 5400 -635
rect 5350 -685 5365 -665
rect 5385 -685 5400 -665
rect 5350 -715 5400 -685
rect 5350 -735 5365 -715
rect 5385 -735 5400 -715
rect 5350 -765 5400 -735
rect 5350 -785 5365 -765
rect 5385 -785 5400 -765
rect 5350 -800 5400 -785
rect 5650 -115 5700 -100
rect 5650 -135 5665 -115
rect 5685 -135 5700 -115
rect 5650 -165 5700 -135
rect 5650 -185 5665 -165
rect 5685 -185 5700 -165
rect 5650 -215 5700 -185
rect 5650 -235 5665 -215
rect 5685 -235 5700 -215
rect 5650 -265 5700 -235
rect 5650 -285 5665 -265
rect 5685 -285 5700 -265
rect 5650 -315 5700 -285
rect 5650 -335 5665 -315
rect 5685 -335 5700 -315
rect 5650 -365 5700 -335
rect 5650 -385 5665 -365
rect 5685 -385 5700 -365
rect 5650 -415 5700 -385
rect 5650 -435 5665 -415
rect 5685 -435 5700 -415
rect 5650 -465 5700 -435
rect 5650 -485 5665 -465
rect 5685 -485 5700 -465
rect 5650 -515 5700 -485
rect 5650 -535 5665 -515
rect 5685 -535 5700 -515
rect 5650 -565 5700 -535
rect 5650 -585 5665 -565
rect 5685 -585 5700 -565
rect 5650 -615 5700 -585
rect 5650 -635 5665 -615
rect 5685 -635 5700 -615
rect 5650 -665 5700 -635
rect 5650 -685 5665 -665
rect 5685 -685 5700 -665
rect 5650 -715 5700 -685
rect 5650 -735 5665 -715
rect 5685 -735 5700 -715
rect 5650 -765 5700 -735
rect 5650 -785 5665 -765
rect 5685 -785 5700 -765
rect 5650 -800 5700 -785
rect 5950 -115 6000 -100
rect 5950 -135 5965 -115
rect 5985 -135 6000 -115
rect 5950 -165 6000 -135
rect 5950 -185 5965 -165
rect 5985 -185 6000 -165
rect 5950 -215 6000 -185
rect 5950 -235 5965 -215
rect 5985 -235 6000 -215
rect 5950 -265 6000 -235
rect 5950 -285 5965 -265
rect 5985 -285 6000 -265
rect 5950 -315 6000 -285
rect 5950 -335 5965 -315
rect 5985 -335 6000 -315
rect 5950 -365 6000 -335
rect 5950 -385 5965 -365
rect 5985 -385 6000 -365
rect 5950 -415 6000 -385
rect 5950 -435 5965 -415
rect 5985 -435 6000 -415
rect 5950 -465 6000 -435
rect 5950 -485 5965 -465
rect 5985 -485 6000 -465
rect 5950 -515 6000 -485
rect 5950 -535 5965 -515
rect 5985 -535 6000 -515
rect 5950 -565 6000 -535
rect 5950 -585 5965 -565
rect 5985 -585 6000 -565
rect 5950 -615 6000 -585
rect 5950 -635 5965 -615
rect 5985 -635 6000 -615
rect 5950 -665 6000 -635
rect 5950 -685 5965 -665
rect 5985 -685 6000 -665
rect 5950 -715 6000 -685
rect 5950 -735 5965 -715
rect 5985 -735 6000 -715
rect 5950 -765 6000 -735
rect 5950 -785 5965 -765
rect 5985 -785 6000 -765
rect 5950 -800 6000 -785
rect 6250 -115 6300 -100
rect 6250 -135 6265 -115
rect 6285 -135 6300 -115
rect 6250 -165 6300 -135
rect 6250 -185 6265 -165
rect 6285 -185 6300 -165
rect 6250 -215 6300 -185
rect 6250 -235 6265 -215
rect 6285 -235 6300 -215
rect 6250 -265 6300 -235
rect 6250 -285 6265 -265
rect 6285 -285 6300 -265
rect 6250 -315 6300 -285
rect 6250 -335 6265 -315
rect 6285 -335 6300 -315
rect 6250 -365 6300 -335
rect 6250 -385 6265 -365
rect 6285 -385 6300 -365
rect 6250 -415 6300 -385
rect 6250 -435 6265 -415
rect 6285 -435 6300 -415
rect 6250 -465 6300 -435
rect 6250 -485 6265 -465
rect 6285 -485 6300 -465
rect 6250 -515 6300 -485
rect 6250 -535 6265 -515
rect 6285 -535 6300 -515
rect 6250 -565 6300 -535
rect 6250 -585 6265 -565
rect 6285 -585 6300 -565
rect 6250 -615 6300 -585
rect 6250 -635 6265 -615
rect 6285 -635 6300 -615
rect 6250 -665 6300 -635
rect 6250 -685 6265 -665
rect 6285 -685 6300 -665
rect 6250 -715 6300 -685
rect 6250 -735 6265 -715
rect 6285 -735 6300 -715
rect 6250 -765 6300 -735
rect 6250 -785 6265 -765
rect 6285 -785 6300 -765
rect 6250 -800 6300 -785
rect 6550 -115 6600 -100
rect 6550 -135 6565 -115
rect 6585 -135 6600 -115
rect 6550 -165 6600 -135
rect 6550 -185 6565 -165
rect 6585 -185 6600 -165
rect 6550 -215 6600 -185
rect 6550 -235 6565 -215
rect 6585 -235 6600 -215
rect 6550 -265 6600 -235
rect 6550 -285 6565 -265
rect 6585 -285 6600 -265
rect 6550 -315 6600 -285
rect 6550 -335 6565 -315
rect 6585 -335 6600 -315
rect 6550 -365 6600 -335
rect 6550 -385 6565 -365
rect 6585 -385 6600 -365
rect 6550 -415 6600 -385
rect 6550 -435 6565 -415
rect 6585 -435 6600 -415
rect 6550 -465 6600 -435
rect 6550 -485 6565 -465
rect 6585 -485 6600 -465
rect 6550 -515 6600 -485
rect 6550 -535 6565 -515
rect 6585 -535 6600 -515
rect 6550 -565 6600 -535
rect 6550 -585 6565 -565
rect 6585 -585 6600 -565
rect 6550 -615 6600 -585
rect 6550 -635 6565 -615
rect 6585 -635 6600 -615
rect 6550 -665 6600 -635
rect 6550 -685 6565 -665
rect 6585 -685 6600 -665
rect 6550 -715 6600 -685
rect 6550 -735 6565 -715
rect 6585 -735 6600 -715
rect 6550 -765 6600 -735
rect 6550 -785 6565 -765
rect 6585 -785 6600 -765
rect 6550 -800 6600 -785
rect 6850 -115 6900 -100
rect 6850 -135 6865 -115
rect 6885 -135 6900 -115
rect 6850 -165 6900 -135
rect 6850 -185 6865 -165
rect 6885 -185 6900 -165
rect 6850 -215 6900 -185
rect 6850 -235 6865 -215
rect 6885 -235 6900 -215
rect 6850 -265 6900 -235
rect 6850 -285 6865 -265
rect 6885 -285 6900 -265
rect 6850 -315 6900 -285
rect 6850 -335 6865 -315
rect 6885 -335 6900 -315
rect 6850 -365 6900 -335
rect 6850 -385 6865 -365
rect 6885 -385 6900 -365
rect 6850 -415 6900 -385
rect 6850 -435 6865 -415
rect 6885 -435 6900 -415
rect 6850 -465 6900 -435
rect 6850 -485 6865 -465
rect 6885 -485 6900 -465
rect 6850 -515 6900 -485
rect 6850 -535 6865 -515
rect 6885 -535 6900 -515
rect 6850 -565 6900 -535
rect 6850 -585 6865 -565
rect 6885 -585 6900 -565
rect 6850 -615 6900 -585
rect 6850 -635 6865 -615
rect 6885 -635 6900 -615
rect 6850 -665 6900 -635
rect 6850 -685 6865 -665
rect 6885 -685 6900 -665
rect 6850 -715 6900 -685
rect 6850 -735 6865 -715
rect 6885 -735 6900 -715
rect 6850 -765 6900 -735
rect 6850 -785 6865 -765
rect 6885 -785 6900 -765
rect 6850 -800 6900 -785
rect 7150 -115 7200 -100
rect 7150 -135 7165 -115
rect 7185 -135 7200 -115
rect 7150 -165 7200 -135
rect 7150 -185 7165 -165
rect 7185 -185 7200 -165
rect 7150 -215 7200 -185
rect 7150 -235 7165 -215
rect 7185 -235 7200 -215
rect 7150 -265 7200 -235
rect 7150 -285 7165 -265
rect 7185 -285 7200 -265
rect 7150 -315 7200 -285
rect 7150 -335 7165 -315
rect 7185 -335 7200 -315
rect 7150 -365 7200 -335
rect 7150 -385 7165 -365
rect 7185 -385 7200 -365
rect 7150 -415 7200 -385
rect 7150 -435 7165 -415
rect 7185 -435 7200 -415
rect 7150 -465 7200 -435
rect 7150 -485 7165 -465
rect 7185 -485 7200 -465
rect 7150 -515 7200 -485
rect 7150 -535 7165 -515
rect 7185 -535 7200 -515
rect 7150 -565 7200 -535
rect 7150 -585 7165 -565
rect 7185 -585 7200 -565
rect 7150 -615 7200 -585
rect 7150 -635 7165 -615
rect 7185 -635 7200 -615
rect 7150 -665 7200 -635
rect 7150 -685 7165 -665
rect 7185 -685 7200 -665
rect 7150 -715 7200 -685
rect 7150 -735 7165 -715
rect 7185 -735 7200 -715
rect 7150 -765 7200 -735
rect 7150 -785 7165 -765
rect 7185 -785 7200 -765
rect 7150 -800 7200 -785
rect 8350 -115 8400 -100
rect 8350 -135 8365 -115
rect 8385 -135 8400 -115
rect 8350 -165 8400 -135
rect 8350 -185 8365 -165
rect 8385 -185 8400 -165
rect 8350 -215 8400 -185
rect 8350 -235 8365 -215
rect 8385 -235 8400 -215
rect 8350 -265 8400 -235
rect 8350 -285 8365 -265
rect 8385 -285 8400 -265
rect 8350 -315 8400 -285
rect 8350 -335 8365 -315
rect 8385 -335 8400 -315
rect 8350 -365 8400 -335
rect 8350 -385 8365 -365
rect 8385 -385 8400 -365
rect 8350 -415 8400 -385
rect 8350 -435 8365 -415
rect 8385 -435 8400 -415
rect 8350 -465 8400 -435
rect 8350 -485 8365 -465
rect 8385 -485 8400 -465
rect 8350 -515 8400 -485
rect 8350 -535 8365 -515
rect 8385 -535 8400 -515
rect 8350 -565 8400 -535
rect 8350 -585 8365 -565
rect 8385 -585 8400 -565
rect 8350 -615 8400 -585
rect 8350 -635 8365 -615
rect 8385 -635 8400 -615
rect 8350 -665 8400 -635
rect 8350 -685 8365 -665
rect 8385 -685 8400 -665
rect 8350 -715 8400 -685
rect 8350 -735 8365 -715
rect 8385 -735 8400 -715
rect 8350 -765 8400 -735
rect 8350 -785 8365 -765
rect 8385 -785 8400 -765
rect 8350 -800 8400 -785
rect 9550 -115 9600 -100
rect 9550 -135 9565 -115
rect 9585 -135 9600 -115
rect 9550 -165 9600 -135
rect 9550 -185 9565 -165
rect 9585 -185 9600 -165
rect 9550 -215 9600 -185
rect 9550 -235 9565 -215
rect 9585 -235 9600 -215
rect 9550 -265 9600 -235
rect 9550 -285 9565 -265
rect 9585 -285 9600 -265
rect 9550 -315 9600 -285
rect 9550 -335 9565 -315
rect 9585 -335 9600 -315
rect 9550 -365 9600 -335
rect 9550 -385 9565 -365
rect 9585 -385 9600 -365
rect 9550 -415 9600 -385
rect 9550 -435 9565 -415
rect 9585 -435 9600 -415
rect 9550 -465 9600 -435
rect 9550 -485 9565 -465
rect 9585 -485 9600 -465
rect 9550 -515 9600 -485
rect 9550 -535 9565 -515
rect 9585 -535 9600 -515
rect 9550 -565 9600 -535
rect 9550 -585 9565 -565
rect 9585 -585 9600 -565
rect 9550 -615 9600 -585
rect 9550 -635 9565 -615
rect 9585 -635 9600 -615
rect 9550 -665 9600 -635
rect 9550 -685 9565 -665
rect 9585 -685 9600 -665
rect 9550 -715 9600 -685
rect 9550 -735 9565 -715
rect 9585 -735 9600 -715
rect 9550 -765 9600 -735
rect 9550 -785 9565 -765
rect 9585 -785 9600 -765
rect 9550 -800 9600 -785
rect 10750 -115 10800 -100
rect 10750 -135 10765 -115
rect 10785 -135 10800 -115
rect 10750 -165 10800 -135
rect 10750 -185 10765 -165
rect 10785 -185 10800 -165
rect 10750 -215 10800 -185
rect 10750 -235 10765 -215
rect 10785 -235 10800 -215
rect 10750 -265 10800 -235
rect 10750 -285 10765 -265
rect 10785 -285 10800 -265
rect 10750 -315 10800 -285
rect 10750 -335 10765 -315
rect 10785 -335 10800 -315
rect 10750 -365 10800 -335
rect 10750 -385 10765 -365
rect 10785 -385 10800 -365
rect 10750 -415 10800 -385
rect 10750 -435 10765 -415
rect 10785 -435 10800 -415
rect 10750 -465 10800 -435
rect 10750 -485 10765 -465
rect 10785 -485 10800 -465
rect 10750 -515 10800 -485
rect 10750 -535 10765 -515
rect 10785 -535 10800 -515
rect 10750 -565 10800 -535
rect 10750 -585 10765 -565
rect 10785 -585 10800 -565
rect 10750 -615 10800 -585
rect 10750 -635 10765 -615
rect 10785 -635 10800 -615
rect 10750 -665 10800 -635
rect 10750 -685 10765 -665
rect 10785 -685 10800 -665
rect 10750 -715 10800 -685
rect 10750 -735 10765 -715
rect 10785 -735 10800 -715
rect 10750 -765 10800 -735
rect 10750 -785 10765 -765
rect 10785 -785 10800 -765
rect 10750 -800 10800 -785
rect 11950 -115 12000 -100
rect 11950 -135 11965 -115
rect 11985 -135 12000 -115
rect 11950 -165 12000 -135
rect 11950 -185 11965 -165
rect 11985 -185 12000 -165
rect 11950 -215 12000 -185
rect 11950 -235 11965 -215
rect 11985 -235 12000 -215
rect 11950 -265 12000 -235
rect 11950 -285 11965 -265
rect 11985 -285 12000 -265
rect 11950 -315 12000 -285
rect 11950 -335 11965 -315
rect 11985 -335 12000 -315
rect 11950 -365 12000 -335
rect 11950 -385 11965 -365
rect 11985 -385 12000 -365
rect 11950 -415 12000 -385
rect 11950 -435 11965 -415
rect 11985 -435 12000 -415
rect 11950 -465 12000 -435
rect 11950 -485 11965 -465
rect 11985 -485 12000 -465
rect 11950 -515 12000 -485
rect 11950 -535 11965 -515
rect 11985 -535 12000 -515
rect 11950 -565 12000 -535
rect 11950 -585 11965 -565
rect 11985 -585 12000 -565
rect 11950 -615 12000 -585
rect 11950 -635 11965 -615
rect 11985 -635 12000 -615
rect 11950 -665 12000 -635
rect 11950 -685 11965 -665
rect 11985 -685 12000 -665
rect 11950 -715 12000 -685
rect 11950 -735 11965 -715
rect 11985 -735 12000 -715
rect 11950 -765 12000 -735
rect 11950 -785 11965 -765
rect 11985 -785 12000 -765
rect 11950 -800 12000 -785
rect 12250 -115 12300 -100
rect 12250 -135 12265 -115
rect 12285 -135 12300 -115
rect 12250 -165 12300 -135
rect 12250 -185 12265 -165
rect 12285 -185 12300 -165
rect 12250 -215 12300 -185
rect 12250 -235 12265 -215
rect 12285 -235 12300 -215
rect 12250 -265 12300 -235
rect 12250 -285 12265 -265
rect 12285 -285 12300 -265
rect 12250 -315 12300 -285
rect 12250 -335 12265 -315
rect 12285 -335 12300 -315
rect 12250 -365 12300 -335
rect 12250 -385 12265 -365
rect 12285 -385 12300 -365
rect 12250 -415 12300 -385
rect 12250 -435 12265 -415
rect 12285 -435 12300 -415
rect 12250 -465 12300 -435
rect 12250 -485 12265 -465
rect 12285 -485 12300 -465
rect 12250 -515 12300 -485
rect 12250 -535 12265 -515
rect 12285 -535 12300 -515
rect 12250 -565 12300 -535
rect 12250 -585 12265 -565
rect 12285 -585 12300 -565
rect 12250 -615 12300 -585
rect 12250 -635 12265 -615
rect 12285 -635 12300 -615
rect 12250 -665 12300 -635
rect 12250 -685 12265 -665
rect 12285 -685 12300 -665
rect 12250 -715 12300 -685
rect 12250 -735 12265 -715
rect 12285 -735 12300 -715
rect 12250 -765 12300 -735
rect 12250 -785 12265 -765
rect 12285 -785 12300 -765
rect 12250 -800 12300 -785
rect 12550 -115 12600 -100
rect 12550 -135 12565 -115
rect 12585 -135 12600 -115
rect 12550 -165 12600 -135
rect 12550 -185 12565 -165
rect 12585 -185 12600 -165
rect 12550 -215 12600 -185
rect 12550 -235 12565 -215
rect 12585 -235 12600 -215
rect 12550 -265 12600 -235
rect 12550 -285 12565 -265
rect 12585 -285 12600 -265
rect 12550 -315 12600 -285
rect 12550 -335 12565 -315
rect 12585 -335 12600 -315
rect 12550 -365 12600 -335
rect 12550 -385 12565 -365
rect 12585 -385 12600 -365
rect 12550 -415 12600 -385
rect 12550 -435 12565 -415
rect 12585 -435 12600 -415
rect 12550 -465 12600 -435
rect 12550 -485 12565 -465
rect 12585 -485 12600 -465
rect 12550 -515 12600 -485
rect 12550 -535 12565 -515
rect 12585 -535 12600 -515
rect 12550 -565 12600 -535
rect 12550 -585 12565 -565
rect 12585 -585 12600 -565
rect 12550 -615 12600 -585
rect 12550 -635 12565 -615
rect 12585 -635 12600 -615
rect 12550 -665 12600 -635
rect 12550 -685 12565 -665
rect 12585 -685 12600 -665
rect 12550 -715 12600 -685
rect 12550 -735 12565 -715
rect 12585 -735 12600 -715
rect 12550 -765 12600 -735
rect 12550 -785 12565 -765
rect 12585 -785 12600 -765
rect 12550 -800 12600 -785
rect 12850 -115 12900 -100
rect 12850 -135 12865 -115
rect 12885 -135 12900 -115
rect 12850 -165 12900 -135
rect 12850 -185 12865 -165
rect 12885 -185 12900 -165
rect 12850 -215 12900 -185
rect 12850 -235 12865 -215
rect 12885 -235 12900 -215
rect 12850 -265 12900 -235
rect 12850 -285 12865 -265
rect 12885 -285 12900 -265
rect 12850 -315 12900 -285
rect 12850 -335 12865 -315
rect 12885 -335 12900 -315
rect 12850 -365 12900 -335
rect 12850 -385 12865 -365
rect 12885 -385 12900 -365
rect 12850 -415 12900 -385
rect 12850 -435 12865 -415
rect 12885 -435 12900 -415
rect 12850 -465 12900 -435
rect 12850 -485 12865 -465
rect 12885 -485 12900 -465
rect 12850 -515 12900 -485
rect 12850 -535 12865 -515
rect 12885 -535 12900 -515
rect 12850 -565 12900 -535
rect 12850 -585 12865 -565
rect 12885 -585 12900 -565
rect 12850 -615 12900 -585
rect 12850 -635 12865 -615
rect 12885 -635 12900 -615
rect 12850 -665 12900 -635
rect 12850 -685 12865 -665
rect 12885 -685 12900 -665
rect 12850 -715 12900 -685
rect 12850 -735 12865 -715
rect 12885 -735 12900 -715
rect 12850 -765 12900 -735
rect 12850 -785 12865 -765
rect 12885 -785 12900 -765
rect 12850 -800 12900 -785
rect 13150 -115 13200 -100
rect 13150 -135 13165 -115
rect 13185 -135 13200 -115
rect 13150 -165 13200 -135
rect 13150 -185 13165 -165
rect 13185 -185 13200 -165
rect 13150 -215 13200 -185
rect 13150 -235 13165 -215
rect 13185 -235 13200 -215
rect 13150 -265 13200 -235
rect 13150 -285 13165 -265
rect 13185 -285 13200 -265
rect 13150 -315 13200 -285
rect 13150 -335 13165 -315
rect 13185 -335 13200 -315
rect 13150 -365 13200 -335
rect 13150 -385 13165 -365
rect 13185 -385 13200 -365
rect 13150 -415 13200 -385
rect 13150 -435 13165 -415
rect 13185 -435 13200 -415
rect 13150 -465 13200 -435
rect 13150 -485 13165 -465
rect 13185 -485 13200 -465
rect 13150 -515 13200 -485
rect 13150 -535 13165 -515
rect 13185 -535 13200 -515
rect 13150 -565 13200 -535
rect 13150 -585 13165 -565
rect 13185 -585 13200 -565
rect 13150 -615 13200 -585
rect 13150 -635 13165 -615
rect 13185 -635 13200 -615
rect 13150 -665 13200 -635
rect 13150 -685 13165 -665
rect 13185 -685 13200 -665
rect 13150 -715 13200 -685
rect 13150 -735 13165 -715
rect 13185 -735 13200 -715
rect 13150 -765 13200 -735
rect 13150 -785 13165 -765
rect 13185 -785 13200 -765
rect 13150 -800 13200 -785
rect 13450 -115 13500 -100
rect 13450 -135 13465 -115
rect 13485 -135 13500 -115
rect 13450 -165 13500 -135
rect 13450 -185 13465 -165
rect 13485 -185 13500 -165
rect 13450 -215 13500 -185
rect 13450 -235 13465 -215
rect 13485 -235 13500 -215
rect 13450 -265 13500 -235
rect 13450 -285 13465 -265
rect 13485 -285 13500 -265
rect 13450 -315 13500 -285
rect 13450 -335 13465 -315
rect 13485 -335 13500 -315
rect 13450 -365 13500 -335
rect 13450 -385 13465 -365
rect 13485 -385 13500 -365
rect 13450 -415 13500 -385
rect 13450 -435 13465 -415
rect 13485 -435 13500 -415
rect 13450 -465 13500 -435
rect 13450 -485 13465 -465
rect 13485 -485 13500 -465
rect 13450 -515 13500 -485
rect 13450 -535 13465 -515
rect 13485 -535 13500 -515
rect 13450 -565 13500 -535
rect 13450 -585 13465 -565
rect 13485 -585 13500 -565
rect 13450 -615 13500 -585
rect 13450 -635 13465 -615
rect 13485 -635 13500 -615
rect 13450 -665 13500 -635
rect 13450 -685 13465 -665
rect 13485 -685 13500 -665
rect 13450 -715 13500 -685
rect 13450 -735 13465 -715
rect 13485 -735 13500 -715
rect 13450 -765 13500 -735
rect 13450 -785 13465 -765
rect 13485 -785 13500 -765
rect 13450 -800 13500 -785
rect 13750 -115 13800 -100
rect 13750 -135 13765 -115
rect 13785 -135 13800 -115
rect 13750 -165 13800 -135
rect 13750 -185 13765 -165
rect 13785 -185 13800 -165
rect 13750 -215 13800 -185
rect 13750 -235 13765 -215
rect 13785 -235 13800 -215
rect 13750 -265 13800 -235
rect 13750 -285 13765 -265
rect 13785 -285 13800 -265
rect 13750 -315 13800 -285
rect 13750 -335 13765 -315
rect 13785 -335 13800 -315
rect 13750 -365 13800 -335
rect 13750 -385 13765 -365
rect 13785 -385 13800 -365
rect 13750 -415 13800 -385
rect 13750 -435 13765 -415
rect 13785 -435 13800 -415
rect 13750 -465 13800 -435
rect 13750 -485 13765 -465
rect 13785 -485 13800 -465
rect 13750 -515 13800 -485
rect 13750 -535 13765 -515
rect 13785 -535 13800 -515
rect 13750 -565 13800 -535
rect 13750 -585 13765 -565
rect 13785 -585 13800 -565
rect 13750 -615 13800 -585
rect 13750 -635 13765 -615
rect 13785 -635 13800 -615
rect 13750 -665 13800 -635
rect 13750 -685 13765 -665
rect 13785 -685 13800 -665
rect 13750 -715 13800 -685
rect 13750 -735 13765 -715
rect 13785 -735 13800 -715
rect 13750 -765 13800 -735
rect 13750 -785 13765 -765
rect 13785 -785 13800 -765
rect 13750 -800 13800 -785
rect 14050 -115 14100 -100
rect 14050 -135 14065 -115
rect 14085 -135 14100 -115
rect 14050 -165 14100 -135
rect 14050 -185 14065 -165
rect 14085 -185 14100 -165
rect 14050 -215 14100 -185
rect 14050 -235 14065 -215
rect 14085 -235 14100 -215
rect 14050 -265 14100 -235
rect 14050 -285 14065 -265
rect 14085 -285 14100 -265
rect 14050 -315 14100 -285
rect 14050 -335 14065 -315
rect 14085 -335 14100 -315
rect 14050 -365 14100 -335
rect 14050 -385 14065 -365
rect 14085 -385 14100 -365
rect 14050 -415 14100 -385
rect 14050 -435 14065 -415
rect 14085 -435 14100 -415
rect 14050 -465 14100 -435
rect 14050 -485 14065 -465
rect 14085 -485 14100 -465
rect 14050 -515 14100 -485
rect 14050 -535 14065 -515
rect 14085 -535 14100 -515
rect 14050 -565 14100 -535
rect 14050 -585 14065 -565
rect 14085 -585 14100 -565
rect 14050 -615 14100 -585
rect 14050 -635 14065 -615
rect 14085 -635 14100 -615
rect 14050 -665 14100 -635
rect 14050 -685 14065 -665
rect 14085 -685 14100 -665
rect 14050 -715 14100 -685
rect 14050 -735 14065 -715
rect 14085 -735 14100 -715
rect 14050 -765 14100 -735
rect 14050 -785 14065 -765
rect 14085 -785 14100 -765
rect 14050 -800 14100 -785
rect 14350 -115 14400 -100
rect 14350 -135 14365 -115
rect 14385 -135 14400 -115
rect 14350 -165 14400 -135
rect 14350 -185 14365 -165
rect 14385 -185 14400 -165
rect 14350 -215 14400 -185
rect 14350 -235 14365 -215
rect 14385 -235 14400 -215
rect 14350 -265 14400 -235
rect 14350 -285 14365 -265
rect 14385 -285 14400 -265
rect 14350 -315 14400 -285
rect 14350 -335 14365 -315
rect 14385 -335 14400 -315
rect 14350 -365 14400 -335
rect 14350 -385 14365 -365
rect 14385 -385 14400 -365
rect 14350 -415 14400 -385
rect 14350 -435 14365 -415
rect 14385 -435 14400 -415
rect 14350 -465 14400 -435
rect 14350 -485 14365 -465
rect 14385 -485 14400 -465
rect 14350 -515 14400 -485
rect 14350 -535 14365 -515
rect 14385 -535 14400 -515
rect 14350 -565 14400 -535
rect 14350 -585 14365 -565
rect 14385 -585 14400 -565
rect 14350 -615 14400 -585
rect 14350 -635 14365 -615
rect 14385 -635 14400 -615
rect 14350 -665 14400 -635
rect 14350 -685 14365 -665
rect 14385 -685 14400 -665
rect 14350 -715 14400 -685
rect 14350 -735 14365 -715
rect 14385 -735 14400 -715
rect 14350 -765 14400 -735
rect 14350 -785 14365 -765
rect 14385 -785 14400 -765
rect 14350 -800 14400 -785
rect 15550 -115 15600 -100
rect 15550 -135 15565 -115
rect 15585 -135 15600 -115
rect 15550 -165 15600 -135
rect 15550 -185 15565 -165
rect 15585 -185 15600 -165
rect 15550 -215 15600 -185
rect 15550 -235 15565 -215
rect 15585 -235 15600 -215
rect 15550 -265 15600 -235
rect 15550 -285 15565 -265
rect 15585 -285 15600 -265
rect 15550 -315 15600 -285
rect 15550 -335 15565 -315
rect 15585 -335 15600 -315
rect 15550 -365 15600 -335
rect 15550 -385 15565 -365
rect 15585 -385 15600 -365
rect 15550 -415 15600 -385
rect 15550 -435 15565 -415
rect 15585 -435 15600 -415
rect 15550 -465 15600 -435
rect 15550 -485 15565 -465
rect 15585 -485 15600 -465
rect 15550 -515 15600 -485
rect 15550 -535 15565 -515
rect 15585 -535 15600 -515
rect 15550 -565 15600 -535
rect 15550 -585 15565 -565
rect 15585 -585 15600 -565
rect 15550 -615 15600 -585
rect 15550 -635 15565 -615
rect 15585 -635 15600 -615
rect 15550 -665 15600 -635
rect 15550 -685 15565 -665
rect 15585 -685 15600 -665
rect 15550 -715 15600 -685
rect 15550 -735 15565 -715
rect 15585 -735 15600 -715
rect 15550 -765 15600 -735
rect 15550 -785 15565 -765
rect 15585 -785 15600 -765
rect 15550 -800 15600 -785
rect 16750 -115 16800 -100
rect 16750 -135 16765 -115
rect 16785 -135 16800 -115
rect 16750 -165 16800 -135
rect 16750 -185 16765 -165
rect 16785 -185 16800 -165
rect 16750 -215 16800 -185
rect 16750 -235 16765 -215
rect 16785 -235 16800 -215
rect 16750 -265 16800 -235
rect 16750 -285 16765 -265
rect 16785 -285 16800 -265
rect 16750 -315 16800 -285
rect 16750 -335 16765 -315
rect 16785 -335 16800 -315
rect 16750 -365 16800 -335
rect 16750 -385 16765 -365
rect 16785 -385 16800 -365
rect 16750 -415 16800 -385
rect 16750 -435 16765 -415
rect 16785 -435 16800 -415
rect 16750 -465 16800 -435
rect 16750 -485 16765 -465
rect 16785 -485 16800 -465
rect 16750 -515 16800 -485
rect 16750 -535 16765 -515
rect 16785 -535 16800 -515
rect 16750 -565 16800 -535
rect 16750 -585 16765 -565
rect 16785 -585 16800 -565
rect 16750 -615 16800 -585
rect 16750 -635 16765 -615
rect 16785 -635 16800 -615
rect 16750 -665 16800 -635
rect 16750 -685 16765 -665
rect 16785 -685 16800 -665
rect 16750 -715 16800 -685
rect 16750 -735 16765 -715
rect 16785 -735 16800 -715
rect 16750 -765 16800 -735
rect 16750 -785 16765 -765
rect 16785 -785 16800 -765
rect 16750 -800 16800 -785
rect 17950 -115 18000 -100
rect 17950 -135 17965 -115
rect 17985 -135 18000 -115
rect 17950 -165 18000 -135
rect 17950 -185 17965 -165
rect 17985 -185 18000 -165
rect 17950 -215 18000 -185
rect 17950 -235 17965 -215
rect 17985 -235 18000 -215
rect 17950 -265 18000 -235
rect 17950 -285 17965 -265
rect 17985 -285 18000 -265
rect 17950 -315 18000 -285
rect 17950 -335 17965 -315
rect 17985 -335 18000 -315
rect 17950 -365 18000 -335
rect 17950 -385 17965 -365
rect 17985 -385 18000 -365
rect 17950 -415 18000 -385
rect 17950 -435 17965 -415
rect 17985 -435 18000 -415
rect 17950 -465 18000 -435
rect 17950 -485 17965 -465
rect 17985 -485 18000 -465
rect 17950 -515 18000 -485
rect 17950 -535 17965 -515
rect 17985 -535 18000 -515
rect 17950 -565 18000 -535
rect 17950 -585 17965 -565
rect 17985 -585 18000 -565
rect 17950 -615 18000 -585
rect 17950 -635 17965 -615
rect 17985 -635 18000 -615
rect 17950 -665 18000 -635
rect 17950 -685 17965 -665
rect 17985 -685 18000 -665
rect 17950 -715 18000 -685
rect 17950 -735 17965 -715
rect 17985 -735 18000 -715
rect 17950 -765 18000 -735
rect 17950 -785 17965 -765
rect 17985 -785 18000 -765
rect 17950 -800 18000 -785
rect 19150 -115 19200 -100
rect 19150 -135 19165 -115
rect 19185 -135 19200 -115
rect 19150 -165 19200 -135
rect 19150 -185 19165 -165
rect 19185 -185 19200 -165
rect 19150 -215 19200 -185
rect 19150 -235 19165 -215
rect 19185 -235 19200 -215
rect 19150 -265 19200 -235
rect 19150 -285 19165 -265
rect 19185 -285 19200 -265
rect 19150 -315 19200 -285
rect 19150 -335 19165 -315
rect 19185 -335 19200 -315
rect 19150 -365 19200 -335
rect 19150 -385 19165 -365
rect 19185 -385 19200 -365
rect 19150 -415 19200 -385
rect 19150 -435 19165 -415
rect 19185 -435 19200 -415
rect 19150 -465 19200 -435
rect 19150 -485 19165 -465
rect 19185 -485 19200 -465
rect 19150 -515 19200 -485
rect 19150 -535 19165 -515
rect 19185 -535 19200 -515
rect 19150 -565 19200 -535
rect 19150 -585 19165 -565
rect 19185 -585 19200 -565
rect 19150 -615 19200 -585
rect 19150 -635 19165 -615
rect 19185 -635 19200 -615
rect 19150 -665 19200 -635
rect 19150 -685 19165 -665
rect 19185 -685 19200 -665
rect 19150 -715 19200 -685
rect 19150 -735 19165 -715
rect 19185 -735 19200 -715
rect 19150 -765 19200 -735
rect 19150 -785 19165 -765
rect 19185 -785 19200 -765
rect 19150 -800 19200 -785
rect 20350 -115 20400 -100
rect 20350 -135 20365 -115
rect 20385 -135 20400 -115
rect 20350 -165 20400 -135
rect 20350 -185 20365 -165
rect 20385 -185 20400 -165
rect 20350 -215 20400 -185
rect 20350 -235 20365 -215
rect 20385 -235 20400 -215
rect 20350 -265 20400 -235
rect 20350 -285 20365 -265
rect 20385 -285 20400 -265
rect 20350 -315 20400 -285
rect 20350 -335 20365 -315
rect 20385 -335 20400 -315
rect 20350 -365 20400 -335
rect 20350 -385 20365 -365
rect 20385 -385 20400 -365
rect 20350 -415 20400 -385
rect 20350 -435 20365 -415
rect 20385 -435 20400 -415
rect 20350 -465 20400 -435
rect 20350 -485 20365 -465
rect 20385 -485 20400 -465
rect 20350 -515 20400 -485
rect 20350 -535 20365 -515
rect 20385 -535 20400 -515
rect 20350 -565 20400 -535
rect 20350 -585 20365 -565
rect 20385 -585 20400 -565
rect 20350 -615 20400 -585
rect 20350 -635 20365 -615
rect 20385 -635 20400 -615
rect 20350 -665 20400 -635
rect 20350 -685 20365 -665
rect 20385 -685 20400 -665
rect 20350 -715 20400 -685
rect 20350 -735 20365 -715
rect 20385 -735 20400 -715
rect 20350 -765 20400 -735
rect 20350 -785 20365 -765
rect 20385 -785 20400 -765
rect 20350 -800 20400 -785
rect -600 -865 -350 -850
rect -600 -885 -585 -865
rect -565 -885 -535 -865
rect -515 -885 -485 -865
rect -465 -885 -435 -865
rect -415 -885 -385 -865
rect -365 -885 -350 -865
rect -600 -900 -350 -885
rect -300 -865 -50 -850
rect -300 -885 -285 -865
rect -265 -885 -235 -865
rect -215 -885 -185 -865
rect -165 -885 -135 -865
rect -115 -885 -85 -865
rect -65 -885 -50 -865
rect -300 -900 -50 -885
rect 0 -865 250 -850
rect 0 -885 15 -865
rect 35 -885 65 -865
rect 85 -885 115 -865
rect 135 -885 165 -865
rect 185 -885 215 -865
rect 235 -885 250 -865
rect 0 -900 250 -885
rect 300 -865 550 -850
rect 300 -885 315 -865
rect 335 -885 365 -865
rect 385 -885 415 -865
rect 435 -885 465 -865
rect 485 -885 515 -865
rect 535 -885 550 -865
rect 300 -900 550 -885
rect 600 -865 850 -850
rect 600 -885 615 -865
rect 635 -885 665 -865
rect 685 -885 715 -865
rect 735 -885 765 -865
rect 785 -885 815 -865
rect 835 -885 850 -865
rect 600 -900 850 -885
rect 900 -865 1150 -850
rect 900 -885 915 -865
rect 935 -885 965 -865
rect 985 -885 1015 -865
rect 1035 -885 1065 -865
rect 1085 -885 1115 -865
rect 1135 -885 1150 -865
rect 900 -900 1150 -885
rect 1200 -865 1450 -850
rect 1200 -885 1215 -865
rect 1235 -885 1265 -865
rect 1285 -885 1315 -865
rect 1335 -885 1365 -865
rect 1385 -885 1415 -865
rect 1435 -885 1450 -865
rect 1200 -900 1450 -885
rect 1500 -865 1750 -850
rect 1500 -885 1515 -865
rect 1535 -885 1565 -865
rect 1585 -885 1615 -865
rect 1635 -885 1665 -865
rect 1685 -885 1715 -865
rect 1735 -885 1750 -865
rect 1500 -900 1750 -885
rect 1800 -865 2050 -850
rect 1800 -885 1815 -865
rect 1835 -885 1865 -865
rect 1885 -885 1915 -865
rect 1935 -885 1965 -865
rect 1985 -885 2015 -865
rect 2035 -885 2050 -865
rect 1800 -900 2050 -885
rect 2100 -865 2350 -850
rect 2100 -885 2115 -865
rect 2135 -885 2165 -865
rect 2185 -885 2215 -865
rect 2235 -885 2265 -865
rect 2285 -885 2315 -865
rect 2335 -885 2350 -865
rect 2100 -900 2350 -885
rect 2400 -865 2650 -850
rect 2400 -885 2415 -865
rect 2435 -885 2465 -865
rect 2485 -885 2515 -865
rect 2535 -885 2565 -865
rect 2585 -885 2615 -865
rect 2635 -885 2650 -865
rect 2400 -900 2650 -885
rect 2700 -865 2950 -850
rect 2700 -885 2715 -865
rect 2735 -885 2765 -865
rect 2785 -885 2815 -865
rect 2835 -885 2865 -865
rect 2885 -885 2915 -865
rect 2935 -885 2950 -865
rect 2700 -900 2950 -885
rect 3000 -865 3250 -850
rect 3000 -885 3015 -865
rect 3035 -885 3065 -865
rect 3085 -885 3115 -865
rect 3135 -885 3165 -865
rect 3185 -885 3215 -865
rect 3235 -885 3250 -865
rect 3000 -900 3250 -885
rect 3300 -865 3550 -850
rect 3300 -885 3315 -865
rect 3335 -885 3365 -865
rect 3385 -885 3415 -865
rect 3435 -885 3465 -865
rect 3485 -885 3515 -865
rect 3535 -885 3550 -865
rect 3300 -900 3550 -885
rect 3600 -865 3850 -850
rect 3600 -885 3615 -865
rect 3635 -885 3665 -865
rect 3685 -885 3715 -865
rect 3735 -885 3765 -865
rect 3785 -885 3815 -865
rect 3835 -885 3850 -865
rect 3600 -900 3850 -885
rect 3900 -865 4150 -850
rect 3900 -885 3915 -865
rect 3935 -885 3965 -865
rect 3985 -885 4015 -865
rect 4035 -885 4065 -865
rect 4085 -885 4115 -865
rect 4135 -885 4150 -865
rect 3900 -900 4150 -885
rect 4200 -865 4450 -850
rect 4200 -885 4215 -865
rect 4235 -885 4265 -865
rect 4285 -885 4315 -865
rect 4335 -885 4365 -865
rect 4385 -885 4415 -865
rect 4435 -885 4450 -865
rect 4200 -900 4450 -885
rect 4500 -865 4750 -850
rect 4500 -885 4515 -865
rect 4535 -885 4565 -865
rect 4585 -885 4615 -865
rect 4635 -885 4665 -865
rect 4685 -885 4715 -865
rect 4735 -885 4750 -865
rect 4500 -900 4750 -885
rect 4800 -865 5050 -850
rect 4800 -885 4815 -865
rect 4835 -885 4865 -865
rect 4885 -885 4915 -865
rect 4935 -885 4965 -865
rect 4985 -885 5015 -865
rect 5035 -885 5050 -865
rect 4800 -900 5050 -885
rect 5100 -865 5350 -850
rect 5100 -885 5115 -865
rect 5135 -885 5165 -865
rect 5185 -885 5215 -865
rect 5235 -885 5265 -865
rect 5285 -885 5315 -865
rect 5335 -885 5350 -865
rect 5100 -900 5350 -885
rect 5400 -865 5650 -850
rect 5400 -885 5415 -865
rect 5435 -885 5465 -865
rect 5485 -885 5515 -865
rect 5535 -885 5565 -865
rect 5585 -885 5615 -865
rect 5635 -885 5650 -865
rect 5400 -900 5650 -885
rect 5700 -865 5950 -850
rect 5700 -885 5715 -865
rect 5735 -885 5765 -865
rect 5785 -885 5815 -865
rect 5835 -885 5865 -865
rect 5885 -885 5915 -865
rect 5935 -885 5950 -865
rect 5700 -900 5950 -885
rect 6000 -865 6250 -850
rect 6000 -885 6015 -865
rect 6035 -885 6065 -865
rect 6085 -885 6115 -865
rect 6135 -885 6165 -865
rect 6185 -885 6215 -865
rect 6235 -885 6250 -865
rect 6000 -900 6250 -885
rect 6300 -865 6550 -850
rect 6300 -885 6315 -865
rect 6335 -885 6365 -865
rect 6385 -885 6415 -865
rect 6435 -885 6465 -865
rect 6485 -885 6515 -865
rect 6535 -885 6550 -865
rect 6300 -900 6550 -885
rect 6600 -865 6850 -850
rect 6600 -885 6615 -865
rect 6635 -885 6665 -865
rect 6685 -885 6715 -865
rect 6735 -885 6765 -865
rect 6785 -885 6815 -865
rect 6835 -885 6850 -865
rect 6600 -900 6850 -885
rect 6900 -865 7150 -850
rect 6900 -885 6915 -865
rect 6935 -885 6965 -865
rect 6985 -885 7015 -865
rect 7035 -885 7065 -865
rect 7085 -885 7115 -865
rect 7135 -885 7150 -865
rect 6900 -900 7150 -885
rect 7200 -865 7450 -850
rect 7200 -885 7215 -865
rect 7235 -885 7265 -865
rect 7285 -885 7315 -865
rect 7335 -885 7365 -865
rect 7385 -885 7415 -865
rect 7435 -885 7450 -865
rect 7200 -900 7450 -885
rect 7500 -865 7750 -850
rect 7500 -885 7515 -865
rect 7535 -885 7565 -865
rect 7585 -885 7615 -865
rect 7635 -885 7665 -865
rect 7685 -885 7715 -865
rect 7735 -885 7750 -865
rect 7500 -900 7750 -885
rect 7800 -865 8050 -850
rect 7800 -885 7815 -865
rect 7835 -885 7865 -865
rect 7885 -885 7915 -865
rect 7935 -885 7965 -865
rect 7985 -885 8015 -865
rect 8035 -885 8050 -865
rect 7800 -900 8050 -885
rect 8100 -865 8350 -850
rect 8100 -885 8115 -865
rect 8135 -885 8165 -865
rect 8185 -885 8215 -865
rect 8235 -885 8265 -865
rect 8285 -885 8315 -865
rect 8335 -885 8350 -865
rect 8100 -900 8350 -885
rect 8400 -865 8650 -850
rect 8400 -885 8415 -865
rect 8435 -885 8465 -865
rect 8485 -885 8515 -865
rect 8535 -885 8565 -865
rect 8585 -885 8615 -865
rect 8635 -885 8650 -865
rect 8400 -900 8650 -885
rect 8700 -865 8950 -850
rect 8700 -885 8715 -865
rect 8735 -885 8765 -865
rect 8785 -885 8815 -865
rect 8835 -885 8865 -865
rect 8885 -885 8915 -865
rect 8935 -885 8950 -865
rect 8700 -900 8950 -885
rect 9000 -865 9250 -850
rect 9000 -885 9015 -865
rect 9035 -885 9065 -865
rect 9085 -885 9115 -865
rect 9135 -885 9165 -865
rect 9185 -885 9215 -865
rect 9235 -885 9250 -865
rect 9000 -900 9250 -885
rect 9300 -865 9550 -850
rect 9300 -885 9315 -865
rect 9335 -885 9365 -865
rect 9385 -885 9415 -865
rect 9435 -885 9465 -865
rect 9485 -885 9515 -865
rect 9535 -885 9550 -865
rect 9300 -900 9550 -885
rect 9600 -865 9850 -850
rect 9600 -885 9615 -865
rect 9635 -885 9665 -865
rect 9685 -885 9715 -865
rect 9735 -885 9765 -865
rect 9785 -885 9815 -865
rect 9835 -885 9850 -865
rect 9600 -900 9850 -885
rect 9900 -865 10150 -850
rect 9900 -885 9915 -865
rect 9935 -885 9965 -865
rect 9985 -885 10015 -865
rect 10035 -885 10065 -865
rect 10085 -885 10115 -865
rect 10135 -885 10150 -865
rect 9900 -900 10150 -885
rect 10200 -865 10450 -850
rect 10200 -885 10215 -865
rect 10235 -885 10265 -865
rect 10285 -885 10315 -865
rect 10335 -885 10365 -865
rect 10385 -885 10415 -865
rect 10435 -885 10450 -865
rect 10200 -900 10450 -885
rect 10500 -865 10750 -850
rect 10500 -885 10515 -865
rect 10535 -885 10565 -865
rect 10585 -885 10615 -865
rect 10635 -885 10665 -865
rect 10685 -885 10715 -865
rect 10735 -885 10750 -865
rect 10500 -900 10750 -885
rect 10800 -865 11050 -850
rect 10800 -885 10815 -865
rect 10835 -885 10865 -865
rect 10885 -885 10915 -865
rect 10935 -885 10965 -865
rect 10985 -885 11015 -865
rect 11035 -885 11050 -865
rect 10800 -900 11050 -885
rect 11100 -865 11350 -850
rect 11100 -885 11115 -865
rect 11135 -885 11165 -865
rect 11185 -885 11215 -865
rect 11235 -885 11265 -865
rect 11285 -885 11315 -865
rect 11335 -885 11350 -865
rect 11100 -900 11350 -885
rect 11400 -865 11650 -850
rect 11400 -885 11415 -865
rect 11435 -885 11465 -865
rect 11485 -885 11515 -865
rect 11535 -885 11565 -865
rect 11585 -885 11615 -865
rect 11635 -885 11650 -865
rect 11400 -900 11650 -885
rect 11700 -865 11950 -850
rect 11700 -885 11715 -865
rect 11735 -885 11765 -865
rect 11785 -885 11815 -865
rect 11835 -885 11865 -865
rect 11885 -885 11915 -865
rect 11935 -885 11950 -865
rect 11700 -900 11950 -885
rect 12000 -865 12250 -850
rect 12000 -885 12015 -865
rect 12035 -885 12065 -865
rect 12085 -885 12115 -865
rect 12135 -885 12165 -865
rect 12185 -885 12215 -865
rect 12235 -885 12250 -865
rect 12000 -900 12250 -885
rect 12300 -865 12550 -850
rect 12300 -885 12315 -865
rect 12335 -885 12365 -865
rect 12385 -885 12415 -865
rect 12435 -885 12465 -865
rect 12485 -885 12515 -865
rect 12535 -885 12550 -865
rect 12300 -900 12550 -885
rect 12600 -865 12850 -850
rect 12600 -885 12615 -865
rect 12635 -885 12665 -865
rect 12685 -885 12715 -865
rect 12735 -885 12765 -865
rect 12785 -885 12815 -865
rect 12835 -885 12850 -865
rect 12600 -900 12850 -885
rect 12900 -865 13150 -850
rect 12900 -885 12915 -865
rect 12935 -885 12965 -865
rect 12985 -885 13015 -865
rect 13035 -885 13065 -865
rect 13085 -885 13115 -865
rect 13135 -885 13150 -865
rect 12900 -900 13150 -885
rect 13200 -865 13450 -850
rect 13200 -885 13215 -865
rect 13235 -885 13265 -865
rect 13285 -885 13315 -865
rect 13335 -885 13365 -865
rect 13385 -885 13415 -865
rect 13435 -885 13450 -865
rect 13200 -900 13450 -885
rect 13500 -865 13750 -850
rect 13500 -885 13515 -865
rect 13535 -885 13565 -865
rect 13585 -885 13615 -865
rect 13635 -885 13665 -865
rect 13685 -885 13715 -865
rect 13735 -885 13750 -865
rect 13500 -900 13750 -885
rect 13800 -865 14050 -850
rect 13800 -885 13815 -865
rect 13835 -885 13865 -865
rect 13885 -885 13915 -865
rect 13935 -885 13965 -865
rect 13985 -885 14015 -865
rect 14035 -885 14050 -865
rect 13800 -900 14050 -885
rect 14100 -865 14350 -850
rect 14100 -885 14115 -865
rect 14135 -885 14165 -865
rect 14185 -885 14215 -865
rect 14235 -885 14265 -865
rect 14285 -885 14315 -865
rect 14335 -885 14350 -865
rect 14100 -900 14350 -885
rect 14400 -865 14650 -850
rect 14400 -885 14415 -865
rect 14435 -885 14465 -865
rect 14485 -885 14515 -865
rect 14535 -885 14565 -865
rect 14585 -885 14615 -865
rect 14635 -885 14650 -865
rect 14400 -900 14650 -885
rect 14700 -865 14950 -850
rect 14700 -885 14715 -865
rect 14735 -885 14765 -865
rect 14785 -885 14815 -865
rect 14835 -885 14865 -865
rect 14885 -885 14915 -865
rect 14935 -885 14950 -865
rect 14700 -900 14950 -885
rect 15000 -865 15250 -850
rect 15000 -885 15015 -865
rect 15035 -885 15065 -865
rect 15085 -885 15115 -865
rect 15135 -885 15165 -865
rect 15185 -885 15215 -865
rect 15235 -885 15250 -865
rect 15000 -900 15250 -885
rect 15300 -865 15550 -850
rect 15300 -885 15315 -865
rect 15335 -885 15365 -865
rect 15385 -885 15415 -865
rect 15435 -885 15465 -865
rect 15485 -885 15515 -865
rect 15535 -885 15550 -865
rect 15300 -900 15550 -885
rect 15600 -865 15850 -850
rect 15600 -885 15615 -865
rect 15635 -885 15665 -865
rect 15685 -885 15715 -865
rect 15735 -885 15765 -865
rect 15785 -885 15815 -865
rect 15835 -885 15850 -865
rect 15600 -900 15850 -885
rect 15900 -865 16150 -850
rect 15900 -885 15915 -865
rect 15935 -885 15965 -865
rect 15985 -885 16015 -865
rect 16035 -885 16065 -865
rect 16085 -885 16115 -865
rect 16135 -885 16150 -865
rect 15900 -900 16150 -885
rect 16200 -865 16450 -850
rect 16200 -885 16215 -865
rect 16235 -885 16265 -865
rect 16285 -885 16315 -865
rect 16335 -885 16365 -865
rect 16385 -885 16415 -865
rect 16435 -885 16450 -865
rect 16200 -900 16450 -885
rect 16500 -865 16750 -850
rect 16500 -885 16515 -865
rect 16535 -885 16565 -865
rect 16585 -885 16615 -865
rect 16635 -885 16665 -865
rect 16685 -885 16715 -865
rect 16735 -885 16750 -865
rect 16500 -900 16750 -885
rect 16800 -865 17050 -850
rect 16800 -885 16815 -865
rect 16835 -885 16865 -865
rect 16885 -885 16915 -865
rect 16935 -885 16965 -865
rect 16985 -885 17015 -865
rect 17035 -885 17050 -865
rect 16800 -900 17050 -885
rect 17100 -865 17350 -850
rect 17100 -885 17115 -865
rect 17135 -885 17165 -865
rect 17185 -885 17215 -865
rect 17235 -885 17265 -865
rect 17285 -885 17315 -865
rect 17335 -885 17350 -865
rect 17100 -900 17350 -885
rect 17400 -865 17650 -850
rect 17400 -885 17415 -865
rect 17435 -885 17465 -865
rect 17485 -885 17515 -865
rect 17535 -885 17565 -865
rect 17585 -885 17615 -865
rect 17635 -885 17650 -865
rect 17400 -900 17650 -885
rect 17700 -865 17950 -850
rect 17700 -885 17715 -865
rect 17735 -885 17765 -865
rect 17785 -885 17815 -865
rect 17835 -885 17865 -865
rect 17885 -885 17915 -865
rect 17935 -885 17950 -865
rect 17700 -900 17950 -885
rect 18000 -865 18250 -850
rect 18000 -885 18015 -865
rect 18035 -885 18065 -865
rect 18085 -885 18115 -865
rect 18135 -885 18165 -865
rect 18185 -885 18215 -865
rect 18235 -885 18250 -865
rect 18000 -900 18250 -885
rect 18300 -865 18550 -850
rect 18300 -885 18315 -865
rect 18335 -885 18365 -865
rect 18385 -885 18415 -865
rect 18435 -885 18465 -865
rect 18485 -885 18515 -865
rect 18535 -885 18550 -865
rect 18300 -900 18550 -885
rect 18600 -865 18850 -850
rect 18600 -885 18615 -865
rect 18635 -885 18665 -865
rect 18685 -885 18715 -865
rect 18735 -885 18765 -865
rect 18785 -885 18815 -865
rect 18835 -885 18850 -865
rect 18600 -900 18850 -885
rect 18900 -865 19150 -850
rect 18900 -885 18915 -865
rect 18935 -885 18965 -865
rect 18985 -885 19015 -865
rect 19035 -885 19065 -865
rect 19085 -885 19115 -865
rect 19135 -885 19150 -865
rect 18900 -900 19150 -885
rect 19200 -865 19450 -850
rect 19200 -885 19215 -865
rect 19235 -885 19265 -865
rect 19285 -885 19315 -865
rect 19335 -885 19365 -865
rect 19385 -885 19415 -865
rect 19435 -885 19450 -865
rect 19200 -900 19450 -885
rect 19500 -865 19750 -850
rect 19500 -885 19515 -865
rect 19535 -885 19565 -865
rect 19585 -885 19615 -865
rect 19635 -885 19665 -865
rect 19685 -885 19715 -865
rect 19735 -885 19750 -865
rect 19500 -900 19750 -885
rect 19800 -865 20050 -850
rect 19800 -885 19815 -865
rect 19835 -885 19865 -865
rect 19885 -885 19915 -865
rect 19935 -885 19965 -865
rect 19985 -885 20015 -865
rect 20035 -885 20050 -865
rect 19800 -900 20050 -885
rect 20100 -865 20350 -850
rect 20100 -885 20115 -865
rect 20135 -885 20165 -865
rect 20185 -885 20215 -865
rect 20235 -885 20265 -865
rect 20285 -885 20315 -865
rect 20335 -885 20350 -865
rect 20100 -900 20350 -885
rect -650 -965 -600 -950
rect -650 -985 -635 -965
rect -615 -985 -600 -965
rect -650 -1015 -600 -985
rect -650 -1035 -635 -1015
rect -615 -1035 -600 -1015
rect -650 -1065 -600 -1035
rect -650 -1085 -635 -1065
rect -615 -1085 -600 -1065
rect -650 -1115 -600 -1085
rect -650 -1135 -635 -1115
rect -615 -1135 -600 -1115
rect -650 -1165 -600 -1135
rect -650 -1185 -635 -1165
rect -615 -1185 -600 -1165
rect -650 -1215 -600 -1185
rect -650 -1235 -635 -1215
rect -615 -1235 -600 -1215
rect -650 -1265 -600 -1235
rect -650 -1285 -635 -1265
rect -615 -1285 -600 -1265
rect -650 -1315 -600 -1285
rect -650 -1335 -635 -1315
rect -615 -1335 -600 -1315
rect -650 -1365 -600 -1335
rect -650 -1385 -635 -1365
rect -615 -1385 -600 -1365
rect -650 -1415 -600 -1385
rect -650 -1435 -635 -1415
rect -615 -1435 -600 -1415
rect -650 -1465 -600 -1435
rect -650 -1485 -635 -1465
rect -615 -1485 -600 -1465
rect -650 -1515 -600 -1485
rect -650 -1535 -635 -1515
rect -615 -1535 -600 -1515
rect -650 -1565 -600 -1535
rect -650 -1585 -635 -1565
rect -615 -1585 -600 -1565
rect -650 -1615 -600 -1585
rect -650 -1635 -635 -1615
rect -615 -1635 -600 -1615
rect -650 -1650 -600 -1635
rect -500 -965 -450 -950
rect -500 -985 -485 -965
rect -465 -985 -450 -965
rect -500 -1015 -450 -985
rect -500 -1035 -485 -1015
rect -465 -1035 -450 -1015
rect -500 -1065 -450 -1035
rect -500 -1085 -485 -1065
rect -465 -1085 -450 -1065
rect -500 -1115 -450 -1085
rect -500 -1135 -485 -1115
rect -465 -1135 -450 -1115
rect -500 -1165 -450 -1135
rect -500 -1185 -485 -1165
rect -465 -1185 -450 -1165
rect -500 -1215 -450 -1185
rect -500 -1235 -485 -1215
rect -465 -1235 -450 -1215
rect -500 -1265 -450 -1235
rect -500 -1285 -485 -1265
rect -465 -1285 -450 -1265
rect -500 -1315 -450 -1285
rect -500 -1335 -485 -1315
rect -465 -1335 -450 -1315
rect -500 -1365 -450 -1335
rect -500 -1385 -485 -1365
rect -465 -1385 -450 -1365
rect -500 -1415 -450 -1385
rect -500 -1435 -485 -1415
rect -465 -1435 -450 -1415
rect -500 -1465 -450 -1435
rect -500 -1485 -485 -1465
rect -465 -1485 -450 -1465
rect -500 -1515 -450 -1485
rect -500 -1535 -485 -1515
rect -465 -1535 -450 -1515
rect -500 -1565 -450 -1535
rect -500 -1585 -485 -1565
rect -465 -1585 -450 -1565
rect -500 -1615 -450 -1585
rect -500 -1635 -485 -1615
rect -465 -1635 -450 -1615
rect -500 -1650 -450 -1635
rect -350 -965 -300 -950
rect -350 -985 -335 -965
rect -315 -985 -300 -965
rect -350 -1015 -300 -985
rect -350 -1035 -335 -1015
rect -315 -1035 -300 -1015
rect -350 -1065 -300 -1035
rect -350 -1085 -335 -1065
rect -315 -1085 -300 -1065
rect -350 -1115 -300 -1085
rect -350 -1135 -335 -1115
rect -315 -1135 -300 -1115
rect -350 -1165 -300 -1135
rect -350 -1185 -335 -1165
rect -315 -1185 -300 -1165
rect -350 -1215 -300 -1185
rect -350 -1235 -335 -1215
rect -315 -1235 -300 -1215
rect -350 -1265 -300 -1235
rect -350 -1285 -335 -1265
rect -315 -1285 -300 -1265
rect -350 -1315 -300 -1285
rect -350 -1335 -335 -1315
rect -315 -1335 -300 -1315
rect -350 -1365 -300 -1335
rect -350 -1385 -335 -1365
rect -315 -1385 -300 -1365
rect -350 -1415 -300 -1385
rect -350 -1435 -335 -1415
rect -315 -1435 -300 -1415
rect -350 -1465 -300 -1435
rect -350 -1485 -335 -1465
rect -315 -1485 -300 -1465
rect -350 -1515 -300 -1485
rect -350 -1535 -335 -1515
rect -315 -1535 -300 -1515
rect -350 -1565 -300 -1535
rect -350 -1585 -335 -1565
rect -315 -1585 -300 -1565
rect -350 -1615 -300 -1585
rect -350 -1635 -335 -1615
rect -315 -1635 -300 -1615
rect -350 -1650 -300 -1635
rect -200 -965 -150 -950
rect -200 -985 -185 -965
rect -165 -985 -150 -965
rect -200 -1015 -150 -985
rect -200 -1035 -185 -1015
rect -165 -1035 -150 -1015
rect -200 -1065 -150 -1035
rect -200 -1085 -185 -1065
rect -165 -1085 -150 -1065
rect -200 -1115 -150 -1085
rect -200 -1135 -185 -1115
rect -165 -1135 -150 -1115
rect -200 -1165 -150 -1135
rect -200 -1185 -185 -1165
rect -165 -1185 -150 -1165
rect -200 -1215 -150 -1185
rect -200 -1235 -185 -1215
rect -165 -1235 -150 -1215
rect -200 -1265 -150 -1235
rect -200 -1285 -185 -1265
rect -165 -1285 -150 -1265
rect -200 -1315 -150 -1285
rect -200 -1335 -185 -1315
rect -165 -1335 -150 -1315
rect -200 -1365 -150 -1335
rect -200 -1385 -185 -1365
rect -165 -1385 -150 -1365
rect -200 -1415 -150 -1385
rect -200 -1435 -185 -1415
rect -165 -1435 -150 -1415
rect -200 -1465 -150 -1435
rect -200 -1485 -185 -1465
rect -165 -1485 -150 -1465
rect -200 -1515 -150 -1485
rect -200 -1535 -185 -1515
rect -165 -1535 -150 -1515
rect -200 -1565 -150 -1535
rect -200 -1585 -185 -1565
rect -165 -1585 -150 -1565
rect -200 -1615 -150 -1585
rect -200 -1635 -185 -1615
rect -165 -1635 -150 -1615
rect -200 -1650 -150 -1635
rect -50 -965 0 -950
rect -50 -985 -35 -965
rect -15 -985 0 -965
rect -50 -1015 0 -985
rect -50 -1035 -35 -1015
rect -15 -1035 0 -1015
rect -50 -1065 0 -1035
rect -50 -1085 -35 -1065
rect -15 -1085 0 -1065
rect -50 -1115 0 -1085
rect -50 -1135 -35 -1115
rect -15 -1135 0 -1115
rect -50 -1165 0 -1135
rect -50 -1185 -35 -1165
rect -15 -1185 0 -1165
rect -50 -1215 0 -1185
rect -50 -1235 -35 -1215
rect -15 -1235 0 -1215
rect -50 -1265 0 -1235
rect -50 -1285 -35 -1265
rect -15 -1285 0 -1265
rect -50 -1315 0 -1285
rect -50 -1335 -35 -1315
rect -15 -1335 0 -1315
rect -50 -1365 0 -1335
rect -50 -1385 -35 -1365
rect -15 -1385 0 -1365
rect -50 -1415 0 -1385
rect -50 -1435 -35 -1415
rect -15 -1435 0 -1415
rect -50 -1465 0 -1435
rect -50 -1485 -35 -1465
rect -15 -1485 0 -1465
rect -50 -1515 0 -1485
rect -50 -1535 -35 -1515
rect -15 -1535 0 -1515
rect -50 -1565 0 -1535
rect -50 -1585 -35 -1565
rect -15 -1585 0 -1565
rect -50 -1615 0 -1585
rect -50 -1635 -35 -1615
rect -15 -1635 0 -1615
rect -50 -1650 0 -1635
rect 1150 -965 1200 -950
rect 1150 -985 1165 -965
rect 1185 -985 1200 -965
rect 1150 -1015 1200 -985
rect 1150 -1035 1165 -1015
rect 1185 -1035 1200 -1015
rect 1150 -1065 1200 -1035
rect 1150 -1085 1165 -1065
rect 1185 -1085 1200 -1065
rect 1150 -1115 1200 -1085
rect 1150 -1135 1165 -1115
rect 1185 -1135 1200 -1115
rect 1150 -1165 1200 -1135
rect 1150 -1185 1165 -1165
rect 1185 -1185 1200 -1165
rect 1150 -1215 1200 -1185
rect 1150 -1235 1165 -1215
rect 1185 -1235 1200 -1215
rect 1150 -1265 1200 -1235
rect 1150 -1285 1165 -1265
rect 1185 -1285 1200 -1265
rect 1150 -1315 1200 -1285
rect 1150 -1335 1165 -1315
rect 1185 -1335 1200 -1315
rect 1150 -1365 1200 -1335
rect 1150 -1385 1165 -1365
rect 1185 -1385 1200 -1365
rect 1150 -1415 1200 -1385
rect 1150 -1435 1165 -1415
rect 1185 -1435 1200 -1415
rect 1150 -1465 1200 -1435
rect 1150 -1485 1165 -1465
rect 1185 -1485 1200 -1465
rect 1150 -1515 1200 -1485
rect 1150 -1535 1165 -1515
rect 1185 -1535 1200 -1515
rect 1150 -1565 1200 -1535
rect 1150 -1585 1165 -1565
rect 1185 -1585 1200 -1565
rect 1150 -1615 1200 -1585
rect 1150 -1635 1165 -1615
rect 1185 -1635 1200 -1615
rect 1150 -1650 1200 -1635
rect 1450 -965 1500 -950
rect 1450 -985 1465 -965
rect 1485 -985 1500 -965
rect 1450 -1015 1500 -985
rect 1450 -1035 1465 -1015
rect 1485 -1035 1500 -1015
rect 1450 -1065 1500 -1035
rect 1450 -1085 1465 -1065
rect 1485 -1085 1500 -1065
rect 1450 -1115 1500 -1085
rect 1450 -1135 1465 -1115
rect 1485 -1135 1500 -1115
rect 1450 -1165 1500 -1135
rect 1450 -1185 1465 -1165
rect 1485 -1185 1500 -1165
rect 1450 -1215 1500 -1185
rect 1450 -1235 1465 -1215
rect 1485 -1235 1500 -1215
rect 1450 -1265 1500 -1235
rect 1450 -1285 1465 -1265
rect 1485 -1285 1500 -1265
rect 1450 -1315 1500 -1285
rect 1450 -1335 1465 -1315
rect 1485 -1335 1500 -1315
rect 1450 -1365 1500 -1335
rect 1450 -1385 1465 -1365
rect 1485 -1385 1500 -1365
rect 1450 -1415 1500 -1385
rect 1450 -1435 1465 -1415
rect 1485 -1435 1500 -1415
rect 1450 -1465 1500 -1435
rect 1450 -1485 1465 -1465
rect 1485 -1485 1500 -1465
rect 1450 -1515 1500 -1485
rect 1450 -1535 1465 -1515
rect 1485 -1535 1500 -1515
rect 1450 -1565 1500 -1535
rect 1450 -1585 1465 -1565
rect 1485 -1585 1500 -1565
rect 1450 -1615 1500 -1585
rect 1450 -1635 1465 -1615
rect 1485 -1635 1500 -1615
rect 1450 -1650 1500 -1635
rect 1750 -965 1800 -950
rect 1750 -985 1765 -965
rect 1785 -985 1800 -965
rect 1750 -1015 1800 -985
rect 1750 -1035 1765 -1015
rect 1785 -1035 1800 -1015
rect 1750 -1065 1800 -1035
rect 1750 -1085 1765 -1065
rect 1785 -1085 1800 -1065
rect 1750 -1115 1800 -1085
rect 1750 -1135 1765 -1115
rect 1785 -1135 1800 -1115
rect 1750 -1165 1800 -1135
rect 1750 -1185 1765 -1165
rect 1785 -1185 1800 -1165
rect 1750 -1215 1800 -1185
rect 1750 -1235 1765 -1215
rect 1785 -1235 1800 -1215
rect 1750 -1265 1800 -1235
rect 1750 -1285 1765 -1265
rect 1785 -1285 1800 -1265
rect 1750 -1315 1800 -1285
rect 1750 -1335 1765 -1315
rect 1785 -1335 1800 -1315
rect 1750 -1365 1800 -1335
rect 1750 -1385 1765 -1365
rect 1785 -1385 1800 -1365
rect 1750 -1415 1800 -1385
rect 1750 -1435 1765 -1415
rect 1785 -1435 1800 -1415
rect 1750 -1465 1800 -1435
rect 1750 -1485 1765 -1465
rect 1785 -1485 1800 -1465
rect 1750 -1515 1800 -1485
rect 1750 -1535 1765 -1515
rect 1785 -1535 1800 -1515
rect 1750 -1565 1800 -1535
rect 1750 -1585 1765 -1565
rect 1785 -1585 1800 -1565
rect 1750 -1615 1800 -1585
rect 1750 -1635 1765 -1615
rect 1785 -1635 1800 -1615
rect 1750 -1650 1800 -1635
rect 2050 -965 2100 -950
rect 2050 -985 2065 -965
rect 2085 -985 2100 -965
rect 2050 -1015 2100 -985
rect 2050 -1035 2065 -1015
rect 2085 -1035 2100 -1015
rect 2050 -1065 2100 -1035
rect 2050 -1085 2065 -1065
rect 2085 -1085 2100 -1065
rect 2050 -1115 2100 -1085
rect 2050 -1135 2065 -1115
rect 2085 -1135 2100 -1115
rect 2050 -1165 2100 -1135
rect 2050 -1185 2065 -1165
rect 2085 -1185 2100 -1165
rect 2050 -1215 2100 -1185
rect 2050 -1235 2065 -1215
rect 2085 -1235 2100 -1215
rect 2050 -1265 2100 -1235
rect 2050 -1285 2065 -1265
rect 2085 -1285 2100 -1265
rect 2050 -1315 2100 -1285
rect 2050 -1335 2065 -1315
rect 2085 -1335 2100 -1315
rect 2050 -1365 2100 -1335
rect 2050 -1385 2065 -1365
rect 2085 -1385 2100 -1365
rect 2050 -1415 2100 -1385
rect 2050 -1435 2065 -1415
rect 2085 -1435 2100 -1415
rect 2050 -1465 2100 -1435
rect 2050 -1485 2065 -1465
rect 2085 -1485 2100 -1465
rect 2050 -1515 2100 -1485
rect 2050 -1535 2065 -1515
rect 2085 -1535 2100 -1515
rect 2050 -1565 2100 -1535
rect 2050 -1585 2065 -1565
rect 2085 -1585 2100 -1565
rect 2050 -1615 2100 -1585
rect 2050 -1635 2065 -1615
rect 2085 -1635 2100 -1615
rect 2050 -1650 2100 -1635
rect 2350 -965 2400 -950
rect 2350 -985 2365 -965
rect 2385 -985 2400 -965
rect 2350 -1015 2400 -985
rect 2350 -1035 2365 -1015
rect 2385 -1035 2400 -1015
rect 2350 -1065 2400 -1035
rect 2350 -1085 2365 -1065
rect 2385 -1085 2400 -1065
rect 2350 -1115 2400 -1085
rect 2350 -1135 2365 -1115
rect 2385 -1135 2400 -1115
rect 2350 -1165 2400 -1135
rect 2350 -1185 2365 -1165
rect 2385 -1185 2400 -1165
rect 2350 -1215 2400 -1185
rect 2350 -1235 2365 -1215
rect 2385 -1235 2400 -1215
rect 2350 -1265 2400 -1235
rect 2350 -1285 2365 -1265
rect 2385 -1285 2400 -1265
rect 2350 -1315 2400 -1285
rect 2350 -1335 2365 -1315
rect 2385 -1335 2400 -1315
rect 2350 -1365 2400 -1335
rect 2350 -1385 2365 -1365
rect 2385 -1385 2400 -1365
rect 2350 -1415 2400 -1385
rect 2350 -1435 2365 -1415
rect 2385 -1435 2400 -1415
rect 2350 -1465 2400 -1435
rect 2350 -1485 2365 -1465
rect 2385 -1485 2400 -1465
rect 2350 -1515 2400 -1485
rect 2350 -1535 2365 -1515
rect 2385 -1535 2400 -1515
rect 2350 -1565 2400 -1535
rect 2350 -1585 2365 -1565
rect 2385 -1585 2400 -1565
rect 2350 -1615 2400 -1585
rect 2350 -1635 2365 -1615
rect 2385 -1635 2400 -1615
rect 2350 -1650 2400 -1635
rect 2650 -965 2700 -950
rect 2650 -985 2665 -965
rect 2685 -985 2700 -965
rect 2650 -1015 2700 -985
rect 2650 -1035 2665 -1015
rect 2685 -1035 2700 -1015
rect 2650 -1065 2700 -1035
rect 2650 -1085 2665 -1065
rect 2685 -1085 2700 -1065
rect 2650 -1115 2700 -1085
rect 2650 -1135 2665 -1115
rect 2685 -1135 2700 -1115
rect 2650 -1165 2700 -1135
rect 2650 -1185 2665 -1165
rect 2685 -1185 2700 -1165
rect 2650 -1215 2700 -1185
rect 2650 -1235 2665 -1215
rect 2685 -1235 2700 -1215
rect 2650 -1265 2700 -1235
rect 2650 -1285 2665 -1265
rect 2685 -1285 2700 -1265
rect 2650 -1315 2700 -1285
rect 2650 -1335 2665 -1315
rect 2685 -1335 2700 -1315
rect 2650 -1365 2700 -1335
rect 2650 -1385 2665 -1365
rect 2685 -1385 2700 -1365
rect 2650 -1415 2700 -1385
rect 2650 -1435 2665 -1415
rect 2685 -1435 2700 -1415
rect 2650 -1465 2700 -1435
rect 2650 -1485 2665 -1465
rect 2685 -1485 2700 -1465
rect 2650 -1515 2700 -1485
rect 2650 -1535 2665 -1515
rect 2685 -1535 2700 -1515
rect 2650 -1565 2700 -1535
rect 2650 -1585 2665 -1565
rect 2685 -1585 2700 -1565
rect 2650 -1615 2700 -1585
rect 2650 -1635 2665 -1615
rect 2685 -1635 2700 -1615
rect 2650 -1650 2700 -1635
rect 2950 -965 3000 -950
rect 2950 -985 2965 -965
rect 2985 -985 3000 -965
rect 2950 -1015 3000 -985
rect 2950 -1035 2965 -1015
rect 2985 -1035 3000 -1015
rect 2950 -1065 3000 -1035
rect 2950 -1085 2965 -1065
rect 2985 -1085 3000 -1065
rect 2950 -1115 3000 -1085
rect 2950 -1135 2965 -1115
rect 2985 -1135 3000 -1115
rect 2950 -1165 3000 -1135
rect 2950 -1185 2965 -1165
rect 2985 -1185 3000 -1165
rect 2950 -1215 3000 -1185
rect 2950 -1235 2965 -1215
rect 2985 -1235 3000 -1215
rect 2950 -1265 3000 -1235
rect 2950 -1285 2965 -1265
rect 2985 -1285 3000 -1265
rect 2950 -1315 3000 -1285
rect 2950 -1335 2965 -1315
rect 2985 -1335 3000 -1315
rect 2950 -1365 3000 -1335
rect 2950 -1385 2965 -1365
rect 2985 -1385 3000 -1365
rect 2950 -1415 3000 -1385
rect 2950 -1435 2965 -1415
rect 2985 -1435 3000 -1415
rect 2950 -1465 3000 -1435
rect 2950 -1485 2965 -1465
rect 2985 -1485 3000 -1465
rect 2950 -1515 3000 -1485
rect 2950 -1535 2965 -1515
rect 2985 -1535 3000 -1515
rect 2950 -1565 3000 -1535
rect 2950 -1585 2965 -1565
rect 2985 -1585 3000 -1565
rect 2950 -1615 3000 -1585
rect 2950 -1635 2965 -1615
rect 2985 -1635 3000 -1615
rect 2950 -1650 3000 -1635
rect 3250 -965 3300 -950
rect 3250 -985 3265 -965
rect 3285 -985 3300 -965
rect 3250 -1015 3300 -985
rect 3250 -1035 3265 -1015
rect 3285 -1035 3300 -1015
rect 3250 -1065 3300 -1035
rect 3250 -1085 3265 -1065
rect 3285 -1085 3300 -1065
rect 3250 -1115 3300 -1085
rect 3250 -1135 3265 -1115
rect 3285 -1135 3300 -1115
rect 3250 -1165 3300 -1135
rect 3250 -1185 3265 -1165
rect 3285 -1185 3300 -1165
rect 3250 -1215 3300 -1185
rect 3250 -1235 3265 -1215
rect 3285 -1235 3300 -1215
rect 3250 -1265 3300 -1235
rect 3250 -1285 3265 -1265
rect 3285 -1285 3300 -1265
rect 3250 -1315 3300 -1285
rect 3250 -1335 3265 -1315
rect 3285 -1335 3300 -1315
rect 3250 -1365 3300 -1335
rect 3250 -1385 3265 -1365
rect 3285 -1385 3300 -1365
rect 3250 -1415 3300 -1385
rect 3250 -1435 3265 -1415
rect 3285 -1435 3300 -1415
rect 3250 -1465 3300 -1435
rect 3250 -1485 3265 -1465
rect 3285 -1485 3300 -1465
rect 3250 -1515 3300 -1485
rect 3250 -1535 3265 -1515
rect 3285 -1535 3300 -1515
rect 3250 -1565 3300 -1535
rect 3250 -1585 3265 -1565
rect 3285 -1585 3300 -1565
rect 3250 -1615 3300 -1585
rect 3250 -1635 3265 -1615
rect 3285 -1635 3300 -1615
rect 3250 -1650 3300 -1635
rect 3550 -965 3600 -950
rect 3550 -985 3565 -965
rect 3585 -985 3600 -965
rect 3550 -1015 3600 -985
rect 3550 -1035 3565 -1015
rect 3585 -1035 3600 -1015
rect 3550 -1065 3600 -1035
rect 3550 -1085 3565 -1065
rect 3585 -1085 3600 -1065
rect 3550 -1115 3600 -1085
rect 3550 -1135 3565 -1115
rect 3585 -1135 3600 -1115
rect 3550 -1165 3600 -1135
rect 3550 -1185 3565 -1165
rect 3585 -1185 3600 -1165
rect 3550 -1215 3600 -1185
rect 3550 -1235 3565 -1215
rect 3585 -1235 3600 -1215
rect 3550 -1265 3600 -1235
rect 3550 -1285 3565 -1265
rect 3585 -1285 3600 -1265
rect 3550 -1315 3600 -1285
rect 3550 -1335 3565 -1315
rect 3585 -1335 3600 -1315
rect 3550 -1365 3600 -1335
rect 3550 -1385 3565 -1365
rect 3585 -1385 3600 -1365
rect 3550 -1415 3600 -1385
rect 3550 -1435 3565 -1415
rect 3585 -1435 3600 -1415
rect 3550 -1465 3600 -1435
rect 3550 -1485 3565 -1465
rect 3585 -1485 3600 -1465
rect 3550 -1515 3600 -1485
rect 3550 -1535 3565 -1515
rect 3585 -1535 3600 -1515
rect 3550 -1565 3600 -1535
rect 3550 -1585 3565 -1565
rect 3585 -1585 3600 -1565
rect 3550 -1615 3600 -1585
rect 3550 -1635 3565 -1615
rect 3585 -1635 3600 -1615
rect 3550 -1650 3600 -1635
rect 3700 -965 3750 -950
rect 3700 -985 3715 -965
rect 3735 -985 3750 -965
rect 3700 -1015 3750 -985
rect 3700 -1035 3715 -1015
rect 3735 -1035 3750 -1015
rect 3700 -1065 3750 -1035
rect 3700 -1085 3715 -1065
rect 3735 -1085 3750 -1065
rect 3700 -1115 3750 -1085
rect 3700 -1135 3715 -1115
rect 3735 -1135 3750 -1115
rect 3700 -1165 3750 -1135
rect 3700 -1185 3715 -1165
rect 3735 -1185 3750 -1165
rect 3700 -1215 3750 -1185
rect 3700 -1235 3715 -1215
rect 3735 -1235 3750 -1215
rect 3700 -1265 3750 -1235
rect 3700 -1285 3715 -1265
rect 3735 -1285 3750 -1265
rect 3700 -1315 3750 -1285
rect 3700 -1335 3715 -1315
rect 3735 -1335 3750 -1315
rect 3700 -1365 3750 -1335
rect 3700 -1385 3715 -1365
rect 3735 -1385 3750 -1365
rect 3700 -1415 3750 -1385
rect 3700 -1435 3715 -1415
rect 3735 -1435 3750 -1415
rect 3700 -1465 3750 -1435
rect 3700 -1485 3715 -1465
rect 3735 -1485 3750 -1465
rect 3700 -1515 3750 -1485
rect 3700 -1535 3715 -1515
rect 3735 -1535 3750 -1515
rect 3700 -1565 3750 -1535
rect 3700 -1585 3715 -1565
rect 3735 -1585 3750 -1565
rect 3700 -1615 3750 -1585
rect 3700 -1635 3715 -1615
rect 3735 -1635 3750 -1615
rect 3700 -1650 3750 -1635
rect 3850 -965 3900 -950
rect 3850 -985 3865 -965
rect 3885 -985 3900 -965
rect 3850 -1015 3900 -985
rect 3850 -1035 3865 -1015
rect 3885 -1035 3900 -1015
rect 3850 -1065 3900 -1035
rect 3850 -1085 3865 -1065
rect 3885 -1085 3900 -1065
rect 3850 -1115 3900 -1085
rect 3850 -1135 3865 -1115
rect 3885 -1135 3900 -1115
rect 3850 -1165 3900 -1135
rect 3850 -1185 3865 -1165
rect 3885 -1185 3900 -1165
rect 3850 -1215 3900 -1185
rect 3850 -1235 3865 -1215
rect 3885 -1235 3900 -1215
rect 3850 -1265 3900 -1235
rect 3850 -1285 3865 -1265
rect 3885 -1285 3900 -1265
rect 3850 -1315 3900 -1285
rect 3850 -1335 3865 -1315
rect 3885 -1335 3900 -1315
rect 3850 -1365 3900 -1335
rect 3850 -1385 3865 -1365
rect 3885 -1385 3900 -1365
rect 3850 -1415 3900 -1385
rect 3850 -1435 3865 -1415
rect 3885 -1435 3900 -1415
rect 3850 -1465 3900 -1435
rect 3850 -1485 3865 -1465
rect 3885 -1485 3900 -1465
rect 3850 -1515 3900 -1485
rect 3850 -1535 3865 -1515
rect 3885 -1535 3900 -1515
rect 3850 -1565 3900 -1535
rect 3850 -1585 3865 -1565
rect 3885 -1585 3900 -1565
rect 3850 -1615 3900 -1585
rect 3850 -1635 3865 -1615
rect 3885 -1635 3900 -1615
rect 3850 -1650 3900 -1635
rect 4000 -965 4050 -950
rect 4000 -985 4015 -965
rect 4035 -985 4050 -965
rect 4000 -1015 4050 -985
rect 4000 -1035 4015 -1015
rect 4035 -1035 4050 -1015
rect 4000 -1065 4050 -1035
rect 4000 -1085 4015 -1065
rect 4035 -1085 4050 -1065
rect 4000 -1115 4050 -1085
rect 4000 -1135 4015 -1115
rect 4035 -1135 4050 -1115
rect 4000 -1165 4050 -1135
rect 4000 -1185 4015 -1165
rect 4035 -1185 4050 -1165
rect 4000 -1215 4050 -1185
rect 4000 -1235 4015 -1215
rect 4035 -1235 4050 -1215
rect 4000 -1265 4050 -1235
rect 4000 -1285 4015 -1265
rect 4035 -1285 4050 -1265
rect 4000 -1315 4050 -1285
rect 4000 -1335 4015 -1315
rect 4035 -1335 4050 -1315
rect 4000 -1365 4050 -1335
rect 4000 -1385 4015 -1365
rect 4035 -1385 4050 -1365
rect 4000 -1415 4050 -1385
rect 4000 -1435 4015 -1415
rect 4035 -1435 4050 -1415
rect 4000 -1465 4050 -1435
rect 4000 -1485 4015 -1465
rect 4035 -1485 4050 -1465
rect 4000 -1515 4050 -1485
rect 4000 -1535 4015 -1515
rect 4035 -1535 4050 -1515
rect 4000 -1565 4050 -1535
rect 4000 -1585 4015 -1565
rect 4035 -1585 4050 -1565
rect 4000 -1615 4050 -1585
rect 4000 -1635 4015 -1615
rect 4035 -1635 4050 -1615
rect 4000 -1650 4050 -1635
rect 4150 -965 4200 -950
rect 4150 -985 4165 -965
rect 4185 -985 4200 -965
rect 4150 -1015 4200 -985
rect 4150 -1035 4165 -1015
rect 4185 -1035 4200 -1015
rect 4150 -1065 4200 -1035
rect 4150 -1085 4165 -1065
rect 4185 -1085 4200 -1065
rect 4150 -1115 4200 -1085
rect 4150 -1135 4165 -1115
rect 4185 -1135 4200 -1115
rect 4150 -1165 4200 -1135
rect 4150 -1185 4165 -1165
rect 4185 -1185 4200 -1165
rect 4150 -1215 4200 -1185
rect 4150 -1235 4165 -1215
rect 4185 -1235 4200 -1215
rect 4150 -1265 4200 -1235
rect 4150 -1285 4165 -1265
rect 4185 -1285 4200 -1265
rect 4150 -1315 4200 -1285
rect 4150 -1335 4165 -1315
rect 4185 -1335 4200 -1315
rect 4150 -1365 4200 -1335
rect 4150 -1385 4165 -1365
rect 4185 -1385 4200 -1365
rect 4150 -1415 4200 -1385
rect 4150 -1435 4165 -1415
rect 4185 -1435 4200 -1415
rect 4150 -1465 4200 -1435
rect 4150 -1485 4165 -1465
rect 4185 -1485 4200 -1465
rect 4150 -1515 4200 -1485
rect 4150 -1535 4165 -1515
rect 4185 -1535 4200 -1515
rect 4150 -1565 4200 -1535
rect 4150 -1585 4165 -1565
rect 4185 -1585 4200 -1565
rect 4150 -1615 4200 -1585
rect 4150 -1635 4165 -1615
rect 4185 -1635 4200 -1615
rect 4150 -1650 4200 -1635
rect 4300 -965 4350 -950
rect 4300 -985 4315 -965
rect 4335 -985 4350 -965
rect 4300 -1015 4350 -985
rect 4300 -1035 4315 -1015
rect 4335 -1035 4350 -1015
rect 4300 -1065 4350 -1035
rect 4300 -1085 4315 -1065
rect 4335 -1085 4350 -1065
rect 4300 -1115 4350 -1085
rect 4300 -1135 4315 -1115
rect 4335 -1135 4350 -1115
rect 4300 -1165 4350 -1135
rect 4300 -1185 4315 -1165
rect 4335 -1185 4350 -1165
rect 4300 -1215 4350 -1185
rect 4300 -1235 4315 -1215
rect 4335 -1235 4350 -1215
rect 4300 -1265 4350 -1235
rect 4300 -1285 4315 -1265
rect 4335 -1285 4350 -1265
rect 4300 -1315 4350 -1285
rect 4300 -1335 4315 -1315
rect 4335 -1335 4350 -1315
rect 4300 -1365 4350 -1335
rect 4300 -1385 4315 -1365
rect 4335 -1385 4350 -1365
rect 4300 -1415 4350 -1385
rect 4300 -1435 4315 -1415
rect 4335 -1435 4350 -1415
rect 4300 -1465 4350 -1435
rect 4300 -1485 4315 -1465
rect 4335 -1485 4350 -1465
rect 4300 -1515 4350 -1485
rect 4300 -1535 4315 -1515
rect 4335 -1535 4350 -1515
rect 4300 -1565 4350 -1535
rect 4300 -1585 4315 -1565
rect 4335 -1585 4350 -1565
rect 4300 -1615 4350 -1585
rect 4300 -1635 4315 -1615
rect 4335 -1635 4350 -1615
rect 4300 -1650 4350 -1635
rect 4450 -965 4500 -950
rect 4450 -985 4465 -965
rect 4485 -985 4500 -965
rect 4450 -1015 4500 -985
rect 4450 -1035 4465 -1015
rect 4485 -1035 4500 -1015
rect 4450 -1065 4500 -1035
rect 4450 -1085 4465 -1065
rect 4485 -1085 4500 -1065
rect 4450 -1115 4500 -1085
rect 4450 -1135 4465 -1115
rect 4485 -1135 4500 -1115
rect 4450 -1165 4500 -1135
rect 4450 -1185 4465 -1165
rect 4485 -1185 4500 -1165
rect 4450 -1215 4500 -1185
rect 4450 -1235 4465 -1215
rect 4485 -1235 4500 -1215
rect 4450 -1265 4500 -1235
rect 4450 -1285 4465 -1265
rect 4485 -1285 4500 -1265
rect 4450 -1315 4500 -1285
rect 4450 -1335 4465 -1315
rect 4485 -1335 4500 -1315
rect 4450 -1365 4500 -1335
rect 4450 -1385 4465 -1365
rect 4485 -1385 4500 -1365
rect 4450 -1415 4500 -1385
rect 4450 -1435 4465 -1415
rect 4485 -1435 4500 -1415
rect 4450 -1465 4500 -1435
rect 4450 -1485 4465 -1465
rect 4485 -1485 4500 -1465
rect 4450 -1515 4500 -1485
rect 4450 -1535 4465 -1515
rect 4485 -1535 4500 -1515
rect 4450 -1565 4500 -1535
rect 4450 -1585 4465 -1565
rect 4485 -1585 4500 -1565
rect 4450 -1615 4500 -1585
rect 4450 -1635 4465 -1615
rect 4485 -1635 4500 -1615
rect 4450 -1650 4500 -1635
rect 4600 -965 4650 -950
rect 4600 -985 4615 -965
rect 4635 -985 4650 -965
rect 4600 -1015 4650 -985
rect 4600 -1035 4615 -1015
rect 4635 -1035 4650 -1015
rect 4600 -1065 4650 -1035
rect 4600 -1085 4615 -1065
rect 4635 -1085 4650 -1065
rect 4600 -1115 4650 -1085
rect 4600 -1135 4615 -1115
rect 4635 -1135 4650 -1115
rect 4600 -1165 4650 -1135
rect 4600 -1185 4615 -1165
rect 4635 -1185 4650 -1165
rect 4600 -1215 4650 -1185
rect 4600 -1235 4615 -1215
rect 4635 -1235 4650 -1215
rect 4600 -1265 4650 -1235
rect 4600 -1285 4615 -1265
rect 4635 -1285 4650 -1265
rect 4600 -1315 4650 -1285
rect 4600 -1335 4615 -1315
rect 4635 -1335 4650 -1315
rect 4600 -1365 4650 -1335
rect 4600 -1385 4615 -1365
rect 4635 -1385 4650 -1365
rect 4600 -1415 4650 -1385
rect 4600 -1435 4615 -1415
rect 4635 -1435 4650 -1415
rect 4600 -1465 4650 -1435
rect 4600 -1485 4615 -1465
rect 4635 -1485 4650 -1465
rect 4600 -1515 4650 -1485
rect 4600 -1535 4615 -1515
rect 4635 -1535 4650 -1515
rect 4600 -1565 4650 -1535
rect 4600 -1585 4615 -1565
rect 4635 -1585 4650 -1565
rect 4600 -1615 4650 -1585
rect 4600 -1635 4615 -1615
rect 4635 -1635 4650 -1615
rect 4600 -1650 4650 -1635
rect 4750 -965 4800 -950
rect 4750 -985 4765 -965
rect 4785 -985 4800 -965
rect 4750 -1015 4800 -985
rect 4750 -1035 4765 -1015
rect 4785 -1035 4800 -1015
rect 4750 -1065 4800 -1035
rect 4750 -1085 4765 -1065
rect 4785 -1085 4800 -1065
rect 4750 -1115 4800 -1085
rect 4750 -1135 4765 -1115
rect 4785 -1135 4800 -1115
rect 4750 -1165 4800 -1135
rect 4750 -1185 4765 -1165
rect 4785 -1185 4800 -1165
rect 4750 -1215 4800 -1185
rect 4750 -1235 4765 -1215
rect 4785 -1235 4800 -1215
rect 4750 -1265 4800 -1235
rect 4750 -1285 4765 -1265
rect 4785 -1285 4800 -1265
rect 4750 -1315 4800 -1285
rect 4750 -1335 4765 -1315
rect 4785 -1335 4800 -1315
rect 4750 -1365 4800 -1335
rect 4750 -1385 4765 -1365
rect 4785 -1385 4800 -1365
rect 4750 -1415 4800 -1385
rect 4750 -1435 4765 -1415
rect 4785 -1435 4800 -1415
rect 4750 -1465 4800 -1435
rect 4750 -1485 4765 -1465
rect 4785 -1485 4800 -1465
rect 4750 -1515 4800 -1485
rect 4750 -1535 4765 -1515
rect 4785 -1535 4800 -1515
rect 4750 -1565 4800 -1535
rect 4750 -1585 4765 -1565
rect 4785 -1585 4800 -1565
rect 4750 -1615 4800 -1585
rect 4750 -1635 4765 -1615
rect 4785 -1635 4800 -1615
rect 4750 -1650 4800 -1635
rect 5050 -965 5100 -950
rect 5050 -985 5065 -965
rect 5085 -985 5100 -965
rect 5050 -1015 5100 -985
rect 5050 -1035 5065 -1015
rect 5085 -1035 5100 -1015
rect 5050 -1065 5100 -1035
rect 5050 -1085 5065 -1065
rect 5085 -1085 5100 -1065
rect 5050 -1115 5100 -1085
rect 5050 -1135 5065 -1115
rect 5085 -1135 5100 -1115
rect 5050 -1165 5100 -1135
rect 5050 -1185 5065 -1165
rect 5085 -1185 5100 -1165
rect 5050 -1215 5100 -1185
rect 5050 -1235 5065 -1215
rect 5085 -1235 5100 -1215
rect 5050 -1265 5100 -1235
rect 5050 -1285 5065 -1265
rect 5085 -1285 5100 -1265
rect 5050 -1315 5100 -1285
rect 5050 -1335 5065 -1315
rect 5085 -1335 5100 -1315
rect 5050 -1365 5100 -1335
rect 5050 -1385 5065 -1365
rect 5085 -1385 5100 -1365
rect 5050 -1415 5100 -1385
rect 5050 -1435 5065 -1415
rect 5085 -1435 5100 -1415
rect 5050 -1465 5100 -1435
rect 5050 -1485 5065 -1465
rect 5085 -1485 5100 -1465
rect 5050 -1515 5100 -1485
rect 5050 -1535 5065 -1515
rect 5085 -1535 5100 -1515
rect 5050 -1565 5100 -1535
rect 5050 -1585 5065 -1565
rect 5085 -1585 5100 -1565
rect 5050 -1615 5100 -1585
rect 5050 -1635 5065 -1615
rect 5085 -1635 5100 -1615
rect 5050 -1650 5100 -1635
rect 5350 -965 5400 -950
rect 5350 -985 5365 -965
rect 5385 -985 5400 -965
rect 5350 -1015 5400 -985
rect 5350 -1035 5365 -1015
rect 5385 -1035 5400 -1015
rect 5350 -1065 5400 -1035
rect 5350 -1085 5365 -1065
rect 5385 -1085 5400 -1065
rect 5350 -1115 5400 -1085
rect 5350 -1135 5365 -1115
rect 5385 -1135 5400 -1115
rect 5350 -1165 5400 -1135
rect 5350 -1185 5365 -1165
rect 5385 -1185 5400 -1165
rect 5350 -1215 5400 -1185
rect 5350 -1235 5365 -1215
rect 5385 -1235 5400 -1215
rect 5350 -1265 5400 -1235
rect 5350 -1285 5365 -1265
rect 5385 -1285 5400 -1265
rect 5350 -1315 5400 -1285
rect 5350 -1335 5365 -1315
rect 5385 -1335 5400 -1315
rect 5350 -1365 5400 -1335
rect 5350 -1385 5365 -1365
rect 5385 -1385 5400 -1365
rect 5350 -1415 5400 -1385
rect 5350 -1435 5365 -1415
rect 5385 -1435 5400 -1415
rect 5350 -1465 5400 -1435
rect 5350 -1485 5365 -1465
rect 5385 -1485 5400 -1465
rect 5350 -1515 5400 -1485
rect 5350 -1535 5365 -1515
rect 5385 -1535 5400 -1515
rect 5350 -1565 5400 -1535
rect 5350 -1585 5365 -1565
rect 5385 -1585 5400 -1565
rect 5350 -1615 5400 -1585
rect 5350 -1635 5365 -1615
rect 5385 -1635 5400 -1615
rect 5350 -1650 5400 -1635
rect 5650 -965 5700 -950
rect 5650 -985 5665 -965
rect 5685 -985 5700 -965
rect 5650 -1015 5700 -985
rect 5650 -1035 5665 -1015
rect 5685 -1035 5700 -1015
rect 5650 -1065 5700 -1035
rect 5650 -1085 5665 -1065
rect 5685 -1085 5700 -1065
rect 5650 -1115 5700 -1085
rect 5650 -1135 5665 -1115
rect 5685 -1135 5700 -1115
rect 5650 -1165 5700 -1135
rect 5650 -1185 5665 -1165
rect 5685 -1185 5700 -1165
rect 5650 -1215 5700 -1185
rect 5650 -1235 5665 -1215
rect 5685 -1235 5700 -1215
rect 5650 -1265 5700 -1235
rect 5650 -1285 5665 -1265
rect 5685 -1285 5700 -1265
rect 5650 -1315 5700 -1285
rect 5650 -1335 5665 -1315
rect 5685 -1335 5700 -1315
rect 5650 -1365 5700 -1335
rect 5650 -1385 5665 -1365
rect 5685 -1385 5700 -1365
rect 5650 -1415 5700 -1385
rect 5650 -1435 5665 -1415
rect 5685 -1435 5700 -1415
rect 5650 -1465 5700 -1435
rect 5650 -1485 5665 -1465
rect 5685 -1485 5700 -1465
rect 5650 -1515 5700 -1485
rect 5650 -1535 5665 -1515
rect 5685 -1535 5700 -1515
rect 5650 -1565 5700 -1535
rect 5650 -1585 5665 -1565
rect 5685 -1585 5700 -1565
rect 5650 -1615 5700 -1585
rect 5650 -1635 5665 -1615
rect 5685 -1635 5700 -1615
rect 5650 -1650 5700 -1635
rect 5950 -965 6000 -950
rect 5950 -985 5965 -965
rect 5985 -985 6000 -965
rect 5950 -1015 6000 -985
rect 5950 -1035 5965 -1015
rect 5985 -1035 6000 -1015
rect 5950 -1065 6000 -1035
rect 5950 -1085 5965 -1065
rect 5985 -1085 6000 -1065
rect 5950 -1115 6000 -1085
rect 5950 -1135 5965 -1115
rect 5985 -1135 6000 -1115
rect 5950 -1165 6000 -1135
rect 5950 -1185 5965 -1165
rect 5985 -1185 6000 -1165
rect 5950 -1215 6000 -1185
rect 5950 -1235 5965 -1215
rect 5985 -1235 6000 -1215
rect 5950 -1265 6000 -1235
rect 5950 -1285 5965 -1265
rect 5985 -1285 6000 -1265
rect 5950 -1315 6000 -1285
rect 5950 -1335 5965 -1315
rect 5985 -1335 6000 -1315
rect 5950 -1365 6000 -1335
rect 5950 -1385 5965 -1365
rect 5985 -1385 6000 -1365
rect 5950 -1415 6000 -1385
rect 5950 -1435 5965 -1415
rect 5985 -1435 6000 -1415
rect 5950 -1465 6000 -1435
rect 5950 -1485 5965 -1465
rect 5985 -1485 6000 -1465
rect 5950 -1515 6000 -1485
rect 5950 -1535 5965 -1515
rect 5985 -1535 6000 -1515
rect 5950 -1565 6000 -1535
rect 5950 -1585 5965 -1565
rect 5985 -1585 6000 -1565
rect 5950 -1615 6000 -1585
rect 5950 -1635 5965 -1615
rect 5985 -1635 6000 -1615
rect 5950 -1650 6000 -1635
rect 6250 -965 6300 -950
rect 6250 -985 6265 -965
rect 6285 -985 6300 -965
rect 6250 -1015 6300 -985
rect 6250 -1035 6265 -1015
rect 6285 -1035 6300 -1015
rect 6250 -1065 6300 -1035
rect 6250 -1085 6265 -1065
rect 6285 -1085 6300 -1065
rect 6250 -1115 6300 -1085
rect 6250 -1135 6265 -1115
rect 6285 -1135 6300 -1115
rect 6250 -1165 6300 -1135
rect 6250 -1185 6265 -1165
rect 6285 -1185 6300 -1165
rect 6250 -1215 6300 -1185
rect 6250 -1235 6265 -1215
rect 6285 -1235 6300 -1215
rect 6250 -1265 6300 -1235
rect 6250 -1285 6265 -1265
rect 6285 -1285 6300 -1265
rect 6250 -1315 6300 -1285
rect 6250 -1335 6265 -1315
rect 6285 -1335 6300 -1315
rect 6250 -1365 6300 -1335
rect 6250 -1385 6265 -1365
rect 6285 -1385 6300 -1365
rect 6250 -1415 6300 -1385
rect 6250 -1435 6265 -1415
rect 6285 -1435 6300 -1415
rect 6250 -1465 6300 -1435
rect 6250 -1485 6265 -1465
rect 6285 -1485 6300 -1465
rect 6250 -1515 6300 -1485
rect 6250 -1535 6265 -1515
rect 6285 -1535 6300 -1515
rect 6250 -1565 6300 -1535
rect 6250 -1585 6265 -1565
rect 6285 -1585 6300 -1565
rect 6250 -1615 6300 -1585
rect 6250 -1635 6265 -1615
rect 6285 -1635 6300 -1615
rect 6250 -1650 6300 -1635
rect 6550 -965 6600 -950
rect 6550 -985 6565 -965
rect 6585 -985 6600 -965
rect 6550 -1015 6600 -985
rect 6550 -1035 6565 -1015
rect 6585 -1035 6600 -1015
rect 6550 -1065 6600 -1035
rect 6550 -1085 6565 -1065
rect 6585 -1085 6600 -1065
rect 6550 -1115 6600 -1085
rect 6550 -1135 6565 -1115
rect 6585 -1135 6600 -1115
rect 6550 -1165 6600 -1135
rect 6550 -1185 6565 -1165
rect 6585 -1185 6600 -1165
rect 6550 -1215 6600 -1185
rect 6550 -1235 6565 -1215
rect 6585 -1235 6600 -1215
rect 6550 -1265 6600 -1235
rect 6550 -1285 6565 -1265
rect 6585 -1285 6600 -1265
rect 6550 -1315 6600 -1285
rect 6550 -1335 6565 -1315
rect 6585 -1335 6600 -1315
rect 6550 -1365 6600 -1335
rect 6550 -1385 6565 -1365
rect 6585 -1385 6600 -1365
rect 6550 -1415 6600 -1385
rect 6550 -1435 6565 -1415
rect 6585 -1435 6600 -1415
rect 6550 -1465 6600 -1435
rect 6550 -1485 6565 -1465
rect 6585 -1485 6600 -1465
rect 6550 -1515 6600 -1485
rect 6550 -1535 6565 -1515
rect 6585 -1535 6600 -1515
rect 6550 -1565 6600 -1535
rect 6550 -1585 6565 -1565
rect 6585 -1585 6600 -1565
rect 6550 -1615 6600 -1585
rect 6550 -1635 6565 -1615
rect 6585 -1635 6600 -1615
rect 6550 -1650 6600 -1635
rect 6850 -965 6900 -950
rect 6850 -985 6865 -965
rect 6885 -985 6900 -965
rect 6850 -1015 6900 -985
rect 6850 -1035 6865 -1015
rect 6885 -1035 6900 -1015
rect 6850 -1065 6900 -1035
rect 6850 -1085 6865 -1065
rect 6885 -1085 6900 -1065
rect 6850 -1115 6900 -1085
rect 6850 -1135 6865 -1115
rect 6885 -1135 6900 -1115
rect 6850 -1165 6900 -1135
rect 6850 -1185 6865 -1165
rect 6885 -1185 6900 -1165
rect 6850 -1215 6900 -1185
rect 6850 -1235 6865 -1215
rect 6885 -1235 6900 -1215
rect 6850 -1265 6900 -1235
rect 6850 -1285 6865 -1265
rect 6885 -1285 6900 -1265
rect 6850 -1315 6900 -1285
rect 6850 -1335 6865 -1315
rect 6885 -1335 6900 -1315
rect 6850 -1365 6900 -1335
rect 6850 -1385 6865 -1365
rect 6885 -1385 6900 -1365
rect 6850 -1415 6900 -1385
rect 6850 -1435 6865 -1415
rect 6885 -1435 6900 -1415
rect 6850 -1465 6900 -1435
rect 6850 -1485 6865 -1465
rect 6885 -1485 6900 -1465
rect 6850 -1515 6900 -1485
rect 6850 -1535 6865 -1515
rect 6885 -1535 6900 -1515
rect 6850 -1565 6900 -1535
rect 6850 -1585 6865 -1565
rect 6885 -1585 6900 -1565
rect 6850 -1615 6900 -1585
rect 6850 -1635 6865 -1615
rect 6885 -1635 6900 -1615
rect 6850 -1650 6900 -1635
rect 7150 -965 7200 -950
rect 7150 -985 7165 -965
rect 7185 -985 7200 -965
rect 7150 -1015 7200 -985
rect 7150 -1035 7165 -1015
rect 7185 -1035 7200 -1015
rect 7150 -1065 7200 -1035
rect 7150 -1085 7165 -1065
rect 7185 -1085 7200 -1065
rect 7150 -1115 7200 -1085
rect 7150 -1135 7165 -1115
rect 7185 -1135 7200 -1115
rect 7150 -1165 7200 -1135
rect 7150 -1185 7165 -1165
rect 7185 -1185 7200 -1165
rect 7150 -1215 7200 -1185
rect 7150 -1235 7165 -1215
rect 7185 -1235 7200 -1215
rect 7150 -1265 7200 -1235
rect 7150 -1285 7165 -1265
rect 7185 -1285 7200 -1265
rect 7150 -1315 7200 -1285
rect 7150 -1335 7165 -1315
rect 7185 -1335 7200 -1315
rect 7150 -1365 7200 -1335
rect 7150 -1385 7165 -1365
rect 7185 -1385 7200 -1365
rect 7150 -1415 7200 -1385
rect 7150 -1435 7165 -1415
rect 7185 -1435 7200 -1415
rect 7150 -1465 7200 -1435
rect 7150 -1485 7165 -1465
rect 7185 -1485 7200 -1465
rect 7150 -1515 7200 -1485
rect 7150 -1535 7165 -1515
rect 7185 -1535 7200 -1515
rect 7150 -1565 7200 -1535
rect 7150 -1585 7165 -1565
rect 7185 -1585 7200 -1565
rect 7150 -1615 7200 -1585
rect 7150 -1635 7165 -1615
rect 7185 -1635 7200 -1615
rect 7150 -1650 7200 -1635
rect 8350 -965 8400 -950
rect 8350 -985 8365 -965
rect 8385 -985 8400 -965
rect 8350 -1015 8400 -985
rect 8350 -1035 8365 -1015
rect 8385 -1035 8400 -1015
rect 8350 -1065 8400 -1035
rect 8350 -1085 8365 -1065
rect 8385 -1085 8400 -1065
rect 8350 -1115 8400 -1085
rect 8350 -1135 8365 -1115
rect 8385 -1135 8400 -1115
rect 8350 -1165 8400 -1135
rect 8350 -1185 8365 -1165
rect 8385 -1185 8400 -1165
rect 8350 -1215 8400 -1185
rect 8350 -1235 8365 -1215
rect 8385 -1235 8400 -1215
rect 8350 -1265 8400 -1235
rect 8350 -1285 8365 -1265
rect 8385 -1285 8400 -1265
rect 8350 -1315 8400 -1285
rect 8350 -1335 8365 -1315
rect 8385 -1335 8400 -1315
rect 8350 -1365 8400 -1335
rect 8350 -1385 8365 -1365
rect 8385 -1385 8400 -1365
rect 8350 -1415 8400 -1385
rect 8350 -1435 8365 -1415
rect 8385 -1435 8400 -1415
rect 8350 -1465 8400 -1435
rect 8350 -1485 8365 -1465
rect 8385 -1485 8400 -1465
rect 8350 -1515 8400 -1485
rect 8350 -1535 8365 -1515
rect 8385 -1535 8400 -1515
rect 8350 -1565 8400 -1535
rect 8350 -1585 8365 -1565
rect 8385 -1585 8400 -1565
rect 8350 -1615 8400 -1585
rect 8350 -1635 8365 -1615
rect 8385 -1635 8400 -1615
rect 8350 -1650 8400 -1635
rect 9550 -965 9600 -950
rect 9550 -985 9565 -965
rect 9585 -985 9600 -965
rect 9550 -1015 9600 -985
rect 9550 -1035 9565 -1015
rect 9585 -1035 9600 -1015
rect 9550 -1065 9600 -1035
rect 9550 -1085 9565 -1065
rect 9585 -1085 9600 -1065
rect 9550 -1115 9600 -1085
rect 9550 -1135 9565 -1115
rect 9585 -1135 9600 -1115
rect 9550 -1165 9600 -1135
rect 9550 -1185 9565 -1165
rect 9585 -1185 9600 -1165
rect 9550 -1215 9600 -1185
rect 9550 -1235 9565 -1215
rect 9585 -1235 9600 -1215
rect 9550 -1265 9600 -1235
rect 9550 -1285 9565 -1265
rect 9585 -1285 9600 -1265
rect 9550 -1315 9600 -1285
rect 9550 -1335 9565 -1315
rect 9585 -1335 9600 -1315
rect 9550 -1365 9600 -1335
rect 9550 -1385 9565 -1365
rect 9585 -1385 9600 -1365
rect 9550 -1415 9600 -1385
rect 9550 -1435 9565 -1415
rect 9585 -1435 9600 -1415
rect 9550 -1465 9600 -1435
rect 9550 -1485 9565 -1465
rect 9585 -1485 9600 -1465
rect 9550 -1515 9600 -1485
rect 9550 -1535 9565 -1515
rect 9585 -1535 9600 -1515
rect 9550 -1565 9600 -1535
rect 9550 -1585 9565 -1565
rect 9585 -1585 9600 -1565
rect 9550 -1615 9600 -1585
rect 9550 -1635 9565 -1615
rect 9585 -1635 9600 -1615
rect 9550 -1650 9600 -1635
rect 10750 -965 10800 -950
rect 10750 -985 10765 -965
rect 10785 -985 10800 -965
rect 10750 -1015 10800 -985
rect 10750 -1035 10765 -1015
rect 10785 -1035 10800 -1015
rect 10750 -1065 10800 -1035
rect 10750 -1085 10765 -1065
rect 10785 -1085 10800 -1065
rect 10750 -1115 10800 -1085
rect 10750 -1135 10765 -1115
rect 10785 -1135 10800 -1115
rect 10750 -1165 10800 -1135
rect 10750 -1185 10765 -1165
rect 10785 -1185 10800 -1165
rect 10750 -1215 10800 -1185
rect 10750 -1235 10765 -1215
rect 10785 -1235 10800 -1215
rect 10750 -1265 10800 -1235
rect 10750 -1285 10765 -1265
rect 10785 -1285 10800 -1265
rect 10750 -1315 10800 -1285
rect 10750 -1335 10765 -1315
rect 10785 -1335 10800 -1315
rect 10750 -1365 10800 -1335
rect 10750 -1385 10765 -1365
rect 10785 -1385 10800 -1365
rect 10750 -1415 10800 -1385
rect 10750 -1435 10765 -1415
rect 10785 -1435 10800 -1415
rect 10750 -1465 10800 -1435
rect 10750 -1485 10765 -1465
rect 10785 -1485 10800 -1465
rect 10750 -1515 10800 -1485
rect 10750 -1535 10765 -1515
rect 10785 -1535 10800 -1515
rect 10750 -1565 10800 -1535
rect 10750 -1585 10765 -1565
rect 10785 -1585 10800 -1565
rect 10750 -1615 10800 -1585
rect 10750 -1635 10765 -1615
rect 10785 -1635 10800 -1615
rect 10750 -1650 10800 -1635
rect 11950 -965 12000 -950
rect 11950 -985 11965 -965
rect 11985 -985 12000 -965
rect 11950 -1015 12000 -985
rect 11950 -1035 11965 -1015
rect 11985 -1035 12000 -1015
rect 11950 -1065 12000 -1035
rect 11950 -1085 11965 -1065
rect 11985 -1085 12000 -1065
rect 11950 -1115 12000 -1085
rect 11950 -1135 11965 -1115
rect 11985 -1135 12000 -1115
rect 11950 -1165 12000 -1135
rect 11950 -1185 11965 -1165
rect 11985 -1185 12000 -1165
rect 11950 -1215 12000 -1185
rect 11950 -1235 11965 -1215
rect 11985 -1235 12000 -1215
rect 11950 -1265 12000 -1235
rect 11950 -1285 11965 -1265
rect 11985 -1285 12000 -1265
rect 11950 -1315 12000 -1285
rect 11950 -1335 11965 -1315
rect 11985 -1335 12000 -1315
rect 11950 -1365 12000 -1335
rect 11950 -1385 11965 -1365
rect 11985 -1385 12000 -1365
rect 11950 -1415 12000 -1385
rect 11950 -1435 11965 -1415
rect 11985 -1435 12000 -1415
rect 11950 -1465 12000 -1435
rect 11950 -1485 11965 -1465
rect 11985 -1485 12000 -1465
rect 11950 -1515 12000 -1485
rect 11950 -1535 11965 -1515
rect 11985 -1535 12000 -1515
rect 11950 -1565 12000 -1535
rect 11950 -1585 11965 -1565
rect 11985 -1585 12000 -1565
rect 11950 -1615 12000 -1585
rect 11950 -1635 11965 -1615
rect 11985 -1635 12000 -1615
rect 11950 -1650 12000 -1635
rect 12250 -965 12300 -950
rect 12250 -985 12265 -965
rect 12285 -985 12300 -965
rect 12250 -1015 12300 -985
rect 12250 -1035 12265 -1015
rect 12285 -1035 12300 -1015
rect 12250 -1065 12300 -1035
rect 12250 -1085 12265 -1065
rect 12285 -1085 12300 -1065
rect 12250 -1115 12300 -1085
rect 12250 -1135 12265 -1115
rect 12285 -1135 12300 -1115
rect 12250 -1165 12300 -1135
rect 12250 -1185 12265 -1165
rect 12285 -1185 12300 -1165
rect 12250 -1215 12300 -1185
rect 12250 -1235 12265 -1215
rect 12285 -1235 12300 -1215
rect 12250 -1265 12300 -1235
rect 12250 -1285 12265 -1265
rect 12285 -1285 12300 -1265
rect 12250 -1315 12300 -1285
rect 12250 -1335 12265 -1315
rect 12285 -1335 12300 -1315
rect 12250 -1365 12300 -1335
rect 12250 -1385 12265 -1365
rect 12285 -1385 12300 -1365
rect 12250 -1415 12300 -1385
rect 12250 -1435 12265 -1415
rect 12285 -1435 12300 -1415
rect 12250 -1465 12300 -1435
rect 12250 -1485 12265 -1465
rect 12285 -1485 12300 -1465
rect 12250 -1515 12300 -1485
rect 12250 -1535 12265 -1515
rect 12285 -1535 12300 -1515
rect 12250 -1565 12300 -1535
rect 12250 -1585 12265 -1565
rect 12285 -1585 12300 -1565
rect 12250 -1615 12300 -1585
rect 12250 -1635 12265 -1615
rect 12285 -1635 12300 -1615
rect 12250 -1650 12300 -1635
rect 12550 -965 12600 -950
rect 12550 -985 12565 -965
rect 12585 -985 12600 -965
rect 12550 -1015 12600 -985
rect 12550 -1035 12565 -1015
rect 12585 -1035 12600 -1015
rect 12550 -1065 12600 -1035
rect 12550 -1085 12565 -1065
rect 12585 -1085 12600 -1065
rect 12550 -1115 12600 -1085
rect 12550 -1135 12565 -1115
rect 12585 -1135 12600 -1115
rect 12550 -1165 12600 -1135
rect 12550 -1185 12565 -1165
rect 12585 -1185 12600 -1165
rect 12550 -1215 12600 -1185
rect 12550 -1235 12565 -1215
rect 12585 -1235 12600 -1215
rect 12550 -1265 12600 -1235
rect 12550 -1285 12565 -1265
rect 12585 -1285 12600 -1265
rect 12550 -1315 12600 -1285
rect 12550 -1335 12565 -1315
rect 12585 -1335 12600 -1315
rect 12550 -1365 12600 -1335
rect 12550 -1385 12565 -1365
rect 12585 -1385 12600 -1365
rect 12550 -1415 12600 -1385
rect 12550 -1435 12565 -1415
rect 12585 -1435 12600 -1415
rect 12550 -1465 12600 -1435
rect 12550 -1485 12565 -1465
rect 12585 -1485 12600 -1465
rect 12550 -1515 12600 -1485
rect 12550 -1535 12565 -1515
rect 12585 -1535 12600 -1515
rect 12550 -1565 12600 -1535
rect 12550 -1585 12565 -1565
rect 12585 -1585 12600 -1565
rect 12550 -1615 12600 -1585
rect 12550 -1635 12565 -1615
rect 12585 -1635 12600 -1615
rect 12550 -1650 12600 -1635
rect 12850 -965 12900 -950
rect 12850 -985 12865 -965
rect 12885 -985 12900 -965
rect 12850 -1015 12900 -985
rect 12850 -1035 12865 -1015
rect 12885 -1035 12900 -1015
rect 12850 -1065 12900 -1035
rect 12850 -1085 12865 -1065
rect 12885 -1085 12900 -1065
rect 12850 -1115 12900 -1085
rect 12850 -1135 12865 -1115
rect 12885 -1135 12900 -1115
rect 12850 -1165 12900 -1135
rect 12850 -1185 12865 -1165
rect 12885 -1185 12900 -1165
rect 12850 -1215 12900 -1185
rect 12850 -1235 12865 -1215
rect 12885 -1235 12900 -1215
rect 12850 -1265 12900 -1235
rect 12850 -1285 12865 -1265
rect 12885 -1285 12900 -1265
rect 12850 -1315 12900 -1285
rect 12850 -1335 12865 -1315
rect 12885 -1335 12900 -1315
rect 12850 -1365 12900 -1335
rect 12850 -1385 12865 -1365
rect 12885 -1385 12900 -1365
rect 12850 -1415 12900 -1385
rect 12850 -1435 12865 -1415
rect 12885 -1435 12900 -1415
rect 12850 -1465 12900 -1435
rect 12850 -1485 12865 -1465
rect 12885 -1485 12900 -1465
rect 12850 -1515 12900 -1485
rect 12850 -1535 12865 -1515
rect 12885 -1535 12900 -1515
rect 12850 -1565 12900 -1535
rect 12850 -1585 12865 -1565
rect 12885 -1585 12900 -1565
rect 12850 -1615 12900 -1585
rect 12850 -1635 12865 -1615
rect 12885 -1635 12900 -1615
rect 12850 -1650 12900 -1635
rect 13150 -965 13200 -950
rect 13150 -985 13165 -965
rect 13185 -985 13200 -965
rect 13150 -1015 13200 -985
rect 13150 -1035 13165 -1015
rect 13185 -1035 13200 -1015
rect 13150 -1065 13200 -1035
rect 13150 -1085 13165 -1065
rect 13185 -1085 13200 -1065
rect 13150 -1115 13200 -1085
rect 13150 -1135 13165 -1115
rect 13185 -1135 13200 -1115
rect 13150 -1165 13200 -1135
rect 13150 -1185 13165 -1165
rect 13185 -1185 13200 -1165
rect 13150 -1215 13200 -1185
rect 13150 -1235 13165 -1215
rect 13185 -1235 13200 -1215
rect 13150 -1265 13200 -1235
rect 13150 -1285 13165 -1265
rect 13185 -1285 13200 -1265
rect 13150 -1315 13200 -1285
rect 13150 -1335 13165 -1315
rect 13185 -1335 13200 -1315
rect 13150 -1365 13200 -1335
rect 13150 -1385 13165 -1365
rect 13185 -1385 13200 -1365
rect 13150 -1415 13200 -1385
rect 13150 -1435 13165 -1415
rect 13185 -1435 13200 -1415
rect 13150 -1465 13200 -1435
rect 13150 -1485 13165 -1465
rect 13185 -1485 13200 -1465
rect 13150 -1515 13200 -1485
rect 13150 -1535 13165 -1515
rect 13185 -1535 13200 -1515
rect 13150 -1565 13200 -1535
rect 13150 -1585 13165 -1565
rect 13185 -1585 13200 -1565
rect 13150 -1615 13200 -1585
rect 13150 -1635 13165 -1615
rect 13185 -1635 13200 -1615
rect 13150 -1650 13200 -1635
rect 13450 -965 13500 -950
rect 13450 -985 13465 -965
rect 13485 -985 13500 -965
rect 13450 -1015 13500 -985
rect 13450 -1035 13465 -1015
rect 13485 -1035 13500 -1015
rect 13450 -1065 13500 -1035
rect 13450 -1085 13465 -1065
rect 13485 -1085 13500 -1065
rect 13450 -1115 13500 -1085
rect 13450 -1135 13465 -1115
rect 13485 -1135 13500 -1115
rect 13450 -1165 13500 -1135
rect 13450 -1185 13465 -1165
rect 13485 -1185 13500 -1165
rect 13450 -1215 13500 -1185
rect 13450 -1235 13465 -1215
rect 13485 -1235 13500 -1215
rect 13450 -1265 13500 -1235
rect 13450 -1285 13465 -1265
rect 13485 -1285 13500 -1265
rect 13450 -1315 13500 -1285
rect 13450 -1335 13465 -1315
rect 13485 -1335 13500 -1315
rect 13450 -1365 13500 -1335
rect 13450 -1385 13465 -1365
rect 13485 -1385 13500 -1365
rect 13450 -1415 13500 -1385
rect 13450 -1435 13465 -1415
rect 13485 -1435 13500 -1415
rect 13450 -1465 13500 -1435
rect 13450 -1485 13465 -1465
rect 13485 -1485 13500 -1465
rect 13450 -1515 13500 -1485
rect 13450 -1535 13465 -1515
rect 13485 -1535 13500 -1515
rect 13450 -1565 13500 -1535
rect 13450 -1585 13465 -1565
rect 13485 -1585 13500 -1565
rect 13450 -1615 13500 -1585
rect 13450 -1635 13465 -1615
rect 13485 -1635 13500 -1615
rect 13450 -1650 13500 -1635
rect 13750 -965 13800 -950
rect 13750 -985 13765 -965
rect 13785 -985 13800 -965
rect 13750 -1015 13800 -985
rect 13750 -1035 13765 -1015
rect 13785 -1035 13800 -1015
rect 13750 -1065 13800 -1035
rect 13750 -1085 13765 -1065
rect 13785 -1085 13800 -1065
rect 13750 -1115 13800 -1085
rect 13750 -1135 13765 -1115
rect 13785 -1135 13800 -1115
rect 13750 -1165 13800 -1135
rect 13750 -1185 13765 -1165
rect 13785 -1185 13800 -1165
rect 13750 -1215 13800 -1185
rect 13750 -1235 13765 -1215
rect 13785 -1235 13800 -1215
rect 13750 -1265 13800 -1235
rect 13750 -1285 13765 -1265
rect 13785 -1285 13800 -1265
rect 13750 -1315 13800 -1285
rect 13750 -1335 13765 -1315
rect 13785 -1335 13800 -1315
rect 13750 -1365 13800 -1335
rect 13750 -1385 13765 -1365
rect 13785 -1385 13800 -1365
rect 13750 -1415 13800 -1385
rect 13750 -1435 13765 -1415
rect 13785 -1435 13800 -1415
rect 13750 -1465 13800 -1435
rect 13750 -1485 13765 -1465
rect 13785 -1485 13800 -1465
rect 13750 -1515 13800 -1485
rect 13750 -1535 13765 -1515
rect 13785 -1535 13800 -1515
rect 13750 -1565 13800 -1535
rect 13750 -1585 13765 -1565
rect 13785 -1585 13800 -1565
rect 13750 -1615 13800 -1585
rect 13750 -1635 13765 -1615
rect 13785 -1635 13800 -1615
rect 13750 -1650 13800 -1635
rect 14050 -965 14100 -950
rect 14050 -985 14065 -965
rect 14085 -985 14100 -965
rect 14050 -1015 14100 -985
rect 14050 -1035 14065 -1015
rect 14085 -1035 14100 -1015
rect 14050 -1065 14100 -1035
rect 14050 -1085 14065 -1065
rect 14085 -1085 14100 -1065
rect 14050 -1115 14100 -1085
rect 14050 -1135 14065 -1115
rect 14085 -1135 14100 -1115
rect 14050 -1165 14100 -1135
rect 14050 -1185 14065 -1165
rect 14085 -1185 14100 -1165
rect 14050 -1215 14100 -1185
rect 14050 -1235 14065 -1215
rect 14085 -1235 14100 -1215
rect 14050 -1265 14100 -1235
rect 14050 -1285 14065 -1265
rect 14085 -1285 14100 -1265
rect 14050 -1315 14100 -1285
rect 14050 -1335 14065 -1315
rect 14085 -1335 14100 -1315
rect 14050 -1365 14100 -1335
rect 14050 -1385 14065 -1365
rect 14085 -1385 14100 -1365
rect 14050 -1415 14100 -1385
rect 14050 -1435 14065 -1415
rect 14085 -1435 14100 -1415
rect 14050 -1465 14100 -1435
rect 14050 -1485 14065 -1465
rect 14085 -1485 14100 -1465
rect 14050 -1515 14100 -1485
rect 14050 -1535 14065 -1515
rect 14085 -1535 14100 -1515
rect 14050 -1565 14100 -1535
rect 14050 -1585 14065 -1565
rect 14085 -1585 14100 -1565
rect 14050 -1615 14100 -1585
rect 14050 -1635 14065 -1615
rect 14085 -1635 14100 -1615
rect 14050 -1650 14100 -1635
rect 14350 -965 14400 -950
rect 14350 -985 14365 -965
rect 14385 -985 14400 -965
rect 14350 -1015 14400 -985
rect 14350 -1035 14365 -1015
rect 14385 -1035 14400 -1015
rect 14350 -1065 14400 -1035
rect 14350 -1085 14365 -1065
rect 14385 -1085 14400 -1065
rect 14350 -1115 14400 -1085
rect 14350 -1135 14365 -1115
rect 14385 -1135 14400 -1115
rect 14350 -1165 14400 -1135
rect 14350 -1185 14365 -1165
rect 14385 -1185 14400 -1165
rect 14350 -1215 14400 -1185
rect 14350 -1235 14365 -1215
rect 14385 -1235 14400 -1215
rect 14350 -1265 14400 -1235
rect 14350 -1285 14365 -1265
rect 14385 -1285 14400 -1265
rect 14350 -1315 14400 -1285
rect 14350 -1335 14365 -1315
rect 14385 -1335 14400 -1315
rect 14350 -1365 14400 -1335
rect 14350 -1385 14365 -1365
rect 14385 -1385 14400 -1365
rect 14350 -1415 14400 -1385
rect 14350 -1435 14365 -1415
rect 14385 -1435 14400 -1415
rect 14350 -1465 14400 -1435
rect 14350 -1485 14365 -1465
rect 14385 -1485 14400 -1465
rect 14350 -1515 14400 -1485
rect 14350 -1535 14365 -1515
rect 14385 -1535 14400 -1515
rect 14350 -1565 14400 -1535
rect 14350 -1585 14365 -1565
rect 14385 -1585 14400 -1565
rect 14350 -1615 14400 -1585
rect 14350 -1635 14365 -1615
rect 14385 -1635 14400 -1615
rect 14350 -1650 14400 -1635
rect 15550 -965 15600 -950
rect 15550 -985 15565 -965
rect 15585 -985 15600 -965
rect 15550 -1015 15600 -985
rect 15550 -1035 15565 -1015
rect 15585 -1035 15600 -1015
rect 15550 -1065 15600 -1035
rect 15550 -1085 15565 -1065
rect 15585 -1085 15600 -1065
rect 15550 -1115 15600 -1085
rect 15550 -1135 15565 -1115
rect 15585 -1135 15600 -1115
rect 15550 -1165 15600 -1135
rect 15550 -1185 15565 -1165
rect 15585 -1185 15600 -1165
rect 15550 -1215 15600 -1185
rect 15550 -1235 15565 -1215
rect 15585 -1235 15600 -1215
rect 15550 -1265 15600 -1235
rect 15550 -1285 15565 -1265
rect 15585 -1285 15600 -1265
rect 15550 -1315 15600 -1285
rect 15550 -1335 15565 -1315
rect 15585 -1335 15600 -1315
rect 15550 -1365 15600 -1335
rect 15550 -1385 15565 -1365
rect 15585 -1385 15600 -1365
rect 15550 -1415 15600 -1385
rect 15550 -1435 15565 -1415
rect 15585 -1435 15600 -1415
rect 15550 -1465 15600 -1435
rect 15550 -1485 15565 -1465
rect 15585 -1485 15600 -1465
rect 15550 -1515 15600 -1485
rect 15550 -1535 15565 -1515
rect 15585 -1535 15600 -1515
rect 15550 -1565 15600 -1535
rect 15550 -1585 15565 -1565
rect 15585 -1585 15600 -1565
rect 15550 -1615 15600 -1585
rect 15550 -1635 15565 -1615
rect 15585 -1635 15600 -1615
rect 15550 -1650 15600 -1635
rect 16750 -965 16800 -950
rect 16750 -985 16765 -965
rect 16785 -985 16800 -965
rect 16750 -1015 16800 -985
rect 16750 -1035 16765 -1015
rect 16785 -1035 16800 -1015
rect 16750 -1065 16800 -1035
rect 16750 -1085 16765 -1065
rect 16785 -1085 16800 -1065
rect 16750 -1115 16800 -1085
rect 16750 -1135 16765 -1115
rect 16785 -1135 16800 -1115
rect 16750 -1165 16800 -1135
rect 16750 -1185 16765 -1165
rect 16785 -1185 16800 -1165
rect 16750 -1215 16800 -1185
rect 16750 -1235 16765 -1215
rect 16785 -1235 16800 -1215
rect 16750 -1265 16800 -1235
rect 16750 -1285 16765 -1265
rect 16785 -1285 16800 -1265
rect 16750 -1315 16800 -1285
rect 16750 -1335 16765 -1315
rect 16785 -1335 16800 -1315
rect 16750 -1365 16800 -1335
rect 16750 -1385 16765 -1365
rect 16785 -1385 16800 -1365
rect 16750 -1415 16800 -1385
rect 16750 -1435 16765 -1415
rect 16785 -1435 16800 -1415
rect 16750 -1465 16800 -1435
rect 16750 -1485 16765 -1465
rect 16785 -1485 16800 -1465
rect 16750 -1515 16800 -1485
rect 16750 -1535 16765 -1515
rect 16785 -1535 16800 -1515
rect 16750 -1565 16800 -1535
rect 16750 -1585 16765 -1565
rect 16785 -1585 16800 -1565
rect 16750 -1615 16800 -1585
rect 16750 -1635 16765 -1615
rect 16785 -1635 16800 -1615
rect 16750 -1650 16800 -1635
rect 17950 -965 18000 -950
rect 17950 -985 17965 -965
rect 17985 -985 18000 -965
rect 17950 -1015 18000 -985
rect 17950 -1035 17965 -1015
rect 17985 -1035 18000 -1015
rect 17950 -1065 18000 -1035
rect 17950 -1085 17965 -1065
rect 17985 -1085 18000 -1065
rect 17950 -1115 18000 -1085
rect 17950 -1135 17965 -1115
rect 17985 -1135 18000 -1115
rect 17950 -1165 18000 -1135
rect 17950 -1185 17965 -1165
rect 17985 -1185 18000 -1165
rect 17950 -1215 18000 -1185
rect 17950 -1235 17965 -1215
rect 17985 -1235 18000 -1215
rect 17950 -1265 18000 -1235
rect 17950 -1285 17965 -1265
rect 17985 -1285 18000 -1265
rect 17950 -1315 18000 -1285
rect 17950 -1335 17965 -1315
rect 17985 -1335 18000 -1315
rect 17950 -1365 18000 -1335
rect 17950 -1385 17965 -1365
rect 17985 -1385 18000 -1365
rect 17950 -1415 18000 -1385
rect 17950 -1435 17965 -1415
rect 17985 -1435 18000 -1415
rect 17950 -1465 18000 -1435
rect 17950 -1485 17965 -1465
rect 17985 -1485 18000 -1465
rect 17950 -1515 18000 -1485
rect 17950 -1535 17965 -1515
rect 17985 -1535 18000 -1515
rect 17950 -1565 18000 -1535
rect 17950 -1585 17965 -1565
rect 17985 -1585 18000 -1565
rect 17950 -1615 18000 -1585
rect 17950 -1635 17965 -1615
rect 17985 -1635 18000 -1615
rect 17950 -1650 18000 -1635
rect 19150 -965 19200 -950
rect 19150 -985 19165 -965
rect 19185 -985 19200 -965
rect 19150 -1015 19200 -985
rect 19150 -1035 19165 -1015
rect 19185 -1035 19200 -1015
rect 19150 -1065 19200 -1035
rect 19150 -1085 19165 -1065
rect 19185 -1085 19200 -1065
rect 19150 -1115 19200 -1085
rect 19150 -1135 19165 -1115
rect 19185 -1135 19200 -1115
rect 19150 -1165 19200 -1135
rect 19150 -1185 19165 -1165
rect 19185 -1185 19200 -1165
rect 19150 -1215 19200 -1185
rect 19150 -1235 19165 -1215
rect 19185 -1235 19200 -1215
rect 19150 -1265 19200 -1235
rect 19150 -1285 19165 -1265
rect 19185 -1285 19200 -1265
rect 19150 -1315 19200 -1285
rect 19150 -1335 19165 -1315
rect 19185 -1335 19200 -1315
rect 19150 -1365 19200 -1335
rect 19150 -1385 19165 -1365
rect 19185 -1385 19200 -1365
rect 19150 -1415 19200 -1385
rect 19150 -1435 19165 -1415
rect 19185 -1435 19200 -1415
rect 19150 -1465 19200 -1435
rect 19150 -1485 19165 -1465
rect 19185 -1485 19200 -1465
rect 19150 -1515 19200 -1485
rect 19150 -1535 19165 -1515
rect 19185 -1535 19200 -1515
rect 19150 -1565 19200 -1535
rect 19150 -1585 19165 -1565
rect 19185 -1585 19200 -1565
rect 19150 -1615 19200 -1585
rect 19150 -1635 19165 -1615
rect 19185 -1635 19200 -1615
rect 19150 -1650 19200 -1635
rect 20350 -965 20400 -950
rect 20350 -985 20365 -965
rect 20385 -985 20400 -965
rect 20350 -1015 20400 -985
rect 20350 -1035 20365 -1015
rect 20385 -1035 20400 -1015
rect 20350 -1065 20400 -1035
rect 20350 -1085 20365 -1065
rect 20385 -1085 20400 -1065
rect 20350 -1115 20400 -1085
rect 20350 -1135 20365 -1115
rect 20385 -1135 20400 -1115
rect 20350 -1165 20400 -1135
rect 20350 -1185 20365 -1165
rect 20385 -1185 20400 -1165
rect 20350 -1215 20400 -1185
rect 20350 -1235 20365 -1215
rect 20385 -1235 20400 -1215
rect 20350 -1265 20400 -1235
rect 20350 -1285 20365 -1265
rect 20385 -1285 20400 -1265
rect 20350 -1315 20400 -1285
rect 20350 -1335 20365 -1315
rect 20385 -1335 20400 -1315
rect 20350 -1365 20400 -1335
rect 20350 -1385 20365 -1365
rect 20385 -1385 20400 -1365
rect 20350 -1415 20400 -1385
rect 20350 -1435 20365 -1415
rect 20385 -1435 20400 -1415
rect 20350 -1465 20400 -1435
rect 20350 -1485 20365 -1465
rect 20385 -1485 20400 -1465
rect 20350 -1515 20400 -1485
rect 20350 -1535 20365 -1515
rect 20385 -1535 20400 -1515
rect 20350 -1565 20400 -1535
rect 20350 -1585 20365 -1565
rect 20385 -1585 20400 -1565
rect 20350 -1615 20400 -1585
rect 20350 -1635 20365 -1615
rect 20385 -1635 20400 -1615
rect 20350 -1650 20400 -1635
rect -650 -1715 20400 -1700
rect -650 -1735 -635 -1715
rect -615 -1735 -585 -1715
rect -565 -1735 -535 -1715
rect -515 -1735 -485 -1715
rect -465 -1735 -435 -1715
rect -415 -1735 -385 -1715
rect -365 -1735 -335 -1715
rect -315 -1735 -285 -1715
rect -265 -1735 -235 -1715
rect -215 -1735 -185 -1715
rect -165 -1735 -135 -1715
rect -115 -1735 -85 -1715
rect -65 -1735 -35 -1715
rect -15 -1735 15 -1715
rect 35 -1735 65 -1715
rect 85 -1735 115 -1715
rect 135 -1735 165 -1715
rect 185 -1735 215 -1715
rect 235 -1735 265 -1715
rect 285 -1735 315 -1715
rect 335 -1735 365 -1715
rect 385 -1735 415 -1715
rect 435 -1735 465 -1715
rect 485 -1735 515 -1715
rect 535 -1735 565 -1715
rect 585 -1735 615 -1715
rect 635 -1735 665 -1715
rect 685 -1735 715 -1715
rect 735 -1735 765 -1715
rect 785 -1735 815 -1715
rect 835 -1735 865 -1715
rect 885 -1735 915 -1715
rect 935 -1735 965 -1715
rect 985 -1735 1015 -1715
rect 1035 -1735 1065 -1715
rect 1085 -1735 1115 -1715
rect 1135 -1735 1165 -1715
rect 1185 -1735 1215 -1715
rect 1235 -1735 1265 -1715
rect 1285 -1735 1315 -1715
rect 1335 -1735 1365 -1715
rect 1385 -1735 1415 -1715
rect 1435 -1735 1465 -1715
rect 1485 -1735 1515 -1715
rect 1535 -1735 1565 -1715
rect 1585 -1735 1615 -1715
rect 1635 -1735 1665 -1715
rect 1685 -1735 1715 -1715
rect 1735 -1735 1765 -1715
rect 1785 -1735 1815 -1715
rect 1835 -1735 1865 -1715
rect 1885 -1735 1915 -1715
rect 1935 -1735 1965 -1715
rect 1985 -1735 2015 -1715
rect 2035 -1735 2065 -1715
rect 2085 -1735 2115 -1715
rect 2135 -1735 2165 -1715
rect 2185 -1735 2215 -1715
rect 2235 -1735 2265 -1715
rect 2285 -1735 2315 -1715
rect 2335 -1735 2365 -1715
rect 2385 -1735 2415 -1715
rect 2435 -1735 2465 -1715
rect 2485 -1735 2515 -1715
rect 2535 -1735 2565 -1715
rect 2585 -1735 2615 -1715
rect 2635 -1735 2665 -1715
rect 2685 -1735 2715 -1715
rect 2735 -1735 2765 -1715
rect 2785 -1735 2815 -1715
rect 2835 -1735 2865 -1715
rect 2885 -1735 2915 -1715
rect 2935 -1735 2965 -1715
rect 2985 -1735 3015 -1715
rect 3035 -1735 3065 -1715
rect 3085 -1735 3115 -1715
rect 3135 -1735 3165 -1715
rect 3185 -1735 3215 -1715
rect 3235 -1735 3265 -1715
rect 3285 -1735 3315 -1715
rect 3335 -1735 3365 -1715
rect 3385 -1735 3415 -1715
rect 3435 -1735 3465 -1715
rect 3485 -1735 3515 -1715
rect 3535 -1735 3565 -1715
rect 3585 -1735 3615 -1715
rect 3635 -1735 3665 -1715
rect 3685 -1735 3715 -1715
rect 3735 -1735 3765 -1715
rect 3785 -1735 3815 -1715
rect 3835 -1735 3865 -1715
rect 3885 -1735 3915 -1715
rect 3935 -1735 3965 -1715
rect 3985 -1735 4015 -1715
rect 4035 -1735 4065 -1715
rect 4085 -1735 4115 -1715
rect 4135 -1735 4165 -1715
rect 4185 -1735 4215 -1715
rect 4235 -1735 4265 -1715
rect 4285 -1735 4315 -1715
rect 4335 -1735 4365 -1715
rect 4385 -1735 4415 -1715
rect 4435 -1735 4465 -1715
rect 4485 -1735 4515 -1715
rect 4535 -1735 4565 -1715
rect 4585 -1735 4615 -1715
rect 4635 -1735 4665 -1715
rect 4685 -1735 4715 -1715
rect 4735 -1735 4765 -1715
rect 4785 -1735 4815 -1715
rect 4835 -1735 4865 -1715
rect 4885 -1735 4915 -1715
rect 4935 -1735 4965 -1715
rect 4985 -1735 5015 -1715
rect 5035 -1735 5065 -1715
rect 5085 -1735 5115 -1715
rect 5135 -1735 5165 -1715
rect 5185 -1735 5215 -1715
rect 5235 -1735 5265 -1715
rect 5285 -1735 5315 -1715
rect 5335 -1735 5365 -1715
rect 5385 -1735 5415 -1715
rect 5435 -1735 5465 -1715
rect 5485 -1735 5515 -1715
rect 5535 -1735 5565 -1715
rect 5585 -1735 5615 -1715
rect 5635 -1735 5665 -1715
rect 5685 -1735 5715 -1715
rect 5735 -1735 5765 -1715
rect 5785 -1735 5815 -1715
rect 5835 -1735 5865 -1715
rect 5885 -1735 5915 -1715
rect 5935 -1735 5965 -1715
rect 5985 -1735 6015 -1715
rect 6035 -1735 6065 -1715
rect 6085 -1735 6115 -1715
rect 6135 -1735 6165 -1715
rect 6185 -1735 6215 -1715
rect 6235 -1735 6265 -1715
rect 6285 -1735 6315 -1715
rect 6335 -1735 6365 -1715
rect 6385 -1735 6415 -1715
rect 6435 -1735 6465 -1715
rect 6485 -1735 6515 -1715
rect 6535 -1735 6565 -1715
rect 6585 -1735 6615 -1715
rect 6635 -1735 6665 -1715
rect 6685 -1735 6715 -1715
rect 6735 -1735 6765 -1715
rect 6785 -1735 6815 -1715
rect 6835 -1735 6865 -1715
rect 6885 -1735 6915 -1715
rect 6935 -1735 6965 -1715
rect 6985 -1735 7015 -1715
rect 7035 -1735 7065 -1715
rect 7085 -1735 7115 -1715
rect 7135 -1735 7165 -1715
rect 7185 -1735 7215 -1715
rect 7235 -1735 7265 -1715
rect 7285 -1735 7315 -1715
rect 7335 -1735 7365 -1715
rect 7385 -1735 7415 -1715
rect 7435 -1735 7465 -1715
rect 7485 -1735 7515 -1715
rect 7535 -1735 7565 -1715
rect 7585 -1735 7615 -1715
rect 7635 -1735 7665 -1715
rect 7685 -1735 7715 -1715
rect 7735 -1735 7765 -1715
rect 7785 -1735 7815 -1715
rect 7835 -1735 7865 -1715
rect 7885 -1735 7915 -1715
rect 7935 -1735 7965 -1715
rect 7985 -1735 8015 -1715
rect 8035 -1735 8065 -1715
rect 8085 -1735 8115 -1715
rect 8135 -1735 8165 -1715
rect 8185 -1735 8215 -1715
rect 8235 -1735 8265 -1715
rect 8285 -1735 8315 -1715
rect 8335 -1735 8365 -1715
rect 8385 -1735 8415 -1715
rect 8435 -1735 8465 -1715
rect 8485 -1735 8515 -1715
rect 8535 -1735 8565 -1715
rect 8585 -1735 8615 -1715
rect 8635 -1735 8665 -1715
rect 8685 -1735 8715 -1715
rect 8735 -1735 8765 -1715
rect 8785 -1735 8815 -1715
rect 8835 -1735 8865 -1715
rect 8885 -1735 8915 -1715
rect 8935 -1735 8965 -1715
rect 8985 -1735 9015 -1715
rect 9035 -1735 9065 -1715
rect 9085 -1735 9115 -1715
rect 9135 -1735 9165 -1715
rect 9185 -1735 9215 -1715
rect 9235 -1735 9265 -1715
rect 9285 -1735 9315 -1715
rect 9335 -1735 9365 -1715
rect 9385 -1735 9415 -1715
rect 9435 -1735 9465 -1715
rect 9485 -1735 9515 -1715
rect 9535 -1735 9565 -1715
rect 9585 -1735 9615 -1715
rect 9635 -1735 9665 -1715
rect 9685 -1735 9715 -1715
rect 9735 -1735 9765 -1715
rect 9785 -1735 9815 -1715
rect 9835 -1735 9865 -1715
rect 9885 -1735 9915 -1715
rect 9935 -1735 9965 -1715
rect 9985 -1735 10015 -1715
rect 10035 -1735 10065 -1715
rect 10085 -1735 10115 -1715
rect 10135 -1735 10165 -1715
rect 10185 -1735 10215 -1715
rect 10235 -1735 10265 -1715
rect 10285 -1735 10315 -1715
rect 10335 -1735 10365 -1715
rect 10385 -1735 10415 -1715
rect 10435 -1735 10465 -1715
rect 10485 -1735 10515 -1715
rect 10535 -1735 10565 -1715
rect 10585 -1735 10615 -1715
rect 10635 -1735 10665 -1715
rect 10685 -1735 10715 -1715
rect 10735 -1735 10765 -1715
rect 10785 -1735 10815 -1715
rect 10835 -1735 10865 -1715
rect 10885 -1735 10915 -1715
rect 10935 -1735 10965 -1715
rect 10985 -1735 11015 -1715
rect 11035 -1735 11065 -1715
rect 11085 -1735 11115 -1715
rect 11135 -1735 11165 -1715
rect 11185 -1735 11215 -1715
rect 11235 -1735 11265 -1715
rect 11285 -1735 11315 -1715
rect 11335 -1735 11365 -1715
rect 11385 -1735 11415 -1715
rect 11435 -1735 11465 -1715
rect 11485 -1735 11515 -1715
rect 11535 -1735 11565 -1715
rect 11585 -1735 11615 -1715
rect 11635 -1735 11665 -1715
rect 11685 -1735 11715 -1715
rect 11735 -1735 11765 -1715
rect 11785 -1735 11815 -1715
rect 11835 -1735 11865 -1715
rect 11885 -1735 11915 -1715
rect 11935 -1735 11965 -1715
rect 11985 -1735 12015 -1715
rect 12035 -1735 12065 -1715
rect 12085 -1735 12115 -1715
rect 12135 -1735 12165 -1715
rect 12185 -1735 12215 -1715
rect 12235 -1735 12265 -1715
rect 12285 -1735 12315 -1715
rect 12335 -1735 12365 -1715
rect 12385 -1735 12415 -1715
rect 12435 -1735 12465 -1715
rect 12485 -1735 12515 -1715
rect 12535 -1735 12565 -1715
rect 12585 -1735 12615 -1715
rect 12635 -1735 12665 -1715
rect 12685 -1735 12715 -1715
rect 12735 -1735 12765 -1715
rect 12785 -1735 12815 -1715
rect 12835 -1735 12865 -1715
rect 12885 -1735 12915 -1715
rect 12935 -1735 12965 -1715
rect 12985 -1735 13015 -1715
rect 13035 -1735 13065 -1715
rect 13085 -1735 13115 -1715
rect 13135 -1735 13165 -1715
rect 13185 -1735 13215 -1715
rect 13235 -1735 13265 -1715
rect 13285 -1735 13315 -1715
rect 13335 -1735 13365 -1715
rect 13385 -1735 13415 -1715
rect 13435 -1735 13465 -1715
rect 13485 -1735 13515 -1715
rect 13535 -1735 13565 -1715
rect 13585 -1735 13615 -1715
rect 13635 -1735 13665 -1715
rect 13685 -1735 13715 -1715
rect 13735 -1735 13765 -1715
rect 13785 -1735 13815 -1715
rect 13835 -1735 13865 -1715
rect 13885 -1735 13915 -1715
rect 13935 -1735 13965 -1715
rect 13985 -1735 14015 -1715
rect 14035 -1735 14065 -1715
rect 14085 -1735 14115 -1715
rect 14135 -1735 14165 -1715
rect 14185 -1735 14215 -1715
rect 14235 -1735 14265 -1715
rect 14285 -1735 14315 -1715
rect 14335 -1735 14365 -1715
rect 14385 -1735 14415 -1715
rect 14435 -1735 14465 -1715
rect 14485 -1735 14515 -1715
rect 14535 -1735 14565 -1715
rect 14585 -1735 14615 -1715
rect 14635 -1735 14665 -1715
rect 14685 -1735 14715 -1715
rect 14735 -1735 14765 -1715
rect 14785 -1735 14815 -1715
rect 14835 -1735 14865 -1715
rect 14885 -1735 14915 -1715
rect 14935 -1735 14965 -1715
rect 14985 -1735 15015 -1715
rect 15035 -1735 15065 -1715
rect 15085 -1735 15115 -1715
rect 15135 -1735 15165 -1715
rect 15185 -1735 15215 -1715
rect 15235 -1735 15265 -1715
rect 15285 -1735 15315 -1715
rect 15335 -1735 15365 -1715
rect 15385 -1735 15415 -1715
rect 15435 -1735 15465 -1715
rect 15485 -1735 15515 -1715
rect 15535 -1735 15565 -1715
rect 15585 -1735 15615 -1715
rect 15635 -1735 15665 -1715
rect 15685 -1735 15715 -1715
rect 15735 -1735 15765 -1715
rect 15785 -1735 15815 -1715
rect 15835 -1735 15865 -1715
rect 15885 -1735 15915 -1715
rect 15935 -1735 15965 -1715
rect 15985 -1735 16015 -1715
rect 16035 -1735 16065 -1715
rect 16085 -1735 16115 -1715
rect 16135 -1735 16165 -1715
rect 16185 -1735 16215 -1715
rect 16235 -1735 16265 -1715
rect 16285 -1735 16315 -1715
rect 16335 -1735 16365 -1715
rect 16385 -1735 16415 -1715
rect 16435 -1735 16465 -1715
rect 16485 -1735 16515 -1715
rect 16535 -1735 16565 -1715
rect 16585 -1735 16615 -1715
rect 16635 -1735 16665 -1715
rect 16685 -1735 16715 -1715
rect 16735 -1735 16765 -1715
rect 16785 -1735 16815 -1715
rect 16835 -1735 16865 -1715
rect 16885 -1735 16915 -1715
rect 16935 -1735 16965 -1715
rect 16985 -1735 17015 -1715
rect 17035 -1735 17065 -1715
rect 17085 -1735 17115 -1715
rect 17135 -1735 17165 -1715
rect 17185 -1735 17215 -1715
rect 17235 -1735 17265 -1715
rect 17285 -1735 17315 -1715
rect 17335 -1735 17365 -1715
rect 17385 -1735 17415 -1715
rect 17435 -1735 17465 -1715
rect 17485 -1735 17515 -1715
rect 17535 -1735 17565 -1715
rect 17585 -1735 17615 -1715
rect 17635 -1735 17665 -1715
rect 17685 -1735 17715 -1715
rect 17735 -1735 17765 -1715
rect 17785 -1735 17815 -1715
rect 17835 -1735 17865 -1715
rect 17885 -1735 17915 -1715
rect 17935 -1735 17965 -1715
rect 17985 -1735 18015 -1715
rect 18035 -1735 18065 -1715
rect 18085 -1735 18115 -1715
rect 18135 -1735 18165 -1715
rect 18185 -1735 18215 -1715
rect 18235 -1735 18265 -1715
rect 18285 -1735 18315 -1715
rect 18335 -1735 18365 -1715
rect 18385 -1735 18415 -1715
rect 18435 -1735 18465 -1715
rect 18485 -1735 18515 -1715
rect 18535 -1735 18565 -1715
rect 18585 -1735 18615 -1715
rect 18635 -1735 18665 -1715
rect 18685 -1735 18715 -1715
rect 18735 -1735 18765 -1715
rect 18785 -1735 18815 -1715
rect 18835 -1735 18865 -1715
rect 18885 -1735 18915 -1715
rect 18935 -1735 18965 -1715
rect 18985 -1735 19015 -1715
rect 19035 -1735 19065 -1715
rect 19085 -1735 19115 -1715
rect 19135 -1735 19165 -1715
rect 19185 -1735 19215 -1715
rect 19235 -1735 19265 -1715
rect 19285 -1735 19315 -1715
rect 19335 -1735 19365 -1715
rect 19385 -1735 19415 -1715
rect 19435 -1735 19465 -1715
rect 19485 -1735 19515 -1715
rect 19535 -1735 19565 -1715
rect 19585 -1735 19615 -1715
rect 19635 -1735 19665 -1715
rect 19685 -1735 19715 -1715
rect 19735 -1735 19765 -1715
rect 19785 -1735 19815 -1715
rect 19835 -1735 19865 -1715
rect 19885 -1735 19915 -1715
rect 19935 -1735 19965 -1715
rect 19985 -1735 20015 -1715
rect 20035 -1735 20065 -1715
rect 20085 -1735 20115 -1715
rect 20135 -1735 20165 -1715
rect 20185 -1735 20215 -1715
rect 20235 -1735 20265 -1715
rect 20285 -1735 20315 -1715
rect 20335 -1735 20365 -1715
rect 20385 -1735 20400 -1715
rect -650 -1750 20400 -1735
rect -650 -1865 20400 -1850
rect -650 -1885 -635 -1865
rect -615 -1885 -585 -1865
rect -565 -1885 -535 -1865
rect -515 -1885 -485 -1865
rect -465 -1885 -435 -1865
rect -415 -1885 -385 -1865
rect -365 -1885 -335 -1865
rect -315 -1885 -285 -1865
rect -265 -1885 -235 -1865
rect -215 -1885 -185 -1865
rect -165 -1885 -135 -1865
rect -115 -1885 -85 -1865
rect -65 -1885 -35 -1865
rect -15 -1885 15 -1865
rect 35 -1885 65 -1865
rect 85 -1885 115 -1865
rect 135 -1885 165 -1865
rect 185 -1885 215 -1865
rect 235 -1885 265 -1865
rect 285 -1885 315 -1865
rect 335 -1885 365 -1865
rect 385 -1885 415 -1865
rect 435 -1885 465 -1865
rect 485 -1885 515 -1865
rect 535 -1885 565 -1865
rect 585 -1885 615 -1865
rect 635 -1885 665 -1865
rect 685 -1885 715 -1865
rect 735 -1885 765 -1865
rect 785 -1885 815 -1865
rect 835 -1885 865 -1865
rect 885 -1885 915 -1865
rect 935 -1885 965 -1865
rect 985 -1885 1015 -1865
rect 1035 -1885 1065 -1865
rect 1085 -1885 1115 -1865
rect 1135 -1885 1165 -1865
rect 1185 -1885 1215 -1865
rect 1235 -1885 1265 -1865
rect 1285 -1885 1315 -1865
rect 1335 -1885 1365 -1865
rect 1385 -1885 1415 -1865
rect 1435 -1885 1465 -1865
rect 1485 -1885 1515 -1865
rect 1535 -1885 1565 -1865
rect 1585 -1885 1615 -1865
rect 1635 -1885 1665 -1865
rect 1685 -1885 1715 -1865
rect 1735 -1885 1765 -1865
rect 1785 -1885 1815 -1865
rect 1835 -1885 1865 -1865
rect 1885 -1885 1915 -1865
rect 1935 -1885 1965 -1865
rect 1985 -1885 2015 -1865
rect 2035 -1885 2065 -1865
rect 2085 -1885 2115 -1865
rect 2135 -1885 2165 -1865
rect 2185 -1885 2215 -1865
rect 2235 -1885 2265 -1865
rect 2285 -1885 2315 -1865
rect 2335 -1885 2365 -1865
rect 2385 -1885 2415 -1865
rect 2435 -1885 2465 -1865
rect 2485 -1885 2515 -1865
rect 2535 -1885 2565 -1865
rect 2585 -1885 2615 -1865
rect 2635 -1885 2665 -1865
rect 2685 -1885 2715 -1865
rect 2735 -1885 2765 -1865
rect 2785 -1885 2815 -1865
rect 2835 -1885 2865 -1865
rect 2885 -1885 2915 -1865
rect 2935 -1885 2965 -1865
rect 2985 -1885 3015 -1865
rect 3035 -1885 3065 -1865
rect 3085 -1885 3115 -1865
rect 3135 -1885 3165 -1865
rect 3185 -1885 3215 -1865
rect 3235 -1885 3265 -1865
rect 3285 -1885 3315 -1865
rect 3335 -1885 3365 -1865
rect 3385 -1885 3415 -1865
rect 3435 -1885 3465 -1865
rect 3485 -1885 3515 -1865
rect 3535 -1885 3565 -1865
rect 3585 -1885 3615 -1865
rect 3635 -1885 3665 -1865
rect 3685 -1885 3715 -1865
rect 3735 -1885 3765 -1865
rect 3785 -1885 3815 -1865
rect 3835 -1885 3865 -1865
rect 3885 -1885 3915 -1865
rect 3935 -1885 3965 -1865
rect 3985 -1885 4015 -1865
rect 4035 -1885 4065 -1865
rect 4085 -1885 4115 -1865
rect 4135 -1885 4165 -1865
rect 4185 -1885 4215 -1865
rect 4235 -1885 4265 -1865
rect 4285 -1885 4315 -1865
rect 4335 -1885 4365 -1865
rect 4385 -1885 4415 -1865
rect 4435 -1885 4465 -1865
rect 4485 -1885 4515 -1865
rect 4535 -1885 4565 -1865
rect 4585 -1885 4615 -1865
rect 4635 -1885 4665 -1865
rect 4685 -1885 4715 -1865
rect 4735 -1885 4765 -1865
rect 4785 -1885 4815 -1865
rect 4835 -1885 4865 -1865
rect 4885 -1885 4915 -1865
rect 4935 -1885 4965 -1865
rect 4985 -1885 5015 -1865
rect 5035 -1885 5065 -1865
rect 5085 -1885 5115 -1865
rect 5135 -1885 5165 -1865
rect 5185 -1885 5215 -1865
rect 5235 -1885 5265 -1865
rect 5285 -1885 5315 -1865
rect 5335 -1885 5365 -1865
rect 5385 -1885 5415 -1865
rect 5435 -1885 5465 -1865
rect 5485 -1885 5515 -1865
rect 5535 -1885 5565 -1865
rect 5585 -1885 5615 -1865
rect 5635 -1885 5665 -1865
rect 5685 -1885 5715 -1865
rect 5735 -1885 5765 -1865
rect 5785 -1885 5815 -1865
rect 5835 -1885 5865 -1865
rect 5885 -1885 5915 -1865
rect 5935 -1885 5965 -1865
rect 5985 -1885 6015 -1865
rect 6035 -1885 6065 -1865
rect 6085 -1885 6115 -1865
rect 6135 -1885 6165 -1865
rect 6185 -1885 6215 -1865
rect 6235 -1885 6265 -1865
rect 6285 -1885 6315 -1865
rect 6335 -1885 6365 -1865
rect 6385 -1885 6415 -1865
rect 6435 -1885 6465 -1865
rect 6485 -1885 6515 -1865
rect 6535 -1885 6565 -1865
rect 6585 -1885 6615 -1865
rect 6635 -1885 6665 -1865
rect 6685 -1885 6715 -1865
rect 6735 -1885 6765 -1865
rect 6785 -1885 6815 -1865
rect 6835 -1885 6865 -1865
rect 6885 -1885 6915 -1865
rect 6935 -1885 6965 -1865
rect 6985 -1885 7015 -1865
rect 7035 -1885 7065 -1865
rect 7085 -1885 7115 -1865
rect 7135 -1885 7165 -1865
rect 7185 -1885 7215 -1865
rect 7235 -1885 7265 -1865
rect 7285 -1885 7315 -1865
rect 7335 -1885 7365 -1865
rect 7385 -1885 7415 -1865
rect 7435 -1885 7465 -1865
rect 7485 -1885 7515 -1865
rect 7535 -1885 7565 -1865
rect 7585 -1885 7615 -1865
rect 7635 -1885 7665 -1865
rect 7685 -1885 7715 -1865
rect 7735 -1885 7765 -1865
rect 7785 -1885 7815 -1865
rect 7835 -1885 7865 -1865
rect 7885 -1885 7915 -1865
rect 7935 -1885 7965 -1865
rect 7985 -1885 8015 -1865
rect 8035 -1885 8065 -1865
rect 8085 -1885 8115 -1865
rect 8135 -1885 8165 -1865
rect 8185 -1885 8215 -1865
rect 8235 -1885 8265 -1865
rect 8285 -1885 8315 -1865
rect 8335 -1885 8365 -1865
rect 8385 -1885 8415 -1865
rect 8435 -1885 8465 -1865
rect 8485 -1885 8515 -1865
rect 8535 -1885 8565 -1865
rect 8585 -1885 8615 -1865
rect 8635 -1885 8665 -1865
rect 8685 -1885 8715 -1865
rect 8735 -1885 8765 -1865
rect 8785 -1885 8815 -1865
rect 8835 -1885 8865 -1865
rect 8885 -1885 8915 -1865
rect 8935 -1885 8965 -1865
rect 8985 -1885 9015 -1865
rect 9035 -1885 9065 -1865
rect 9085 -1885 9115 -1865
rect 9135 -1885 9165 -1865
rect 9185 -1885 9215 -1865
rect 9235 -1885 9265 -1865
rect 9285 -1885 9315 -1865
rect 9335 -1885 9365 -1865
rect 9385 -1885 9415 -1865
rect 9435 -1885 9465 -1865
rect 9485 -1885 9515 -1865
rect 9535 -1885 9565 -1865
rect 9585 -1885 9615 -1865
rect 9635 -1885 9665 -1865
rect 9685 -1885 9715 -1865
rect 9735 -1885 9765 -1865
rect 9785 -1885 9815 -1865
rect 9835 -1885 9865 -1865
rect 9885 -1885 9915 -1865
rect 9935 -1885 9965 -1865
rect 9985 -1885 10015 -1865
rect 10035 -1885 10065 -1865
rect 10085 -1885 10115 -1865
rect 10135 -1885 10165 -1865
rect 10185 -1885 10215 -1865
rect 10235 -1885 10265 -1865
rect 10285 -1885 10315 -1865
rect 10335 -1885 10365 -1865
rect 10385 -1885 10415 -1865
rect 10435 -1885 10465 -1865
rect 10485 -1885 10515 -1865
rect 10535 -1885 10565 -1865
rect 10585 -1885 10615 -1865
rect 10635 -1885 10665 -1865
rect 10685 -1885 10715 -1865
rect 10735 -1885 10765 -1865
rect 10785 -1885 10815 -1865
rect 10835 -1885 10865 -1865
rect 10885 -1885 10915 -1865
rect 10935 -1885 10965 -1865
rect 10985 -1885 11015 -1865
rect 11035 -1885 11065 -1865
rect 11085 -1885 11115 -1865
rect 11135 -1885 11165 -1865
rect 11185 -1885 11215 -1865
rect 11235 -1885 11265 -1865
rect 11285 -1885 11315 -1865
rect 11335 -1885 11365 -1865
rect 11385 -1885 11415 -1865
rect 11435 -1885 11465 -1865
rect 11485 -1885 11515 -1865
rect 11535 -1885 11565 -1865
rect 11585 -1885 11615 -1865
rect 11635 -1885 11665 -1865
rect 11685 -1885 11715 -1865
rect 11735 -1885 11765 -1865
rect 11785 -1885 11815 -1865
rect 11835 -1885 11865 -1865
rect 11885 -1885 11915 -1865
rect 11935 -1885 11965 -1865
rect 11985 -1885 12015 -1865
rect 12035 -1885 12065 -1865
rect 12085 -1885 12115 -1865
rect 12135 -1885 12165 -1865
rect 12185 -1885 12215 -1865
rect 12235 -1885 12265 -1865
rect 12285 -1885 12315 -1865
rect 12335 -1885 12365 -1865
rect 12385 -1885 12415 -1865
rect 12435 -1885 12465 -1865
rect 12485 -1885 12515 -1865
rect 12535 -1885 12565 -1865
rect 12585 -1885 12615 -1865
rect 12635 -1885 12665 -1865
rect 12685 -1885 12715 -1865
rect 12735 -1885 12765 -1865
rect 12785 -1885 12815 -1865
rect 12835 -1885 12865 -1865
rect 12885 -1885 12915 -1865
rect 12935 -1885 12965 -1865
rect 12985 -1885 13015 -1865
rect 13035 -1885 13065 -1865
rect 13085 -1885 13115 -1865
rect 13135 -1885 13165 -1865
rect 13185 -1885 13215 -1865
rect 13235 -1885 13265 -1865
rect 13285 -1885 13315 -1865
rect 13335 -1885 13365 -1865
rect 13385 -1885 13415 -1865
rect 13435 -1885 13465 -1865
rect 13485 -1885 13515 -1865
rect 13535 -1885 13565 -1865
rect 13585 -1885 13615 -1865
rect 13635 -1885 13665 -1865
rect 13685 -1885 13715 -1865
rect 13735 -1885 13765 -1865
rect 13785 -1885 13815 -1865
rect 13835 -1885 13865 -1865
rect 13885 -1885 13915 -1865
rect 13935 -1885 13965 -1865
rect 13985 -1885 14015 -1865
rect 14035 -1885 14065 -1865
rect 14085 -1885 14115 -1865
rect 14135 -1885 14165 -1865
rect 14185 -1885 14215 -1865
rect 14235 -1885 14265 -1865
rect 14285 -1885 14315 -1865
rect 14335 -1885 14365 -1865
rect 14385 -1885 14415 -1865
rect 14435 -1885 14465 -1865
rect 14485 -1885 14515 -1865
rect 14535 -1885 14565 -1865
rect 14585 -1885 14615 -1865
rect 14635 -1885 14665 -1865
rect 14685 -1885 14715 -1865
rect 14735 -1885 14765 -1865
rect 14785 -1885 14815 -1865
rect 14835 -1885 14865 -1865
rect 14885 -1885 14915 -1865
rect 14935 -1885 14965 -1865
rect 14985 -1885 15015 -1865
rect 15035 -1885 15065 -1865
rect 15085 -1885 15115 -1865
rect 15135 -1885 15165 -1865
rect 15185 -1885 15215 -1865
rect 15235 -1885 15265 -1865
rect 15285 -1885 15315 -1865
rect 15335 -1885 15365 -1865
rect 15385 -1885 15415 -1865
rect 15435 -1885 15465 -1865
rect 15485 -1885 15515 -1865
rect 15535 -1885 15565 -1865
rect 15585 -1885 15615 -1865
rect 15635 -1885 15665 -1865
rect 15685 -1885 15715 -1865
rect 15735 -1885 15765 -1865
rect 15785 -1885 15815 -1865
rect 15835 -1885 15865 -1865
rect 15885 -1885 15915 -1865
rect 15935 -1885 15965 -1865
rect 15985 -1885 16015 -1865
rect 16035 -1885 16065 -1865
rect 16085 -1885 16115 -1865
rect 16135 -1885 16165 -1865
rect 16185 -1885 16215 -1865
rect 16235 -1885 16265 -1865
rect 16285 -1885 16315 -1865
rect 16335 -1885 16365 -1865
rect 16385 -1885 16415 -1865
rect 16435 -1885 16465 -1865
rect 16485 -1885 16515 -1865
rect 16535 -1885 16565 -1865
rect 16585 -1885 16615 -1865
rect 16635 -1885 16665 -1865
rect 16685 -1885 16715 -1865
rect 16735 -1885 16765 -1865
rect 16785 -1885 16815 -1865
rect 16835 -1885 16865 -1865
rect 16885 -1885 16915 -1865
rect 16935 -1885 16965 -1865
rect 16985 -1885 17015 -1865
rect 17035 -1885 17065 -1865
rect 17085 -1885 17115 -1865
rect 17135 -1885 17165 -1865
rect 17185 -1885 17215 -1865
rect 17235 -1885 17265 -1865
rect 17285 -1885 17315 -1865
rect 17335 -1885 17365 -1865
rect 17385 -1885 17415 -1865
rect 17435 -1885 17465 -1865
rect 17485 -1885 17515 -1865
rect 17535 -1885 17565 -1865
rect 17585 -1885 17615 -1865
rect 17635 -1885 17665 -1865
rect 17685 -1885 17715 -1865
rect 17735 -1885 17765 -1865
rect 17785 -1885 17815 -1865
rect 17835 -1885 17865 -1865
rect 17885 -1885 17915 -1865
rect 17935 -1885 17965 -1865
rect 17985 -1885 18015 -1865
rect 18035 -1885 18065 -1865
rect 18085 -1885 18115 -1865
rect 18135 -1885 18165 -1865
rect 18185 -1885 18215 -1865
rect 18235 -1885 18265 -1865
rect 18285 -1885 18315 -1865
rect 18335 -1885 18365 -1865
rect 18385 -1885 18415 -1865
rect 18435 -1885 18465 -1865
rect 18485 -1885 18515 -1865
rect 18535 -1885 18565 -1865
rect 18585 -1885 18615 -1865
rect 18635 -1885 18665 -1865
rect 18685 -1885 18715 -1865
rect 18735 -1885 18765 -1865
rect 18785 -1885 18815 -1865
rect 18835 -1885 18865 -1865
rect 18885 -1885 18915 -1865
rect 18935 -1885 18965 -1865
rect 18985 -1885 19015 -1865
rect 19035 -1885 19065 -1865
rect 19085 -1885 19115 -1865
rect 19135 -1885 19165 -1865
rect 19185 -1885 19215 -1865
rect 19235 -1885 19265 -1865
rect 19285 -1885 19315 -1865
rect 19335 -1885 19365 -1865
rect 19385 -1885 19415 -1865
rect 19435 -1885 19465 -1865
rect 19485 -1885 19515 -1865
rect 19535 -1885 19565 -1865
rect 19585 -1885 19615 -1865
rect 19635 -1885 19665 -1865
rect 19685 -1885 19715 -1865
rect 19735 -1885 19765 -1865
rect 19785 -1885 19815 -1865
rect 19835 -1885 19865 -1865
rect 19885 -1885 19915 -1865
rect 19935 -1885 19965 -1865
rect 19985 -1885 20015 -1865
rect 20035 -1885 20065 -1865
rect 20085 -1885 20115 -1865
rect 20135 -1885 20165 -1865
rect 20185 -1885 20215 -1865
rect 20235 -1885 20265 -1865
rect 20285 -1885 20315 -1865
rect 20335 -1885 20365 -1865
rect 20385 -1885 20400 -1865
rect -650 -1900 20400 -1885
<< viali >>
rect -635 5165 -615 5185
rect 8365 5165 8385 5185
rect 8665 5165 8685 5185
rect 8965 5165 8985 5185
rect 9265 5165 9285 5185
rect 9565 5165 9585 5185
rect 9865 5165 9885 5185
rect 10165 5165 10185 5185
rect 10465 5165 10485 5185
rect 10765 5165 10785 5185
rect 11965 5165 11985 5185
rect 13165 5165 13185 5185
rect 14365 5165 14385 5185
rect 15565 5165 15585 5185
rect 17965 5165 17985 5185
rect 20365 5165 20385 5185
rect -635 5065 -615 5085
rect -635 5015 -615 5035
rect -635 4965 -615 4985
rect -635 4915 -615 4935
rect -635 4865 -615 4885
rect -635 4815 -615 4835
rect -635 4765 -615 4785
rect -635 4715 -615 4735
rect -635 4665 -615 4685
rect -635 4615 -615 4635
rect -485 5065 -465 5085
rect -485 5015 -465 5035
rect -485 4965 -465 4985
rect -485 4915 -465 4935
rect -485 4865 -465 4885
rect -485 4815 -465 4835
rect -485 4765 -465 4785
rect -485 4715 -465 4735
rect -485 4665 -465 4685
rect -485 4615 -465 4635
rect -335 5065 -315 5085
rect -335 5015 -315 5035
rect -335 4965 -315 4985
rect -335 4915 -315 4935
rect -335 4865 -315 4885
rect -335 4815 -315 4835
rect -335 4765 -315 4785
rect -335 4715 -315 4735
rect -185 5065 -165 5085
rect -185 5015 -165 5035
rect -185 4965 -165 4985
rect -185 4915 -165 4935
rect -185 4865 -165 4885
rect -185 4815 -165 4835
rect -185 4765 -165 4785
rect -185 4715 -165 4735
rect -185 4665 -165 4685
rect -185 4615 -165 4635
rect -35 5065 -15 5085
rect -35 5015 -15 5035
rect -35 4965 -15 4985
rect -35 4915 -15 4935
rect -35 4865 -15 4885
rect -35 4815 -15 4835
rect -35 4765 -15 4785
rect -35 4715 -15 4735
rect 565 5065 585 5085
rect 565 5015 585 5035
rect 565 4965 585 4985
rect 565 4915 585 4935
rect 565 4865 585 4885
rect 565 4815 585 4835
rect 565 4765 585 4785
rect 565 4715 585 4735
rect 565 4665 585 4685
rect 565 4615 585 4635
rect 715 4965 735 4985
rect 715 4915 735 4935
rect 715 4865 735 4885
rect 715 4815 735 4835
rect 715 4765 735 4785
rect 715 4715 735 4735
rect 715 4665 735 4685
rect 715 4615 735 4635
rect 865 5065 885 5085
rect 865 5015 885 5035
rect 865 4965 885 4985
rect 865 4915 885 4935
rect 865 4865 885 4885
rect 865 4815 885 4835
rect 865 4765 885 4785
rect 865 4715 885 4735
rect 1015 4965 1035 4985
rect 1015 4915 1035 4935
rect 1015 4865 1035 4885
rect 1015 4815 1035 4835
rect 1015 4765 1035 4785
rect 1015 4715 1035 4735
rect 1015 4665 1035 4685
rect 1165 5065 1185 5085
rect 1165 5015 1185 5035
rect 1165 4965 1185 4985
rect 1165 4915 1185 4935
rect 1165 4865 1185 4885
rect 1165 4815 1185 4835
rect 1165 4765 1185 4785
rect 1165 4715 1185 4735
rect 1315 4965 1335 4985
rect 1315 4915 1335 4935
rect 1315 4865 1335 4885
rect 1315 4815 1335 4835
rect 1315 4765 1335 4785
rect 1315 4715 1335 4735
rect 1315 4665 1335 4685
rect 1465 5065 1485 5085
rect 1465 5015 1485 5035
rect 1465 4965 1485 4985
rect 1465 4915 1485 4935
rect 1465 4865 1485 4885
rect 1465 4815 1485 4835
rect 1465 4765 1485 4785
rect 1465 4715 1485 4735
rect 1615 4965 1635 4985
rect 1615 4915 1635 4935
rect 1615 4865 1635 4885
rect 1615 4815 1635 4835
rect 1615 4765 1635 4785
rect 1615 4715 1635 4735
rect 1615 4665 1635 4685
rect 1765 5065 1785 5085
rect 1765 5015 1785 5035
rect 1765 4965 1785 4985
rect 1765 4915 1785 4935
rect 1765 4865 1785 4885
rect 1765 4815 1785 4835
rect 1765 4765 1785 4785
rect 1765 4715 1785 4735
rect 1765 4665 1785 4685
rect 1765 4615 1785 4635
rect 1915 4965 1935 4985
rect 1915 4915 1935 4935
rect 1915 4865 1935 4885
rect 1915 4815 1935 4835
rect 1915 4765 1935 4785
rect 1915 4715 1935 4735
rect 1915 4665 1935 4685
rect 1915 4615 1935 4635
rect 2065 5065 2085 5085
rect 2065 5015 2085 5035
rect 2065 4965 2085 4985
rect 2065 4915 2085 4935
rect 2065 4865 2085 4885
rect 2065 4815 2085 4835
rect 2065 4765 2085 4785
rect 2065 4715 2085 4735
rect 2215 4965 2235 4985
rect 2215 4915 2235 4935
rect 2215 4865 2235 4885
rect 2215 4815 2235 4835
rect 2215 4765 2235 4785
rect 2215 4715 2235 4735
rect 2215 4665 2235 4685
rect 2215 4615 2235 4635
rect 2365 5065 2385 5085
rect 2365 5015 2385 5035
rect 2365 4965 2385 4985
rect 2365 4915 2385 4935
rect 2365 4865 2385 4885
rect 2365 4815 2385 4835
rect 2365 4765 2385 4785
rect 2365 4715 2385 4735
rect 2365 4665 2385 4685
rect 2365 4615 2385 4635
rect 2515 4965 2535 4985
rect 2515 4915 2535 4935
rect 2515 4865 2535 4885
rect 2515 4815 2535 4835
rect 2515 4765 2535 4785
rect 2515 4715 2535 4735
rect 2515 4665 2535 4685
rect 2665 5065 2685 5085
rect 2665 5015 2685 5035
rect 2665 4965 2685 4985
rect 2665 4915 2685 4935
rect 2665 4865 2685 4885
rect 2665 4815 2685 4835
rect 2665 4765 2685 4785
rect 2665 4715 2685 4735
rect 2815 4965 2835 4985
rect 2815 4915 2835 4935
rect 2815 4865 2835 4885
rect 2815 4815 2835 4835
rect 2815 4765 2835 4785
rect 2815 4715 2835 4735
rect 2815 4665 2835 4685
rect 2965 5065 2985 5085
rect 2965 5015 2985 5035
rect 2965 4965 2985 4985
rect 2965 4915 2985 4935
rect 2965 4865 2985 4885
rect 2965 4815 2985 4835
rect 2965 4765 2985 4785
rect 2965 4715 2985 4735
rect 3115 4965 3135 4985
rect 3115 4915 3135 4935
rect 3115 4865 3135 4885
rect 3115 4815 3135 4835
rect 3115 4765 3135 4785
rect 3115 4715 3135 4735
rect 3115 4665 3135 4685
rect 3265 5065 3285 5085
rect 3265 5015 3285 5035
rect 3265 4965 3285 4985
rect 3265 4915 3285 4935
rect 3265 4865 3285 4885
rect 3265 4815 3285 4835
rect 3265 4765 3285 4785
rect 3265 4715 3285 4735
rect 3415 4965 3435 4985
rect 3415 4915 3435 4935
rect 3415 4865 3435 4885
rect 3415 4815 3435 4835
rect 3415 4765 3435 4785
rect 3415 4715 3435 4735
rect 3415 4665 3435 4685
rect 3415 4615 3435 4635
rect 3565 5065 3585 5085
rect 3565 5015 3585 5035
rect 3565 4965 3585 4985
rect 3565 4915 3585 4935
rect 3565 4865 3585 4885
rect 3565 4815 3585 4835
rect 3565 4765 3585 4785
rect 3565 4715 3585 4735
rect 3565 4665 3585 4685
rect 3565 4615 3585 4635
rect 4165 5065 4185 5085
rect 4165 5015 4185 5035
rect 4165 4965 4185 4985
rect 4165 4915 4185 4935
rect 4165 4865 4185 4885
rect 4165 4815 4185 4835
rect 4165 4765 4185 4785
rect 4165 4715 4185 4735
rect 4765 5065 4785 5085
rect 4765 5015 4785 5035
rect 4765 4965 4785 4985
rect 4765 4915 4785 4935
rect 4765 4865 4785 4885
rect 4765 4815 4785 4835
rect 4765 4765 4785 4785
rect 4765 4715 4785 4735
rect 4765 4665 4785 4685
rect 4765 4615 4785 4635
rect 4915 4965 4935 4985
rect 4915 4915 4935 4935
rect 4915 4865 4935 4885
rect 4915 4815 4935 4835
rect 4915 4765 4935 4785
rect 4915 4715 4935 4735
rect 4915 4665 4935 4685
rect 4915 4615 4935 4635
rect 5065 5065 5085 5085
rect 5065 5015 5085 5035
rect 5065 4965 5085 4985
rect 5065 4915 5085 4935
rect 5065 4865 5085 4885
rect 5065 4815 5085 4835
rect 5065 4765 5085 4785
rect 5065 4715 5085 4735
rect 5215 4965 5235 4985
rect 5215 4915 5235 4935
rect 5215 4865 5235 4885
rect 5215 4815 5235 4835
rect 5215 4765 5235 4785
rect 5215 4715 5235 4735
rect 5215 4665 5235 4685
rect 5365 5065 5385 5085
rect 5365 5015 5385 5035
rect 5365 4965 5385 4985
rect 5365 4915 5385 4935
rect 5365 4865 5385 4885
rect 5365 4815 5385 4835
rect 5365 4765 5385 4785
rect 5365 4715 5385 4735
rect 5515 4965 5535 4985
rect 5515 4915 5535 4935
rect 5515 4865 5535 4885
rect 5515 4815 5535 4835
rect 5515 4765 5535 4785
rect 5515 4715 5535 4735
rect 5515 4665 5535 4685
rect 5665 5065 5685 5085
rect 5665 5015 5685 5035
rect 5665 4965 5685 4985
rect 5665 4915 5685 4935
rect 5665 4865 5685 4885
rect 5665 4815 5685 4835
rect 5665 4765 5685 4785
rect 5665 4715 5685 4735
rect 5815 4965 5835 4985
rect 5815 4915 5835 4935
rect 5815 4865 5835 4885
rect 5815 4815 5835 4835
rect 5815 4765 5835 4785
rect 5815 4715 5835 4735
rect 5815 4665 5835 4685
rect 5965 5065 5985 5085
rect 5965 5015 5985 5035
rect 5965 4965 5985 4985
rect 5965 4915 5985 4935
rect 5965 4865 5985 4885
rect 5965 4815 5985 4835
rect 5965 4765 5985 4785
rect 5965 4715 5985 4735
rect 5965 4665 5985 4685
rect 5965 4615 5985 4635
rect 6115 4965 6135 4985
rect 6115 4915 6135 4935
rect 6115 4865 6135 4885
rect 6115 4815 6135 4835
rect 6115 4765 6135 4785
rect 6115 4715 6135 4735
rect 6115 4665 6135 4685
rect 6115 4615 6135 4635
rect 6265 5065 6285 5085
rect 6265 5015 6285 5035
rect 6265 4965 6285 4985
rect 6265 4915 6285 4935
rect 6265 4865 6285 4885
rect 6265 4815 6285 4835
rect 6265 4765 6285 4785
rect 6265 4715 6285 4735
rect 6415 4965 6435 4985
rect 6415 4915 6435 4935
rect 6415 4865 6435 4885
rect 6415 4815 6435 4835
rect 6415 4765 6435 4785
rect 6415 4715 6435 4735
rect 6415 4665 6435 4685
rect 6415 4615 6435 4635
rect 6565 5065 6585 5085
rect 6565 5015 6585 5035
rect 6565 4965 6585 4985
rect 6565 4915 6585 4935
rect 6565 4865 6585 4885
rect 6565 4815 6585 4835
rect 6565 4765 6585 4785
rect 6565 4715 6585 4735
rect 6565 4665 6585 4685
rect 6565 4615 6585 4635
rect 6715 4965 6735 4985
rect 6715 4915 6735 4935
rect 6715 4865 6735 4885
rect 6715 4815 6735 4835
rect 6715 4765 6735 4785
rect 6715 4715 6735 4735
rect 6715 4665 6735 4685
rect 6865 5065 6885 5085
rect 6865 5015 6885 5035
rect 6865 4965 6885 4985
rect 6865 4915 6885 4935
rect 6865 4865 6885 4885
rect 6865 4815 6885 4835
rect 6865 4765 6885 4785
rect 6865 4715 6885 4735
rect 7015 4965 7035 4985
rect 7015 4915 7035 4935
rect 7015 4865 7035 4885
rect 7015 4815 7035 4835
rect 7015 4765 7035 4785
rect 7015 4715 7035 4735
rect 7015 4665 7035 4685
rect 7165 5065 7185 5085
rect 7165 5015 7185 5035
rect 7165 4965 7185 4985
rect 7165 4915 7185 4935
rect 7165 4865 7185 4885
rect 7165 4815 7185 4835
rect 7165 4765 7185 4785
rect 7165 4715 7185 4735
rect 7315 4965 7335 4985
rect 7315 4915 7335 4935
rect 7315 4865 7335 4885
rect 7315 4815 7335 4835
rect 7315 4765 7335 4785
rect 7315 4715 7335 4735
rect 7315 4665 7335 4685
rect 7465 5065 7485 5085
rect 7465 5015 7485 5035
rect 7465 4965 7485 4985
rect 7465 4915 7485 4935
rect 7465 4865 7485 4885
rect 7465 4815 7485 4835
rect 7465 4765 7485 4785
rect 7465 4715 7485 4735
rect 7615 4965 7635 4985
rect 7615 4915 7635 4935
rect 7615 4865 7635 4885
rect 7615 4815 7635 4835
rect 7615 4765 7635 4785
rect 7615 4715 7635 4735
rect 7615 4665 7635 4685
rect 7615 4615 7635 4635
rect 7765 5065 7785 5085
rect 7765 5015 7785 5035
rect 7765 4965 7785 4985
rect 7765 4915 7785 4935
rect 7765 4865 7785 4885
rect 7765 4815 7785 4835
rect 7765 4765 7785 4785
rect 7765 4715 7785 4735
rect 7765 4665 7785 4685
rect 7765 4615 7785 4635
rect 8365 5065 8385 5085
rect 8365 5015 8385 5035
rect 8365 4965 8385 4985
rect 8365 4915 8385 4935
rect 8365 4865 8385 4885
rect 8365 4815 8385 4835
rect 8365 4765 8385 4785
rect 8365 4715 8385 4735
rect 8365 4665 8385 4685
rect 8365 4615 8385 4635
rect 8515 5065 8535 5085
rect 8515 5015 8535 5035
rect 8515 4965 8535 4985
rect 8515 4915 8535 4935
rect 8515 4865 8535 4885
rect 8515 4815 8535 4835
rect 8515 4765 8535 4785
rect 8515 4715 8535 4735
rect 8515 4665 8535 4685
rect 8515 4615 8535 4635
rect 8665 5065 8685 5085
rect 8665 5015 8685 5035
rect 8665 4965 8685 4985
rect 8665 4915 8685 4935
rect 8665 4865 8685 4885
rect 8665 4815 8685 4835
rect 8665 4765 8685 4785
rect 8665 4715 8685 4735
rect 8665 4665 8685 4685
rect 8665 4615 8685 4635
rect 8815 5065 8835 5085
rect 8815 5015 8835 5035
rect 8815 4965 8835 4985
rect 8815 4915 8835 4935
rect 8815 4865 8835 4885
rect 8815 4815 8835 4835
rect 8815 4765 8835 4785
rect 8815 4715 8835 4735
rect 8815 4665 8835 4685
rect 8815 4615 8835 4635
rect 8965 5065 8985 5085
rect 8965 5015 8985 5035
rect 8965 4965 8985 4985
rect 8965 4915 8985 4935
rect 8965 4865 8985 4885
rect 8965 4815 8985 4835
rect 8965 4765 8985 4785
rect 8965 4715 8985 4735
rect 8965 4665 8985 4685
rect 8965 4615 8985 4635
rect 9115 5065 9135 5085
rect 9115 5015 9135 5035
rect 9115 4965 9135 4985
rect 9115 4915 9135 4935
rect 9115 4865 9135 4885
rect 9115 4815 9135 4835
rect 9115 4765 9135 4785
rect 9115 4715 9135 4735
rect 9115 4665 9135 4685
rect 9115 4615 9135 4635
rect 9265 5065 9285 5085
rect 9265 5015 9285 5035
rect 9265 4965 9285 4985
rect 9265 4915 9285 4935
rect 9265 4865 9285 4885
rect 9265 4815 9285 4835
rect 9265 4765 9285 4785
rect 9265 4715 9285 4735
rect 9265 4665 9285 4685
rect 9265 4615 9285 4635
rect 9415 5065 9435 5085
rect 9415 5015 9435 5035
rect 9415 4965 9435 4985
rect 9415 4915 9435 4935
rect 9415 4865 9435 4885
rect 9415 4815 9435 4835
rect 9415 4765 9435 4785
rect 9415 4715 9435 4735
rect 9415 4665 9435 4685
rect 9415 4615 9435 4635
rect 9565 5065 9585 5085
rect 9565 5015 9585 5035
rect 9565 4965 9585 4985
rect 9565 4915 9585 4935
rect 9565 4865 9585 4885
rect 9565 4815 9585 4835
rect 9565 4765 9585 4785
rect 9565 4715 9585 4735
rect 9565 4665 9585 4685
rect 9565 4615 9585 4635
rect 9715 5065 9735 5085
rect 9715 5015 9735 5035
rect 9715 4965 9735 4985
rect 9715 4915 9735 4935
rect 9715 4865 9735 4885
rect 9715 4815 9735 4835
rect 9715 4765 9735 4785
rect 9715 4715 9735 4735
rect 9715 4665 9735 4685
rect 9715 4615 9735 4635
rect 9865 5065 9885 5085
rect 9865 5015 9885 5035
rect 9865 4965 9885 4985
rect 9865 4915 9885 4935
rect 9865 4865 9885 4885
rect 9865 4815 9885 4835
rect 9865 4765 9885 4785
rect 9865 4715 9885 4735
rect 9865 4665 9885 4685
rect 9865 4615 9885 4635
rect 10015 5065 10035 5085
rect 10015 5015 10035 5035
rect 10015 4965 10035 4985
rect 10015 4915 10035 4935
rect 10015 4865 10035 4885
rect 10015 4815 10035 4835
rect 10015 4765 10035 4785
rect 10015 4715 10035 4735
rect 10015 4665 10035 4685
rect 10015 4615 10035 4635
rect 10165 5065 10185 5085
rect 10165 5015 10185 5035
rect 10165 4965 10185 4985
rect 10165 4915 10185 4935
rect 10165 4865 10185 4885
rect 10165 4815 10185 4835
rect 10165 4765 10185 4785
rect 10165 4715 10185 4735
rect 10165 4665 10185 4685
rect 10165 4615 10185 4635
rect 10315 5065 10335 5085
rect 10315 5015 10335 5035
rect 10315 4965 10335 4985
rect 10315 4915 10335 4935
rect 10315 4865 10335 4885
rect 10315 4815 10335 4835
rect 10315 4765 10335 4785
rect 10315 4715 10335 4735
rect 10315 4665 10335 4685
rect 10315 4615 10335 4635
rect 10465 5065 10485 5085
rect 10465 5015 10485 5035
rect 10465 4965 10485 4985
rect 10465 4915 10485 4935
rect 10465 4865 10485 4885
rect 10465 4815 10485 4835
rect 10465 4765 10485 4785
rect 10465 4715 10485 4735
rect 10465 4665 10485 4685
rect 10465 4615 10485 4635
rect 10615 5065 10635 5085
rect 10615 5015 10635 5035
rect 10615 4965 10635 4985
rect 10615 4915 10635 4935
rect 10615 4865 10635 4885
rect 10615 4815 10635 4835
rect 10615 4765 10635 4785
rect 10615 4715 10635 4735
rect 10615 4665 10635 4685
rect 10615 4615 10635 4635
rect 10765 5065 10785 5085
rect 10765 5015 10785 5035
rect 10765 4965 10785 4985
rect 10765 4915 10785 4935
rect 10765 4865 10785 4885
rect 10765 4815 10785 4835
rect 10765 4765 10785 4785
rect 10765 4715 10785 4735
rect 10765 4665 10785 4685
rect 10765 4615 10785 4635
rect 11365 5065 11385 5085
rect 11365 5015 11385 5035
rect 11365 4965 11385 4985
rect 11365 4915 11385 4935
rect 11365 4865 11385 4885
rect 11365 4815 11385 4835
rect 11365 4765 11385 4785
rect 11365 4715 11385 4735
rect 11365 4665 11385 4685
rect 11365 4615 11385 4635
rect 11965 5065 11985 5085
rect 11965 5015 11985 5035
rect 11965 4965 11985 4985
rect 11965 4915 11985 4935
rect 11965 4865 11985 4885
rect 11965 4815 11985 4835
rect 11965 4765 11985 4785
rect 11965 4715 11985 4735
rect 11965 4665 11985 4685
rect 11965 4615 11985 4635
rect 12565 5065 12585 5085
rect 12565 5015 12585 5035
rect 12565 4965 12585 4985
rect 12565 4915 12585 4935
rect 12565 4865 12585 4885
rect 12565 4815 12585 4835
rect 12565 4765 12585 4785
rect 12565 4715 12585 4735
rect 12565 4665 12585 4685
rect 12565 4615 12585 4635
rect 13165 5065 13185 5085
rect 13165 5015 13185 5035
rect 13165 4965 13185 4985
rect 13165 4915 13185 4935
rect 13165 4865 13185 4885
rect 13165 4815 13185 4835
rect 13165 4765 13185 4785
rect 13165 4715 13185 4735
rect 13165 4665 13185 4685
rect 13165 4615 13185 4635
rect 13765 5065 13785 5085
rect 13765 5015 13785 5035
rect 13765 4965 13785 4985
rect 13765 4915 13785 4935
rect 13765 4865 13785 4885
rect 13765 4815 13785 4835
rect 13765 4765 13785 4785
rect 13765 4715 13785 4735
rect 13765 4665 13785 4685
rect 13765 4615 13785 4635
rect 14365 5065 14385 5085
rect 14365 5015 14385 5035
rect 14365 4965 14385 4985
rect 14365 4915 14385 4935
rect 14365 4865 14385 4885
rect 14365 4815 14385 4835
rect 14365 4765 14385 4785
rect 14365 4715 14385 4735
rect 14365 4665 14385 4685
rect 14365 4615 14385 4635
rect 14965 5065 14985 5085
rect 14965 5015 14985 5035
rect 14965 4965 14985 4985
rect 14965 4915 14985 4935
rect 14965 4865 14985 4885
rect 14965 4815 14985 4835
rect 14965 4765 14985 4785
rect 14965 4715 14985 4735
rect 14965 4665 14985 4685
rect 14965 4615 14985 4635
rect 15565 5065 15585 5085
rect 15565 5015 15585 5035
rect 15565 4965 15585 4985
rect 15565 4915 15585 4935
rect 15565 4865 15585 4885
rect 15565 4815 15585 4835
rect 15565 4765 15585 4785
rect 15565 4715 15585 4735
rect 15565 4665 15585 4685
rect 15565 4615 15585 4635
rect 16165 5065 16185 5085
rect 16165 5015 16185 5035
rect 16165 4965 16185 4985
rect 16165 4915 16185 4935
rect 16165 4865 16185 4885
rect 16165 4815 16185 4835
rect 16165 4765 16185 4785
rect 16165 4715 16185 4735
rect 16165 4665 16185 4685
rect 16165 4615 16185 4635
rect 16315 4965 16335 4985
rect 16315 4915 16335 4935
rect 16315 4865 16335 4885
rect 16315 4815 16335 4835
rect 16315 4765 16335 4785
rect 16315 4715 16335 4735
rect 16315 4665 16335 4685
rect 16315 4615 16335 4635
rect 16465 5065 16485 5085
rect 16465 5015 16485 5035
rect 16465 4965 16485 4985
rect 16465 4915 16485 4935
rect 16465 4865 16485 4885
rect 16465 4815 16485 4835
rect 16465 4765 16485 4785
rect 16465 4715 16485 4735
rect 16615 4965 16635 4985
rect 16615 4915 16635 4935
rect 16615 4865 16635 4885
rect 16615 4815 16635 4835
rect 16615 4765 16635 4785
rect 16615 4715 16635 4735
rect 16615 4665 16635 4685
rect 16615 4615 16635 4635
rect 16765 5065 16785 5085
rect 16765 5015 16785 5035
rect 16765 4965 16785 4985
rect 16765 4915 16785 4935
rect 16765 4865 16785 4885
rect 16765 4815 16785 4835
rect 16765 4765 16785 4785
rect 16765 4715 16785 4735
rect 16915 4965 16935 4985
rect 16915 4915 16935 4935
rect 16915 4865 16935 4885
rect 16915 4815 16935 4835
rect 16915 4765 16935 4785
rect 16915 4715 16935 4735
rect 16915 4665 16935 4685
rect 16915 4615 16935 4635
rect 17065 5065 17085 5085
rect 17065 5015 17085 5035
rect 17065 4965 17085 4985
rect 17065 4915 17085 4935
rect 17065 4865 17085 4885
rect 17065 4815 17085 4835
rect 17065 4765 17085 4785
rect 17065 4715 17085 4735
rect 17215 4965 17235 4985
rect 17215 4915 17235 4935
rect 17215 4865 17235 4885
rect 17215 4815 17235 4835
rect 17215 4765 17235 4785
rect 17215 4715 17235 4735
rect 17215 4665 17235 4685
rect 17215 4615 17235 4635
rect 17365 5065 17385 5085
rect 17365 5015 17385 5035
rect 17365 4965 17385 4985
rect 17365 4915 17385 4935
rect 17365 4865 17385 4885
rect 17365 4815 17385 4835
rect 17365 4765 17385 4785
rect 17365 4715 17385 4735
rect 17365 4665 17385 4685
rect 17365 4615 17385 4635
rect 17965 4965 17985 4985
rect 17965 4915 17985 4935
rect 17965 4865 17985 4885
rect 17965 4815 17985 4835
rect 17965 4765 17985 4785
rect 17965 4715 17985 4735
rect 17965 4665 17985 4685
rect 17965 4615 17985 4635
rect 18565 5065 18585 5085
rect 18565 5015 18585 5035
rect 18565 4965 18585 4985
rect 18565 4915 18585 4935
rect 18565 4865 18585 4885
rect 18565 4815 18585 4835
rect 18565 4765 18585 4785
rect 18565 4715 18585 4735
rect 18565 4665 18585 4685
rect 18565 4615 18585 4635
rect 18715 4965 18735 4985
rect 18715 4915 18735 4935
rect 18715 4865 18735 4885
rect 18715 4815 18735 4835
rect 18715 4765 18735 4785
rect 18715 4715 18735 4735
rect 18715 4665 18735 4685
rect 18715 4615 18735 4635
rect 18865 5065 18885 5085
rect 18865 5015 18885 5035
rect 18865 4965 18885 4985
rect 18865 4915 18885 4935
rect 18865 4865 18885 4885
rect 18865 4815 18885 4835
rect 18865 4765 18885 4785
rect 18865 4715 18885 4735
rect 19015 4965 19035 4985
rect 19015 4915 19035 4935
rect 19015 4865 19035 4885
rect 19015 4815 19035 4835
rect 19015 4765 19035 4785
rect 19015 4715 19035 4735
rect 19015 4665 19035 4685
rect 19015 4615 19035 4635
rect 19165 5065 19185 5085
rect 19165 5015 19185 5035
rect 19165 4965 19185 4985
rect 19165 4915 19185 4935
rect 19165 4865 19185 4885
rect 19165 4815 19185 4835
rect 19165 4765 19185 4785
rect 19165 4715 19185 4735
rect 19315 4965 19335 4985
rect 19315 4915 19335 4935
rect 19315 4865 19335 4885
rect 19315 4815 19335 4835
rect 19315 4765 19335 4785
rect 19315 4715 19335 4735
rect 19315 4665 19335 4685
rect 19315 4615 19335 4635
rect 19465 5065 19485 5085
rect 19465 5015 19485 5035
rect 19465 4965 19485 4985
rect 19465 4915 19485 4935
rect 19465 4865 19485 4885
rect 19465 4815 19485 4835
rect 19465 4765 19485 4785
rect 19465 4715 19485 4735
rect 19615 4965 19635 4985
rect 19615 4915 19635 4935
rect 19615 4865 19635 4885
rect 19615 4815 19635 4835
rect 19615 4765 19635 4785
rect 19615 4715 19635 4735
rect 19615 4665 19635 4685
rect 19615 4615 19635 4635
rect 19765 5065 19785 5085
rect 19765 5015 19785 5035
rect 19765 4965 19785 4985
rect 19765 4915 19785 4935
rect 19765 4865 19785 4885
rect 19765 4815 19785 4835
rect 19765 4765 19785 4785
rect 19765 4715 19785 4735
rect 19765 4665 19785 4685
rect 19765 4615 19785 4635
rect 20365 5065 20385 5085
rect 20365 5015 20385 5035
rect 20365 4965 20385 4985
rect 20365 4915 20385 4935
rect 20365 4865 20385 4885
rect 20365 4815 20385 4835
rect 20365 4765 20385 4785
rect 20365 4715 20385 4735
rect 20365 4665 20385 4685
rect 20365 4615 20385 4635
rect -485 4515 -465 4535
rect -185 4515 -165 4535
rect 115 4515 135 4535
rect 415 4515 435 4535
rect 715 4515 735 4535
rect 1015 4515 1035 4535
rect 1315 4515 1335 4535
rect 1615 4515 1635 4535
rect 1915 4515 1935 4535
rect 2215 4515 2235 4535
rect 2515 4515 2535 4535
rect 2815 4515 2835 4535
rect 3115 4515 3135 4535
rect 3415 4515 3435 4535
rect 3715 4515 3735 4535
rect 4015 4515 4035 4535
rect 4315 4515 4335 4535
rect 4615 4515 4635 4535
rect 4915 4515 4935 4535
rect 5215 4515 5235 4535
rect 5515 4515 5535 4535
rect 5815 4515 5835 4535
rect 6115 4515 6135 4535
rect 6415 4515 6435 4535
rect 6715 4515 6735 4535
rect 7015 4515 7035 4535
rect 7315 4515 7335 4535
rect 7615 4515 7635 4535
rect 7915 4515 7935 4535
rect 8215 4515 8235 4535
rect 8515 4515 8535 4535
rect 8815 4515 8835 4535
rect 9115 4515 9135 4535
rect 9415 4515 9435 4535
rect 9715 4515 9735 4535
rect 10015 4515 10035 4535
rect 10315 4515 10335 4535
rect 10615 4515 10635 4535
rect 10915 4515 10935 4535
rect 11215 4515 11235 4535
rect 11515 4515 11535 4535
rect 11815 4515 11835 4535
rect 12115 4515 12135 4535
rect 12415 4515 12435 4535
rect 12715 4515 12735 4535
rect 13015 4515 13035 4535
rect 13315 4515 13335 4535
rect 13615 4515 13635 4535
rect 13915 4515 13935 4535
rect 14215 4515 14235 4535
rect 14515 4515 14535 4535
rect 14815 4515 14835 4535
rect 15115 4515 15135 4535
rect 15415 4515 15435 4535
rect 15715 4515 15735 4535
rect 16015 4515 16035 4535
rect 16315 4515 16335 4535
rect 16615 4515 16635 4535
rect 16915 4515 16935 4535
rect 17215 4515 17235 4535
rect 17515 4515 17535 4535
rect 17815 4515 17835 4535
rect 18115 4515 18135 4535
rect 18415 4515 18435 4535
rect 18715 4515 18735 4535
rect 19015 4515 19035 4535
rect 19315 4515 19335 4535
rect 19615 4515 19635 4535
rect 19915 4515 19935 4535
rect 20215 4515 20235 4535
rect -635 4415 -615 4435
rect -635 4365 -615 4385
rect -635 4315 -615 4335
rect -635 4265 -615 4285
rect -635 4215 -615 4235
rect -635 4165 -615 4185
rect -635 4115 -615 4135
rect -635 4065 -615 4085
rect -635 4015 -615 4035
rect -635 3965 -615 3985
rect -485 4415 -465 4435
rect -485 4365 -465 4385
rect -485 4315 -465 4335
rect -485 4265 -465 4285
rect -485 4215 -465 4235
rect -485 4165 -465 4185
rect -485 4115 -465 4135
rect -485 4065 -465 4085
rect -485 4015 -465 4035
rect -485 3965 -465 3985
rect -335 4315 -315 4335
rect -335 4265 -315 4285
rect -335 4215 -315 4235
rect -335 4165 -315 4185
rect -335 4115 -315 4135
rect -335 4065 -315 4085
rect -335 4015 -315 4035
rect -335 3965 -315 3985
rect -185 4415 -165 4435
rect -185 4365 -165 4385
rect -185 4315 -165 4335
rect -185 4265 -165 4285
rect -185 4215 -165 4235
rect -185 4165 -165 4185
rect -185 4115 -165 4135
rect -185 4065 -165 4085
rect -185 4015 -165 4035
rect -185 3965 -165 3985
rect -35 4315 -15 4335
rect -35 4265 -15 4285
rect -35 4215 -15 4235
rect -35 4165 -15 4185
rect -35 4115 -15 4135
rect -35 4065 -15 4085
rect -35 4015 -15 4035
rect -35 3965 -15 3985
rect 565 4415 585 4435
rect 565 4365 585 4385
rect 565 4315 585 4335
rect 565 4265 585 4285
rect 565 4215 585 4235
rect 565 4165 585 4185
rect 565 4115 585 4135
rect 565 4065 585 4085
rect 565 4015 585 4035
rect 565 3965 585 3985
rect 715 4415 735 4435
rect 715 4365 735 4385
rect 715 4315 735 4335
rect 715 4265 735 4285
rect 715 4215 735 4235
rect 715 4165 735 4185
rect 715 4115 735 4135
rect 715 4065 735 4085
rect 865 4315 885 4335
rect 865 4265 885 4285
rect 865 4215 885 4235
rect 865 4165 885 4185
rect 865 4115 885 4135
rect 865 4065 885 4085
rect 865 4015 885 4035
rect 865 3965 885 3985
rect 1015 4365 1035 4385
rect 1015 4315 1035 4335
rect 1015 4265 1035 4285
rect 1015 4215 1035 4235
rect 1015 4165 1035 4185
rect 1015 4115 1035 4135
rect 1015 4065 1035 4085
rect 1165 4315 1185 4335
rect 1165 4265 1185 4285
rect 1165 4215 1185 4235
rect 1165 4165 1185 4185
rect 1165 4115 1185 4135
rect 1165 4065 1185 4085
rect 1165 4015 1185 4035
rect 1165 3965 1185 3985
rect 1315 4365 1335 4385
rect 1315 4315 1335 4335
rect 1315 4265 1335 4285
rect 1315 4215 1335 4235
rect 1315 4165 1335 4185
rect 1315 4115 1335 4135
rect 1315 4065 1335 4085
rect 1465 4315 1485 4335
rect 1465 4265 1485 4285
rect 1465 4215 1485 4235
rect 1465 4165 1485 4185
rect 1465 4115 1485 4135
rect 1465 4065 1485 4085
rect 1465 4015 1485 4035
rect 1465 3965 1485 3985
rect 1615 4365 1635 4385
rect 1615 4315 1635 4335
rect 1615 4265 1635 4285
rect 1615 4215 1635 4235
rect 1615 4165 1635 4185
rect 1615 4115 1635 4135
rect 1615 4065 1635 4085
rect 1765 4415 1785 4435
rect 1765 4365 1785 4385
rect 1765 4315 1785 4335
rect 1765 4265 1785 4285
rect 1765 4215 1785 4235
rect 1765 4165 1785 4185
rect 1765 4115 1785 4135
rect 1765 4065 1785 4085
rect 1765 4015 1785 4035
rect 1765 3965 1785 3985
rect 1915 4415 1935 4435
rect 1915 4365 1935 4385
rect 1915 4315 1935 4335
rect 1915 4265 1935 4285
rect 1915 4215 1935 4235
rect 1915 4165 1935 4185
rect 1915 4115 1935 4135
rect 1915 4065 1935 4085
rect 2065 4315 2085 4335
rect 2065 4265 2085 4285
rect 2065 4215 2085 4235
rect 2065 4165 2085 4185
rect 2065 4115 2085 4135
rect 2065 4065 2085 4085
rect 2065 4015 2085 4035
rect 2065 3965 2085 3985
rect 2215 4415 2235 4435
rect 2215 4365 2235 4385
rect 2215 4315 2235 4335
rect 2215 4265 2235 4285
rect 2215 4215 2235 4235
rect 2215 4165 2235 4185
rect 2215 4115 2235 4135
rect 2215 4065 2235 4085
rect 2365 4415 2385 4435
rect 2365 4365 2385 4385
rect 2365 4315 2385 4335
rect 2365 4265 2385 4285
rect 2365 4215 2385 4235
rect 2365 4165 2385 4185
rect 2365 4115 2385 4135
rect 2365 4065 2385 4085
rect 2365 4015 2385 4035
rect 2365 3965 2385 3985
rect 2515 4365 2535 4385
rect 2515 4315 2535 4335
rect 2515 4265 2535 4285
rect 2515 4215 2535 4235
rect 2515 4165 2535 4185
rect 2515 4115 2535 4135
rect 2515 4065 2535 4085
rect 2665 4315 2685 4335
rect 2665 4265 2685 4285
rect 2665 4215 2685 4235
rect 2665 4165 2685 4185
rect 2665 4115 2685 4135
rect 2665 4065 2685 4085
rect 2665 4015 2685 4035
rect 2665 3965 2685 3985
rect 2815 4365 2835 4385
rect 2815 4315 2835 4335
rect 2815 4265 2835 4285
rect 2815 4215 2835 4235
rect 2815 4165 2835 4185
rect 2815 4115 2835 4135
rect 2815 4065 2835 4085
rect 2965 4315 2985 4335
rect 2965 4265 2985 4285
rect 2965 4215 2985 4235
rect 2965 4165 2985 4185
rect 2965 4115 2985 4135
rect 2965 4065 2985 4085
rect 2965 4015 2985 4035
rect 2965 3965 2985 3985
rect 3115 4365 3135 4385
rect 3115 4315 3135 4335
rect 3115 4265 3135 4285
rect 3115 4215 3135 4235
rect 3115 4165 3135 4185
rect 3115 4115 3135 4135
rect 3115 4065 3135 4085
rect 3265 4315 3285 4335
rect 3265 4265 3285 4285
rect 3265 4215 3285 4235
rect 3265 4165 3285 4185
rect 3265 4115 3285 4135
rect 3265 4065 3285 4085
rect 3265 4015 3285 4035
rect 3265 3965 3285 3985
rect 3415 4415 3435 4435
rect 3415 4365 3435 4385
rect 3415 4315 3435 4335
rect 3415 4265 3435 4285
rect 3415 4215 3435 4235
rect 3415 4165 3435 4185
rect 3415 4115 3435 4135
rect 3415 4065 3435 4085
rect 3565 4415 3585 4435
rect 3565 4365 3585 4385
rect 3565 4315 3585 4335
rect 3565 4265 3585 4285
rect 3565 4215 3585 4235
rect 3565 4165 3585 4185
rect 3565 4115 3585 4135
rect 3565 4065 3585 4085
rect 3565 4015 3585 4035
rect 3565 3965 3585 3985
rect 4165 4315 4185 4335
rect 4165 4265 4185 4285
rect 4165 4215 4185 4235
rect 4165 4165 4185 4185
rect 4165 4115 4185 4135
rect 4165 4065 4185 4085
rect 4165 4015 4185 4035
rect 4165 3965 4185 3985
rect 4765 4415 4785 4435
rect 4765 4365 4785 4385
rect 4765 4315 4785 4335
rect 4765 4265 4785 4285
rect 4765 4215 4785 4235
rect 4765 4165 4785 4185
rect 4765 4115 4785 4135
rect 4765 4065 4785 4085
rect 4765 4015 4785 4035
rect 4765 3965 4785 3985
rect 4915 4415 4935 4435
rect 4915 4365 4935 4385
rect 4915 4315 4935 4335
rect 4915 4265 4935 4285
rect 4915 4215 4935 4235
rect 4915 4165 4935 4185
rect 4915 4115 4935 4135
rect 4915 4065 4935 4085
rect 5065 4315 5085 4335
rect 5065 4265 5085 4285
rect 5065 4215 5085 4235
rect 5065 4165 5085 4185
rect 5065 4115 5085 4135
rect 5065 4065 5085 4085
rect 5065 4015 5085 4035
rect 5065 3965 5085 3985
rect 5215 4365 5235 4385
rect 5215 4315 5235 4335
rect 5215 4265 5235 4285
rect 5215 4215 5235 4235
rect 5215 4165 5235 4185
rect 5215 4115 5235 4135
rect 5215 4065 5235 4085
rect 5365 4315 5385 4335
rect 5365 4265 5385 4285
rect 5365 4215 5385 4235
rect 5365 4165 5385 4185
rect 5365 4115 5385 4135
rect 5365 4065 5385 4085
rect 5365 4015 5385 4035
rect 5365 3965 5385 3985
rect 5515 4365 5535 4385
rect 5515 4315 5535 4335
rect 5515 4265 5535 4285
rect 5515 4215 5535 4235
rect 5515 4165 5535 4185
rect 5515 4115 5535 4135
rect 5515 4065 5535 4085
rect 5665 4315 5685 4335
rect 5665 4265 5685 4285
rect 5665 4215 5685 4235
rect 5665 4165 5685 4185
rect 5665 4115 5685 4135
rect 5665 4065 5685 4085
rect 5665 4015 5685 4035
rect 5665 3965 5685 3985
rect 5815 4365 5835 4385
rect 5815 4315 5835 4335
rect 5815 4265 5835 4285
rect 5815 4215 5835 4235
rect 5815 4165 5835 4185
rect 5815 4115 5835 4135
rect 5815 4065 5835 4085
rect 5965 4415 5985 4435
rect 5965 4365 5985 4385
rect 5965 4315 5985 4335
rect 5965 4265 5985 4285
rect 5965 4215 5985 4235
rect 5965 4165 5985 4185
rect 5965 4115 5985 4135
rect 5965 4065 5985 4085
rect 5965 4015 5985 4035
rect 5965 3965 5985 3985
rect 6115 4415 6135 4435
rect 6115 4365 6135 4385
rect 6115 4315 6135 4335
rect 6115 4265 6135 4285
rect 6115 4215 6135 4235
rect 6115 4165 6135 4185
rect 6115 4115 6135 4135
rect 6115 4065 6135 4085
rect 6265 4315 6285 4335
rect 6265 4265 6285 4285
rect 6265 4215 6285 4235
rect 6265 4165 6285 4185
rect 6265 4115 6285 4135
rect 6265 4065 6285 4085
rect 6265 4015 6285 4035
rect 6265 3965 6285 3985
rect 6415 4415 6435 4435
rect 6415 4365 6435 4385
rect 6415 4315 6435 4335
rect 6415 4265 6435 4285
rect 6415 4215 6435 4235
rect 6415 4165 6435 4185
rect 6415 4115 6435 4135
rect 6415 4065 6435 4085
rect 6565 4415 6585 4435
rect 6565 4365 6585 4385
rect 6565 4315 6585 4335
rect 6565 4265 6585 4285
rect 6565 4215 6585 4235
rect 6565 4165 6585 4185
rect 6565 4115 6585 4135
rect 6565 4065 6585 4085
rect 6565 4015 6585 4035
rect 6565 3965 6585 3985
rect 6715 4365 6735 4385
rect 6715 4315 6735 4335
rect 6715 4265 6735 4285
rect 6715 4215 6735 4235
rect 6715 4165 6735 4185
rect 6715 4115 6735 4135
rect 6715 4065 6735 4085
rect 6865 4315 6885 4335
rect 6865 4265 6885 4285
rect 6865 4215 6885 4235
rect 6865 4165 6885 4185
rect 6865 4115 6885 4135
rect 6865 4065 6885 4085
rect 6865 4015 6885 4035
rect 6865 3965 6885 3985
rect 7015 4365 7035 4385
rect 7015 4315 7035 4335
rect 7015 4265 7035 4285
rect 7015 4215 7035 4235
rect 7015 4165 7035 4185
rect 7015 4115 7035 4135
rect 7015 4065 7035 4085
rect 7165 4315 7185 4335
rect 7165 4265 7185 4285
rect 7165 4215 7185 4235
rect 7165 4165 7185 4185
rect 7165 4115 7185 4135
rect 7165 4065 7185 4085
rect 7165 4015 7185 4035
rect 7165 3965 7185 3985
rect 7315 4365 7335 4385
rect 7315 4315 7335 4335
rect 7315 4265 7335 4285
rect 7315 4215 7335 4235
rect 7315 4165 7335 4185
rect 7315 4115 7335 4135
rect 7315 4065 7335 4085
rect 7465 4315 7485 4335
rect 7465 4265 7485 4285
rect 7465 4215 7485 4235
rect 7465 4165 7485 4185
rect 7465 4115 7485 4135
rect 7465 4065 7485 4085
rect 7465 4015 7485 4035
rect 7465 3965 7485 3985
rect 7615 4415 7635 4435
rect 7615 4365 7635 4385
rect 7615 4315 7635 4335
rect 7615 4265 7635 4285
rect 7615 4215 7635 4235
rect 7615 4165 7635 4185
rect 7615 4115 7635 4135
rect 7615 4065 7635 4085
rect 7765 4415 7785 4435
rect 7765 4365 7785 4385
rect 7765 4315 7785 4335
rect 7765 4265 7785 4285
rect 7765 4215 7785 4235
rect 7765 4165 7785 4185
rect 7765 4115 7785 4135
rect 7765 4065 7785 4085
rect 7765 4015 7785 4035
rect 7765 3965 7785 3985
rect 8365 4415 8385 4435
rect 8365 4365 8385 4385
rect 8365 4315 8385 4335
rect 8365 4265 8385 4285
rect 8365 4215 8385 4235
rect 8365 4165 8385 4185
rect 8365 4115 8385 4135
rect 8365 4065 8385 4085
rect 8365 4015 8385 4035
rect 8365 3965 8385 3985
rect 8515 4415 8535 4435
rect 8515 4365 8535 4385
rect 8515 4315 8535 4335
rect 8515 4265 8535 4285
rect 8515 4215 8535 4235
rect 8515 4165 8535 4185
rect 8515 4115 8535 4135
rect 8515 4065 8535 4085
rect 8515 4015 8535 4035
rect 8515 3965 8535 3985
rect 8665 4415 8685 4435
rect 8665 4365 8685 4385
rect 8665 4315 8685 4335
rect 8665 4265 8685 4285
rect 8665 4215 8685 4235
rect 8665 4165 8685 4185
rect 8665 4115 8685 4135
rect 8665 4065 8685 4085
rect 8665 4015 8685 4035
rect 8665 3965 8685 3985
rect 8815 4415 8835 4435
rect 8815 4365 8835 4385
rect 8815 4315 8835 4335
rect 8815 4265 8835 4285
rect 8815 4215 8835 4235
rect 8815 4165 8835 4185
rect 8815 4115 8835 4135
rect 8815 4065 8835 4085
rect 8815 4015 8835 4035
rect 8815 3965 8835 3985
rect 8965 4415 8985 4435
rect 8965 4365 8985 4385
rect 8965 4315 8985 4335
rect 8965 4265 8985 4285
rect 8965 4215 8985 4235
rect 8965 4165 8985 4185
rect 8965 4115 8985 4135
rect 8965 4065 8985 4085
rect 8965 4015 8985 4035
rect 8965 3965 8985 3985
rect 9115 4415 9135 4435
rect 9115 4365 9135 4385
rect 9115 4315 9135 4335
rect 9115 4265 9135 4285
rect 9115 4215 9135 4235
rect 9115 4165 9135 4185
rect 9115 4115 9135 4135
rect 9115 4065 9135 4085
rect 9115 4015 9135 4035
rect 9115 3965 9135 3985
rect 9265 4415 9285 4435
rect 9265 4365 9285 4385
rect 9265 4315 9285 4335
rect 9265 4265 9285 4285
rect 9265 4215 9285 4235
rect 9265 4165 9285 4185
rect 9265 4115 9285 4135
rect 9265 4065 9285 4085
rect 9265 4015 9285 4035
rect 9265 3965 9285 3985
rect 9415 4415 9435 4435
rect 9415 4365 9435 4385
rect 9415 4315 9435 4335
rect 9415 4265 9435 4285
rect 9415 4215 9435 4235
rect 9415 4165 9435 4185
rect 9415 4115 9435 4135
rect 9415 4065 9435 4085
rect 9415 4015 9435 4035
rect 9415 3965 9435 3985
rect 9565 4415 9585 4435
rect 9565 4365 9585 4385
rect 9565 4315 9585 4335
rect 9565 4265 9585 4285
rect 9565 4215 9585 4235
rect 9565 4165 9585 4185
rect 9565 4115 9585 4135
rect 9565 4065 9585 4085
rect 9565 4015 9585 4035
rect 9565 3965 9585 3985
rect 9715 4415 9735 4435
rect 9715 4365 9735 4385
rect 9715 4315 9735 4335
rect 9715 4265 9735 4285
rect 9715 4215 9735 4235
rect 9715 4165 9735 4185
rect 9715 4115 9735 4135
rect 9715 4065 9735 4085
rect 9715 4015 9735 4035
rect 9715 3965 9735 3985
rect 9865 4415 9885 4435
rect 9865 4365 9885 4385
rect 9865 4315 9885 4335
rect 9865 4265 9885 4285
rect 9865 4215 9885 4235
rect 9865 4165 9885 4185
rect 9865 4115 9885 4135
rect 9865 4065 9885 4085
rect 9865 4015 9885 4035
rect 9865 3965 9885 3985
rect 10015 4415 10035 4435
rect 10015 4365 10035 4385
rect 10015 4315 10035 4335
rect 10015 4265 10035 4285
rect 10015 4215 10035 4235
rect 10015 4165 10035 4185
rect 10015 4115 10035 4135
rect 10015 4065 10035 4085
rect 10015 4015 10035 4035
rect 10015 3965 10035 3985
rect 10165 4415 10185 4435
rect 10165 4365 10185 4385
rect 10165 4315 10185 4335
rect 10165 4265 10185 4285
rect 10165 4215 10185 4235
rect 10165 4165 10185 4185
rect 10165 4115 10185 4135
rect 10165 4065 10185 4085
rect 10165 4015 10185 4035
rect 10165 3965 10185 3985
rect 10315 4415 10335 4435
rect 10315 4365 10335 4385
rect 10315 4315 10335 4335
rect 10315 4265 10335 4285
rect 10315 4215 10335 4235
rect 10315 4165 10335 4185
rect 10315 4115 10335 4135
rect 10315 4065 10335 4085
rect 10315 4015 10335 4035
rect 10315 3965 10335 3985
rect 10465 4415 10485 4435
rect 10465 4365 10485 4385
rect 10465 4315 10485 4335
rect 10465 4265 10485 4285
rect 10465 4215 10485 4235
rect 10465 4165 10485 4185
rect 10465 4115 10485 4135
rect 10465 4065 10485 4085
rect 10465 4015 10485 4035
rect 10465 3965 10485 3985
rect 10615 4415 10635 4435
rect 10615 4365 10635 4385
rect 10615 4315 10635 4335
rect 10615 4265 10635 4285
rect 10615 4215 10635 4235
rect 10615 4165 10635 4185
rect 10615 4115 10635 4135
rect 10615 4065 10635 4085
rect 10615 4015 10635 4035
rect 10615 3965 10635 3985
rect 10765 4415 10785 4435
rect 10765 4365 10785 4385
rect 10765 4315 10785 4335
rect 10765 4265 10785 4285
rect 10765 4215 10785 4235
rect 10765 4165 10785 4185
rect 10765 4115 10785 4135
rect 10765 4065 10785 4085
rect 10765 4015 10785 4035
rect 10765 3965 10785 3985
rect 11365 4415 11385 4435
rect 11365 4365 11385 4385
rect 11365 4315 11385 4335
rect 11365 4265 11385 4285
rect 11365 4215 11385 4235
rect 11365 4165 11385 4185
rect 11365 4115 11385 4135
rect 11365 4065 11385 4085
rect 11365 4015 11385 4035
rect 11365 3965 11385 3985
rect 11965 4415 11985 4435
rect 11965 4365 11985 4385
rect 11965 4315 11985 4335
rect 11965 4265 11985 4285
rect 11965 4215 11985 4235
rect 11965 4165 11985 4185
rect 11965 4115 11985 4135
rect 11965 4065 11985 4085
rect 11965 4015 11985 4035
rect 11965 3965 11985 3985
rect 12565 4415 12585 4435
rect 12565 4365 12585 4385
rect 12565 4315 12585 4335
rect 12565 4265 12585 4285
rect 12565 4215 12585 4235
rect 12565 4165 12585 4185
rect 12565 4115 12585 4135
rect 12565 4065 12585 4085
rect 12565 4015 12585 4035
rect 12565 3965 12585 3985
rect 13165 4415 13185 4435
rect 13165 4365 13185 4385
rect 13165 4315 13185 4335
rect 13165 4265 13185 4285
rect 13165 4215 13185 4235
rect 13165 4165 13185 4185
rect 13165 4115 13185 4135
rect 13165 4065 13185 4085
rect 13165 4015 13185 4035
rect 13165 3965 13185 3985
rect 13765 4415 13785 4435
rect 13765 4365 13785 4385
rect 13765 4315 13785 4335
rect 13765 4265 13785 4285
rect 13765 4215 13785 4235
rect 13765 4165 13785 4185
rect 13765 4115 13785 4135
rect 13765 4065 13785 4085
rect 13765 4015 13785 4035
rect 13765 3965 13785 3985
rect 14365 4415 14385 4435
rect 14365 4365 14385 4385
rect 14365 4315 14385 4335
rect 14365 4265 14385 4285
rect 14365 4215 14385 4235
rect 14365 4165 14385 4185
rect 14365 4115 14385 4135
rect 14365 4065 14385 4085
rect 14365 4015 14385 4035
rect 14365 3965 14385 3985
rect 14965 4415 14985 4435
rect 14965 4365 14985 4385
rect 14965 4315 14985 4335
rect 14965 4265 14985 4285
rect 14965 4215 14985 4235
rect 14965 4165 14985 4185
rect 14965 4115 14985 4135
rect 14965 4065 14985 4085
rect 14965 4015 14985 4035
rect 14965 3965 14985 3985
rect 15565 4415 15585 4435
rect 15565 4365 15585 4385
rect 15565 4315 15585 4335
rect 15565 4265 15585 4285
rect 15565 4215 15585 4235
rect 15565 4165 15585 4185
rect 15565 4115 15585 4135
rect 15565 4065 15585 4085
rect 15565 4015 15585 4035
rect 15565 3965 15585 3985
rect 16165 4415 16185 4435
rect 16165 4365 16185 4385
rect 16165 4315 16185 4335
rect 16165 4265 16185 4285
rect 16165 4215 16185 4235
rect 16165 4165 16185 4185
rect 16165 4115 16185 4135
rect 16165 4065 16185 4085
rect 16165 4015 16185 4035
rect 16165 3965 16185 3985
rect 16315 4415 16335 4435
rect 16315 4365 16335 4385
rect 16315 4315 16335 4335
rect 16315 4265 16335 4285
rect 16315 4215 16335 4235
rect 16315 4165 16335 4185
rect 16315 4115 16335 4135
rect 16315 4065 16335 4085
rect 16465 4315 16485 4335
rect 16465 4265 16485 4285
rect 16465 4215 16485 4235
rect 16465 4165 16485 4185
rect 16465 4115 16485 4135
rect 16465 4065 16485 4085
rect 16465 4015 16485 4035
rect 16465 3965 16485 3985
rect 16615 4415 16635 4435
rect 16615 4365 16635 4385
rect 16615 4315 16635 4335
rect 16615 4265 16635 4285
rect 16615 4215 16635 4235
rect 16615 4165 16635 4185
rect 16615 4115 16635 4135
rect 16615 4065 16635 4085
rect 16765 4315 16785 4335
rect 16765 4265 16785 4285
rect 16765 4215 16785 4235
rect 16765 4165 16785 4185
rect 16765 4115 16785 4135
rect 16765 4065 16785 4085
rect 16765 4015 16785 4035
rect 16765 3965 16785 3985
rect 16915 4415 16935 4435
rect 16915 4365 16935 4385
rect 16915 4315 16935 4335
rect 16915 4265 16935 4285
rect 16915 4215 16935 4235
rect 16915 4165 16935 4185
rect 16915 4115 16935 4135
rect 16915 4065 16935 4085
rect 17065 4315 17085 4335
rect 17065 4265 17085 4285
rect 17065 4215 17085 4235
rect 17065 4165 17085 4185
rect 17065 4115 17085 4135
rect 17065 4065 17085 4085
rect 17065 4015 17085 4035
rect 17065 3965 17085 3985
rect 17215 4415 17235 4435
rect 17215 4365 17235 4385
rect 17215 4315 17235 4335
rect 17215 4265 17235 4285
rect 17215 4215 17235 4235
rect 17215 4165 17235 4185
rect 17215 4115 17235 4135
rect 17215 4065 17235 4085
rect 17365 4415 17385 4435
rect 17365 4365 17385 4385
rect 17365 4315 17385 4335
rect 17365 4265 17385 4285
rect 17365 4215 17385 4235
rect 17365 4165 17385 4185
rect 17365 4115 17385 4135
rect 17365 4065 17385 4085
rect 17365 4015 17385 4035
rect 17365 3965 17385 3985
rect 17965 4415 17985 4435
rect 17965 4365 17985 4385
rect 17965 4315 17985 4335
rect 17965 4265 17985 4285
rect 17965 4215 17985 4235
rect 17965 4165 17985 4185
rect 17965 4115 17985 4135
rect 17965 4065 17985 4085
rect 18565 4415 18585 4435
rect 18565 4365 18585 4385
rect 18565 4315 18585 4335
rect 18565 4265 18585 4285
rect 18565 4215 18585 4235
rect 18565 4165 18585 4185
rect 18565 4115 18585 4135
rect 18565 4065 18585 4085
rect 18565 4015 18585 4035
rect 18565 3965 18585 3985
rect 18715 4415 18735 4435
rect 18715 4365 18735 4385
rect 18715 4315 18735 4335
rect 18715 4265 18735 4285
rect 18715 4215 18735 4235
rect 18715 4165 18735 4185
rect 18715 4115 18735 4135
rect 18715 4065 18735 4085
rect 18865 4315 18885 4335
rect 18865 4265 18885 4285
rect 18865 4215 18885 4235
rect 18865 4165 18885 4185
rect 18865 4115 18885 4135
rect 18865 4065 18885 4085
rect 18865 4015 18885 4035
rect 18865 3965 18885 3985
rect 19015 4415 19035 4435
rect 19015 4365 19035 4385
rect 19015 4315 19035 4335
rect 19015 4265 19035 4285
rect 19015 4215 19035 4235
rect 19015 4165 19035 4185
rect 19015 4115 19035 4135
rect 19015 4065 19035 4085
rect 19165 4315 19185 4335
rect 19165 4265 19185 4285
rect 19165 4215 19185 4235
rect 19165 4165 19185 4185
rect 19165 4115 19185 4135
rect 19165 4065 19185 4085
rect 19165 4015 19185 4035
rect 19165 3965 19185 3985
rect 19315 4415 19335 4435
rect 19315 4365 19335 4385
rect 19315 4315 19335 4335
rect 19315 4265 19335 4285
rect 19315 4215 19335 4235
rect 19315 4165 19335 4185
rect 19315 4115 19335 4135
rect 19315 4065 19335 4085
rect 19465 4315 19485 4335
rect 19465 4265 19485 4285
rect 19465 4215 19485 4235
rect 19465 4165 19485 4185
rect 19465 4115 19485 4135
rect 19465 4065 19485 4085
rect 19465 4015 19485 4035
rect 19465 3965 19485 3985
rect 19615 4415 19635 4435
rect 19615 4365 19635 4385
rect 19615 4315 19635 4335
rect 19615 4265 19635 4285
rect 19615 4215 19635 4235
rect 19615 4165 19635 4185
rect 19615 4115 19635 4135
rect 19615 4065 19635 4085
rect 19765 4415 19785 4435
rect 19765 4365 19785 4385
rect 19765 4315 19785 4335
rect 19765 4265 19785 4285
rect 19765 4215 19785 4235
rect 19765 4165 19785 4185
rect 19765 4115 19785 4135
rect 19765 4065 19785 4085
rect 19765 4015 19785 4035
rect 19765 3965 19785 3985
rect 20365 4415 20385 4435
rect 20365 4365 20385 4385
rect 20365 4315 20385 4335
rect 20365 4265 20385 4285
rect 20365 4215 20385 4235
rect 20365 4165 20385 4185
rect 20365 4115 20385 4135
rect 20365 4065 20385 4085
rect 20365 4015 20385 4035
rect 20365 3965 20385 3985
rect -635 3865 -615 3885
rect -35 3865 -15 3885
rect 4165 3865 4185 3885
rect 8365 3865 8385 3885
rect 8665 3865 8685 3885
rect 8965 3865 8985 3885
rect 9265 3865 9285 3885
rect 9565 3865 9585 3885
rect 9865 3865 9885 3885
rect 10165 3865 10185 3885
rect 10465 3865 10485 3885
rect 10765 3865 10785 3885
rect 11965 3865 11985 3885
rect 13165 3865 13185 3885
rect 14365 3865 14385 3885
rect 15565 3865 15585 3885
rect 20365 3865 20385 3885
rect -635 3765 -615 3785
rect -635 3715 -615 3735
rect -635 3665 -615 3685
rect -635 3615 -615 3635
rect -635 3565 -615 3585
rect -635 3515 -615 3535
rect -635 3465 -615 3485
rect -635 3415 -615 3435
rect -635 3365 -615 3385
rect -635 3315 -615 3335
rect -485 3765 -465 3785
rect -485 3715 -465 3735
rect -485 3665 -465 3685
rect -485 3615 -465 3635
rect -485 3565 -465 3585
rect -485 3515 -465 3535
rect -485 3465 -465 3485
rect -485 3415 -465 3435
rect -485 3365 -465 3385
rect -485 3315 -465 3335
rect -335 3765 -315 3785
rect -335 3715 -315 3735
rect -335 3665 -315 3685
rect -335 3615 -315 3635
rect -335 3565 -315 3585
rect -335 3515 -315 3535
rect -335 3465 -315 3485
rect -335 3415 -315 3435
rect -185 3765 -165 3785
rect -185 3715 -165 3735
rect -185 3665 -165 3685
rect -185 3615 -165 3635
rect -185 3565 -165 3585
rect -185 3515 -165 3535
rect -185 3465 -165 3485
rect -185 3415 -165 3435
rect -185 3365 -165 3385
rect -185 3315 -165 3335
rect -35 3765 -15 3785
rect -35 3715 -15 3735
rect -35 3665 -15 3685
rect -35 3615 -15 3635
rect -35 3565 -15 3585
rect -35 3515 -15 3535
rect -35 3465 -15 3485
rect -35 3415 -15 3435
rect 565 3765 585 3785
rect 565 3715 585 3735
rect 565 3665 585 3685
rect 565 3615 585 3635
rect 565 3565 585 3585
rect 565 3515 585 3535
rect 565 3465 585 3485
rect 565 3415 585 3435
rect 565 3365 585 3385
rect 565 3315 585 3335
rect 715 3665 735 3685
rect 715 3615 735 3635
rect 715 3565 735 3585
rect 715 3515 735 3535
rect 715 3465 735 3485
rect 715 3415 735 3435
rect 715 3365 735 3385
rect 715 3315 735 3335
rect 865 3765 885 3785
rect 865 3715 885 3735
rect 865 3665 885 3685
rect 865 3615 885 3635
rect 865 3565 885 3585
rect 865 3515 885 3535
rect 865 3465 885 3485
rect 865 3415 885 3435
rect 1015 3665 1035 3685
rect 1015 3615 1035 3635
rect 1015 3565 1035 3585
rect 1015 3515 1035 3535
rect 1015 3465 1035 3485
rect 1015 3415 1035 3435
rect 1015 3365 1035 3385
rect 1165 3765 1185 3785
rect 1165 3715 1185 3735
rect 1165 3665 1185 3685
rect 1165 3615 1185 3635
rect 1165 3565 1185 3585
rect 1165 3515 1185 3535
rect 1165 3465 1185 3485
rect 1165 3415 1185 3435
rect 1315 3665 1335 3685
rect 1315 3615 1335 3635
rect 1315 3565 1335 3585
rect 1315 3515 1335 3535
rect 1315 3465 1335 3485
rect 1315 3415 1335 3435
rect 1315 3365 1335 3385
rect 1465 3765 1485 3785
rect 1465 3715 1485 3735
rect 1465 3665 1485 3685
rect 1465 3615 1485 3635
rect 1465 3565 1485 3585
rect 1465 3515 1485 3535
rect 1465 3465 1485 3485
rect 1465 3415 1485 3435
rect 1615 3665 1635 3685
rect 1615 3615 1635 3635
rect 1615 3565 1635 3585
rect 1615 3515 1635 3535
rect 1615 3465 1635 3485
rect 1615 3415 1635 3435
rect 1615 3365 1635 3385
rect 1765 3765 1785 3785
rect 1765 3715 1785 3735
rect 1765 3665 1785 3685
rect 1765 3615 1785 3635
rect 1765 3565 1785 3585
rect 1765 3515 1785 3535
rect 1765 3465 1785 3485
rect 1765 3415 1785 3435
rect 1765 3365 1785 3385
rect 1765 3315 1785 3335
rect 1915 3665 1935 3685
rect 1915 3615 1935 3635
rect 1915 3565 1935 3585
rect 1915 3515 1935 3535
rect 1915 3465 1935 3485
rect 1915 3415 1935 3435
rect 1915 3365 1935 3385
rect 1915 3315 1935 3335
rect 2065 3765 2085 3785
rect 2065 3715 2085 3735
rect 2065 3665 2085 3685
rect 2065 3615 2085 3635
rect 2065 3565 2085 3585
rect 2065 3515 2085 3535
rect 2065 3465 2085 3485
rect 2065 3415 2085 3435
rect 2215 3665 2235 3685
rect 2215 3615 2235 3635
rect 2215 3565 2235 3585
rect 2215 3515 2235 3535
rect 2215 3465 2235 3485
rect 2215 3415 2235 3435
rect 2215 3365 2235 3385
rect 2215 3315 2235 3335
rect 2365 3765 2385 3785
rect 2365 3715 2385 3735
rect 2365 3665 2385 3685
rect 2365 3615 2385 3635
rect 2365 3565 2385 3585
rect 2365 3515 2385 3535
rect 2365 3465 2385 3485
rect 2365 3415 2385 3435
rect 2365 3365 2385 3385
rect 2365 3315 2385 3335
rect 2515 3665 2535 3685
rect 2515 3615 2535 3635
rect 2515 3565 2535 3585
rect 2515 3515 2535 3535
rect 2515 3465 2535 3485
rect 2515 3415 2535 3435
rect 2515 3365 2535 3385
rect 2665 3765 2685 3785
rect 2665 3715 2685 3735
rect 2665 3665 2685 3685
rect 2665 3615 2685 3635
rect 2665 3565 2685 3585
rect 2665 3515 2685 3535
rect 2665 3465 2685 3485
rect 2665 3415 2685 3435
rect 2815 3665 2835 3685
rect 2815 3615 2835 3635
rect 2815 3565 2835 3585
rect 2815 3515 2835 3535
rect 2815 3465 2835 3485
rect 2815 3415 2835 3435
rect 2815 3365 2835 3385
rect 2965 3765 2985 3785
rect 2965 3715 2985 3735
rect 2965 3665 2985 3685
rect 2965 3615 2985 3635
rect 2965 3565 2985 3585
rect 2965 3515 2985 3535
rect 2965 3465 2985 3485
rect 2965 3415 2985 3435
rect 3115 3665 3135 3685
rect 3115 3615 3135 3635
rect 3115 3565 3135 3585
rect 3115 3515 3135 3535
rect 3115 3465 3135 3485
rect 3115 3415 3135 3435
rect 3115 3365 3135 3385
rect 3265 3765 3285 3785
rect 3265 3715 3285 3735
rect 3265 3665 3285 3685
rect 3265 3615 3285 3635
rect 3265 3565 3285 3585
rect 3265 3515 3285 3535
rect 3265 3465 3285 3485
rect 3265 3415 3285 3435
rect 3415 3665 3435 3685
rect 3415 3615 3435 3635
rect 3415 3565 3435 3585
rect 3415 3515 3435 3535
rect 3415 3465 3435 3485
rect 3415 3415 3435 3435
rect 3415 3365 3435 3385
rect 3415 3315 3435 3335
rect 3565 3765 3585 3785
rect 3565 3715 3585 3735
rect 3565 3665 3585 3685
rect 3565 3615 3585 3635
rect 3565 3565 3585 3585
rect 3565 3515 3585 3535
rect 3565 3465 3585 3485
rect 3565 3415 3585 3435
rect 3565 3365 3585 3385
rect 3565 3315 3585 3335
rect 4165 3765 4185 3785
rect 4165 3715 4185 3735
rect 4165 3665 4185 3685
rect 4165 3615 4185 3635
rect 4165 3565 4185 3585
rect 4165 3515 4185 3535
rect 4165 3465 4185 3485
rect 4165 3415 4185 3435
rect 4765 3765 4785 3785
rect 4765 3715 4785 3735
rect 4765 3665 4785 3685
rect 4765 3615 4785 3635
rect 4765 3565 4785 3585
rect 4765 3515 4785 3535
rect 4765 3465 4785 3485
rect 4765 3415 4785 3435
rect 4765 3365 4785 3385
rect 4765 3315 4785 3335
rect 4915 3665 4935 3685
rect 4915 3615 4935 3635
rect 4915 3565 4935 3585
rect 4915 3515 4935 3535
rect 4915 3465 4935 3485
rect 4915 3415 4935 3435
rect 4915 3365 4935 3385
rect 4915 3315 4935 3335
rect 5065 3765 5085 3785
rect 5065 3715 5085 3735
rect 5065 3665 5085 3685
rect 5065 3615 5085 3635
rect 5065 3565 5085 3585
rect 5065 3515 5085 3535
rect 5065 3465 5085 3485
rect 5065 3415 5085 3435
rect 5215 3665 5235 3685
rect 5215 3615 5235 3635
rect 5215 3565 5235 3585
rect 5215 3515 5235 3535
rect 5215 3465 5235 3485
rect 5215 3415 5235 3435
rect 5215 3365 5235 3385
rect 5365 3765 5385 3785
rect 5365 3715 5385 3735
rect 5365 3665 5385 3685
rect 5365 3615 5385 3635
rect 5365 3565 5385 3585
rect 5365 3515 5385 3535
rect 5365 3465 5385 3485
rect 5365 3415 5385 3435
rect 5515 3665 5535 3685
rect 5515 3615 5535 3635
rect 5515 3565 5535 3585
rect 5515 3515 5535 3535
rect 5515 3465 5535 3485
rect 5515 3415 5535 3435
rect 5515 3365 5535 3385
rect 5665 3765 5685 3785
rect 5665 3715 5685 3735
rect 5665 3665 5685 3685
rect 5665 3615 5685 3635
rect 5665 3565 5685 3585
rect 5665 3515 5685 3535
rect 5665 3465 5685 3485
rect 5665 3415 5685 3435
rect 5815 3665 5835 3685
rect 5815 3615 5835 3635
rect 5815 3565 5835 3585
rect 5815 3515 5835 3535
rect 5815 3465 5835 3485
rect 5815 3415 5835 3435
rect 5815 3365 5835 3385
rect 5965 3765 5985 3785
rect 5965 3715 5985 3735
rect 5965 3665 5985 3685
rect 5965 3615 5985 3635
rect 5965 3565 5985 3585
rect 5965 3515 5985 3535
rect 5965 3465 5985 3485
rect 5965 3415 5985 3435
rect 5965 3365 5985 3385
rect 5965 3315 5985 3335
rect 6115 3665 6135 3685
rect 6115 3615 6135 3635
rect 6115 3565 6135 3585
rect 6115 3515 6135 3535
rect 6115 3465 6135 3485
rect 6115 3415 6135 3435
rect 6115 3365 6135 3385
rect 6115 3315 6135 3335
rect 6265 3765 6285 3785
rect 6265 3715 6285 3735
rect 6265 3665 6285 3685
rect 6265 3615 6285 3635
rect 6265 3565 6285 3585
rect 6265 3515 6285 3535
rect 6265 3465 6285 3485
rect 6265 3415 6285 3435
rect 6415 3665 6435 3685
rect 6415 3615 6435 3635
rect 6415 3565 6435 3585
rect 6415 3515 6435 3535
rect 6415 3465 6435 3485
rect 6415 3415 6435 3435
rect 6415 3365 6435 3385
rect 6415 3315 6435 3335
rect 6565 3765 6585 3785
rect 6565 3715 6585 3735
rect 6565 3665 6585 3685
rect 6565 3615 6585 3635
rect 6565 3565 6585 3585
rect 6565 3515 6585 3535
rect 6565 3465 6585 3485
rect 6565 3415 6585 3435
rect 6565 3365 6585 3385
rect 6565 3315 6585 3335
rect 6715 3665 6735 3685
rect 6715 3615 6735 3635
rect 6715 3565 6735 3585
rect 6715 3515 6735 3535
rect 6715 3465 6735 3485
rect 6715 3415 6735 3435
rect 6715 3365 6735 3385
rect 6865 3765 6885 3785
rect 6865 3715 6885 3735
rect 6865 3665 6885 3685
rect 6865 3615 6885 3635
rect 6865 3565 6885 3585
rect 6865 3515 6885 3535
rect 6865 3465 6885 3485
rect 6865 3415 6885 3435
rect 7015 3665 7035 3685
rect 7015 3615 7035 3635
rect 7015 3565 7035 3585
rect 7015 3515 7035 3535
rect 7015 3465 7035 3485
rect 7015 3415 7035 3435
rect 7015 3365 7035 3385
rect 7165 3765 7185 3785
rect 7165 3715 7185 3735
rect 7165 3665 7185 3685
rect 7165 3615 7185 3635
rect 7165 3565 7185 3585
rect 7165 3515 7185 3535
rect 7165 3465 7185 3485
rect 7165 3415 7185 3435
rect 7315 3665 7335 3685
rect 7315 3615 7335 3635
rect 7315 3565 7335 3585
rect 7315 3515 7335 3535
rect 7315 3465 7335 3485
rect 7315 3415 7335 3435
rect 7315 3365 7335 3385
rect 7465 3765 7485 3785
rect 7465 3715 7485 3735
rect 7465 3665 7485 3685
rect 7465 3615 7485 3635
rect 7465 3565 7485 3585
rect 7465 3515 7485 3535
rect 7465 3465 7485 3485
rect 7465 3415 7485 3435
rect 7615 3665 7635 3685
rect 7615 3615 7635 3635
rect 7615 3565 7635 3585
rect 7615 3515 7635 3535
rect 7615 3465 7635 3485
rect 7615 3415 7635 3435
rect 7615 3365 7635 3385
rect 7615 3315 7635 3335
rect 7765 3765 7785 3785
rect 7765 3715 7785 3735
rect 7765 3665 7785 3685
rect 7765 3615 7785 3635
rect 7765 3565 7785 3585
rect 7765 3515 7785 3535
rect 7765 3465 7785 3485
rect 7765 3415 7785 3435
rect 7765 3365 7785 3385
rect 7765 3315 7785 3335
rect 8365 3765 8385 3785
rect 8365 3715 8385 3735
rect 8365 3665 8385 3685
rect 8365 3615 8385 3635
rect 8365 3565 8385 3585
rect 8365 3515 8385 3535
rect 8365 3465 8385 3485
rect 8365 3415 8385 3435
rect 8365 3365 8385 3385
rect 8365 3315 8385 3335
rect 8515 3765 8535 3785
rect 8515 3715 8535 3735
rect 8515 3665 8535 3685
rect 8515 3615 8535 3635
rect 8515 3565 8535 3585
rect 8515 3515 8535 3535
rect 8515 3465 8535 3485
rect 8515 3415 8535 3435
rect 8515 3365 8535 3385
rect 8515 3315 8535 3335
rect 8665 3765 8685 3785
rect 8665 3715 8685 3735
rect 8665 3665 8685 3685
rect 8665 3615 8685 3635
rect 8665 3565 8685 3585
rect 8665 3515 8685 3535
rect 8665 3465 8685 3485
rect 8665 3415 8685 3435
rect 8665 3365 8685 3385
rect 8665 3315 8685 3335
rect 8815 3765 8835 3785
rect 8815 3715 8835 3735
rect 8815 3665 8835 3685
rect 8815 3615 8835 3635
rect 8815 3565 8835 3585
rect 8815 3515 8835 3535
rect 8815 3465 8835 3485
rect 8815 3415 8835 3435
rect 8815 3365 8835 3385
rect 8815 3315 8835 3335
rect 8965 3765 8985 3785
rect 8965 3715 8985 3735
rect 8965 3665 8985 3685
rect 8965 3615 8985 3635
rect 8965 3565 8985 3585
rect 8965 3515 8985 3535
rect 8965 3465 8985 3485
rect 8965 3415 8985 3435
rect 8965 3365 8985 3385
rect 8965 3315 8985 3335
rect 9115 3765 9135 3785
rect 9115 3715 9135 3735
rect 9115 3665 9135 3685
rect 9115 3615 9135 3635
rect 9115 3565 9135 3585
rect 9115 3515 9135 3535
rect 9115 3465 9135 3485
rect 9115 3415 9135 3435
rect 9115 3365 9135 3385
rect 9115 3315 9135 3335
rect 9265 3765 9285 3785
rect 9265 3715 9285 3735
rect 9265 3665 9285 3685
rect 9265 3615 9285 3635
rect 9265 3565 9285 3585
rect 9265 3515 9285 3535
rect 9265 3465 9285 3485
rect 9265 3415 9285 3435
rect 9265 3365 9285 3385
rect 9265 3315 9285 3335
rect 9415 3765 9435 3785
rect 9415 3715 9435 3735
rect 9415 3665 9435 3685
rect 9415 3615 9435 3635
rect 9415 3565 9435 3585
rect 9415 3515 9435 3535
rect 9415 3465 9435 3485
rect 9415 3415 9435 3435
rect 9415 3365 9435 3385
rect 9415 3315 9435 3335
rect 9565 3765 9585 3785
rect 9565 3715 9585 3735
rect 9565 3665 9585 3685
rect 9565 3615 9585 3635
rect 9565 3565 9585 3585
rect 9565 3515 9585 3535
rect 9565 3465 9585 3485
rect 9565 3415 9585 3435
rect 9565 3365 9585 3385
rect 9565 3315 9585 3335
rect 9715 3765 9735 3785
rect 9715 3715 9735 3735
rect 9715 3665 9735 3685
rect 9715 3615 9735 3635
rect 9715 3565 9735 3585
rect 9715 3515 9735 3535
rect 9715 3465 9735 3485
rect 9715 3415 9735 3435
rect 9715 3365 9735 3385
rect 9715 3315 9735 3335
rect 9865 3765 9885 3785
rect 9865 3715 9885 3735
rect 9865 3665 9885 3685
rect 9865 3615 9885 3635
rect 9865 3565 9885 3585
rect 9865 3515 9885 3535
rect 9865 3465 9885 3485
rect 9865 3415 9885 3435
rect 9865 3365 9885 3385
rect 9865 3315 9885 3335
rect 10015 3765 10035 3785
rect 10015 3715 10035 3735
rect 10015 3665 10035 3685
rect 10015 3615 10035 3635
rect 10015 3565 10035 3585
rect 10015 3515 10035 3535
rect 10015 3465 10035 3485
rect 10015 3415 10035 3435
rect 10015 3365 10035 3385
rect 10015 3315 10035 3335
rect 10165 3765 10185 3785
rect 10165 3715 10185 3735
rect 10165 3665 10185 3685
rect 10165 3615 10185 3635
rect 10165 3565 10185 3585
rect 10165 3515 10185 3535
rect 10165 3465 10185 3485
rect 10165 3415 10185 3435
rect 10165 3365 10185 3385
rect 10165 3315 10185 3335
rect 10315 3765 10335 3785
rect 10315 3715 10335 3735
rect 10315 3665 10335 3685
rect 10315 3615 10335 3635
rect 10315 3565 10335 3585
rect 10315 3515 10335 3535
rect 10315 3465 10335 3485
rect 10315 3415 10335 3435
rect 10315 3365 10335 3385
rect 10315 3315 10335 3335
rect 10465 3765 10485 3785
rect 10465 3715 10485 3735
rect 10465 3665 10485 3685
rect 10465 3615 10485 3635
rect 10465 3565 10485 3585
rect 10465 3515 10485 3535
rect 10465 3465 10485 3485
rect 10465 3415 10485 3435
rect 10465 3365 10485 3385
rect 10465 3315 10485 3335
rect 10615 3765 10635 3785
rect 10615 3715 10635 3735
rect 10615 3665 10635 3685
rect 10615 3615 10635 3635
rect 10615 3565 10635 3585
rect 10615 3515 10635 3535
rect 10615 3465 10635 3485
rect 10615 3415 10635 3435
rect 10615 3365 10635 3385
rect 10615 3315 10635 3335
rect 10765 3765 10785 3785
rect 10765 3715 10785 3735
rect 10765 3665 10785 3685
rect 10765 3615 10785 3635
rect 10765 3565 10785 3585
rect 10765 3515 10785 3535
rect 10765 3465 10785 3485
rect 10765 3415 10785 3435
rect 10765 3365 10785 3385
rect 10765 3315 10785 3335
rect 11365 3765 11385 3785
rect 11365 3715 11385 3735
rect 11365 3665 11385 3685
rect 11365 3615 11385 3635
rect 11365 3565 11385 3585
rect 11365 3515 11385 3535
rect 11365 3465 11385 3485
rect 11365 3415 11385 3435
rect 11365 3365 11385 3385
rect 11365 3315 11385 3335
rect 11965 3765 11985 3785
rect 11965 3715 11985 3735
rect 11965 3665 11985 3685
rect 11965 3615 11985 3635
rect 11965 3565 11985 3585
rect 11965 3515 11985 3535
rect 11965 3465 11985 3485
rect 11965 3415 11985 3435
rect 11965 3365 11985 3385
rect 11965 3315 11985 3335
rect 12565 3765 12585 3785
rect 12565 3715 12585 3735
rect 12565 3665 12585 3685
rect 12565 3615 12585 3635
rect 12565 3565 12585 3585
rect 12565 3515 12585 3535
rect 12565 3465 12585 3485
rect 12565 3415 12585 3435
rect 12565 3365 12585 3385
rect 12565 3315 12585 3335
rect 13165 3765 13185 3785
rect 13165 3715 13185 3735
rect 13165 3665 13185 3685
rect 13165 3615 13185 3635
rect 13165 3565 13185 3585
rect 13165 3515 13185 3535
rect 13165 3465 13185 3485
rect 13165 3415 13185 3435
rect 13165 3365 13185 3385
rect 13165 3315 13185 3335
rect 13765 3765 13785 3785
rect 13765 3715 13785 3735
rect 13765 3665 13785 3685
rect 13765 3615 13785 3635
rect 13765 3565 13785 3585
rect 13765 3515 13785 3535
rect 13765 3465 13785 3485
rect 13765 3415 13785 3435
rect 13765 3365 13785 3385
rect 13765 3315 13785 3335
rect 14365 3765 14385 3785
rect 14365 3715 14385 3735
rect 14365 3665 14385 3685
rect 14365 3615 14385 3635
rect 14365 3565 14385 3585
rect 14365 3515 14385 3535
rect 14365 3465 14385 3485
rect 14365 3415 14385 3435
rect 14365 3365 14385 3385
rect 14365 3315 14385 3335
rect 14965 3765 14985 3785
rect 14965 3715 14985 3735
rect 14965 3665 14985 3685
rect 14965 3615 14985 3635
rect 14965 3565 14985 3585
rect 14965 3515 14985 3535
rect 14965 3465 14985 3485
rect 14965 3415 14985 3435
rect 14965 3365 14985 3385
rect 14965 3315 14985 3335
rect 15565 3765 15585 3785
rect 15565 3715 15585 3735
rect 15565 3665 15585 3685
rect 15565 3615 15585 3635
rect 15565 3565 15585 3585
rect 15565 3515 15585 3535
rect 15565 3465 15585 3485
rect 15565 3415 15585 3435
rect 15565 3365 15585 3385
rect 15565 3315 15585 3335
rect 16165 3765 16185 3785
rect 16165 3715 16185 3735
rect 16165 3665 16185 3685
rect 16165 3615 16185 3635
rect 16165 3565 16185 3585
rect 16165 3515 16185 3535
rect 16165 3465 16185 3485
rect 16165 3415 16185 3435
rect 16165 3365 16185 3385
rect 16165 3315 16185 3335
rect 16315 3665 16335 3685
rect 16315 3615 16335 3635
rect 16315 3565 16335 3585
rect 16315 3515 16335 3535
rect 16315 3465 16335 3485
rect 16315 3415 16335 3435
rect 16315 3365 16335 3385
rect 16315 3315 16335 3335
rect 16465 3765 16485 3785
rect 16465 3715 16485 3735
rect 16465 3665 16485 3685
rect 16465 3615 16485 3635
rect 16465 3565 16485 3585
rect 16465 3515 16485 3535
rect 16465 3465 16485 3485
rect 16465 3415 16485 3435
rect 16615 3665 16635 3685
rect 16615 3615 16635 3635
rect 16615 3565 16635 3585
rect 16615 3515 16635 3535
rect 16615 3465 16635 3485
rect 16615 3415 16635 3435
rect 16615 3365 16635 3385
rect 16615 3315 16635 3335
rect 16765 3765 16785 3785
rect 16765 3715 16785 3735
rect 16765 3665 16785 3685
rect 16765 3615 16785 3635
rect 16765 3565 16785 3585
rect 16765 3515 16785 3535
rect 16765 3465 16785 3485
rect 16765 3415 16785 3435
rect 16915 3665 16935 3685
rect 16915 3615 16935 3635
rect 16915 3565 16935 3585
rect 16915 3515 16935 3535
rect 16915 3465 16935 3485
rect 16915 3415 16935 3435
rect 16915 3365 16935 3385
rect 16915 3315 16935 3335
rect 17065 3765 17085 3785
rect 17065 3715 17085 3735
rect 17065 3665 17085 3685
rect 17065 3615 17085 3635
rect 17065 3565 17085 3585
rect 17065 3515 17085 3535
rect 17065 3465 17085 3485
rect 17065 3415 17085 3435
rect 17215 3665 17235 3685
rect 17215 3615 17235 3635
rect 17215 3565 17235 3585
rect 17215 3515 17235 3535
rect 17215 3465 17235 3485
rect 17215 3415 17235 3435
rect 17215 3365 17235 3385
rect 17215 3315 17235 3335
rect 17365 3765 17385 3785
rect 17365 3715 17385 3735
rect 17365 3665 17385 3685
rect 17365 3615 17385 3635
rect 17365 3565 17385 3585
rect 17365 3515 17385 3535
rect 17365 3465 17385 3485
rect 17365 3415 17385 3435
rect 17365 3365 17385 3385
rect 17365 3315 17385 3335
rect 17965 3665 17985 3685
rect 17965 3615 17985 3635
rect 17965 3565 17985 3585
rect 17965 3515 17985 3535
rect 17965 3465 17985 3485
rect 17965 3415 17985 3435
rect 17965 3365 17985 3385
rect 17965 3315 17985 3335
rect 18565 3765 18585 3785
rect 18565 3715 18585 3735
rect 18565 3665 18585 3685
rect 18565 3615 18585 3635
rect 18565 3565 18585 3585
rect 18565 3515 18585 3535
rect 18565 3465 18585 3485
rect 18565 3415 18585 3435
rect 18565 3365 18585 3385
rect 18565 3315 18585 3335
rect 18715 3665 18735 3685
rect 18715 3615 18735 3635
rect 18715 3565 18735 3585
rect 18715 3515 18735 3535
rect 18715 3465 18735 3485
rect 18715 3415 18735 3435
rect 18715 3365 18735 3385
rect 18715 3315 18735 3335
rect 18865 3765 18885 3785
rect 18865 3715 18885 3735
rect 18865 3665 18885 3685
rect 18865 3615 18885 3635
rect 18865 3565 18885 3585
rect 18865 3515 18885 3535
rect 18865 3465 18885 3485
rect 18865 3415 18885 3435
rect 19015 3665 19035 3685
rect 19015 3615 19035 3635
rect 19015 3565 19035 3585
rect 19015 3515 19035 3535
rect 19015 3465 19035 3485
rect 19015 3415 19035 3435
rect 19015 3365 19035 3385
rect 19015 3315 19035 3335
rect 19165 3765 19185 3785
rect 19165 3715 19185 3735
rect 19165 3665 19185 3685
rect 19165 3615 19185 3635
rect 19165 3565 19185 3585
rect 19165 3515 19185 3535
rect 19165 3465 19185 3485
rect 19165 3415 19185 3435
rect 19315 3665 19335 3685
rect 19315 3615 19335 3635
rect 19315 3565 19335 3585
rect 19315 3515 19335 3535
rect 19315 3465 19335 3485
rect 19315 3415 19335 3435
rect 19315 3365 19335 3385
rect 19315 3315 19335 3335
rect 19465 3765 19485 3785
rect 19465 3715 19485 3735
rect 19465 3665 19485 3685
rect 19465 3615 19485 3635
rect 19465 3565 19485 3585
rect 19465 3515 19485 3535
rect 19465 3465 19485 3485
rect 19465 3415 19485 3435
rect 19615 3665 19635 3685
rect 19615 3615 19635 3635
rect 19615 3565 19635 3585
rect 19615 3515 19635 3535
rect 19615 3465 19635 3485
rect 19615 3415 19635 3435
rect 19615 3365 19635 3385
rect 19615 3315 19635 3335
rect 19765 3765 19785 3785
rect 19765 3715 19785 3735
rect 19765 3665 19785 3685
rect 19765 3615 19785 3635
rect 19765 3565 19785 3585
rect 19765 3515 19785 3535
rect 19765 3465 19785 3485
rect 19765 3415 19785 3435
rect 19765 3365 19785 3385
rect 19765 3315 19785 3335
rect 20365 3765 20385 3785
rect 20365 3715 20385 3735
rect 20365 3665 20385 3685
rect 20365 3615 20385 3635
rect 20365 3565 20385 3585
rect 20365 3515 20385 3535
rect 20365 3465 20385 3485
rect 20365 3415 20385 3435
rect 20365 3365 20385 3385
rect 20365 3315 20385 3335
rect -485 3215 -465 3235
rect -185 3215 -165 3235
rect 115 3215 135 3235
rect 415 3215 435 3235
rect 715 3215 735 3235
rect 1015 3215 1035 3235
rect 1315 3215 1335 3235
rect 1615 3215 1635 3235
rect 1915 3215 1935 3235
rect 2215 3215 2235 3235
rect 2515 3215 2535 3235
rect 2815 3215 2835 3235
rect 3115 3215 3135 3235
rect 3415 3215 3435 3235
rect 3715 3215 3735 3235
rect 4015 3215 4035 3235
rect 4315 3215 4335 3235
rect 4615 3215 4635 3235
rect 4915 3215 4935 3235
rect 5215 3215 5235 3235
rect 5515 3215 5535 3235
rect 5815 3215 5835 3235
rect 6115 3215 6135 3235
rect 6415 3215 6435 3235
rect 6715 3215 6735 3235
rect 7015 3215 7035 3235
rect 7315 3215 7335 3235
rect 7615 3215 7635 3235
rect 7915 3215 7935 3235
rect 8215 3215 8235 3235
rect 8515 3215 8535 3235
rect 8815 3215 8835 3235
rect 9115 3215 9135 3235
rect 9415 3215 9435 3235
rect 9715 3215 9735 3235
rect 10015 3215 10035 3235
rect 10315 3215 10335 3235
rect 10615 3215 10635 3235
rect 10915 3215 10935 3235
rect 11215 3215 11235 3235
rect 11515 3215 11535 3235
rect 11815 3215 11835 3235
rect 12115 3215 12135 3235
rect 12415 3215 12435 3235
rect 12715 3215 12735 3235
rect 13015 3215 13035 3235
rect 13315 3215 13335 3235
rect 13615 3215 13635 3235
rect 13915 3215 13935 3235
rect 14215 3215 14235 3235
rect 14515 3215 14535 3235
rect 14815 3215 14835 3235
rect 15115 3215 15135 3235
rect 15415 3215 15435 3235
rect 15715 3215 15735 3235
rect 16015 3215 16035 3235
rect 16315 3215 16335 3235
rect 16615 3215 16635 3235
rect 16915 3215 16935 3235
rect 17215 3215 17235 3235
rect 17515 3215 17535 3235
rect 17815 3215 17835 3235
rect 18115 3215 18135 3235
rect 18415 3215 18435 3235
rect 18715 3215 18735 3235
rect 19015 3215 19035 3235
rect 19315 3215 19335 3235
rect 19615 3215 19635 3235
rect 19915 3215 19935 3235
rect 20215 3215 20235 3235
rect -635 3115 -615 3135
rect -635 3065 -615 3085
rect -635 3015 -615 3035
rect -635 2965 -615 2985
rect -635 2915 -615 2935
rect -635 2865 -615 2885
rect -635 2815 -615 2835
rect -635 2765 -615 2785
rect -635 2715 -615 2735
rect -635 2665 -615 2685
rect -485 3115 -465 3135
rect -485 3065 -465 3085
rect -485 3015 -465 3035
rect -485 2965 -465 2985
rect -485 2915 -465 2935
rect -485 2865 -465 2885
rect -485 2815 -465 2835
rect -485 2765 -465 2785
rect -485 2715 -465 2735
rect -485 2665 -465 2685
rect -335 3015 -315 3035
rect -335 2965 -315 2985
rect -335 2915 -315 2935
rect -335 2865 -315 2885
rect -335 2815 -315 2835
rect -335 2765 -315 2785
rect -335 2715 -315 2735
rect -335 2665 -315 2685
rect -185 3115 -165 3135
rect -185 3065 -165 3085
rect -185 3015 -165 3035
rect -185 2965 -165 2985
rect -185 2915 -165 2935
rect -185 2865 -165 2885
rect -185 2815 -165 2835
rect -185 2765 -165 2785
rect -185 2715 -165 2735
rect -185 2665 -165 2685
rect -35 3015 -15 3035
rect -35 2965 -15 2985
rect -35 2915 -15 2935
rect -35 2865 -15 2885
rect -35 2815 -15 2835
rect -35 2765 -15 2785
rect -35 2715 -15 2735
rect -35 2665 -15 2685
rect 565 3115 585 3135
rect 565 3065 585 3085
rect 565 3015 585 3035
rect 565 2965 585 2985
rect 565 2915 585 2935
rect 565 2865 585 2885
rect 565 2815 585 2835
rect 565 2765 585 2785
rect 565 2715 585 2735
rect 565 2665 585 2685
rect 715 3115 735 3135
rect 715 3065 735 3085
rect 715 3015 735 3035
rect 715 2965 735 2985
rect 715 2915 735 2935
rect 715 2865 735 2885
rect 715 2815 735 2835
rect 715 2765 735 2785
rect 865 3015 885 3035
rect 865 2965 885 2985
rect 865 2915 885 2935
rect 865 2865 885 2885
rect 865 2815 885 2835
rect 865 2765 885 2785
rect 865 2715 885 2735
rect 865 2665 885 2685
rect 1015 3115 1035 3135
rect 1015 3065 1035 3085
rect 1015 3015 1035 3035
rect 1015 2965 1035 2985
rect 1015 2915 1035 2935
rect 1015 2865 1035 2885
rect 1015 2815 1035 2835
rect 1015 2765 1035 2785
rect 1165 3015 1185 3035
rect 1165 2965 1185 2985
rect 1165 2915 1185 2935
rect 1165 2865 1185 2885
rect 1165 2815 1185 2835
rect 1165 2765 1185 2785
rect 1165 2715 1185 2735
rect 1165 2665 1185 2685
rect 1315 3115 1335 3135
rect 1315 3065 1335 3085
rect 1315 3015 1335 3035
rect 1315 2965 1335 2985
rect 1315 2915 1335 2935
rect 1315 2865 1335 2885
rect 1315 2815 1335 2835
rect 1315 2765 1335 2785
rect 1465 3015 1485 3035
rect 1465 2965 1485 2985
rect 1465 2915 1485 2935
rect 1465 2865 1485 2885
rect 1465 2815 1485 2835
rect 1465 2765 1485 2785
rect 1465 2715 1485 2735
rect 1465 2665 1485 2685
rect 1615 3115 1635 3135
rect 1615 3065 1635 3085
rect 1615 3015 1635 3035
rect 1615 2965 1635 2985
rect 1615 2915 1635 2935
rect 1615 2865 1635 2885
rect 1615 2815 1635 2835
rect 1615 2765 1635 2785
rect 1765 3115 1785 3135
rect 1765 3065 1785 3085
rect 1765 3015 1785 3035
rect 1765 2965 1785 2985
rect 1765 2915 1785 2935
rect 1765 2865 1785 2885
rect 1765 2815 1785 2835
rect 1765 2765 1785 2785
rect 1765 2715 1785 2735
rect 1765 2665 1785 2685
rect 1915 3115 1935 3135
rect 1915 3065 1935 3085
rect 1915 3015 1935 3035
rect 1915 2965 1935 2985
rect 1915 2915 1935 2935
rect 1915 2865 1935 2885
rect 1915 2815 1935 2835
rect 1915 2765 1935 2785
rect 2065 3015 2085 3035
rect 2065 2965 2085 2985
rect 2065 2915 2085 2935
rect 2065 2865 2085 2885
rect 2065 2815 2085 2835
rect 2065 2765 2085 2785
rect 2065 2715 2085 2735
rect 2065 2665 2085 2685
rect 2215 3115 2235 3135
rect 2215 3065 2235 3085
rect 2215 3015 2235 3035
rect 2215 2965 2235 2985
rect 2215 2915 2235 2935
rect 2215 2865 2235 2885
rect 2215 2815 2235 2835
rect 2215 2765 2235 2785
rect 2365 3115 2385 3135
rect 2365 3065 2385 3085
rect 2365 3015 2385 3035
rect 2365 2965 2385 2985
rect 2365 2915 2385 2935
rect 2365 2865 2385 2885
rect 2365 2815 2385 2835
rect 2365 2765 2385 2785
rect 2365 2715 2385 2735
rect 2365 2665 2385 2685
rect 2515 3115 2535 3135
rect 2515 3065 2535 3085
rect 2515 3015 2535 3035
rect 2515 2965 2535 2985
rect 2515 2915 2535 2935
rect 2515 2865 2535 2885
rect 2515 2815 2535 2835
rect 2515 2765 2535 2785
rect 2665 3015 2685 3035
rect 2665 2965 2685 2985
rect 2665 2915 2685 2935
rect 2665 2865 2685 2885
rect 2665 2815 2685 2835
rect 2665 2765 2685 2785
rect 2665 2715 2685 2735
rect 2665 2665 2685 2685
rect 2815 3115 2835 3135
rect 2815 3065 2835 3085
rect 2815 3015 2835 3035
rect 2815 2965 2835 2985
rect 2815 2915 2835 2935
rect 2815 2865 2835 2885
rect 2815 2815 2835 2835
rect 2815 2765 2835 2785
rect 2965 3015 2985 3035
rect 2965 2965 2985 2985
rect 2965 2915 2985 2935
rect 2965 2865 2985 2885
rect 2965 2815 2985 2835
rect 2965 2765 2985 2785
rect 2965 2715 2985 2735
rect 2965 2665 2985 2685
rect 3115 3115 3135 3135
rect 3115 3065 3135 3085
rect 3115 3015 3135 3035
rect 3115 2965 3135 2985
rect 3115 2915 3135 2935
rect 3115 2865 3135 2885
rect 3115 2815 3135 2835
rect 3115 2765 3135 2785
rect 3265 3015 3285 3035
rect 3265 2965 3285 2985
rect 3265 2915 3285 2935
rect 3265 2865 3285 2885
rect 3265 2815 3285 2835
rect 3265 2765 3285 2785
rect 3265 2715 3285 2735
rect 3265 2665 3285 2685
rect 3415 3115 3435 3135
rect 3415 3065 3435 3085
rect 3415 3015 3435 3035
rect 3415 2965 3435 2985
rect 3415 2915 3435 2935
rect 3415 2865 3435 2885
rect 3415 2815 3435 2835
rect 3415 2765 3435 2785
rect 3565 3115 3585 3135
rect 3565 3065 3585 3085
rect 3565 3015 3585 3035
rect 3565 2965 3585 2985
rect 3565 2915 3585 2935
rect 3565 2865 3585 2885
rect 3565 2815 3585 2835
rect 3565 2765 3585 2785
rect 3565 2715 3585 2735
rect 3565 2665 3585 2685
rect 4165 3015 4185 3035
rect 4165 2965 4185 2985
rect 4165 2915 4185 2935
rect 4165 2865 4185 2885
rect 4165 2815 4185 2835
rect 4165 2765 4185 2785
rect 4165 2715 4185 2735
rect 4165 2665 4185 2685
rect 4765 3115 4785 3135
rect 4765 3065 4785 3085
rect 4765 3015 4785 3035
rect 4765 2965 4785 2985
rect 4765 2915 4785 2935
rect 4765 2865 4785 2885
rect 4765 2815 4785 2835
rect 4765 2765 4785 2785
rect 4765 2715 4785 2735
rect 4765 2665 4785 2685
rect 4915 3115 4935 3135
rect 4915 3065 4935 3085
rect 4915 3015 4935 3035
rect 4915 2965 4935 2985
rect 4915 2915 4935 2935
rect 4915 2865 4935 2885
rect 4915 2815 4935 2835
rect 4915 2765 4935 2785
rect 5065 3015 5085 3035
rect 5065 2965 5085 2985
rect 5065 2915 5085 2935
rect 5065 2865 5085 2885
rect 5065 2815 5085 2835
rect 5065 2765 5085 2785
rect 5065 2715 5085 2735
rect 5065 2665 5085 2685
rect 5215 3115 5235 3135
rect 5215 3065 5235 3085
rect 5215 3015 5235 3035
rect 5215 2965 5235 2985
rect 5215 2915 5235 2935
rect 5215 2865 5235 2885
rect 5215 2815 5235 2835
rect 5215 2765 5235 2785
rect 5365 3015 5385 3035
rect 5365 2965 5385 2985
rect 5365 2915 5385 2935
rect 5365 2865 5385 2885
rect 5365 2815 5385 2835
rect 5365 2765 5385 2785
rect 5365 2715 5385 2735
rect 5365 2665 5385 2685
rect 5515 3115 5535 3135
rect 5515 3065 5535 3085
rect 5515 3015 5535 3035
rect 5515 2965 5535 2985
rect 5515 2915 5535 2935
rect 5515 2865 5535 2885
rect 5515 2815 5535 2835
rect 5515 2765 5535 2785
rect 5665 3015 5685 3035
rect 5665 2965 5685 2985
rect 5665 2915 5685 2935
rect 5665 2865 5685 2885
rect 5665 2815 5685 2835
rect 5665 2765 5685 2785
rect 5665 2715 5685 2735
rect 5665 2665 5685 2685
rect 5815 3115 5835 3135
rect 5815 3065 5835 3085
rect 5815 3015 5835 3035
rect 5815 2965 5835 2985
rect 5815 2915 5835 2935
rect 5815 2865 5835 2885
rect 5815 2815 5835 2835
rect 5815 2765 5835 2785
rect 5965 3115 5985 3135
rect 5965 3065 5985 3085
rect 5965 3015 5985 3035
rect 5965 2965 5985 2985
rect 5965 2915 5985 2935
rect 5965 2865 5985 2885
rect 5965 2815 5985 2835
rect 5965 2765 5985 2785
rect 5965 2715 5985 2735
rect 5965 2665 5985 2685
rect 6115 3115 6135 3135
rect 6115 3065 6135 3085
rect 6115 3015 6135 3035
rect 6115 2965 6135 2985
rect 6115 2915 6135 2935
rect 6115 2865 6135 2885
rect 6115 2815 6135 2835
rect 6115 2765 6135 2785
rect 6265 3015 6285 3035
rect 6265 2965 6285 2985
rect 6265 2915 6285 2935
rect 6265 2865 6285 2885
rect 6265 2815 6285 2835
rect 6265 2765 6285 2785
rect 6265 2715 6285 2735
rect 6265 2665 6285 2685
rect 6415 3115 6435 3135
rect 6415 3065 6435 3085
rect 6415 3015 6435 3035
rect 6415 2965 6435 2985
rect 6415 2915 6435 2935
rect 6415 2865 6435 2885
rect 6415 2815 6435 2835
rect 6415 2765 6435 2785
rect 6565 3115 6585 3135
rect 6565 3065 6585 3085
rect 6565 3015 6585 3035
rect 6565 2965 6585 2985
rect 6565 2915 6585 2935
rect 6565 2865 6585 2885
rect 6565 2815 6585 2835
rect 6565 2765 6585 2785
rect 6565 2715 6585 2735
rect 6565 2665 6585 2685
rect 6715 3115 6735 3135
rect 6715 3065 6735 3085
rect 6715 3015 6735 3035
rect 6715 2965 6735 2985
rect 6715 2915 6735 2935
rect 6715 2865 6735 2885
rect 6715 2815 6735 2835
rect 6715 2765 6735 2785
rect 6865 3015 6885 3035
rect 6865 2965 6885 2985
rect 6865 2915 6885 2935
rect 6865 2865 6885 2885
rect 6865 2815 6885 2835
rect 6865 2765 6885 2785
rect 6865 2715 6885 2735
rect 6865 2665 6885 2685
rect 7015 3115 7035 3135
rect 7015 3065 7035 3085
rect 7015 3015 7035 3035
rect 7015 2965 7035 2985
rect 7015 2915 7035 2935
rect 7015 2865 7035 2885
rect 7015 2815 7035 2835
rect 7015 2765 7035 2785
rect 7165 3015 7185 3035
rect 7165 2965 7185 2985
rect 7165 2915 7185 2935
rect 7165 2865 7185 2885
rect 7165 2815 7185 2835
rect 7165 2765 7185 2785
rect 7165 2715 7185 2735
rect 7165 2665 7185 2685
rect 7315 3115 7335 3135
rect 7315 3065 7335 3085
rect 7315 3015 7335 3035
rect 7315 2965 7335 2985
rect 7315 2915 7335 2935
rect 7315 2865 7335 2885
rect 7315 2815 7335 2835
rect 7315 2765 7335 2785
rect 7465 3015 7485 3035
rect 7465 2965 7485 2985
rect 7465 2915 7485 2935
rect 7465 2865 7485 2885
rect 7465 2815 7485 2835
rect 7465 2765 7485 2785
rect 7465 2715 7485 2735
rect 7465 2665 7485 2685
rect 7615 3115 7635 3135
rect 7615 3065 7635 3085
rect 7615 3015 7635 3035
rect 7615 2965 7635 2985
rect 7615 2915 7635 2935
rect 7615 2865 7635 2885
rect 7615 2815 7635 2835
rect 7615 2765 7635 2785
rect 7765 3115 7785 3135
rect 7765 3065 7785 3085
rect 7765 3015 7785 3035
rect 7765 2965 7785 2985
rect 7765 2915 7785 2935
rect 7765 2865 7785 2885
rect 7765 2815 7785 2835
rect 7765 2765 7785 2785
rect 7765 2715 7785 2735
rect 7765 2665 7785 2685
rect 8365 3115 8385 3135
rect 8365 3065 8385 3085
rect 8365 3015 8385 3035
rect 8365 2965 8385 2985
rect 8365 2915 8385 2935
rect 8365 2865 8385 2885
rect 8365 2815 8385 2835
rect 8365 2765 8385 2785
rect 8365 2715 8385 2735
rect 8365 2665 8385 2685
rect 8515 3115 8535 3135
rect 8515 3065 8535 3085
rect 8515 3015 8535 3035
rect 8515 2965 8535 2985
rect 8515 2915 8535 2935
rect 8515 2865 8535 2885
rect 8515 2815 8535 2835
rect 8515 2765 8535 2785
rect 8515 2715 8535 2735
rect 8515 2665 8535 2685
rect 8665 3115 8685 3135
rect 8665 3065 8685 3085
rect 8665 3015 8685 3035
rect 8665 2965 8685 2985
rect 8665 2915 8685 2935
rect 8665 2865 8685 2885
rect 8665 2815 8685 2835
rect 8665 2765 8685 2785
rect 8665 2715 8685 2735
rect 8665 2665 8685 2685
rect 8815 3115 8835 3135
rect 8815 3065 8835 3085
rect 8815 3015 8835 3035
rect 8815 2965 8835 2985
rect 8815 2915 8835 2935
rect 8815 2865 8835 2885
rect 8815 2815 8835 2835
rect 8815 2765 8835 2785
rect 8815 2715 8835 2735
rect 8815 2665 8835 2685
rect 8965 3115 8985 3135
rect 8965 3065 8985 3085
rect 8965 3015 8985 3035
rect 8965 2965 8985 2985
rect 8965 2915 8985 2935
rect 8965 2865 8985 2885
rect 8965 2815 8985 2835
rect 8965 2765 8985 2785
rect 8965 2715 8985 2735
rect 8965 2665 8985 2685
rect 9115 3115 9135 3135
rect 9115 3065 9135 3085
rect 9115 3015 9135 3035
rect 9115 2965 9135 2985
rect 9115 2915 9135 2935
rect 9115 2865 9135 2885
rect 9115 2815 9135 2835
rect 9115 2765 9135 2785
rect 9115 2715 9135 2735
rect 9115 2665 9135 2685
rect 9265 3115 9285 3135
rect 9265 3065 9285 3085
rect 9265 3015 9285 3035
rect 9265 2965 9285 2985
rect 9265 2915 9285 2935
rect 9265 2865 9285 2885
rect 9265 2815 9285 2835
rect 9265 2765 9285 2785
rect 9265 2715 9285 2735
rect 9265 2665 9285 2685
rect 9415 3115 9435 3135
rect 9415 3065 9435 3085
rect 9415 3015 9435 3035
rect 9415 2965 9435 2985
rect 9415 2915 9435 2935
rect 9415 2865 9435 2885
rect 9415 2815 9435 2835
rect 9415 2765 9435 2785
rect 9415 2715 9435 2735
rect 9415 2665 9435 2685
rect 9565 3115 9585 3135
rect 9565 3065 9585 3085
rect 9565 3015 9585 3035
rect 9565 2965 9585 2985
rect 9565 2915 9585 2935
rect 9565 2865 9585 2885
rect 9565 2815 9585 2835
rect 9565 2765 9585 2785
rect 9565 2715 9585 2735
rect 9565 2665 9585 2685
rect 9715 3115 9735 3135
rect 9715 3065 9735 3085
rect 9715 3015 9735 3035
rect 9715 2965 9735 2985
rect 9715 2915 9735 2935
rect 9715 2865 9735 2885
rect 9715 2815 9735 2835
rect 9715 2765 9735 2785
rect 9715 2715 9735 2735
rect 9715 2665 9735 2685
rect 9865 3115 9885 3135
rect 9865 3065 9885 3085
rect 9865 3015 9885 3035
rect 9865 2965 9885 2985
rect 9865 2915 9885 2935
rect 9865 2865 9885 2885
rect 9865 2815 9885 2835
rect 9865 2765 9885 2785
rect 9865 2715 9885 2735
rect 9865 2665 9885 2685
rect 10015 3115 10035 3135
rect 10015 3065 10035 3085
rect 10015 3015 10035 3035
rect 10015 2965 10035 2985
rect 10015 2915 10035 2935
rect 10015 2865 10035 2885
rect 10015 2815 10035 2835
rect 10015 2765 10035 2785
rect 10015 2715 10035 2735
rect 10015 2665 10035 2685
rect 10165 3115 10185 3135
rect 10165 3065 10185 3085
rect 10165 3015 10185 3035
rect 10165 2965 10185 2985
rect 10165 2915 10185 2935
rect 10165 2865 10185 2885
rect 10165 2815 10185 2835
rect 10165 2765 10185 2785
rect 10165 2715 10185 2735
rect 10165 2665 10185 2685
rect 10315 3115 10335 3135
rect 10315 3065 10335 3085
rect 10315 3015 10335 3035
rect 10315 2965 10335 2985
rect 10315 2915 10335 2935
rect 10315 2865 10335 2885
rect 10315 2815 10335 2835
rect 10315 2765 10335 2785
rect 10315 2715 10335 2735
rect 10315 2665 10335 2685
rect 10465 3115 10485 3135
rect 10465 3065 10485 3085
rect 10465 3015 10485 3035
rect 10465 2965 10485 2985
rect 10465 2915 10485 2935
rect 10465 2865 10485 2885
rect 10465 2815 10485 2835
rect 10465 2765 10485 2785
rect 10465 2715 10485 2735
rect 10465 2665 10485 2685
rect 10615 3115 10635 3135
rect 10615 3065 10635 3085
rect 10615 3015 10635 3035
rect 10615 2965 10635 2985
rect 10615 2915 10635 2935
rect 10615 2865 10635 2885
rect 10615 2815 10635 2835
rect 10615 2765 10635 2785
rect 10615 2715 10635 2735
rect 10615 2665 10635 2685
rect 10765 3115 10785 3135
rect 10765 3065 10785 3085
rect 10765 3015 10785 3035
rect 10765 2965 10785 2985
rect 10765 2915 10785 2935
rect 10765 2865 10785 2885
rect 10765 2815 10785 2835
rect 10765 2765 10785 2785
rect 10765 2715 10785 2735
rect 10765 2665 10785 2685
rect 11365 3115 11385 3135
rect 11365 3065 11385 3085
rect 11365 3015 11385 3035
rect 11365 2965 11385 2985
rect 11365 2915 11385 2935
rect 11365 2865 11385 2885
rect 11365 2815 11385 2835
rect 11365 2765 11385 2785
rect 11365 2715 11385 2735
rect 11365 2665 11385 2685
rect 11965 3115 11985 3135
rect 11965 3065 11985 3085
rect 11965 3015 11985 3035
rect 11965 2965 11985 2985
rect 11965 2915 11985 2935
rect 11965 2865 11985 2885
rect 11965 2815 11985 2835
rect 11965 2765 11985 2785
rect 11965 2715 11985 2735
rect 11965 2665 11985 2685
rect 12565 3115 12585 3135
rect 12565 3065 12585 3085
rect 12565 3015 12585 3035
rect 12565 2965 12585 2985
rect 12565 2915 12585 2935
rect 12565 2865 12585 2885
rect 12565 2815 12585 2835
rect 12565 2765 12585 2785
rect 12565 2715 12585 2735
rect 12565 2665 12585 2685
rect 13165 3115 13185 3135
rect 13165 3065 13185 3085
rect 13165 3015 13185 3035
rect 13165 2965 13185 2985
rect 13165 2915 13185 2935
rect 13165 2865 13185 2885
rect 13165 2815 13185 2835
rect 13165 2765 13185 2785
rect 13165 2715 13185 2735
rect 13165 2665 13185 2685
rect 13765 3115 13785 3135
rect 13765 3065 13785 3085
rect 13765 3015 13785 3035
rect 13765 2965 13785 2985
rect 13765 2915 13785 2935
rect 13765 2865 13785 2885
rect 13765 2815 13785 2835
rect 13765 2765 13785 2785
rect 13765 2715 13785 2735
rect 13765 2665 13785 2685
rect 14365 3115 14385 3135
rect 14365 3065 14385 3085
rect 14365 3015 14385 3035
rect 14365 2965 14385 2985
rect 14365 2915 14385 2935
rect 14365 2865 14385 2885
rect 14365 2815 14385 2835
rect 14365 2765 14385 2785
rect 14365 2715 14385 2735
rect 14365 2665 14385 2685
rect 14965 3115 14985 3135
rect 14965 3065 14985 3085
rect 14965 3015 14985 3035
rect 14965 2965 14985 2985
rect 14965 2915 14985 2935
rect 14965 2865 14985 2885
rect 14965 2815 14985 2835
rect 14965 2765 14985 2785
rect 14965 2715 14985 2735
rect 14965 2665 14985 2685
rect 15565 3115 15585 3135
rect 15565 3065 15585 3085
rect 15565 3015 15585 3035
rect 15565 2965 15585 2985
rect 15565 2915 15585 2935
rect 15565 2865 15585 2885
rect 15565 2815 15585 2835
rect 15565 2765 15585 2785
rect 15565 2715 15585 2735
rect 15565 2665 15585 2685
rect 16165 3115 16185 3135
rect 16165 3065 16185 3085
rect 16165 3015 16185 3035
rect 16165 2965 16185 2985
rect 16165 2915 16185 2935
rect 16165 2865 16185 2885
rect 16165 2815 16185 2835
rect 16165 2765 16185 2785
rect 16165 2715 16185 2735
rect 16165 2665 16185 2685
rect 16315 3115 16335 3135
rect 16315 3065 16335 3085
rect 16315 3015 16335 3035
rect 16315 2965 16335 2985
rect 16315 2915 16335 2935
rect 16315 2865 16335 2885
rect 16315 2815 16335 2835
rect 16315 2765 16335 2785
rect 16465 3015 16485 3035
rect 16465 2965 16485 2985
rect 16465 2915 16485 2935
rect 16465 2865 16485 2885
rect 16465 2815 16485 2835
rect 16465 2765 16485 2785
rect 16465 2715 16485 2735
rect 16465 2665 16485 2685
rect 16615 3115 16635 3135
rect 16615 3065 16635 3085
rect 16615 3015 16635 3035
rect 16615 2965 16635 2985
rect 16615 2915 16635 2935
rect 16615 2865 16635 2885
rect 16615 2815 16635 2835
rect 16615 2765 16635 2785
rect 16765 3015 16785 3035
rect 16765 2965 16785 2985
rect 16765 2915 16785 2935
rect 16765 2865 16785 2885
rect 16765 2815 16785 2835
rect 16765 2765 16785 2785
rect 16765 2715 16785 2735
rect 16765 2665 16785 2685
rect 16915 3115 16935 3135
rect 16915 3065 16935 3085
rect 16915 3015 16935 3035
rect 16915 2965 16935 2985
rect 16915 2915 16935 2935
rect 16915 2865 16935 2885
rect 16915 2815 16935 2835
rect 16915 2765 16935 2785
rect 17065 3015 17085 3035
rect 17065 2965 17085 2985
rect 17065 2915 17085 2935
rect 17065 2865 17085 2885
rect 17065 2815 17085 2835
rect 17065 2765 17085 2785
rect 17065 2715 17085 2735
rect 17065 2665 17085 2685
rect 17215 3115 17235 3135
rect 17215 3065 17235 3085
rect 17215 3015 17235 3035
rect 17215 2965 17235 2985
rect 17215 2915 17235 2935
rect 17215 2865 17235 2885
rect 17215 2815 17235 2835
rect 17215 2765 17235 2785
rect 17365 3115 17385 3135
rect 17365 3065 17385 3085
rect 17365 3015 17385 3035
rect 17365 2965 17385 2985
rect 17365 2915 17385 2935
rect 17365 2865 17385 2885
rect 17365 2815 17385 2835
rect 17365 2765 17385 2785
rect 17365 2715 17385 2735
rect 17365 2665 17385 2685
rect 17965 3115 17985 3135
rect 17965 3065 17985 3085
rect 17965 3015 17985 3035
rect 17965 2965 17985 2985
rect 17965 2915 17985 2935
rect 17965 2865 17985 2885
rect 17965 2815 17985 2835
rect 17965 2765 17985 2785
rect 18565 3115 18585 3135
rect 18565 3065 18585 3085
rect 18565 3015 18585 3035
rect 18565 2965 18585 2985
rect 18565 2915 18585 2935
rect 18565 2865 18585 2885
rect 18565 2815 18585 2835
rect 18565 2765 18585 2785
rect 18565 2715 18585 2735
rect 18565 2665 18585 2685
rect 18715 3115 18735 3135
rect 18715 3065 18735 3085
rect 18715 3015 18735 3035
rect 18715 2965 18735 2985
rect 18715 2915 18735 2935
rect 18715 2865 18735 2885
rect 18715 2815 18735 2835
rect 18715 2765 18735 2785
rect 18865 3015 18885 3035
rect 18865 2965 18885 2985
rect 18865 2915 18885 2935
rect 18865 2865 18885 2885
rect 18865 2815 18885 2835
rect 18865 2765 18885 2785
rect 18865 2715 18885 2735
rect 18865 2665 18885 2685
rect 19015 3115 19035 3135
rect 19015 3065 19035 3085
rect 19015 3015 19035 3035
rect 19015 2965 19035 2985
rect 19015 2915 19035 2935
rect 19015 2865 19035 2885
rect 19015 2815 19035 2835
rect 19015 2765 19035 2785
rect 19165 3015 19185 3035
rect 19165 2965 19185 2985
rect 19165 2915 19185 2935
rect 19165 2865 19185 2885
rect 19165 2815 19185 2835
rect 19165 2765 19185 2785
rect 19165 2715 19185 2735
rect 19165 2665 19185 2685
rect 19315 3115 19335 3135
rect 19315 3065 19335 3085
rect 19315 3015 19335 3035
rect 19315 2965 19335 2985
rect 19315 2915 19335 2935
rect 19315 2865 19335 2885
rect 19315 2815 19335 2835
rect 19315 2765 19335 2785
rect 19465 3015 19485 3035
rect 19465 2965 19485 2985
rect 19465 2915 19485 2935
rect 19465 2865 19485 2885
rect 19465 2815 19485 2835
rect 19465 2765 19485 2785
rect 19465 2715 19485 2735
rect 19465 2665 19485 2685
rect 19615 3115 19635 3135
rect 19615 3065 19635 3085
rect 19615 3015 19635 3035
rect 19615 2965 19635 2985
rect 19615 2915 19635 2935
rect 19615 2865 19635 2885
rect 19615 2815 19635 2835
rect 19615 2765 19635 2785
rect 19765 3115 19785 3135
rect 19765 3065 19785 3085
rect 19765 3015 19785 3035
rect 19765 2965 19785 2985
rect 19765 2915 19785 2935
rect 19765 2865 19785 2885
rect 19765 2815 19785 2835
rect 19765 2765 19785 2785
rect 19765 2715 19785 2735
rect 19765 2665 19785 2685
rect 20365 3115 20385 3135
rect 20365 3065 20385 3085
rect 20365 3015 20385 3035
rect 20365 2965 20385 2985
rect 20365 2915 20385 2935
rect 20365 2865 20385 2885
rect 20365 2815 20385 2835
rect 20365 2765 20385 2785
rect 20365 2715 20385 2735
rect 20365 2665 20385 2685
rect -635 2565 -615 2585
rect -35 2565 -15 2585
rect 4165 2565 4185 2585
rect 8365 2565 8385 2585
rect 8665 2565 8685 2585
rect 8965 2565 8985 2585
rect 9265 2565 9285 2585
rect 9565 2565 9585 2585
rect 9865 2565 9885 2585
rect 10165 2565 10185 2585
rect 10465 2565 10485 2585
rect 10765 2565 10785 2585
rect 11965 2565 11985 2585
rect 13165 2565 13185 2585
rect 14365 2565 14385 2585
rect 15565 2565 15585 2585
rect 17965 2565 17985 2585
rect 20365 2565 20385 2585
rect -635 1665 -615 1685
rect -35 1665 -15 1685
rect 8365 1665 8385 1685
rect 10765 1665 10785 1685
rect 15565 1665 15585 1685
rect 17965 1665 17985 1685
rect 20365 1665 20385 1685
rect -635 1565 -615 1585
rect -635 1515 -615 1535
rect -635 1465 -615 1485
rect -635 1415 -615 1435
rect -635 1365 -615 1385
rect -635 1315 -615 1335
rect -635 1265 -615 1285
rect -635 1215 -615 1235
rect -635 1165 -615 1185
rect -635 1115 -615 1135
rect -635 1065 -615 1085
rect -635 1015 -615 1035
rect -635 965 -615 985
rect -635 915 -615 935
rect -485 1565 -465 1585
rect -485 1515 -465 1535
rect -485 1465 -465 1485
rect -485 1415 -465 1435
rect -485 1365 -465 1385
rect -485 1315 -465 1335
rect -485 1265 -465 1285
rect -485 1215 -465 1235
rect -485 1165 -465 1185
rect -485 1115 -465 1135
rect -485 1065 -465 1085
rect -485 1015 -465 1035
rect -485 965 -465 985
rect -485 915 -465 935
rect -335 1565 -315 1585
rect -335 1515 -315 1535
rect -335 1465 -315 1485
rect -335 1415 -315 1435
rect -335 1365 -315 1385
rect -335 1315 -315 1335
rect -335 1265 -315 1285
rect -335 1215 -315 1235
rect -335 1165 -315 1185
rect -335 1115 -315 1135
rect -335 1065 -315 1085
rect -335 1015 -315 1035
rect -335 965 -315 985
rect -335 915 -315 935
rect -185 1565 -165 1585
rect -185 1515 -165 1535
rect -185 1465 -165 1485
rect -185 1415 -165 1435
rect -185 1365 -165 1385
rect -185 1315 -165 1335
rect -185 1265 -165 1285
rect -185 1215 -165 1235
rect -185 1165 -165 1185
rect -185 1115 -165 1135
rect -185 1065 -165 1085
rect -185 1015 -165 1035
rect -185 965 -165 985
rect -185 915 -165 935
rect -35 1565 -15 1585
rect -35 1515 -15 1535
rect -35 1465 -15 1485
rect -35 1415 -15 1435
rect -35 1365 -15 1385
rect -35 1315 -15 1335
rect -35 1265 -15 1285
rect -35 1215 -15 1235
rect -35 1165 -15 1185
rect -35 1115 -15 1135
rect -35 1065 -15 1085
rect -35 1015 -15 1035
rect -35 965 -15 985
rect -35 915 -15 935
rect 1165 1565 1185 1585
rect 1165 1515 1185 1535
rect 1165 1465 1185 1485
rect 1165 1415 1185 1435
rect 1165 1365 1185 1385
rect 1165 1315 1185 1335
rect 1165 1265 1185 1285
rect 1165 1215 1185 1235
rect 1165 1165 1185 1185
rect 1165 1115 1185 1135
rect 1165 1065 1185 1085
rect 1165 1015 1185 1035
rect 1165 965 1185 985
rect 1165 915 1185 935
rect 1465 1465 1485 1485
rect 1465 1415 1485 1435
rect 1465 1365 1485 1385
rect 1465 1315 1485 1335
rect 1465 1265 1485 1285
rect 1465 1215 1485 1235
rect 1465 1165 1485 1185
rect 1465 1115 1485 1135
rect 1465 1065 1485 1085
rect 1465 1015 1485 1035
rect 1465 965 1485 985
rect 1465 915 1485 935
rect 1765 1565 1785 1585
rect 1765 1515 1785 1535
rect 1765 1465 1785 1485
rect 1765 1415 1785 1435
rect 1765 1365 1785 1385
rect 1765 1315 1785 1335
rect 1765 1265 1785 1285
rect 1765 1215 1785 1235
rect 1765 1165 1785 1185
rect 1765 1115 1785 1135
rect 1765 1065 1785 1085
rect 1765 1015 1785 1035
rect 2065 1465 2085 1485
rect 2065 1415 2085 1435
rect 2065 1365 2085 1385
rect 2065 1315 2085 1335
rect 2065 1265 2085 1285
rect 2065 1215 2085 1235
rect 2065 1165 2085 1185
rect 2065 1115 2085 1135
rect 2065 1065 2085 1085
rect 2065 1015 2085 1035
rect 2065 965 2085 985
rect 2065 915 2085 935
rect 2365 1565 2385 1585
rect 2365 1515 2385 1535
rect 2365 1465 2385 1485
rect 2365 1415 2385 1435
rect 2365 1365 2385 1385
rect 2365 1315 2385 1335
rect 2365 1265 2385 1285
rect 2365 1215 2385 1235
rect 2365 1165 2385 1185
rect 2365 1115 2385 1135
rect 2365 1065 2385 1085
rect 2365 1015 2385 1035
rect 2665 1465 2685 1485
rect 2665 1415 2685 1435
rect 2665 1365 2685 1385
rect 2665 1315 2685 1335
rect 2665 1265 2685 1285
rect 2665 1215 2685 1235
rect 2665 1165 2685 1185
rect 2665 1115 2685 1135
rect 2665 1065 2685 1085
rect 2665 1015 2685 1035
rect 2665 965 2685 985
rect 2665 915 2685 935
rect 2965 1565 2985 1585
rect 2965 1515 2985 1535
rect 2965 1465 2985 1485
rect 2965 1415 2985 1435
rect 2965 1365 2985 1385
rect 2965 1315 2985 1335
rect 2965 1265 2985 1285
rect 2965 1215 2985 1235
rect 2965 1165 2985 1185
rect 2965 1115 2985 1135
rect 2965 1065 2985 1085
rect 2965 1015 2985 1035
rect 3265 1465 3285 1485
rect 3265 1415 3285 1435
rect 3265 1365 3285 1385
rect 3265 1315 3285 1335
rect 3265 1265 3285 1285
rect 3265 1215 3285 1235
rect 3265 1165 3285 1185
rect 3265 1115 3285 1135
rect 3265 1065 3285 1085
rect 3265 1015 3285 1035
rect 3265 965 3285 985
rect 3265 915 3285 935
rect 3565 1565 3585 1585
rect 3565 1515 3585 1535
rect 3565 1465 3585 1485
rect 3565 1415 3585 1435
rect 3565 1365 3585 1385
rect 3565 1315 3585 1335
rect 3565 1265 3585 1285
rect 3565 1215 3585 1235
rect 3565 1165 3585 1185
rect 3565 1115 3585 1135
rect 3565 1065 3585 1085
rect 3565 1015 3585 1035
rect 3565 965 3585 985
rect 3565 915 3585 935
rect 3715 1465 3735 1485
rect 3715 1415 3735 1435
rect 3715 1365 3735 1385
rect 3715 1315 3735 1335
rect 3715 1265 3735 1285
rect 3715 1215 3735 1235
rect 3715 1165 3735 1185
rect 3715 1115 3735 1135
rect 3715 1065 3735 1085
rect 3715 1015 3735 1035
rect 3715 965 3735 985
rect 3715 915 3735 935
rect 3865 1565 3885 1585
rect 3865 1515 3885 1535
rect 3865 1465 3885 1485
rect 3865 1415 3885 1435
rect 3865 1365 3885 1385
rect 3865 1315 3885 1335
rect 3865 1265 3885 1285
rect 3865 1215 3885 1235
rect 3865 1165 3885 1185
rect 3865 1115 3885 1135
rect 3865 1065 3885 1085
rect 3865 1015 3885 1035
rect 4015 1465 4035 1485
rect 4015 1415 4035 1435
rect 4015 1365 4035 1385
rect 4015 1315 4035 1335
rect 4015 1265 4035 1285
rect 4015 1215 4035 1235
rect 4015 1165 4035 1185
rect 4015 1115 4035 1135
rect 4015 1065 4035 1085
rect 4015 1015 4035 1035
rect 4015 965 4035 985
rect 4015 915 4035 935
rect 4165 1565 4185 1585
rect 4165 1515 4185 1535
rect 4165 1465 4185 1485
rect 4165 1415 4185 1435
rect 4165 1365 4185 1385
rect 4165 1315 4185 1335
rect 4165 1265 4185 1285
rect 4165 1215 4185 1235
rect 4165 1165 4185 1185
rect 4165 1115 4185 1135
rect 4165 1065 4185 1085
rect 4165 1015 4185 1035
rect 4165 965 4185 985
rect 4165 915 4185 935
rect 4315 1465 4335 1485
rect 4315 1415 4335 1435
rect 4315 1365 4335 1385
rect 4315 1315 4335 1335
rect 4315 1265 4335 1285
rect 4315 1215 4335 1235
rect 4315 1165 4335 1185
rect 4315 1115 4335 1135
rect 4315 1065 4335 1085
rect 4315 1015 4335 1035
rect 4315 965 4335 985
rect 4315 915 4335 935
rect 4465 1565 4485 1585
rect 4465 1515 4485 1535
rect 4465 1465 4485 1485
rect 4465 1415 4485 1435
rect 4465 1365 4485 1385
rect 4465 1315 4485 1335
rect 4465 1265 4485 1285
rect 4465 1215 4485 1235
rect 4465 1165 4485 1185
rect 4465 1115 4485 1135
rect 4465 1065 4485 1085
rect 4465 1015 4485 1035
rect 4615 1465 4635 1485
rect 4615 1415 4635 1435
rect 4615 1365 4635 1385
rect 4615 1315 4635 1335
rect 4615 1265 4635 1285
rect 4615 1215 4635 1235
rect 4615 1165 4635 1185
rect 4615 1115 4635 1135
rect 4615 1065 4635 1085
rect 4615 1015 4635 1035
rect 4615 965 4635 985
rect 4615 915 4635 935
rect 4765 1565 4785 1585
rect 4765 1515 4785 1535
rect 4765 1465 4785 1485
rect 4765 1415 4785 1435
rect 4765 1365 4785 1385
rect 4765 1315 4785 1335
rect 4765 1265 4785 1285
rect 4765 1215 4785 1235
rect 4765 1165 4785 1185
rect 4765 1115 4785 1135
rect 4765 1065 4785 1085
rect 4765 1015 4785 1035
rect 4765 965 4785 985
rect 4765 915 4785 935
rect 5065 1465 5085 1485
rect 5065 1415 5085 1435
rect 5065 1365 5085 1385
rect 5065 1315 5085 1335
rect 5065 1265 5085 1285
rect 5065 1215 5085 1235
rect 5065 1165 5085 1185
rect 5065 1115 5085 1135
rect 5065 1065 5085 1085
rect 5065 1015 5085 1035
rect 5065 965 5085 985
rect 5065 915 5085 935
rect 5365 1565 5385 1585
rect 5365 1515 5385 1535
rect 5365 1465 5385 1485
rect 5365 1415 5385 1435
rect 5365 1365 5385 1385
rect 5365 1315 5385 1335
rect 5365 1265 5385 1285
rect 5365 1215 5385 1235
rect 5365 1165 5385 1185
rect 5365 1115 5385 1135
rect 5365 1065 5385 1085
rect 5365 1015 5385 1035
rect 5665 1465 5685 1485
rect 5665 1415 5685 1435
rect 5665 1365 5685 1385
rect 5665 1315 5685 1335
rect 5665 1265 5685 1285
rect 5665 1215 5685 1235
rect 5665 1165 5685 1185
rect 5665 1115 5685 1135
rect 5665 1065 5685 1085
rect 5665 1015 5685 1035
rect 5665 965 5685 985
rect 5665 915 5685 935
rect 5965 1565 5985 1585
rect 5965 1515 5985 1535
rect 5965 1465 5985 1485
rect 5965 1415 5985 1435
rect 5965 1365 5985 1385
rect 5965 1315 5985 1335
rect 5965 1265 5985 1285
rect 5965 1215 5985 1235
rect 5965 1165 5985 1185
rect 5965 1115 5985 1135
rect 5965 1065 5985 1085
rect 5965 1015 5985 1035
rect 6265 1465 6285 1485
rect 6265 1415 6285 1435
rect 6265 1365 6285 1385
rect 6265 1315 6285 1335
rect 6265 1265 6285 1285
rect 6265 1215 6285 1235
rect 6265 1165 6285 1185
rect 6265 1115 6285 1135
rect 6265 1065 6285 1085
rect 6265 1015 6285 1035
rect 6265 965 6285 985
rect 6265 915 6285 935
rect 6565 1565 6585 1585
rect 6565 1515 6585 1535
rect 6565 1465 6585 1485
rect 6565 1415 6585 1435
rect 6565 1365 6585 1385
rect 6565 1315 6585 1335
rect 6565 1265 6585 1285
rect 6565 1215 6585 1235
rect 6565 1165 6585 1185
rect 6565 1115 6585 1135
rect 6565 1065 6585 1085
rect 6565 1015 6585 1035
rect 6865 1465 6885 1485
rect 6865 1415 6885 1435
rect 6865 1365 6885 1385
rect 6865 1315 6885 1335
rect 6865 1265 6885 1285
rect 6865 1215 6885 1235
rect 6865 1165 6885 1185
rect 6865 1115 6885 1135
rect 6865 1065 6885 1085
rect 6865 1015 6885 1035
rect 6865 965 6885 985
rect 6865 915 6885 935
rect 7165 1565 7185 1585
rect 7165 1515 7185 1535
rect 7165 1465 7185 1485
rect 7165 1415 7185 1435
rect 7165 1365 7185 1385
rect 7165 1315 7185 1335
rect 7165 1265 7185 1285
rect 7165 1215 7185 1235
rect 7165 1165 7185 1185
rect 7165 1115 7185 1135
rect 7165 1065 7185 1085
rect 7165 1015 7185 1035
rect 7165 965 7185 985
rect 7165 915 7185 935
rect 8365 1565 8385 1585
rect 8365 1515 8385 1535
rect 8365 1465 8385 1485
rect 8365 1415 8385 1435
rect 8365 1365 8385 1385
rect 8365 1315 8385 1335
rect 8365 1265 8385 1285
rect 8365 1215 8385 1235
rect 8365 1165 8385 1185
rect 8365 1115 8385 1135
rect 8365 1065 8385 1085
rect 8365 1015 8385 1035
rect 8365 965 8385 985
rect 8365 915 8385 935
rect 9565 1565 9585 1585
rect 9565 1515 9585 1535
rect 9565 1465 9585 1485
rect 9565 1415 9585 1435
rect 9565 1365 9585 1385
rect 9565 1315 9585 1335
rect 9565 1265 9585 1285
rect 9565 1215 9585 1235
rect 9565 1165 9585 1185
rect 9565 1115 9585 1135
rect 9565 1065 9585 1085
rect 9565 1015 9585 1035
rect 9565 965 9585 985
rect 9565 915 9585 935
rect 10765 1565 10785 1585
rect 10765 1515 10785 1535
rect 10765 1465 10785 1485
rect 10765 1415 10785 1435
rect 10765 1365 10785 1385
rect 10765 1315 10785 1335
rect 10765 1265 10785 1285
rect 10765 1215 10785 1235
rect 10765 1165 10785 1185
rect 10765 1115 10785 1135
rect 10765 1065 10785 1085
rect 10765 1015 10785 1035
rect 10765 965 10785 985
rect 10765 915 10785 935
rect 11965 1565 11985 1585
rect 11965 1515 11985 1535
rect 11965 1465 11985 1485
rect 11965 1415 11985 1435
rect 11965 1365 11985 1385
rect 11965 1315 11985 1335
rect 11965 1265 11985 1285
rect 11965 1215 11985 1235
rect 11965 1165 11985 1185
rect 11965 1115 11985 1135
rect 11965 1065 11985 1085
rect 11965 1015 11985 1035
rect 11965 965 11985 985
rect 11965 915 11985 935
rect 12265 1465 12285 1485
rect 12265 1415 12285 1435
rect 12265 1365 12285 1385
rect 12265 1315 12285 1335
rect 12265 1265 12285 1285
rect 12265 1215 12285 1235
rect 12265 1165 12285 1185
rect 12265 1115 12285 1135
rect 12265 1065 12285 1085
rect 12265 1015 12285 1035
rect 12265 965 12285 985
rect 12265 915 12285 935
rect 12565 1565 12585 1585
rect 12565 1515 12585 1535
rect 12565 1465 12585 1485
rect 12565 1415 12585 1435
rect 12565 1365 12585 1385
rect 12565 1315 12585 1335
rect 12565 1265 12585 1285
rect 12565 1215 12585 1235
rect 12565 1165 12585 1185
rect 12565 1115 12585 1135
rect 12565 1065 12585 1085
rect 12565 1015 12585 1035
rect 12865 1465 12885 1485
rect 12865 1415 12885 1435
rect 12865 1365 12885 1385
rect 12865 1315 12885 1335
rect 12865 1265 12885 1285
rect 12865 1215 12885 1235
rect 12865 1165 12885 1185
rect 12865 1115 12885 1135
rect 12865 1065 12885 1085
rect 12865 1015 12885 1035
rect 12865 965 12885 985
rect 12865 915 12885 935
rect 13165 1565 13185 1585
rect 13165 1515 13185 1535
rect 13165 1465 13185 1485
rect 13165 1415 13185 1435
rect 13165 1365 13185 1385
rect 13165 1315 13185 1335
rect 13165 1265 13185 1285
rect 13165 1215 13185 1235
rect 13165 1165 13185 1185
rect 13165 1115 13185 1135
rect 13165 1065 13185 1085
rect 13165 1015 13185 1035
rect 13465 1465 13485 1485
rect 13465 1415 13485 1435
rect 13465 1365 13485 1385
rect 13465 1315 13485 1335
rect 13465 1265 13485 1285
rect 13465 1215 13485 1235
rect 13465 1165 13485 1185
rect 13465 1115 13485 1135
rect 13465 1065 13485 1085
rect 13465 1015 13485 1035
rect 13465 965 13485 985
rect 13465 915 13485 935
rect 13765 1565 13785 1585
rect 13765 1515 13785 1535
rect 13765 1465 13785 1485
rect 13765 1415 13785 1435
rect 13765 1365 13785 1385
rect 13765 1315 13785 1335
rect 13765 1265 13785 1285
rect 13765 1215 13785 1235
rect 13765 1165 13785 1185
rect 13765 1115 13785 1135
rect 13765 1065 13785 1085
rect 13765 1015 13785 1035
rect 14065 1465 14085 1485
rect 14065 1415 14085 1435
rect 14065 1365 14085 1385
rect 14065 1315 14085 1335
rect 14065 1265 14085 1285
rect 14065 1215 14085 1235
rect 14065 1165 14085 1185
rect 14065 1115 14085 1135
rect 14065 1065 14085 1085
rect 14065 1015 14085 1035
rect 14065 965 14085 985
rect 14065 915 14085 935
rect 14365 1565 14385 1585
rect 14365 1515 14385 1535
rect 14365 1465 14385 1485
rect 14365 1415 14385 1435
rect 14365 1365 14385 1385
rect 14365 1315 14385 1335
rect 14365 1265 14385 1285
rect 14365 1215 14385 1235
rect 14365 1165 14385 1185
rect 14365 1115 14385 1135
rect 14365 1065 14385 1085
rect 14365 1015 14385 1035
rect 14365 965 14385 985
rect 14365 915 14385 935
rect 15565 1565 15585 1585
rect 15565 1515 15585 1535
rect 15565 1465 15585 1485
rect 15565 1415 15585 1435
rect 15565 1365 15585 1385
rect 15565 1315 15585 1335
rect 15565 1265 15585 1285
rect 15565 1215 15585 1235
rect 15565 1165 15585 1185
rect 15565 1115 15585 1135
rect 15565 1065 15585 1085
rect 15565 1015 15585 1035
rect 15565 965 15585 985
rect 15565 915 15585 935
rect 16765 1565 16785 1585
rect 16765 1515 16785 1535
rect 16765 1465 16785 1485
rect 16765 1415 16785 1435
rect 16765 1365 16785 1385
rect 16765 1315 16785 1335
rect 16765 1265 16785 1285
rect 16765 1215 16785 1235
rect 16765 1165 16785 1185
rect 16765 1115 16785 1135
rect 16765 1065 16785 1085
rect 16765 1015 16785 1035
rect 16765 965 16785 985
rect 16765 915 16785 935
rect 17965 1565 17985 1585
rect 17965 1515 17985 1535
rect 17965 1465 17985 1485
rect 17965 1415 17985 1435
rect 17965 1365 17985 1385
rect 17965 1315 17985 1335
rect 17965 1265 17985 1285
rect 17965 1215 17985 1235
rect 17965 1165 17985 1185
rect 17965 1115 17985 1135
rect 17965 1065 17985 1085
rect 17965 1015 17985 1035
rect 17965 965 17985 985
rect 17965 915 17985 935
rect 19165 1565 19185 1585
rect 19165 1515 19185 1535
rect 19165 1465 19185 1485
rect 19165 1415 19185 1435
rect 19165 1365 19185 1385
rect 19165 1315 19185 1335
rect 19165 1265 19185 1285
rect 19165 1215 19185 1235
rect 19165 1165 19185 1185
rect 19165 1115 19185 1135
rect 19165 1065 19185 1085
rect 19165 1015 19185 1035
rect 19165 965 19185 985
rect 19165 915 19185 935
rect 20365 1565 20385 1585
rect 20365 1515 20385 1535
rect 20365 1465 20385 1485
rect 20365 1415 20385 1435
rect 20365 1365 20385 1385
rect 20365 1315 20385 1335
rect 20365 1265 20385 1285
rect 20365 1215 20385 1235
rect 20365 1165 20385 1185
rect 20365 1115 20385 1135
rect 20365 1065 20385 1085
rect 20365 1015 20385 1035
rect 20365 965 20385 985
rect 20365 915 20385 935
rect -485 815 -465 835
rect -185 815 -165 835
rect 115 815 135 835
rect 415 815 435 835
rect 715 815 735 835
rect 1015 815 1035 835
rect 1315 815 1335 835
rect 1615 815 1635 835
rect 1915 815 1935 835
rect 2215 815 2235 835
rect 2515 815 2535 835
rect 2815 815 2835 835
rect 3115 815 3135 835
rect 3415 815 3435 835
rect 3715 815 3735 835
rect 4015 815 4035 835
rect 4315 815 4335 835
rect 4615 815 4635 835
rect 4915 815 4935 835
rect 5215 815 5235 835
rect 5515 815 5535 835
rect 5815 815 5835 835
rect 6115 815 6135 835
rect 6415 815 6435 835
rect 6715 815 6735 835
rect 7015 815 7035 835
rect 7315 815 7335 835
rect 7615 815 7635 835
rect 7915 815 7935 835
rect 8215 815 8235 835
rect 8515 815 8535 835
rect 8815 815 8835 835
rect 9115 815 9135 835
rect 9415 815 9435 835
rect 9715 815 9735 835
rect 10015 815 10035 835
rect 10315 815 10335 835
rect 10615 815 10635 835
rect 10915 815 10935 835
rect 11215 815 11235 835
rect 11515 815 11535 835
rect 11815 815 11835 835
rect 12115 815 12135 835
rect 12415 815 12435 835
rect 12715 815 12735 835
rect 13015 815 13035 835
rect 13315 815 13335 835
rect 13615 815 13635 835
rect 13915 815 13935 835
rect 14215 815 14235 835
rect 14515 815 14535 835
rect 14815 815 14835 835
rect 15115 815 15135 835
rect 15415 815 15435 835
rect 15715 815 15735 835
rect 16015 815 16035 835
rect 16315 815 16335 835
rect 16615 815 16635 835
rect 16915 815 16935 835
rect 17215 815 17235 835
rect 17515 815 17535 835
rect 17815 815 17835 835
rect 18115 815 18135 835
rect 18415 815 18435 835
rect 18715 815 18735 835
rect 19015 815 19035 835
rect 19315 815 19335 835
rect 19615 815 19635 835
rect 19915 815 19935 835
rect 20215 815 20235 835
rect -635 715 -615 735
rect -635 665 -615 685
rect -635 615 -615 635
rect -635 565 -615 585
rect -635 515 -615 535
rect -635 465 -615 485
rect -635 415 -615 435
rect -635 365 -615 385
rect -635 315 -615 335
rect -635 265 -615 285
rect -635 215 -615 235
rect -635 165 -615 185
rect -635 115 -615 135
rect -635 65 -615 85
rect -485 715 -465 735
rect -485 665 -465 685
rect -485 615 -465 635
rect -485 565 -465 585
rect -485 515 -465 535
rect -485 465 -465 485
rect -485 415 -465 435
rect -485 365 -465 385
rect -485 315 -465 335
rect -485 265 -465 285
rect -485 215 -465 235
rect -485 165 -465 185
rect -485 115 -465 135
rect -485 65 -465 85
rect -335 715 -315 735
rect -335 665 -315 685
rect -335 615 -315 635
rect -335 565 -315 585
rect -335 515 -315 535
rect -335 465 -315 485
rect -335 415 -315 435
rect -335 365 -315 385
rect -335 315 -315 335
rect -335 265 -315 285
rect -335 215 -315 235
rect -335 165 -315 185
rect -335 115 -315 135
rect -335 65 -315 85
rect -185 715 -165 735
rect -185 665 -165 685
rect -185 615 -165 635
rect -185 565 -165 585
rect -185 515 -165 535
rect -185 465 -165 485
rect -185 415 -165 435
rect -185 365 -165 385
rect -185 315 -165 335
rect -185 265 -165 285
rect -185 215 -165 235
rect -185 165 -165 185
rect -185 115 -165 135
rect -185 65 -165 85
rect -35 715 -15 735
rect -35 665 -15 685
rect -35 615 -15 635
rect -35 565 -15 585
rect -35 515 -15 535
rect -35 465 -15 485
rect -35 415 -15 435
rect -35 365 -15 385
rect -35 315 -15 335
rect -35 265 -15 285
rect -35 215 -15 235
rect -35 165 -15 185
rect -35 115 -15 135
rect -35 65 -15 85
rect 1165 715 1185 735
rect 1165 665 1185 685
rect 1165 615 1185 635
rect 1165 565 1185 585
rect 1165 515 1185 535
rect 1165 465 1185 485
rect 1165 415 1185 435
rect 1165 365 1185 385
rect 1165 315 1185 335
rect 1165 265 1185 285
rect 1165 215 1185 235
rect 1165 165 1185 185
rect 1165 115 1185 135
rect 1165 65 1185 85
rect 1465 715 1485 735
rect 1465 665 1485 685
rect 1465 615 1485 635
rect 1465 565 1485 585
rect 1465 515 1485 535
rect 1465 465 1485 485
rect 1465 415 1485 435
rect 1465 365 1485 385
rect 1465 315 1485 335
rect 1465 265 1485 285
rect 1465 215 1485 235
rect 1465 165 1485 185
rect 1765 615 1785 635
rect 1765 565 1785 585
rect 1765 515 1785 535
rect 1765 465 1785 485
rect 1765 415 1785 435
rect 1765 365 1785 385
rect 1765 315 1785 335
rect 1765 265 1785 285
rect 1765 215 1785 235
rect 1765 165 1785 185
rect 1765 115 1785 135
rect 1765 65 1785 85
rect 2065 715 2085 735
rect 2065 665 2085 685
rect 2065 615 2085 635
rect 2065 565 2085 585
rect 2065 515 2085 535
rect 2065 465 2085 485
rect 2065 415 2085 435
rect 2065 365 2085 385
rect 2065 315 2085 335
rect 2065 265 2085 285
rect 2065 215 2085 235
rect 2065 165 2085 185
rect 2365 615 2385 635
rect 2365 565 2385 585
rect 2365 515 2385 535
rect 2365 465 2385 485
rect 2365 415 2385 435
rect 2365 365 2385 385
rect 2365 315 2385 335
rect 2365 265 2385 285
rect 2365 215 2385 235
rect 2365 165 2385 185
rect 2365 115 2385 135
rect 2365 65 2385 85
rect 2665 715 2685 735
rect 2665 665 2685 685
rect 2665 615 2685 635
rect 2665 565 2685 585
rect 2665 515 2685 535
rect 2665 465 2685 485
rect 2665 415 2685 435
rect 2665 365 2685 385
rect 2665 315 2685 335
rect 2665 265 2685 285
rect 2665 215 2685 235
rect 2665 165 2685 185
rect 2965 615 2985 635
rect 2965 565 2985 585
rect 2965 515 2985 535
rect 2965 465 2985 485
rect 2965 415 2985 435
rect 2965 365 2985 385
rect 2965 315 2985 335
rect 2965 265 2985 285
rect 2965 215 2985 235
rect 2965 165 2985 185
rect 2965 115 2985 135
rect 2965 65 2985 85
rect 3265 715 3285 735
rect 3265 665 3285 685
rect 3265 615 3285 635
rect 3265 565 3285 585
rect 3265 515 3285 535
rect 3265 465 3285 485
rect 3265 415 3285 435
rect 3265 365 3285 385
rect 3265 315 3285 335
rect 3265 265 3285 285
rect 3265 215 3285 235
rect 3265 165 3285 185
rect 3565 715 3585 735
rect 3565 665 3585 685
rect 3565 615 3585 635
rect 3565 565 3585 585
rect 3565 515 3585 535
rect 3565 465 3585 485
rect 3565 415 3585 435
rect 3565 365 3585 385
rect 3565 315 3585 335
rect 3565 265 3585 285
rect 3565 215 3585 235
rect 3565 165 3585 185
rect 3565 115 3585 135
rect 3565 65 3585 85
rect 3715 715 3735 735
rect 3715 665 3735 685
rect 3715 615 3735 635
rect 3715 565 3735 585
rect 3715 515 3735 535
rect 3715 465 3735 485
rect 3715 415 3735 435
rect 3715 365 3735 385
rect 3715 315 3735 335
rect 3715 265 3735 285
rect 3715 215 3735 235
rect 3715 165 3735 185
rect 3865 615 3885 635
rect 3865 565 3885 585
rect 3865 515 3885 535
rect 3865 465 3885 485
rect 3865 415 3885 435
rect 3865 365 3885 385
rect 3865 315 3885 335
rect 3865 265 3885 285
rect 3865 215 3885 235
rect 3865 165 3885 185
rect 3865 115 3885 135
rect 3865 65 3885 85
rect 4015 715 4035 735
rect 4015 665 4035 685
rect 4015 615 4035 635
rect 4015 565 4035 585
rect 4015 515 4035 535
rect 4015 465 4035 485
rect 4015 415 4035 435
rect 4015 365 4035 385
rect 4015 315 4035 335
rect 4015 265 4035 285
rect 4015 215 4035 235
rect 4015 165 4035 185
rect 4165 715 4185 735
rect 4165 665 4185 685
rect 4165 615 4185 635
rect 4165 565 4185 585
rect 4165 515 4185 535
rect 4165 465 4185 485
rect 4165 415 4185 435
rect 4165 365 4185 385
rect 4165 315 4185 335
rect 4165 265 4185 285
rect 4165 215 4185 235
rect 4165 165 4185 185
rect 4165 115 4185 135
rect 4165 65 4185 85
rect 4315 715 4335 735
rect 4315 665 4335 685
rect 4315 615 4335 635
rect 4315 565 4335 585
rect 4315 515 4335 535
rect 4315 465 4335 485
rect 4315 415 4335 435
rect 4315 365 4335 385
rect 4315 315 4335 335
rect 4315 265 4335 285
rect 4315 215 4335 235
rect 4315 165 4335 185
rect 4465 615 4485 635
rect 4465 565 4485 585
rect 4465 515 4485 535
rect 4465 465 4485 485
rect 4465 415 4485 435
rect 4465 365 4485 385
rect 4465 315 4485 335
rect 4465 265 4485 285
rect 4465 215 4485 235
rect 4465 165 4485 185
rect 4465 115 4485 135
rect 4465 65 4485 85
rect 4615 715 4635 735
rect 4615 665 4635 685
rect 4615 615 4635 635
rect 4615 565 4635 585
rect 4615 515 4635 535
rect 4615 465 4635 485
rect 4615 415 4635 435
rect 4615 365 4635 385
rect 4615 315 4635 335
rect 4615 265 4635 285
rect 4615 215 4635 235
rect 4615 165 4635 185
rect 4765 715 4785 735
rect 4765 665 4785 685
rect 4765 615 4785 635
rect 4765 565 4785 585
rect 4765 515 4785 535
rect 4765 465 4785 485
rect 4765 415 4785 435
rect 4765 365 4785 385
rect 4765 315 4785 335
rect 4765 265 4785 285
rect 4765 215 4785 235
rect 4765 165 4785 185
rect 4765 115 4785 135
rect 4765 65 4785 85
rect 5065 715 5085 735
rect 5065 665 5085 685
rect 5065 615 5085 635
rect 5065 565 5085 585
rect 5065 515 5085 535
rect 5065 465 5085 485
rect 5065 415 5085 435
rect 5065 365 5085 385
rect 5065 315 5085 335
rect 5065 265 5085 285
rect 5065 215 5085 235
rect 5065 165 5085 185
rect 5365 615 5385 635
rect 5365 565 5385 585
rect 5365 515 5385 535
rect 5365 465 5385 485
rect 5365 415 5385 435
rect 5365 365 5385 385
rect 5365 315 5385 335
rect 5365 265 5385 285
rect 5365 215 5385 235
rect 5365 165 5385 185
rect 5365 115 5385 135
rect 5365 65 5385 85
rect 5665 715 5685 735
rect 5665 665 5685 685
rect 5665 615 5685 635
rect 5665 565 5685 585
rect 5665 515 5685 535
rect 5665 465 5685 485
rect 5665 415 5685 435
rect 5665 365 5685 385
rect 5665 315 5685 335
rect 5665 265 5685 285
rect 5665 215 5685 235
rect 5665 165 5685 185
rect 5965 615 5985 635
rect 5965 565 5985 585
rect 5965 515 5985 535
rect 5965 465 5985 485
rect 5965 415 5985 435
rect 5965 365 5985 385
rect 5965 315 5985 335
rect 5965 265 5985 285
rect 5965 215 5985 235
rect 5965 165 5985 185
rect 5965 115 5985 135
rect 5965 65 5985 85
rect 6265 715 6285 735
rect 6265 665 6285 685
rect 6265 615 6285 635
rect 6265 565 6285 585
rect 6265 515 6285 535
rect 6265 465 6285 485
rect 6265 415 6285 435
rect 6265 365 6285 385
rect 6265 315 6285 335
rect 6265 265 6285 285
rect 6265 215 6285 235
rect 6265 165 6285 185
rect 6565 615 6585 635
rect 6565 565 6585 585
rect 6565 515 6585 535
rect 6565 465 6585 485
rect 6565 415 6585 435
rect 6565 365 6585 385
rect 6565 315 6585 335
rect 6565 265 6585 285
rect 6565 215 6585 235
rect 6565 165 6585 185
rect 6565 115 6585 135
rect 6565 65 6585 85
rect 6865 715 6885 735
rect 6865 665 6885 685
rect 6865 615 6885 635
rect 6865 565 6885 585
rect 6865 515 6885 535
rect 6865 465 6885 485
rect 6865 415 6885 435
rect 6865 365 6885 385
rect 6865 315 6885 335
rect 6865 265 6885 285
rect 6865 215 6885 235
rect 6865 165 6885 185
rect 7165 715 7185 735
rect 7165 665 7185 685
rect 7165 615 7185 635
rect 7165 565 7185 585
rect 7165 515 7185 535
rect 7165 465 7185 485
rect 7165 415 7185 435
rect 7165 365 7185 385
rect 7165 315 7185 335
rect 7165 265 7185 285
rect 7165 215 7185 235
rect 7165 165 7185 185
rect 7165 115 7185 135
rect 7165 65 7185 85
rect 8365 715 8385 735
rect 8365 665 8385 685
rect 8365 615 8385 635
rect 8365 565 8385 585
rect 8365 515 8385 535
rect 8365 465 8385 485
rect 8365 415 8385 435
rect 8365 365 8385 385
rect 8365 315 8385 335
rect 8365 265 8385 285
rect 8365 215 8385 235
rect 8365 165 8385 185
rect 8365 115 8385 135
rect 8365 65 8385 85
rect 9565 715 9585 735
rect 9565 665 9585 685
rect 9565 615 9585 635
rect 9565 565 9585 585
rect 9565 515 9585 535
rect 9565 465 9585 485
rect 9565 415 9585 435
rect 9565 365 9585 385
rect 9565 315 9585 335
rect 9565 265 9585 285
rect 9565 215 9585 235
rect 9565 165 9585 185
rect 9565 115 9585 135
rect 9565 65 9585 85
rect 10765 715 10785 735
rect 10765 665 10785 685
rect 10765 615 10785 635
rect 10765 565 10785 585
rect 10765 515 10785 535
rect 10765 465 10785 485
rect 10765 415 10785 435
rect 10765 365 10785 385
rect 10765 315 10785 335
rect 10765 265 10785 285
rect 10765 215 10785 235
rect 10765 165 10785 185
rect 10765 115 10785 135
rect 10765 65 10785 85
rect 11965 715 11985 735
rect 11965 665 11985 685
rect 11965 615 11985 635
rect 11965 565 11985 585
rect 11965 515 11985 535
rect 11965 465 11985 485
rect 11965 415 11985 435
rect 11965 365 11985 385
rect 11965 315 11985 335
rect 11965 265 11985 285
rect 11965 215 11985 235
rect 11965 165 11985 185
rect 11965 115 11985 135
rect 11965 65 11985 85
rect 12265 715 12285 735
rect 12265 665 12285 685
rect 12265 615 12285 635
rect 12265 565 12285 585
rect 12265 515 12285 535
rect 12265 465 12285 485
rect 12265 415 12285 435
rect 12265 365 12285 385
rect 12265 315 12285 335
rect 12265 265 12285 285
rect 12265 215 12285 235
rect 12265 165 12285 185
rect 12565 615 12585 635
rect 12565 565 12585 585
rect 12565 515 12585 535
rect 12565 465 12585 485
rect 12565 415 12585 435
rect 12565 365 12585 385
rect 12565 315 12585 335
rect 12565 265 12585 285
rect 12565 215 12585 235
rect 12565 165 12585 185
rect 12565 115 12585 135
rect 12565 65 12585 85
rect 12865 715 12885 735
rect 12865 665 12885 685
rect 12865 615 12885 635
rect 12865 565 12885 585
rect 12865 515 12885 535
rect 12865 465 12885 485
rect 12865 415 12885 435
rect 12865 365 12885 385
rect 12865 315 12885 335
rect 12865 265 12885 285
rect 12865 215 12885 235
rect 12865 165 12885 185
rect 13165 615 13185 635
rect 13165 565 13185 585
rect 13165 515 13185 535
rect 13165 465 13185 485
rect 13165 415 13185 435
rect 13165 365 13185 385
rect 13165 315 13185 335
rect 13165 265 13185 285
rect 13165 215 13185 235
rect 13165 165 13185 185
rect 13165 115 13185 135
rect 13165 65 13185 85
rect 13465 715 13485 735
rect 13465 665 13485 685
rect 13465 615 13485 635
rect 13465 565 13485 585
rect 13465 515 13485 535
rect 13465 465 13485 485
rect 13465 415 13485 435
rect 13465 365 13485 385
rect 13465 315 13485 335
rect 13465 265 13485 285
rect 13465 215 13485 235
rect 13465 165 13485 185
rect 13765 615 13785 635
rect 13765 565 13785 585
rect 13765 515 13785 535
rect 13765 465 13785 485
rect 13765 415 13785 435
rect 13765 365 13785 385
rect 13765 315 13785 335
rect 13765 265 13785 285
rect 13765 215 13785 235
rect 13765 165 13785 185
rect 13765 115 13785 135
rect 13765 65 13785 85
rect 14065 715 14085 735
rect 14065 665 14085 685
rect 14065 615 14085 635
rect 14065 565 14085 585
rect 14065 515 14085 535
rect 14065 465 14085 485
rect 14065 415 14085 435
rect 14065 365 14085 385
rect 14065 315 14085 335
rect 14065 265 14085 285
rect 14065 215 14085 235
rect 14065 165 14085 185
rect 14365 715 14385 735
rect 14365 665 14385 685
rect 14365 615 14385 635
rect 14365 565 14385 585
rect 14365 515 14385 535
rect 14365 465 14385 485
rect 14365 415 14385 435
rect 14365 365 14385 385
rect 14365 315 14385 335
rect 14365 265 14385 285
rect 14365 215 14385 235
rect 14365 165 14385 185
rect 14365 115 14385 135
rect 14365 65 14385 85
rect 15565 715 15585 735
rect 15565 665 15585 685
rect 15565 615 15585 635
rect 15565 565 15585 585
rect 15565 515 15585 535
rect 15565 465 15585 485
rect 15565 415 15585 435
rect 15565 365 15585 385
rect 15565 315 15585 335
rect 15565 265 15585 285
rect 15565 215 15585 235
rect 15565 165 15585 185
rect 15565 115 15585 135
rect 15565 65 15585 85
rect 16765 715 16785 735
rect 16765 665 16785 685
rect 16765 615 16785 635
rect 16765 565 16785 585
rect 16765 515 16785 535
rect 16765 465 16785 485
rect 16765 415 16785 435
rect 16765 365 16785 385
rect 16765 315 16785 335
rect 16765 265 16785 285
rect 16765 215 16785 235
rect 16765 165 16785 185
rect 16765 115 16785 135
rect 16765 65 16785 85
rect 17965 715 17985 735
rect 17965 665 17985 685
rect 17965 615 17985 635
rect 17965 565 17985 585
rect 17965 515 17985 535
rect 17965 465 17985 485
rect 17965 415 17985 435
rect 17965 365 17985 385
rect 17965 315 17985 335
rect 17965 265 17985 285
rect 17965 215 17985 235
rect 17965 165 17985 185
rect 17965 115 17985 135
rect 17965 65 17985 85
rect 19165 715 19185 735
rect 19165 665 19185 685
rect 19165 615 19185 635
rect 19165 565 19185 585
rect 19165 515 19185 535
rect 19165 465 19185 485
rect 19165 415 19185 435
rect 19165 365 19185 385
rect 19165 315 19185 335
rect 19165 265 19185 285
rect 19165 215 19185 235
rect 19165 165 19185 185
rect 19165 115 19185 135
rect 19165 65 19185 85
rect 20365 715 20385 735
rect 20365 665 20385 685
rect 20365 615 20385 635
rect 20365 565 20385 585
rect 20365 515 20385 535
rect 20365 465 20385 485
rect 20365 415 20385 435
rect 20365 365 20385 385
rect 20365 315 20385 335
rect 20365 265 20385 285
rect 20365 215 20385 235
rect 20365 165 20385 185
rect 20365 115 20385 135
rect 20365 65 20385 85
rect -635 -35 -615 -15
rect -35 -35 -15 -15
rect 8365 -35 8385 -15
rect 10765 -35 10785 -15
rect 15565 -35 15585 -15
rect 17965 -35 17985 -15
rect 20365 -35 20385 -15
rect -635 -135 -615 -115
rect -635 -185 -615 -165
rect -635 -235 -615 -215
rect -635 -285 -615 -265
rect -635 -335 -615 -315
rect -635 -385 -615 -365
rect -635 -435 -615 -415
rect -635 -485 -615 -465
rect -635 -535 -615 -515
rect -635 -585 -615 -565
rect -635 -635 -615 -615
rect -635 -685 -615 -665
rect -635 -735 -615 -715
rect -635 -785 -615 -765
rect -485 -135 -465 -115
rect -485 -185 -465 -165
rect -485 -235 -465 -215
rect -485 -285 -465 -265
rect -485 -335 -465 -315
rect -485 -385 -465 -365
rect -485 -435 -465 -415
rect -485 -485 -465 -465
rect -485 -535 -465 -515
rect -485 -585 -465 -565
rect -485 -635 -465 -615
rect -485 -685 -465 -665
rect -485 -735 -465 -715
rect -485 -785 -465 -765
rect -335 -135 -315 -115
rect -335 -185 -315 -165
rect -335 -235 -315 -215
rect -335 -285 -315 -265
rect -335 -335 -315 -315
rect -335 -385 -315 -365
rect -335 -435 -315 -415
rect -335 -485 -315 -465
rect -335 -535 -315 -515
rect -335 -585 -315 -565
rect -335 -635 -315 -615
rect -335 -685 -315 -665
rect -335 -735 -315 -715
rect -335 -785 -315 -765
rect -185 -135 -165 -115
rect -185 -185 -165 -165
rect -185 -235 -165 -215
rect -185 -285 -165 -265
rect -185 -335 -165 -315
rect -185 -385 -165 -365
rect -185 -435 -165 -415
rect -185 -485 -165 -465
rect -185 -535 -165 -515
rect -185 -585 -165 -565
rect -185 -635 -165 -615
rect -185 -685 -165 -665
rect -185 -735 -165 -715
rect -185 -785 -165 -765
rect -35 -135 -15 -115
rect -35 -185 -15 -165
rect -35 -235 -15 -215
rect -35 -285 -15 -265
rect -35 -335 -15 -315
rect -35 -385 -15 -365
rect -35 -435 -15 -415
rect -35 -485 -15 -465
rect -35 -535 -15 -515
rect -35 -585 -15 -565
rect -35 -635 -15 -615
rect -35 -685 -15 -665
rect -35 -735 -15 -715
rect -35 -785 -15 -765
rect 1165 -135 1185 -115
rect 1165 -185 1185 -165
rect 1165 -235 1185 -215
rect 1165 -285 1185 -265
rect 1165 -335 1185 -315
rect 1165 -385 1185 -365
rect 1165 -435 1185 -415
rect 1165 -485 1185 -465
rect 1165 -535 1185 -515
rect 1165 -585 1185 -565
rect 1165 -635 1185 -615
rect 1165 -685 1185 -665
rect 1165 -735 1185 -715
rect 1165 -785 1185 -765
rect 1465 -235 1485 -215
rect 1465 -285 1485 -265
rect 1465 -335 1485 -315
rect 1465 -385 1485 -365
rect 1465 -435 1485 -415
rect 1465 -485 1485 -465
rect 1465 -535 1485 -515
rect 1465 -585 1485 -565
rect 1465 -635 1485 -615
rect 1465 -685 1485 -665
rect 1465 -735 1485 -715
rect 1465 -785 1485 -765
rect 1765 -135 1785 -115
rect 1765 -185 1785 -165
rect 1765 -235 1785 -215
rect 1765 -285 1785 -265
rect 1765 -335 1785 -315
rect 1765 -385 1785 -365
rect 1765 -435 1785 -415
rect 1765 -485 1785 -465
rect 1765 -535 1785 -515
rect 1765 -585 1785 -565
rect 1765 -635 1785 -615
rect 1765 -685 1785 -665
rect 2065 -235 2085 -215
rect 2065 -285 2085 -265
rect 2065 -335 2085 -315
rect 2065 -385 2085 -365
rect 2065 -435 2085 -415
rect 2065 -485 2085 -465
rect 2065 -535 2085 -515
rect 2065 -585 2085 -565
rect 2065 -635 2085 -615
rect 2065 -685 2085 -665
rect 2065 -735 2085 -715
rect 2065 -785 2085 -765
rect 2365 -135 2385 -115
rect 2365 -185 2385 -165
rect 2365 -235 2385 -215
rect 2365 -285 2385 -265
rect 2365 -335 2385 -315
rect 2365 -385 2385 -365
rect 2365 -435 2385 -415
rect 2365 -485 2385 -465
rect 2365 -535 2385 -515
rect 2365 -585 2385 -565
rect 2365 -635 2385 -615
rect 2365 -685 2385 -665
rect 2665 -235 2685 -215
rect 2665 -285 2685 -265
rect 2665 -335 2685 -315
rect 2665 -385 2685 -365
rect 2665 -435 2685 -415
rect 2665 -485 2685 -465
rect 2665 -535 2685 -515
rect 2665 -585 2685 -565
rect 2665 -635 2685 -615
rect 2665 -685 2685 -665
rect 2665 -735 2685 -715
rect 2665 -785 2685 -765
rect 2965 -135 2985 -115
rect 2965 -185 2985 -165
rect 2965 -235 2985 -215
rect 2965 -285 2985 -265
rect 2965 -335 2985 -315
rect 2965 -385 2985 -365
rect 2965 -435 2985 -415
rect 2965 -485 2985 -465
rect 2965 -535 2985 -515
rect 2965 -585 2985 -565
rect 2965 -635 2985 -615
rect 2965 -685 2985 -665
rect 3265 -235 3285 -215
rect 3265 -285 3285 -265
rect 3265 -335 3285 -315
rect 3265 -385 3285 -365
rect 3265 -435 3285 -415
rect 3265 -485 3285 -465
rect 3265 -535 3285 -515
rect 3265 -585 3285 -565
rect 3265 -635 3285 -615
rect 3265 -685 3285 -665
rect 3265 -735 3285 -715
rect 3265 -785 3285 -765
rect 3565 -135 3585 -115
rect 3565 -185 3585 -165
rect 3565 -235 3585 -215
rect 3565 -285 3585 -265
rect 3565 -335 3585 -315
rect 3565 -385 3585 -365
rect 3565 -435 3585 -415
rect 3565 -485 3585 -465
rect 3565 -535 3585 -515
rect 3565 -585 3585 -565
rect 3565 -635 3585 -615
rect 3565 -685 3585 -665
rect 3565 -735 3585 -715
rect 3565 -785 3585 -765
rect 3715 -235 3735 -215
rect 3715 -285 3735 -265
rect 3715 -335 3735 -315
rect 3715 -385 3735 -365
rect 3715 -435 3735 -415
rect 3715 -485 3735 -465
rect 3715 -535 3735 -515
rect 3715 -585 3735 -565
rect 3715 -635 3735 -615
rect 3715 -685 3735 -665
rect 3715 -735 3735 -715
rect 3715 -785 3735 -765
rect 3865 -135 3885 -115
rect 3865 -185 3885 -165
rect 3865 -235 3885 -215
rect 3865 -285 3885 -265
rect 3865 -335 3885 -315
rect 3865 -385 3885 -365
rect 3865 -435 3885 -415
rect 3865 -485 3885 -465
rect 3865 -535 3885 -515
rect 3865 -585 3885 -565
rect 3865 -635 3885 -615
rect 3865 -685 3885 -665
rect 4015 -235 4035 -215
rect 4015 -285 4035 -265
rect 4015 -335 4035 -315
rect 4015 -385 4035 -365
rect 4015 -435 4035 -415
rect 4015 -485 4035 -465
rect 4015 -535 4035 -515
rect 4015 -585 4035 -565
rect 4015 -635 4035 -615
rect 4015 -685 4035 -665
rect 4015 -735 4035 -715
rect 4015 -785 4035 -765
rect 4165 -135 4185 -115
rect 4165 -185 4185 -165
rect 4165 -235 4185 -215
rect 4165 -285 4185 -265
rect 4165 -335 4185 -315
rect 4165 -385 4185 -365
rect 4165 -435 4185 -415
rect 4165 -485 4185 -465
rect 4165 -535 4185 -515
rect 4165 -585 4185 -565
rect 4165 -635 4185 -615
rect 4165 -685 4185 -665
rect 4165 -735 4185 -715
rect 4165 -785 4185 -765
rect 4315 -235 4335 -215
rect 4315 -285 4335 -265
rect 4315 -335 4335 -315
rect 4315 -385 4335 -365
rect 4315 -435 4335 -415
rect 4315 -485 4335 -465
rect 4315 -535 4335 -515
rect 4315 -585 4335 -565
rect 4315 -635 4335 -615
rect 4315 -685 4335 -665
rect 4315 -735 4335 -715
rect 4315 -785 4335 -765
rect 4465 -135 4485 -115
rect 4465 -185 4485 -165
rect 4465 -235 4485 -215
rect 4465 -285 4485 -265
rect 4465 -335 4485 -315
rect 4465 -385 4485 -365
rect 4465 -435 4485 -415
rect 4465 -485 4485 -465
rect 4465 -535 4485 -515
rect 4465 -585 4485 -565
rect 4465 -635 4485 -615
rect 4465 -685 4485 -665
rect 4615 -235 4635 -215
rect 4615 -285 4635 -265
rect 4615 -335 4635 -315
rect 4615 -385 4635 -365
rect 4615 -435 4635 -415
rect 4615 -485 4635 -465
rect 4615 -535 4635 -515
rect 4615 -585 4635 -565
rect 4615 -635 4635 -615
rect 4615 -685 4635 -665
rect 4615 -735 4635 -715
rect 4615 -785 4635 -765
rect 4765 -135 4785 -115
rect 4765 -185 4785 -165
rect 4765 -235 4785 -215
rect 4765 -285 4785 -265
rect 4765 -335 4785 -315
rect 4765 -385 4785 -365
rect 4765 -435 4785 -415
rect 4765 -485 4785 -465
rect 4765 -535 4785 -515
rect 4765 -585 4785 -565
rect 4765 -635 4785 -615
rect 4765 -685 4785 -665
rect 4765 -735 4785 -715
rect 4765 -785 4785 -765
rect 5065 -235 5085 -215
rect 5065 -285 5085 -265
rect 5065 -335 5085 -315
rect 5065 -385 5085 -365
rect 5065 -435 5085 -415
rect 5065 -485 5085 -465
rect 5065 -535 5085 -515
rect 5065 -585 5085 -565
rect 5065 -635 5085 -615
rect 5065 -685 5085 -665
rect 5065 -735 5085 -715
rect 5065 -785 5085 -765
rect 5365 -135 5385 -115
rect 5365 -185 5385 -165
rect 5365 -235 5385 -215
rect 5365 -285 5385 -265
rect 5365 -335 5385 -315
rect 5365 -385 5385 -365
rect 5365 -435 5385 -415
rect 5365 -485 5385 -465
rect 5365 -535 5385 -515
rect 5365 -585 5385 -565
rect 5365 -635 5385 -615
rect 5365 -685 5385 -665
rect 5665 -235 5685 -215
rect 5665 -285 5685 -265
rect 5665 -335 5685 -315
rect 5665 -385 5685 -365
rect 5665 -435 5685 -415
rect 5665 -485 5685 -465
rect 5665 -535 5685 -515
rect 5665 -585 5685 -565
rect 5665 -635 5685 -615
rect 5665 -685 5685 -665
rect 5665 -735 5685 -715
rect 5665 -785 5685 -765
rect 5965 -135 5985 -115
rect 5965 -185 5985 -165
rect 5965 -235 5985 -215
rect 5965 -285 5985 -265
rect 5965 -335 5985 -315
rect 5965 -385 5985 -365
rect 5965 -435 5985 -415
rect 5965 -485 5985 -465
rect 5965 -535 5985 -515
rect 5965 -585 5985 -565
rect 5965 -635 5985 -615
rect 5965 -685 5985 -665
rect 6265 -235 6285 -215
rect 6265 -285 6285 -265
rect 6265 -335 6285 -315
rect 6265 -385 6285 -365
rect 6265 -435 6285 -415
rect 6265 -485 6285 -465
rect 6265 -535 6285 -515
rect 6265 -585 6285 -565
rect 6265 -635 6285 -615
rect 6265 -685 6285 -665
rect 6265 -735 6285 -715
rect 6265 -785 6285 -765
rect 6565 -135 6585 -115
rect 6565 -185 6585 -165
rect 6565 -235 6585 -215
rect 6565 -285 6585 -265
rect 6565 -335 6585 -315
rect 6565 -385 6585 -365
rect 6565 -435 6585 -415
rect 6565 -485 6585 -465
rect 6565 -535 6585 -515
rect 6565 -585 6585 -565
rect 6565 -635 6585 -615
rect 6565 -685 6585 -665
rect 6865 -235 6885 -215
rect 6865 -285 6885 -265
rect 6865 -335 6885 -315
rect 6865 -385 6885 -365
rect 6865 -435 6885 -415
rect 6865 -485 6885 -465
rect 6865 -535 6885 -515
rect 6865 -585 6885 -565
rect 6865 -635 6885 -615
rect 6865 -685 6885 -665
rect 6865 -735 6885 -715
rect 6865 -785 6885 -765
rect 7165 -135 7185 -115
rect 7165 -185 7185 -165
rect 7165 -235 7185 -215
rect 7165 -285 7185 -265
rect 7165 -335 7185 -315
rect 7165 -385 7185 -365
rect 7165 -435 7185 -415
rect 7165 -485 7185 -465
rect 7165 -535 7185 -515
rect 7165 -585 7185 -565
rect 7165 -635 7185 -615
rect 7165 -685 7185 -665
rect 7165 -735 7185 -715
rect 7165 -785 7185 -765
rect 8365 -135 8385 -115
rect 8365 -185 8385 -165
rect 8365 -235 8385 -215
rect 8365 -285 8385 -265
rect 8365 -335 8385 -315
rect 8365 -385 8385 -365
rect 8365 -435 8385 -415
rect 8365 -485 8385 -465
rect 8365 -535 8385 -515
rect 8365 -585 8385 -565
rect 8365 -635 8385 -615
rect 8365 -685 8385 -665
rect 8365 -735 8385 -715
rect 8365 -785 8385 -765
rect 9565 -135 9585 -115
rect 9565 -185 9585 -165
rect 9565 -235 9585 -215
rect 9565 -285 9585 -265
rect 9565 -335 9585 -315
rect 9565 -385 9585 -365
rect 9565 -435 9585 -415
rect 9565 -485 9585 -465
rect 9565 -535 9585 -515
rect 9565 -585 9585 -565
rect 9565 -635 9585 -615
rect 9565 -685 9585 -665
rect 9565 -735 9585 -715
rect 9565 -785 9585 -765
rect 10765 -135 10785 -115
rect 10765 -185 10785 -165
rect 10765 -235 10785 -215
rect 10765 -285 10785 -265
rect 10765 -335 10785 -315
rect 10765 -385 10785 -365
rect 10765 -435 10785 -415
rect 10765 -485 10785 -465
rect 10765 -535 10785 -515
rect 10765 -585 10785 -565
rect 10765 -635 10785 -615
rect 10765 -685 10785 -665
rect 10765 -735 10785 -715
rect 10765 -785 10785 -765
rect 11965 -135 11985 -115
rect 11965 -185 11985 -165
rect 11965 -235 11985 -215
rect 11965 -285 11985 -265
rect 11965 -335 11985 -315
rect 11965 -385 11985 -365
rect 11965 -435 11985 -415
rect 11965 -485 11985 -465
rect 11965 -535 11985 -515
rect 11965 -585 11985 -565
rect 11965 -635 11985 -615
rect 11965 -685 11985 -665
rect 11965 -735 11985 -715
rect 11965 -785 11985 -765
rect 12265 -235 12285 -215
rect 12265 -285 12285 -265
rect 12265 -335 12285 -315
rect 12265 -385 12285 -365
rect 12265 -435 12285 -415
rect 12265 -485 12285 -465
rect 12265 -535 12285 -515
rect 12265 -585 12285 -565
rect 12265 -635 12285 -615
rect 12265 -685 12285 -665
rect 12265 -735 12285 -715
rect 12265 -785 12285 -765
rect 12565 -135 12585 -115
rect 12565 -185 12585 -165
rect 12565 -235 12585 -215
rect 12565 -285 12585 -265
rect 12565 -335 12585 -315
rect 12565 -385 12585 -365
rect 12565 -435 12585 -415
rect 12565 -485 12585 -465
rect 12565 -535 12585 -515
rect 12565 -585 12585 -565
rect 12565 -635 12585 -615
rect 12565 -685 12585 -665
rect 12865 -235 12885 -215
rect 12865 -285 12885 -265
rect 12865 -335 12885 -315
rect 12865 -385 12885 -365
rect 12865 -435 12885 -415
rect 12865 -485 12885 -465
rect 12865 -535 12885 -515
rect 12865 -585 12885 -565
rect 12865 -635 12885 -615
rect 12865 -685 12885 -665
rect 12865 -735 12885 -715
rect 12865 -785 12885 -765
rect 13165 -135 13185 -115
rect 13165 -185 13185 -165
rect 13165 -235 13185 -215
rect 13165 -285 13185 -265
rect 13165 -335 13185 -315
rect 13165 -385 13185 -365
rect 13165 -435 13185 -415
rect 13165 -485 13185 -465
rect 13165 -535 13185 -515
rect 13165 -585 13185 -565
rect 13165 -635 13185 -615
rect 13165 -685 13185 -665
rect 13465 -235 13485 -215
rect 13465 -285 13485 -265
rect 13465 -335 13485 -315
rect 13465 -385 13485 -365
rect 13465 -435 13485 -415
rect 13465 -485 13485 -465
rect 13465 -535 13485 -515
rect 13465 -585 13485 -565
rect 13465 -635 13485 -615
rect 13465 -685 13485 -665
rect 13465 -735 13485 -715
rect 13465 -785 13485 -765
rect 13765 -135 13785 -115
rect 13765 -185 13785 -165
rect 13765 -235 13785 -215
rect 13765 -285 13785 -265
rect 13765 -335 13785 -315
rect 13765 -385 13785 -365
rect 13765 -435 13785 -415
rect 13765 -485 13785 -465
rect 13765 -535 13785 -515
rect 13765 -585 13785 -565
rect 13765 -635 13785 -615
rect 13765 -685 13785 -665
rect 14065 -235 14085 -215
rect 14065 -285 14085 -265
rect 14065 -335 14085 -315
rect 14065 -385 14085 -365
rect 14065 -435 14085 -415
rect 14065 -485 14085 -465
rect 14065 -535 14085 -515
rect 14065 -585 14085 -565
rect 14065 -635 14085 -615
rect 14065 -685 14085 -665
rect 14065 -735 14085 -715
rect 14065 -785 14085 -765
rect 14365 -135 14385 -115
rect 14365 -185 14385 -165
rect 14365 -235 14385 -215
rect 14365 -285 14385 -265
rect 14365 -335 14385 -315
rect 14365 -385 14385 -365
rect 14365 -435 14385 -415
rect 14365 -485 14385 -465
rect 14365 -535 14385 -515
rect 14365 -585 14385 -565
rect 14365 -635 14385 -615
rect 14365 -685 14385 -665
rect 14365 -735 14385 -715
rect 14365 -785 14385 -765
rect 15565 -135 15585 -115
rect 15565 -185 15585 -165
rect 15565 -235 15585 -215
rect 15565 -285 15585 -265
rect 15565 -335 15585 -315
rect 15565 -385 15585 -365
rect 15565 -435 15585 -415
rect 15565 -485 15585 -465
rect 15565 -535 15585 -515
rect 15565 -585 15585 -565
rect 15565 -635 15585 -615
rect 15565 -685 15585 -665
rect 15565 -735 15585 -715
rect 15565 -785 15585 -765
rect 16765 -135 16785 -115
rect 16765 -185 16785 -165
rect 16765 -235 16785 -215
rect 16765 -285 16785 -265
rect 16765 -335 16785 -315
rect 16765 -385 16785 -365
rect 16765 -435 16785 -415
rect 16765 -485 16785 -465
rect 16765 -535 16785 -515
rect 16765 -585 16785 -565
rect 16765 -635 16785 -615
rect 16765 -685 16785 -665
rect 16765 -735 16785 -715
rect 16765 -785 16785 -765
rect 17965 -135 17985 -115
rect 17965 -185 17985 -165
rect 17965 -235 17985 -215
rect 17965 -285 17985 -265
rect 17965 -335 17985 -315
rect 17965 -385 17985 -365
rect 17965 -435 17985 -415
rect 17965 -485 17985 -465
rect 17965 -535 17985 -515
rect 17965 -585 17985 -565
rect 17965 -635 17985 -615
rect 17965 -685 17985 -665
rect 17965 -735 17985 -715
rect 17965 -785 17985 -765
rect 19165 -135 19185 -115
rect 19165 -185 19185 -165
rect 19165 -235 19185 -215
rect 19165 -285 19185 -265
rect 19165 -335 19185 -315
rect 19165 -385 19185 -365
rect 19165 -435 19185 -415
rect 19165 -485 19185 -465
rect 19165 -535 19185 -515
rect 19165 -585 19185 -565
rect 19165 -635 19185 -615
rect 19165 -685 19185 -665
rect 19165 -735 19185 -715
rect 19165 -785 19185 -765
rect 20365 -135 20385 -115
rect 20365 -185 20385 -165
rect 20365 -235 20385 -215
rect 20365 -285 20385 -265
rect 20365 -335 20385 -315
rect 20365 -385 20385 -365
rect 20365 -435 20385 -415
rect 20365 -485 20385 -465
rect 20365 -535 20385 -515
rect 20365 -585 20385 -565
rect 20365 -635 20385 -615
rect 20365 -685 20385 -665
rect 20365 -735 20385 -715
rect 20365 -785 20385 -765
rect -485 -885 -465 -865
rect -185 -885 -165 -865
rect 115 -885 135 -865
rect 415 -885 435 -865
rect 715 -885 735 -865
rect 1015 -885 1035 -865
rect 1315 -885 1335 -865
rect 1615 -885 1635 -865
rect 1915 -885 1935 -865
rect 2215 -885 2235 -865
rect 2515 -885 2535 -865
rect 2815 -885 2835 -865
rect 3115 -885 3135 -865
rect 3415 -885 3435 -865
rect 3715 -885 3735 -865
rect 4015 -885 4035 -865
rect 4315 -885 4335 -865
rect 4615 -885 4635 -865
rect 4915 -885 4935 -865
rect 5215 -885 5235 -865
rect 5515 -885 5535 -865
rect 5815 -885 5835 -865
rect 6115 -885 6135 -865
rect 6415 -885 6435 -865
rect 6715 -885 6735 -865
rect 7015 -885 7035 -865
rect 7315 -885 7335 -865
rect 7615 -885 7635 -865
rect 7915 -885 7935 -865
rect 8215 -885 8235 -865
rect 8515 -885 8535 -865
rect 8815 -885 8835 -865
rect 9115 -885 9135 -865
rect 9415 -885 9435 -865
rect 9715 -885 9735 -865
rect 10015 -885 10035 -865
rect 10315 -885 10335 -865
rect 10615 -885 10635 -865
rect 10915 -885 10935 -865
rect 11215 -885 11235 -865
rect 11515 -885 11535 -865
rect 11815 -885 11835 -865
rect 12115 -885 12135 -865
rect 12415 -885 12435 -865
rect 12715 -885 12735 -865
rect 13015 -885 13035 -865
rect 13315 -885 13335 -865
rect 13615 -885 13635 -865
rect 13915 -885 13935 -865
rect 14215 -885 14235 -865
rect 14515 -885 14535 -865
rect 14815 -885 14835 -865
rect 15115 -885 15135 -865
rect 15415 -885 15435 -865
rect 15715 -885 15735 -865
rect 16015 -885 16035 -865
rect 16315 -885 16335 -865
rect 16615 -885 16635 -865
rect 16915 -885 16935 -865
rect 17215 -885 17235 -865
rect 17515 -885 17535 -865
rect 17815 -885 17835 -865
rect 18115 -885 18135 -865
rect 18415 -885 18435 -865
rect 18715 -885 18735 -865
rect 19015 -885 19035 -865
rect 19315 -885 19335 -865
rect 19615 -885 19635 -865
rect 19915 -885 19935 -865
rect 20215 -885 20235 -865
rect -635 -985 -615 -965
rect -635 -1035 -615 -1015
rect -635 -1085 -615 -1065
rect -635 -1135 -615 -1115
rect -635 -1185 -615 -1165
rect -635 -1235 -615 -1215
rect -635 -1285 -615 -1265
rect -635 -1335 -615 -1315
rect -635 -1385 -615 -1365
rect -635 -1435 -615 -1415
rect -635 -1485 -615 -1465
rect -635 -1535 -615 -1515
rect -635 -1585 -615 -1565
rect -635 -1635 -615 -1615
rect -485 -985 -465 -965
rect -485 -1035 -465 -1015
rect -485 -1085 -465 -1065
rect -485 -1135 -465 -1115
rect -485 -1185 -465 -1165
rect -485 -1235 -465 -1215
rect -485 -1285 -465 -1265
rect -485 -1335 -465 -1315
rect -485 -1385 -465 -1365
rect -485 -1435 -465 -1415
rect -485 -1485 -465 -1465
rect -485 -1535 -465 -1515
rect -485 -1585 -465 -1565
rect -485 -1635 -465 -1615
rect -335 -985 -315 -965
rect -335 -1035 -315 -1015
rect -335 -1085 -315 -1065
rect -335 -1135 -315 -1115
rect -335 -1185 -315 -1165
rect -335 -1235 -315 -1215
rect -335 -1285 -315 -1265
rect -335 -1335 -315 -1315
rect -335 -1385 -315 -1365
rect -335 -1435 -315 -1415
rect -335 -1485 -315 -1465
rect -335 -1535 -315 -1515
rect -335 -1585 -315 -1565
rect -335 -1635 -315 -1615
rect -185 -985 -165 -965
rect -185 -1035 -165 -1015
rect -185 -1085 -165 -1065
rect -185 -1135 -165 -1115
rect -185 -1185 -165 -1165
rect -185 -1235 -165 -1215
rect -185 -1285 -165 -1265
rect -185 -1335 -165 -1315
rect -185 -1385 -165 -1365
rect -185 -1435 -165 -1415
rect -185 -1485 -165 -1465
rect -185 -1535 -165 -1515
rect -185 -1585 -165 -1565
rect -185 -1635 -165 -1615
rect -35 -985 -15 -965
rect -35 -1035 -15 -1015
rect -35 -1085 -15 -1065
rect -35 -1135 -15 -1115
rect -35 -1185 -15 -1165
rect -35 -1235 -15 -1215
rect -35 -1285 -15 -1265
rect -35 -1335 -15 -1315
rect -35 -1385 -15 -1365
rect -35 -1435 -15 -1415
rect -35 -1485 -15 -1465
rect -35 -1535 -15 -1515
rect -35 -1585 -15 -1565
rect -35 -1635 -15 -1615
rect 1165 -985 1185 -965
rect 1165 -1035 1185 -1015
rect 1165 -1085 1185 -1065
rect 1165 -1135 1185 -1115
rect 1165 -1185 1185 -1165
rect 1165 -1235 1185 -1215
rect 1165 -1285 1185 -1265
rect 1165 -1335 1185 -1315
rect 1165 -1385 1185 -1365
rect 1165 -1435 1185 -1415
rect 1165 -1485 1185 -1465
rect 1165 -1535 1185 -1515
rect 1165 -1585 1185 -1565
rect 1165 -1635 1185 -1615
rect 1465 -985 1485 -965
rect 1465 -1035 1485 -1015
rect 1465 -1085 1485 -1065
rect 1465 -1135 1485 -1115
rect 1465 -1185 1485 -1165
rect 1465 -1235 1485 -1215
rect 1465 -1285 1485 -1265
rect 1465 -1335 1485 -1315
rect 1465 -1385 1485 -1365
rect 1465 -1435 1485 -1415
rect 1465 -1485 1485 -1465
rect 1465 -1535 1485 -1515
rect 1765 -1085 1785 -1065
rect 1765 -1135 1785 -1115
rect 1765 -1185 1785 -1165
rect 1765 -1235 1785 -1215
rect 1765 -1285 1785 -1265
rect 1765 -1335 1785 -1315
rect 1765 -1385 1785 -1365
rect 1765 -1435 1785 -1415
rect 1765 -1485 1785 -1465
rect 1765 -1535 1785 -1515
rect 1765 -1585 1785 -1565
rect 1765 -1635 1785 -1615
rect 2065 -985 2085 -965
rect 2065 -1035 2085 -1015
rect 2065 -1085 2085 -1065
rect 2065 -1135 2085 -1115
rect 2065 -1185 2085 -1165
rect 2065 -1235 2085 -1215
rect 2065 -1285 2085 -1265
rect 2065 -1335 2085 -1315
rect 2065 -1385 2085 -1365
rect 2065 -1435 2085 -1415
rect 2065 -1485 2085 -1465
rect 2065 -1535 2085 -1515
rect 2365 -1085 2385 -1065
rect 2365 -1135 2385 -1115
rect 2365 -1185 2385 -1165
rect 2365 -1235 2385 -1215
rect 2365 -1285 2385 -1265
rect 2365 -1335 2385 -1315
rect 2365 -1385 2385 -1365
rect 2365 -1435 2385 -1415
rect 2365 -1485 2385 -1465
rect 2365 -1535 2385 -1515
rect 2365 -1585 2385 -1565
rect 2365 -1635 2385 -1615
rect 2665 -985 2685 -965
rect 2665 -1035 2685 -1015
rect 2665 -1085 2685 -1065
rect 2665 -1135 2685 -1115
rect 2665 -1185 2685 -1165
rect 2665 -1235 2685 -1215
rect 2665 -1285 2685 -1265
rect 2665 -1335 2685 -1315
rect 2665 -1385 2685 -1365
rect 2665 -1435 2685 -1415
rect 2665 -1485 2685 -1465
rect 2665 -1535 2685 -1515
rect 2965 -1085 2985 -1065
rect 2965 -1135 2985 -1115
rect 2965 -1185 2985 -1165
rect 2965 -1235 2985 -1215
rect 2965 -1285 2985 -1265
rect 2965 -1335 2985 -1315
rect 2965 -1385 2985 -1365
rect 2965 -1435 2985 -1415
rect 2965 -1485 2985 -1465
rect 2965 -1535 2985 -1515
rect 2965 -1585 2985 -1565
rect 2965 -1635 2985 -1615
rect 3265 -985 3285 -965
rect 3265 -1035 3285 -1015
rect 3265 -1085 3285 -1065
rect 3265 -1135 3285 -1115
rect 3265 -1185 3285 -1165
rect 3265 -1235 3285 -1215
rect 3265 -1285 3285 -1265
rect 3265 -1335 3285 -1315
rect 3265 -1385 3285 -1365
rect 3265 -1435 3285 -1415
rect 3265 -1485 3285 -1465
rect 3265 -1535 3285 -1515
rect 3565 -985 3585 -965
rect 3565 -1035 3585 -1015
rect 3565 -1085 3585 -1065
rect 3565 -1135 3585 -1115
rect 3565 -1185 3585 -1165
rect 3565 -1235 3585 -1215
rect 3565 -1285 3585 -1265
rect 3565 -1335 3585 -1315
rect 3565 -1385 3585 -1365
rect 3565 -1435 3585 -1415
rect 3565 -1485 3585 -1465
rect 3565 -1535 3585 -1515
rect 3565 -1585 3585 -1565
rect 3565 -1635 3585 -1615
rect 3715 -985 3735 -965
rect 3715 -1035 3735 -1015
rect 3715 -1085 3735 -1065
rect 3715 -1135 3735 -1115
rect 3715 -1185 3735 -1165
rect 3715 -1235 3735 -1215
rect 3715 -1285 3735 -1265
rect 3715 -1335 3735 -1315
rect 3715 -1385 3735 -1365
rect 3715 -1435 3735 -1415
rect 3715 -1485 3735 -1465
rect 3715 -1535 3735 -1515
rect 3865 -1085 3885 -1065
rect 3865 -1135 3885 -1115
rect 3865 -1185 3885 -1165
rect 3865 -1235 3885 -1215
rect 3865 -1285 3885 -1265
rect 3865 -1335 3885 -1315
rect 3865 -1385 3885 -1365
rect 3865 -1435 3885 -1415
rect 3865 -1485 3885 -1465
rect 3865 -1535 3885 -1515
rect 3865 -1585 3885 -1565
rect 3865 -1635 3885 -1615
rect 4015 -985 4035 -965
rect 4015 -1035 4035 -1015
rect 4015 -1085 4035 -1065
rect 4015 -1135 4035 -1115
rect 4015 -1185 4035 -1165
rect 4015 -1235 4035 -1215
rect 4015 -1285 4035 -1265
rect 4015 -1335 4035 -1315
rect 4015 -1385 4035 -1365
rect 4015 -1435 4035 -1415
rect 4015 -1485 4035 -1465
rect 4015 -1535 4035 -1515
rect 4165 -985 4185 -965
rect 4165 -1035 4185 -1015
rect 4165 -1085 4185 -1065
rect 4165 -1135 4185 -1115
rect 4165 -1185 4185 -1165
rect 4165 -1235 4185 -1215
rect 4165 -1285 4185 -1265
rect 4165 -1335 4185 -1315
rect 4165 -1385 4185 -1365
rect 4165 -1435 4185 -1415
rect 4165 -1485 4185 -1465
rect 4165 -1535 4185 -1515
rect 4165 -1585 4185 -1565
rect 4165 -1635 4185 -1615
rect 4315 -985 4335 -965
rect 4315 -1035 4335 -1015
rect 4315 -1085 4335 -1065
rect 4315 -1135 4335 -1115
rect 4315 -1185 4335 -1165
rect 4315 -1235 4335 -1215
rect 4315 -1285 4335 -1265
rect 4315 -1335 4335 -1315
rect 4315 -1385 4335 -1365
rect 4315 -1435 4335 -1415
rect 4315 -1485 4335 -1465
rect 4315 -1535 4335 -1515
rect 4465 -1085 4485 -1065
rect 4465 -1135 4485 -1115
rect 4465 -1185 4485 -1165
rect 4465 -1235 4485 -1215
rect 4465 -1285 4485 -1265
rect 4465 -1335 4485 -1315
rect 4465 -1385 4485 -1365
rect 4465 -1435 4485 -1415
rect 4465 -1485 4485 -1465
rect 4465 -1535 4485 -1515
rect 4465 -1585 4485 -1565
rect 4465 -1635 4485 -1615
rect 4615 -985 4635 -965
rect 4615 -1035 4635 -1015
rect 4615 -1085 4635 -1065
rect 4615 -1135 4635 -1115
rect 4615 -1185 4635 -1165
rect 4615 -1235 4635 -1215
rect 4615 -1285 4635 -1265
rect 4615 -1335 4635 -1315
rect 4615 -1385 4635 -1365
rect 4615 -1435 4635 -1415
rect 4615 -1485 4635 -1465
rect 4615 -1535 4635 -1515
rect 4765 -985 4785 -965
rect 4765 -1035 4785 -1015
rect 4765 -1085 4785 -1065
rect 4765 -1135 4785 -1115
rect 4765 -1185 4785 -1165
rect 4765 -1235 4785 -1215
rect 4765 -1285 4785 -1265
rect 4765 -1335 4785 -1315
rect 4765 -1385 4785 -1365
rect 4765 -1435 4785 -1415
rect 4765 -1485 4785 -1465
rect 4765 -1535 4785 -1515
rect 4765 -1585 4785 -1565
rect 4765 -1635 4785 -1615
rect 5065 -985 5085 -965
rect 5065 -1035 5085 -1015
rect 5065 -1085 5085 -1065
rect 5065 -1135 5085 -1115
rect 5065 -1185 5085 -1165
rect 5065 -1235 5085 -1215
rect 5065 -1285 5085 -1265
rect 5065 -1335 5085 -1315
rect 5065 -1385 5085 -1365
rect 5065 -1435 5085 -1415
rect 5065 -1485 5085 -1465
rect 5065 -1535 5085 -1515
rect 5365 -1085 5385 -1065
rect 5365 -1135 5385 -1115
rect 5365 -1185 5385 -1165
rect 5365 -1235 5385 -1215
rect 5365 -1285 5385 -1265
rect 5365 -1335 5385 -1315
rect 5365 -1385 5385 -1365
rect 5365 -1435 5385 -1415
rect 5365 -1485 5385 -1465
rect 5365 -1535 5385 -1515
rect 5365 -1585 5385 -1565
rect 5365 -1635 5385 -1615
rect 5665 -985 5685 -965
rect 5665 -1035 5685 -1015
rect 5665 -1085 5685 -1065
rect 5665 -1135 5685 -1115
rect 5665 -1185 5685 -1165
rect 5665 -1235 5685 -1215
rect 5665 -1285 5685 -1265
rect 5665 -1335 5685 -1315
rect 5665 -1385 5685 -1365
rect 5665 -1435 5685 -1415
rect 5665 -1485 5685 -1465
rect 5665 -1535 5685 -1515
rect 5965 -1085 5985 -1065
rect 5965 -1135 5985 -1115
rect 5965 -1185 5985 -1165
rect 5965 -1235 5985 -1215
rect 5965 -1285 5985 -1265
rect 5965 -1335 5985 -1315
rect 5965 -1385 5985 -1365
rect 5965 -1435 5985 -1415
rect 5965 -1485 5985 -1465
rect 5965 -1535 5985 -1515
rect 5965 -1585 5985 -1565
rect 5965 -1635 5985 -1615
rect 6265 -985 6285 -965
rect 6265 -1035 6285 -1015
rect 6265 -1085 6285 -1065
rect 6265 -1135 6285 -1115
rect 6265 -1185 6285 -1165
rect 6265 -1235 6285 -1215
rect 6265 -1285 6285 -1265
rect 6265 -1335 6285 -1315
rect 6265 -1385 6285 -1365
rect 6265 -1435 6285 -1415
rect 6265 -1485 6285 -1465
rect 6265 -1535 6285 -1515
rect 6565 -1085 6585 -1065
rect 6565 -1135 6585 -1115
rect 6565 -1185 6585 -1165
rect 6565 -1235 6585 -1215
rect 6565 -1285 6585 -1265
rect 6565 -1335 6585 -1315
rect 6565 -1385 6585 -1365
rect 6565 -1435 6585 -1415
rect 6565 -1485 6585 -1465
rect 6565 -1535 6585 -1515
rect 6565 -1585 6585 -1565
rect 6565 -1635 6585 -1615
rect 6865 -985 6885 -965
rect 6865 -1035 6885 -1015
rect 6865 -1085 6885 -1065
rect 6865 -1135 6885 -1115
rect 6865 -1185 6885 -1165
rect 6865 -1235 6885 -1215
rect 6865 -1285 6885 -1265
rect 6865 -1335 6885 -1315
rect 6865 -1385 6885 -1365
rect 6865 -1435 6885 -1415
rect 6865 -1485 6885 -1465
rect 6865 -1535 6885 -1515
rect 7165 -985 7185 -965
rect 7165 -1035 7185 -1015
rect 7165 -1085 7185 -1065
rect 7165 -1135 7185 -1115
rect 7165 -1185 7185 -1165
rect 7165 -1235 7185 -1215
rect 7165 -1285 7185 -1265
rect 7165 -1335 7185 -1315
rect 7165 -1385 7185 -1365
rect 7165 -1435 7185 -1415
rect 7165 -1485 7185 -1465
rect 7165 -1535 7185 -1515
rect 7165 -1585 7185 -1565
rect 7165 -1635 7185 -1615
rect 8365 -985 8385 -965
rect 8365 -1035 8385 -1015
rect 8365 -1085 8385 -1065
rect 8365 -1135 8385 -1115
rect 8365 -1185 8385 -1165
rect 8365 -1235 8385 -1215
rect 8365 -1285 8385 -1265
rect 8365 -1335 8385 -1315
rect 8365 -1385 8385 -1365
rect 8365 -1435 8385 -1415
rect 8365 -1485 8385 -1465
rect 8365 -1535 8385 -1515
rect 8365 -1585 8385 -1565
rect 8365 -1635 8385 -1615
rect 9565 -985 9585 -965
rect 9565 -1035 9585 -1015
rect 9565 -1085 9585 -1065
rect 9565 -1135 9585 -1115
rect 9565 -1185 9585 -1165
rect 9565 -1235 9585 -1215
rect 9565 -1285 9585 -1265
rect 9565 -1335 9585 -1315
rect 9565 -1385 9585 -1365
rect 9565 -1435 9585 -1415
rect 9565 -1485 9585 -1465
rect 9565 -1535 9585 -1515
rect 9565 -1585 9585 -1565
rect 9565 -1635 9585 -1615
rect 10765 -985 10785 -965
rect 10765 -1035 10785 -1015
rect 10765 -1085 10785 -1065
rect 10765 -1135 10785 -1115
rect 10765 -1185 10785 -1165
rect 10765 -1235 10785 -1215
rect 10765 -1285 10785 -1265
rect 10765 -1335 10785 -1315
rect 10765 -1385 10785 -1365
rect 10765 -1435 10785 -1415
rect 10765 -1485 10785 -1465
rect 10765 -1535 10785 -1515
rect 10765 -1585 10785 -1565
rect 10765 -1635 10785 -1615
rect 11965 -985 11985 -965
rect 11965 -1035 11985 -1015
rect 11965 -1085 11985 -1065
rect 11965 -1135 11985 -1115
rect 11965 -1185 11985 -1165
rect 11965 -1235 11985 -1215
rect 11965 -1285 11985 -1265
rect 11965 -1335 11985 -1315
rect 11965 -1385 11985 -1365
rect 11965 -1435 11985 -1415
rect 11965 -1485 11985 -1465
rect 11965 -1535 11985 -1515
rect 11965 -1585 11985 -1565
rect 11965 -1635 11985 -1615
rect 12265 -985 12285 -965
rect 12265 -1035 12285 -1015
rect 12265 -1085 12285 -1065
rect 12265 -1135 12285 -1115
rect 12265 -1185 12285 -1165
rect 12265 -1235 12285 -1215
rect 12265 -1285 12285 -1265
rect 12265 -1335 12285 -1315
rect 12265 -1385 12285 -1365
rect 12265 -1435 12285 -1415
rect 12265 -1485 12285 -1465
rect 12265 -1535 12285 -1515
rect 12565 -1085 12585 -1065
rect 12565 -1135 12585 -1115
rect 12565 -1185 12585 -1165
rect 12565 -1235 12585 -1215
rect 12565 -1285 12585 -1265
rect 12565 -1335 12585 -1315
rect 12565 -1385 12585 -1365
rect 12565 -1435 12585 -1415
rect 12565 -1485 12585 -1465
rect 12565 -1535 12585 -1515
rect 12565 -1585 12585 -1565
rect 12565 -1635 12585 -1615
rect 12865 -985 12885 -965
rect 12865 -1035 12885 -1015
rect 12865 -1085 12885 -1065
rect 12865 -1135 12885 -1115
rect 12865 -1185 12885 -1165
rect 12865 -1235 12885 -1215
rect 12865 -1285 12885 -1265
rect 12865 -1335 12885 -1315
rect 12865 -1385 12885 -1365
rect 12865 -1435 12885 -1415
rect 12865 -1485 12885 -1465
rect 12865 -1535 12885 -1515
rect 13165 -1085 13185 -1065
rect 13165 -1135 13185 -1115
rect 13165 -1185 13185 -1165
rect 13165 -1235 13185 -1215
rect 13165 -1285 13185 -1265
rect 13165 -1335 13185 -1315
rect 13165 -1385 13185 -1365
rect 13165 -1435 13185 -1415
rect 13165 -1485 13185 -1465
rect 13165 -1535 13185 -1515
rect 13165 -1585 13185 -1565
rect 13165 -1635 13185 -1615
rect 13465 -985 13485 -965
rect 13465 -1035 13485 -1015
rect 13465 -1085 13485 -1065
rect 13465 -1135 13485 -1115
rect 13465 -1185 13485 -1165
rect 13465 -1235 13485 -1215
rect 13465 -1285 13485 -1265
rect 13465 -1335 13485 -1315
rect 13465 -1385 13485 -1365
rect 13465 -1435 13485 -1415
rect 13465 -1485 13485 -1465
rect 13465 -1535 13485 -1515
rect 13765 -1085 13785 -1065
rect 13765 -1135 13785 -1115
rect 13765 -1185 13785 -1165
rect 13765 -1235 13785 -1215
rect 13765 -1285 13785 -1265
rect 13765 -1335 13785 -1315
rect 13765 -1385 13785 -1365
rect 13765 -1435 13785 -1415
rect 13765 -1485 13785 -1465
rect 13765 -1535 13785 -1515
rect 13765 -1585 13785 -1565
rect 13765 -1635 13785 -1615
rect 14065 -985 14085 -965
rect 14065 -1035 14085 -1015
rect 14065 -1085 14085 -1065
rect 14065 -1135 14085 -1115
rect 14065 -1185 14085 -1165
rect 14065 -1235 14085 -1215
rect 14065 -1285 14085 -1265
rect 14065 -1335 14085 -1315
rect 14065 -1385 14085 -1365
rect 14065 -1435 14085 -1415
rect 14065 -1485 14085 -1465
rect 14065 -1535 14085 -1515
rect 14365 -985 14385 -965
rect 14365 -1035 14385 -1015
rect 14365 -1085 14385 -1065
rect 14365 -1135 14385 -1115
rect 14365 -1185 14385 -1165
rect 14365 -1235 14385 -1215
rect 14365 -1285 14385 -1265
rect 14365 -1335 14385 -1315
rect 14365 -1385 14385 -1365
rect 14365 -1435 14385 -1415
rect 14365 -1485 14385 -1465
rect 14365 -1535 14385 -1515
rect 14365 -1585 14385 -1565
rect 14365 -1635 14385 -1615
rect 15565 -985 15585 -965
rect 15565 -1035 15585 -1015
rect 15565 -1085 15585 -1065
rect 15565 -1135 15585 -1115
rect 15565 -1185 15585 -1165
rect 15565 -1235 15585 -1215
rect 15565 -1285 15585 -1265
rect 15565 -1335 15585 -1315
rect 15565 -1385 15585 -1365
rect 15565 -1435 15585 -1415
rect 15565 -1485 15585 -1465
rect 15565 -1535 15585 -1515
rect 15565 -1585 15585 -1565
rect 15565 -1635 15585 -1615
rect 16765 -985 16785 -965
rect 16765 -1035 16785 -1015
rect 16765 -1085 16785 -1065
rect 16765 -1135 16785 -1115
rect 16765 -1185 16785 -1165
rect 16765 -1235 16785 -1215
rect 16765 -1285 16785 -1265
rect 16765 -1335 16785 -1315
rect 16765 -1385 16785 -1365
rect 16765 -1435 16785 -1415
rect 16765 -1485 16785 -1465
rect 16765 -1535 16785 -1515
rect 16765 -1585 16785 -1565
rect 16765 -1635 16785 -1615
rect 17965 -985 17985 -965
rect 17965 -1035 17985 -1015
rect 17965 -1085 17985 -1065
rect 17965 -1135 17985 -1115
rect 17965 -1185 17985 -1165
rect 17965 -1235 17985 -1215
rect 17965 -1285 17985 -1265
rect 17965 -1335 17985 -1315
rect 17965 -1385 17985 -1365
rect 17965 -1435 17985 -1415
rect 17965 -1485 17985 -1465
rect 17965 -1535 17985 -1515
rect 17965 -1585 17985 -1565
rect 17965 -1635 17985 -1615
rect 19165 -985 19185 -965
rect 19165 -1035 19185 -1015
rect 19165 -1085 19185 -1065
rect 19165 -1135 19185 -1115
rect 19165 -1185 19185 -1165
rect 19165 -1235 19185 -1215
rect 19165 -1285 19185 -1265
rect 19165 -1335 19185 -1315
rect 19165 -1385 19185 -1365
rect 19165 -1435 19185 -1415
rect 19165 -1485 19185 -1465
rect 19165 -1535 19185 -1515
rect 19165 -1585 19185 -1565
rect 19165 -1635 19185 -1615
rect 20365 -985 20385 -965
rect 20365 -1035 20385 -1015
rect 20365 -1085 20385 -1065
rect 20365 -1135 20385 -1115
rect 20365 -1185 20385 -1165
rect 20365 -1235 20385 -1215
rect 20365 -1285 20385 -1265
rect 20365 -1335 20385 -1315
rect 20365 -1385 20385 -1365
rect 20365 -1435 20385 -1415
rect 20365 -1485 20385 -1465
rect 20365 -1535 20385 -1515
rect 20365 -1585 20385 -1565
rect 20365 -1635 20385 -1615
rect -635 -1735 -615 -1715
rect -35 -1735 -15 -1715
rect 8365 -1735 8385 -1715
rect 10765 -1735 10785 -1715
rect 15565 -1735 15585 -1715
rect 17965 -1735 17985 -1715
rect 20365 -1735 20385 -1715
<< metal1 >>
rect -650 5190 -600 5200
rect -650 5160 -640 5190
rect -610 5160 -600 5190
rect -650 5085 -600 5160
rect -50 5190 0 5200
rect -50 5160 -40 5190
rect -10 5160 0 5190
rect -650 5065 -635 5085
rect -615 5065 -600 5085
rect -650 5040 -600 5065
rect -650 5010 -640 5040
rect -610 5010 -600 5040
rect -650 4985 -600 5010
rect -650 4965 -635 4985
rect -615 4965 -600 4985
rect -650 4940 -600 4965
rect -650 4910 -640 4940
rect -610 4910 -600 4940
rect -650 4885 -600 4910
rect -650 4865 -635 4885
rect -615 4865 -600 4885
rect -650 4840 -600 4865
rect -650 4810 -640 4840
rect -610 4810 -600 4840
rect -650 4785 -600 4810
rect -650 4765 -635 4785
rect -615 4765 -600 4785
rect -650 4740 -600 4765
rect -650 4710 -640 4740
rect -610 4710 -600 4740
rect -650 4685 -600 4710
rect -650 4665 -635 4685
rect -615 4665 -600 4685
rect -650 4640 -600 4665
rect -650 4610 -640 4640
rect -610 4610 -600 4640
rect -650 4440 -600 4610
rect -500 5085 -450 5100
rect -500 5065 -485 5085
rect -465 5065 -450 5085
rect -500 5035 -450 5065
rect -500 5015 -485 5035
rect -465 5015 -450 5035
rect -500 4985 -450 5015
rect -500 4965 -485 4985
rect -465 4965 -450 4985
rect -500 4935 -450 4965
rect -500 4915 -485 4935
rect -465 4915 -450 4935
rect -500 4885 -450 4915
rect -500 4865 -485 4885
rect -465 4865 -450 4885
rect -500 4835 -450 4865
rect -500 4815 -485 4835
rect -465 4815 -450 4835
rect -500 4785 -450 4815
rect -500 4765 -485 4785
rect -465 4765 -450 4785
rect -500 4735 -450 4765
rect -500 4715 -485 4735
rect -465 4715 -450 4735
rect -500 4685 -450 4715
rect -350 5085 -300 5100
rect -350 5065 -335 5085
rect -315 5065 -300 5085
rect -350 5035 -300 5065
rect -350 5015 -335 5035
rect -315 5015 -300 5035
rect -350 4985 -300 5015
rect -350 4965 -335 4985
rect -315 4965 -300 4985
rect -350 4935 -300 4965
rect -350 4915 -335 4935
rect -315 4915 -300 4935
rect -350 4885 -300 4915
rect -350 4865 -335 4885
rect -315 4865 -300 4885
rect -350 4835 -300 4865
rect -350 4815 -335 4835
rect -315 4815 -300 4835
rect -350 4785 -300 4815
rect -350 4765 -335 4785
rect -315 4765 -300 4785
rect -350 4735 -300 4765
rect -350 4715 -335 4735
rect -315 4715 -300 4735
rect -350 4700 -300 4715
rect -200 5085 -150 5100
rect -200 5065 -185 5085
rect -165 5065 -150 5085
rect -200 5035 -150 5065
rect -200 5015 -185 5035
rect -165 5015 -150 5035
rect -200 4985 -150 5015
rect -200 4965 -185 4985
rect -165 4965 -150 4985
rect -200 4935 -150 4965
rect -200 4915 -185 4935
rect -165 4915 -150 4935
rect -200 4885 -150 4915
rect -200 4865 -185 4885
rect -165 4865 -150 4885
rect -200 4835 -150 4865
rect -200 4815 -185 4835
rect -165 4815 -150 4835
rect -200 4785 -150 4815
rect -200 4765 -185 4785
rect -165 4765 -150 4785
rect -200 4735 -150 4765
rect -200 4715 -185 4735
rect -165 4715 -150 4735
rect -500 4665 -485 4685
rect -465 4665 -450 4685
rect -500 4650 -450 4665
rect -200 4685 -150 4715
rect -200 4665 -185 4685
rect -165 4665 -150 4685
rect -200 4650 -150 4665
rect -500 4635 -150 4650
rect -500 4615 -485 4635
rect -465 4615 -185 4635
rect -165 4615 -150 4635
rect -500 4600 -150 4615
rect -50 5085 0 5160
rect 4150 5190 4200 5200
rect 4150 5160 4160 5190
rect 4190 5160 4200 5190
rect -50 5065 -35 5085
rect -15 5065 0 5085
rect -50 5035 0 5065
rect -50 5015 -35 5035
rect -15 5015 0 5035
rect -50 4985 0 5015
rect -50 4965 -35 4985
rect -15 4965 0 4985
rect -50 4935 0 4965
rect -50 4915 -35 4935
rect -15 4915 0 4935
rect -50 4885 0 4915
rect -50 4865 -35 4885
rect -15 4865 0 4885
rect -50 4835 0 4865
rect -50 4815 -35 4835
rect -15 4815 0 4835
rect -50 4785 0 4815
rect -50 4765 -35 4785
rect -15 4765 0 4785
rect -50 4735 0 4765
rect -50 4715 -35 4735
rect -15 4715 0 4735
rect -500 4540 -450 4550
rect -500 4510 -490 4540
rect -460 4510 -450 4540
rect -500 4500 -450 4510
rect -350 4540 -300 4600
rect -350 4510 -340 4540
rect -310 4510 -300 4540
rect -350 4450 -300 4510
rect -200 4540 -150 4550
rect -200 4510 -190 4540
rect -160 4510 -150 4540
rect -200 4500 -150 4510
rect -650 4410 -640 4440
rect -610 4410 -600 4440
rect -650 4385 -600 4410
rect -650 4365 -635 4385
rect -615 4365 -600 4385
rect -650 4340 -600 4365
rect -650 4310 -640 4340
rect -610 4310 -600 4340
rect -650 4285 -600 4310
rect -650 4265 -635 4285
rect -615 4265 -600 4285
rect -650 4240 -600 4265
rect -650 4210 -640 4240
rect -610 4210 -600 4240
rect -650 4185 -600 4210
rect -650 4165 -635 4185
rect -615 4165 -600 4185
rect -650 4140 -600 4165
rect -650 4110 -640 4140
rect -610 4110 -600 4140
rect -650 4085 -600 4110
rect -650 4065 -635 4085
rect -615 4065 -600 4085
rect -650 4040 -600 4065
rect -650 4010 -640 4040
rect -610 4010 -600 4040
rect -650 3985 -600 4010
rect -650 3965 -635 3985
rect -615 3965 -600 3985
rect -650 3890 -600 3965
rect -500 4435 -150 4450
rect -500 4415 -485 4435
rect -465 4415 -185 4435
rect -165 4415 -150 4435
rect -500 4400 -150 4415
rect -500 4385 -450 4400
rect -500 4365 -485 4385
rect -465 4365 -450 4385
rect -500 4335 -450 4365
rect -200 4385 -150 4400
rect -200 4365 -185 4385
rect -165 4365 -150 4385
rect -500 4315 -485 4335
rect -465 4315 -450 4335
rect -500 4285 -450 4315
rect -500 4265 -485 4285
rect -465 4265 -450 4285
rect -500 4235 -450 4265
rect -500 4215 -485 4235
rect -465 4215 -450 4235
rect -500 4185 -450 4215
rect -500 4165 -485 4185
rect -465 4165 -450 4185
rect -500 4135 -450 4165
rect -500 4115 -485 4135
rect -465 4115 -450 4135
rect -500 4085 -450 4115
rect -500 4065 -485 4085
rect -465 4065 -450 4085
rect -500 4035 -450 4065
rect -500 4015 -485 4035
rect -465 4015 -450 4035
rect -500 3985 -450 4015
rect -500 3965 -485 3985
rect -465 3965 -450 3985
rect -500 3950 -450 3965
rect -350 4335 -300 4350
rect -350 4315 -335 4335
rect -315 4315 -300 4335
rect -350 4285 -300 4315
rect -350 4265 -335 4285
rect -315 4265 -300 4285
rect -350 4235 -300 4265
rect -350 4215 -335 4235
rect -315 4215 -300 4235
rect -350 4185 -300 4215
rect -350 4165 -335 4185
rect -315 4165 -300 4185
rect -350 4135 -300 4165
rect -350 4115 -335 4135
rect -315 4115 -300 4135
rect -350 4085 -300 4115
rect -350 4065 -335 4085
rect -315 4065 -300 4085
rect -350 4035 -300 4065
rect -350 4015 -335 4035
rect -315 4015 -300 4035
rect -350 3985 -300 4015
rect -350 3965 -335 3985
rect -315 3965 -300 3985
rect -350 3950 -300 3965
rect -200 4335 -150 4365
rect -200 4315 -185 4335
rect -165 4315 -150 4335
rect -200 4285 -150 4315
rect -200 4265 -185 4285
rect -165 4265 -150 4285
rect -200 4235 -150 4265
rect -200 4215 -185 4235
rect -165 4215 -150 4235
rect -200 4185 -150 4215
rect -200 4165 -185 4185
rect -165 4165 -150 4185
rect -200 4135 -150 4165
rect -200 4115 -185 4135
rect -165 4115 -150 4135
rect -200 4085 -150 4115
rect -200 4065 -185 4085
rect -165 4065 -150 4085
rect -200 4035 -150 4065
rect -200 4015 -185 4035
rect -165 4015 -150 4035
rect -200 3985 -150 4015
rect -200 3965 -185 3985
rect -165 3965 -150 3985
rect -200 3950 -150 3965
rect -50 4440 0 4715
rect 550 5085 3600 5100
rect 550 5065 565 5085
rect 585 5065 865 5085
rect 885 5065 1165 5085
rect 1185 5065 1465 5085
rect 1485 5065 1765 5085
rect 1785 5065 2065 5085
rect 2085 5065 2365 5085
rect 2385 5065 2665 5085
rect 2685 5065 2965 5085
rect 2985 5065 3265 5085
rect 3285 5065 3565 5085
rect 3585 5065 3600 5085
rect 550 5050 3600 5065
rect 550 5035 600 5050
rect 550 5015 565 5035
rect 585 5015 600 5035
rect 550 4985 600 5015
rect 850 5035 900 5050
rect 850 5015 865 5035
rect 885 5015 900 5035
rect 550 4965 565 4985
rect 585 4965 600 4985
rect 550 4935 600 4965
rect 550 4915 565 4935
rect 585 4915 600 4935
rect 550 4885 600 4915
rect 550 4865 565 4885
rect 585 4865 600 4885
rect 550 4835 600 4865
rect 550 4815 565 4835
rect 585 4815 600 4835
rect 550 4785 600 4815
rect 550 4765 565 4785
rect 585 4765 600 4785
rect 550 4735 600 4765
rect 550 4715 565 4735
rect 585 4715 600 4735
rect 550 4685 600 4715
rect 550 4665 565 4685
rect 585 4665 600 4685
rect 550 4635 600 4665
rect 550 4615 565 4635
rect 585 4615 600 4635
rect 550 4600 600 4615
rect 700 4985 750 5000
rect 700 4965 715 4985
rect 735 4965 750 4985
rect 700 4935 750 4965
rect 700 4915 715 4935
rect 735 4915 750 4935
rect 700 4885 750 4915
rect 700 4865 715 4885
rect 735 4865 750 4885
rect 700 4835 750 4865
rect 700 4815 715 4835
rect 735 4815 750 4835
rect 700 4785 750 4815
rect 700 4765 715 4785
rect 735 4765 750 4785
rect 700 4735 750 4765
rect 700 4715 715 4735
rect 735 4715 750 4735
rect 700 4685 750 4715
rect 850 4985 900 5015
rect 1150 5035 1200 5050
rect 1150 5015 1165 5035
rect 1185 5015 1200 5035
rect 850 4965 865 4985
rect 885 4965 900 4985
rect 850 4935 900 4965
rect 850 4915 865 4935
rect 885 4915 900 4935
rect 850 4885 900 4915
rect 850 4865 865 4885
rect 885 4865 900 4885
rect 850 4835 900 4865
rect 850 4815 865 4835
rect 885 4815 900 4835
rect 850 4785 900 4815
rect 850 4765 865 4785
rect 885 4765 900 4785
rect 850 4735 900 4765
rect 850 4715 865 4735
rect 885 4715 900 4735
rect 850 4700 900 4715
rect 1000 4985 1050 5000
rect 1000 4965 1015 4985
rect 1035 4965 1050 4985
rect 1000 4935 1050 4965
rect 1000 4915 1015 4935
rect 1035 4915 1050 4935
rect 1000 4885 1050 4915
rect 1000 4865 1015 4885
rect 1035 4865 1050 4885
rect 1000 4835 1050 4865
rect 1000 4815 1015 4835
rect 1035 4815 1050 4835
rect 1000 4785 1050 4815
rect 1000 4765 1015 4785
rect 1035 4765 1050 4785
rect 1000 4735 1050 4765
rect 1000 4715 1015 4735
rect 1035 4715 1050 4735
rect 700 4665 715 4685
rect 735 4665 750 4685
rect 700 4650 750 4665
rect 1000 4685 1050 4715
rect 1150 4985 1200 5015
rect 1450 5035 1500 5050
rect 1450 5015 1465 5035
rect 1485 5015 1500 5035
rect 1150 4965 1165 4985
rect 1185 4965 1200 4985
rect 1150 4935 1200 4965
rect 1150 4915 1165 4935
rect 1185 4915 1200 4935
rect 1150 4885 1200 4915
rect 1150 4865 1165 4885
rect 1185 4865 1200 4885
rect 1150 4835 1200 4865
rect 1150 4815 1165 4835
rect 1185 4815 1200 4835
rect 1150 4785 1200 4815
rect 1150 4765 1165 4785
rect 1185 4765 1200 4785
rect 1150 4735 1200 4765
rect 1150 4715 1165 4735
rect 1185 4715 1200 4735
rect 1150 4700 1200 4715
rect 1300 4985 1350 5000
rect 1300 4965 1315 4985
rect 1335 4965 1350 4985
rect 1300 4935 1350 4965
rect 1300 4915 1315 4935
rect 1335 4915 1350 4935
rect 1300 4885 1350 4915
rect 1300 4865 1315 4885
rect 1335 4865 1350 4885
rect 1300 4835 1350 4865
rect 1300 4815 1315 4835
rect 1335 4815 1350 4835
rect 1300 4785 1350 4815
rect 1300 4765 1315 4785
rect 1335 4765 1350 4785
rect 1300 4735 1350 4765
rect 1300 4715 1315 4735
rect 1335 4715 1350 4735
rect 1000 4665 1015 4685
rect 1035 4665 1050 4685
rect 1000 4650 1050 4665
rect 1300 4685 1350 4715
rect 1450 4985 1500 5015
rect 1750 5035 1800 5050
rect 1750 5015 1765 5035
rect 1785 5015 1800 5035
rect 1450 4965 1465 4985
rect 1485 4965 1500 4985
rect 1450 4935 1500 4965
rect 1450 4915 1465 4935
rect 1485 4915 1500 4935
rect 1450 4885 1500 4915
rect 1450 4865 1465 4885
rect 1485 4865 1500 4885
rect 1450 4835 1500 4865
rect 1450 4815 1465 4835
rect 1485 4815 1500 4835
rect 1450 4785 1500 4815
rect 1450 4765 1465 4785
rect 1485 4765 1500 4785
rect 1450 4735 1500 4765
rect 1450 4715 1465 4735
rect 1485 4715 1500 4735
rect 1450 4700 1500 4715
rect 1600 4985 1650 5000
rect 1600 4965 1615 4985
rect 1635 4965 1650 4985
rect 1600 4935 1650 4965
rect 1600 4915 1615 4935
rect 1635 4915 1650 4935
rect 1600 4885 1650 4915
rect 1600 4865 1615 4885
rect 1635 4865 1650 4885
rect 1600 4835 1650 4865
rect 1600 4815 1615 4835
rect 1635 4815 1650 4835
rect 1600 4785 1650 4815
rect 1600 4765 1615 4785
rect 1635 4765 1650 4785
rect 1600 4735 1650 4765
rect 1600 4715 1615 4735
rect 1635 4715 1650 4735
rect 1300 4665 1315 4685
rect 1335 4665 1350 4685
rect 1300 4650 1350 4665
rect 1600 4685 1650 4715
rect 1600 4665 1615 4685
rect 1635 4665 1650 4685
rect 1600 4650 1650 4665
rect 700 4635 1650 4650
rect 700 4615 715 4635
rect 735 4615 1650 4635
rect 700 4600 1650 4615
rect 1750 4985 1800 5015
rect 2050 5035 2100 5050
rect 2050 5015 2065 5035
rect 2085 5015 2100 5035
rect 1750 4965 1765 4985
rect 1785 4965 1800 4985
rect 1750 4935 1800 4965
rect 1750 4915 1765 4935
rect 1785 4915 1800 4935
rect 1750 4885 1800 4915
rect 1750 4865 1765 4885
rect 1785 4865 1800 4885
rect 1750 4835 1800 4865
rect 1750 4815 1765 4835
rect 1785 4815 1800 4835
rect 1750 4785 1800 4815
rect 1750 4765 1765 4785
rect 1785 4765 1800 4785
rect 1750 4735 1800 4765
rect 1750 4715 1765 4735
rect 1785 4715 1800 4735
rect 1750 4685 1800 4715
rect 1750 4665 1765 4685
rect 1785 4665 1800 4685
rect 1750 4635 1800 4665
rect 1750 4615 1765 4635
rect 1785 4615 1800 4635
rect 100 4540 150 4550
rect 100 4510 110 4540
rect 140 4510 150 4540
rect 100 4500 150 4510
rect 400 4540 450 4550
rect 400 4510 410 4540
rect 440 4510 450 4540
rect 400 4500 450 4510
rect 700 4540 750 4550
rect 700 4510 710 4540
rect 740 4510 750 4540
rect 700 4500 750 4510
rect 1000 4540 1050 4550
rect 1000 4510 1010 4540
rect 1040 4510 1050 4540
rect 1000 4500 1050 4510
rect 1150 4540 1200 4550
rect 1150 4510 1160 4540
rect 1190 4510 1200 4540
rect 1150 4500 1200 4510
rect 1300 4540 1350 4550
rect 1300 4510 1310 4540
rect 1340 4510 1350 4540
rect 1300 4500 1350 4510
rect 1600 4540 1650 4550
rect 1600 4510 1610 4540
rect 1640 4510 1650 4540
rect 1600 4500 1650 4510
rect -50 4410 -40 4440
rect -10 4410 0 4440
rect -50 4340 0 4410
rect -50 4310 -40 4340
rect -10 4310 0 4340
rect -50 4285 0 4310
rect -50 4265 -35 4285
rect -15 4265 0 4285
rect -50 4240 0 4265
rect -50 4210 -40 4240
rect -10 4210 0 4240
rect -50 4185 0 4210
rect -50 4165 -35 4185
rect -15 4165 0 4185
rect -50 4140 0 4165
rect -50 4110 -40 4140
rect -10 4110 0 4140
rect -50 4085 0 4110
rect -50 4065 -35 4085
rect -15 4065 0 4085
rect -50 4040 0 4065
rect -50 4010 -40 4040
rect -10 4010 0 4040
rect -50 3985 0 4010
rect -50 3965 -35 3985
rect -15 3965 0 3985
rect -650 3860 -640 3890
rect -610 3860 -600 3890
rect -650 3785 -600 3860
rect -50 3890 0 3965
rect 550 4435 600 4450
rect 550 4415 565 4435
rect 585 4415 600 4435
rect 550 4385 600 4415
rect 550 4365 565 4385
rect 585 4365 600 4385
rect 550 4335 600 4365
rect 550 4315 565 4335
rect 585 4315 600 4335
rect 550 4285 600 4315
rect 550 4265 565 4285
rect 585 4265 600 4285
rect 550 4235 600 4265
rect 550 4215 565 4235
rect 585 4215 600 4235
rect 550 4185 600 4215
rect 550 4165 565 4185
rect 585 4165 600 4185
rect 550 4135 600 4165
rect 550 4115 565 4135
rect 585 4115 600 4135
rect 550 4085 600 4115
rect 550 4065 565 4085
rect 585 4065 600 4085
rect 550 4035 600 4065
rect 700 4435 1650 4450
rect 700 4415 715 4435
rect 735 4415 1650 4435
rect 700 4400 1650 4415
rect 700 4385 750 4400
rect 700 4365 715 4385
rect 735 4365 750 4385
rect 700 4335 750 4365
rect 1000 4385 1050 4400
rect 1000 4365 1015 4385
rect 1035 4365 1050 4385
rect 700 4315 715 4335
rect 735 4315 750 4335
rect 700 4285 750 4315
rect 700 4265 715 4285
rect 735 4265 750 4285
rect 700 4235 750 4265
rect 700 4215 715 4235
rect 735 4215 750 4235
rect 700 4185 750 4215
rect 700 4165 715 4185
rect 735 4165 750 4185
rect 700 4135 750 4165
rect 700 4115 715 4135
rect 735 4115 750 4135
rect 700 4085 750 4115
rect 700 4065 715 4085
rect 735 4065 750 4085
rect 700 4050 750 4065
rect 850 4335 900 4350
rect 850 4315 865 4335
rect 885 4315 900 4335
rect 850 4285 900 4315
rect 850 4265 865 4285
rect 885 4265 900 4285
rect 850 4235 900 4265
rect 850 4215 865 4235
rect 885 4215 900 4235
rect 850 4185 900 4215
rect 850 4165 865 4185
rect 885 4165 900 4185
rect 850 4135 900 4165
rect 850 4115 865 4135
rect 885 4115 900 4135
rect 850 4085 900 4115
rect 850 4065 865 4085
rect 885 4065 900 4085
rect 550 4015 565 4035
rect 585 4015 600 4035
rect 550 4000 600 4015
rect 850 4035 900 4065
rect 1000 4335 1050 4365
rect 1300 4385 1350 4400
rect 1300 4365 1315 4385
rect 1335 4365 1350 4385
rect 1000 4315 1015 4335
rect 1035 4315 1050 4335
rect 1000 4285 1050 4315
rect 1000 4265 1015 4285
rect 1035 4265 1050 4285
rect 1000 4235 1050 4265
rect 1000 4215 1015 4235
rect 1035 4215 1050 4235
rect 1000 4185 1050 4215
rect 1000 4165 1015 4185
rect 1035 4165 1050 4185
rect 1000 4135 1050 4165
rect 1000 4115 1015 4135
rect 1035 4115 1050 4135
rect 1000 4085 1050 4115
rect 1000 4065 1015 4085
rect 1035 4065 1050 4085
rect 1000 4050 1050 4065
rect 1150 4335 1200 4350
rect 1150 4315 1165 4335
rect 1185 4315 1200 4335
rect 1150 4285 1200 4315
rect 1150 4265 1165 4285
rect 1185 4265 1200 4285
rect 1150 4235 1200 4265
rect 1150 4215 1165 4235
rect 1185 4215 1200 4235
rect 1150 4185 1200 4215
rect 1150 4165 1165 4185
rect 1185 4165 1200 4185
rect 1150 4135 1200 4165
rect 1150 4115 1165 4135
rect 1185 4115 1200 4135
rect 1150 4085 1200 4115
rect 1150 4065 1165 4085
rect 1185 4065 1200 4085
rect 850 4015 865 4035
rect 885 4015 900 4035
rect 850 4000 900 4015
rect 1150 4035 1200 4065
rect 1300 4335 1350 4365
rect 1600 4385 1650 4400
rect 1600 4365 1615 4385
rect 1635 4365 1650 4385
rect 1300 4315 1315 4335
rect 1335 4315 1350 4335
rect 1300 4285 1350 4315
rect 1300 4265 1315 4285
rect 1335 4265 1350 4285
rect 1300 4235 1350 4265
rect 1300 4215 1315 4235
rect 1335 4215 1350 4235
rect 1300 4185 1350 4215
rect 1300 4165 1315 4185
rect 1335 4165 1350 4185
rect 1300 4135 1350 4165
rect 1300 4115 1315 4135
rect 1335 4115 1350 4135
rect 1300 4085 1350 4115
rect 1300 4065 1315 4085
rect 1335 4065 1350 4085
rect 1300 4050 1350 4065
rect 1450 4335 1500 4350
rect 1450 4315 1465 4335
rect 1485 4315 1500 4335
rect 1450 4285 1500 4315
rect 1450 4265 1465 4285
rect 1485 4265 1500 4285
rect 1450 4235 1500 4265
rect 1450 4215 1465 4235
rect 1485 4215 1500 4235
rect 1450 4185 1500 4215
rect 1450 4165 1465 4185
rect 1485 4165 1500 4185
rect 1450 4135 1500 4165
rect 1450 4115 1465 4135
rect 1485 4115 1500 4135
rect 1450 4085 1500 4115
rect 1450 4065 1465 4085
rect 1485 4065 1500 4085
rect 1150 4015 1165 4035
rect 1185 4015 1200 4035
rect 1150 4000 1200 4015
rect 1450 4035 1500 4065
rect 1600 4335 1650 4365
rect 1600 4315 1615 4335
rect 1635 4315 1650 4335
rect 1600 4285 1650 4315
rect 1600 4265 1615 4285
rect 1635 4265 1650 4285
rect 1600 4235 1650 4265
rect 1600 4215 1615 4235
rect 1635 4215 1650 4235
rect 1600 4185 1650 4215
rect 1600 4165 1615 4185
rect 1635 4165 1650 4185
rect 1600 4135 1650 4165
rect 1600 4115 1615 4135
rect 1635 4115 1650 4135
rect 1600 4085 1650 4115
rect 1600 4065 1615 4085
rect 1635 4065 1650 4085
rect 1600 4050 1650 4065
rect 1750 4435 1800 4615
rect 1900 4985 1950 5000
rect 1900 4965 1915 4985
rect 1935 4965 1950 4985
rect 1900 4935 1950 4965
rect 1900 4915 1915 4935
rect 1935 4915 1950 4935
rect 1900 4885 1950 4915
rect 1900 4865 1915 4885
rect 1935 4865 1950 4885
rect 1900 4835 1950 4865
rect 1900 4815 1915 4835
rect 1935 4815 1950 4835
rect 1900 4785 1950 4815
rect 1900 4765 1915 4785
rect 1935 4765 1950 4785
rect 1900 4735 1950 4765
rect 1900 4715 1915 4735
rect 1935 4715 1950 4735
rect 1900 4685 1950 4715
rect 2050 4985 2100 5015
rect 2350 5035 2400 5050
rect 2350 5015 2365 5035
rect 2385 5015 2400 5035
rect 2050 4965 2065 4985
rect 2085 4965 2100 4985
rect 2050 4935 2100 4965
rect 2050 4915 2065 4935
rect 2085 4915 2100 4935
rect 2050 4885 2100 4915
rect 2050 4865 2065 4885
rect 2085 4865 2100 4885
rect 2050 4835 2100 4865
rect 2050 4815 2065 4835
rect 2085 4815 2100 4835
rect 2050 4785 2100 4815
rect 2050 4765 2065 4785
rect 2085 4765 2100 4785
rect 2050 4735 2100 4765
rect 2050 4715 2065 4735
rect 2085 4715 2100 4735
rect 2050 4700 2100 4715
rect 2200 4985 2250 5000
rect 2200 4965 2215 4985
rect 2235 4965 2250 4985
rect 2200 4935 2250 4965
rect 2200 4915 2215 4935
rect 2235 4915 2250 4935
rect 2200 4885 2250 4915
rect 2200 4865 2215 4885
rect 2235 4865 2250 4885
rect 2200 4835 2250 4865
rect 2200 4815 2215 4835
rect 2235 4815 2250 4835
rect 2200 4785 2250 4815
rect 2200 4765 2215 4785
rect 2235 4765 2250 4785
rect 2200 4735 2250 4765
rect 2200 4715 2215 4735
rect 2235 4715 2250 4735
rect 1900 4665 1915 4685
rect 1935 4665 1950 4685
rect 1900 4650 1950 4665
rect 2200 4685 2250 4715
rect 2200 4665 2215 4685
rect 2235 4665 2250 4685
rect 2200 4650 2250 4665
rect 1900 4635 2250 4650
rect 1900 4615 1915 4635
rect 1935 4615 2215 4635
rect 2235 4615 2250 4635
rect 1900 4600 2250 4615
rect 2350 4985 2400 5015
rect 2650 5035 2700 5050
rect 2650 5015 2665 5035
rect 2685 5015 2700 5035
rect 2350 4965 2365 4985
rect 2385 4965 2400 4985
rect 2350 4935 2400 4965
rect 2350 4915 2365 4935
rect 2385 4915 2400 4935
rect 2350 4885 2400 4915
rect 2350 4865 2365 4885
rect 2385 4865 2400 4885
rect 2350 4835 2400 4865
rect 2350 4815 2365 4835
rect 2385 4815 2400 4835
rect 2350 4785 2400 4815
rect 2350 4765 2365 4785
rect 2385 4765 2400 4785
rect 2350 4735 2400 4765
rect 2350 4715 2365 4735
rect 2385 4715 2400 4735
rect 2350 4685 2400 4715
rect 2350 4665 2365 4685
rect 2385 4665 2400 4685
rect 2350 4635 2400 4665
rect 2350 4615 2365 4635
rect 2385 4615 2400 4635
rect 1900 4540 1950 4550
rect 1900 4510 1910 4540
rect 1940 4510 1950 4540
rect 1900 4500 1950 4510
rect 2050 4540 2100 4600
rect 2050 4510 2060 4540
rect 2090 4510 2100 4540
rect 2050 4450 2100 4510
rect 2200 4540 2250 4550
rect 2200 4510 2210 4540
rect 2240 4510 2250 4540
rect 2200 4500 2250 4510
rect 1750 4415 1765 4435
rect 1785 4415 1800 4435
rect 1750 4385 1800 4415
rect 1750 4365 1765 4385
rect 1785 4365 1800 4385
rect 1750 4335 1800 4365
rect 1750 4315 1765 4335
rect 1785 4315 1800 4335
rect 1750 4285 1800 4315
rect 1750 4265 1765 4285
rect 1785 4265 1800 4285
rect 1750 4235 1800 4265
rect 1750 4215 1765 4235
rect 1785 4215 1800 4235
rect 1750 4185 1800 4215
rect 1750 4165 1765 4185
rect 1785 4165 1800 4185
rect 1750 4135 1800 4165
rect 1750 4115 1765 4135
rect 1785 4115 1800 4135
rect 1750 4085 1800 4115
rect 1750 4065 1765 4085
rect 1785 4065 1800 4085
rect 1450 4015 1465 4035
rect 1485 4015 1500 4035
rect 1450 4000 1500 4015
rect 1750 4035 1800 4065
rect 1900 4435 2250 4450
rect 1900 4415 1915 4435
rect 1935 4415 2215 4435
rect 2235 4415 2250 4435
rect 1900 4400 2250 4415
rect 1900 4385 1950 4400
rect 1900 4365 1915 4385
rect 1935 4365 1950 4385
rect 1900 4335 1950 4365
rect 2200 4385 2250 4400
rect 2200 4365 2215 4385
rect 2235 4365 2250 4385
rect 1900 4315 1915 4335
rect 1935 4315 1950 4335
rect 1900 4285 1950 4315
rect 1900 4265 1915 4285
rect 1935 4265 1950 4285
rect 1900 4235 1950 4265
rect 1900 4215 1915 4235
rect 1935 4215 1950 4235
rect 1900 4185 1950 4215
rect 1900 4165 1915 4185
rect 1935 4165 1950 4185
rect 1900 4135 1950 4165
rect 1900 4115 1915 4135
rect 1935 4115 1950 4135
rect 1900 4085 1950 4115
rect 1900 4065 1915 4085
rect 1935 4065 1950 4085
rect 1900 4050 1950 4065
rect 2050 4335 2100 4350
rect 2050 4315 2065 4335
rect 2085 4315 2100 4335
rect 2050 4285 2100 4315
rect 2050 4265 2065 4285
rect 2085 4265 2100 4285
rect 2050 4235 2100 4265
rect 2050 4215 2065 4235
rect 2085 4215 2100 4235
rect 2050 4185 2100 4215
rect 2050 4165 2065 4185
rect 2085 4165 2100 4185
rect 2050 4135 2100 4165
rect 2050 4115 2065 4135
rect 2085 4115 2100 4135
rect 2050 4085 2100 4115
rect 2050 4065 2065 4085
rect 2085 4065 2100 4085
rect 1750 4015 1765 4035
rect 1785 4015 1800 4035
rect 1750 4000 1800 4015
rect 2050 4035 2100 4065
rect 2200 4335 2250 4365
rect 2200 4315 2215 4335
rect 2235 4315 2250 4335
rect 2200 4285 2250 4315
rect 2200 4265 2215 4285
rect 2235 4265 2250 4285
rect 2200 4235 2250 4265
rect 2200 4215 2215 4235
rect 2235 4215 2250 4235
rect 2200 4185 2250 4215
rect 2200 4165 2215 4185
rect 2235 4165 2250 4185
rect 2200 4135 2250 4165
rect 2200 4115 2215 4135
rect 2235 4115 2250 4135
rect 2200 4085 2250 4115
rect 2200 4065 2215 4085
rect 2235 4065 2250 4085
rect 2200 4050 2250 4065
rect 2350 4435 2400 4615
rect 2500 4985 2550 5000
rect 2500 4965 2515 4985
rect 2535 4965 2550 4985
rect 2500 4935 2550 4965
rect 2500 4915 2515 4935
rect 2535 4915 2550 4935
rect 2500 4885 2550 4915
rect 2500 4865 2515 4885
rect 2535 4865 2550 4885
rect 2500 4835 2550 4865
rect 2500 4815 2515 4835
rect 2535 4815 2550 4835
rect 2500 4785 2550 4815
rect 2500 4765 2515 4785
rect 2535 4765 2550 4785
rect 2500 4735 2550 4765
rect 2500 4715 2515 4735
rect 2535 4715 2550 4735
rect 2500 4685 2550 4715
rect 2650 4985 2700 5015
rect 2950 5035 3000 5050
rect 2950 5015 2965 5035
rect 2985 5015 3000 5035
rect 2650 4965 2665 4985
rect 2685 4965 2700 4985
rect 2650 4935 2700 4965
rect 2650 4915 2665 4935
rect 2685 4915 2700 4935
rect 2650 4885 2700 4915
rect 2650 4865 2665 4885
rect 2685 4865 2700 4885
rect 2650 4835 2700 4865
rect 2650 4815 2665 4835
rect 2685 4815 2700 4835
rect 2650 4785 2700 4815
rect 2650 4765 2665 4785
rect 2685 4765 2700 4785
rect 2650 4735 2700 4765
rect 2650 4715 2665 4735
rect 2685 4715 2700 4735
rect 2650 4700 2700 4715
rect 2800 4985 2850 5000
rect 2800 4965 2815 4985
rect 2835 4965 2850 4985
rect 2800 4935 2850 4965
rect 2800 4915 2815 4935
rect 2835 4915 2850 4935
rect 2800 4885 2850 4915
rect 2800 4865 2815 4885
rect 2835 4865 2850 4885
rect 2800 4835 2850 4865
rect 2800 4815 2815 4835
rect 2835 4815 2850 4835
rect 2800 4785 2850 4815
rect 2800 4765 2815 4785
rect 2835 4765 2850 4785
rect 2800 4735 2850 4765
rect 2800 4715 2815 4735
rect 2835 4715 2850 4735
rect 2500 4665 2515 4685
rect 2535 4665 2550 4685
rect 2500 4650 2550 4665
rect 2800 4685 2850 4715
rect 2950 4985 3000 5015
rect 3250 5035 3300 5050
rect 3250 5015 3265 5035
rect 3285 5015 3300 5035
rect 2950 4965 2965 4985
rect 2985 4965 3000 4985
rect 2950 4935 3000 4965
rect 2950 4915 2965 4935
rect 2985 4915 3000 4935
rect 2950 4885 3000 4915
rect 2950 4865 2965 4885
rect 2985 4865 3000 4885
rect 2950 4835 3000 4865
rect 2950 4815 2965 4835
rect 2985 4815 3000 4835
rect 2950 4785 3000 4815
rect 2950 4765 2965 4785
rect 2985 4765 3000 4785
rect 2950 4735 3000 4765
rect 2950 4715 2965 4735
rect 2985 4715 3000 4735
rect 2950 4700 3000 4715
rect 3100 4985 3150 5000
rect 3100 4965 3115 4985
rect 3135 4965 3150 4985
rect 3100 4935 3150 4965
rect 3100 4915 3115 4935
rect 3135 4915 3150 4935
rect 3100 4885 3150 4915
rect 3100 4865 3115 4885
rect 3135 4865 3150 4885
rect 3100 4835 3150 4865
rect 3100 4815 3115 4835
rect 3135 4815 3150 4835
rect 3100 4785 3150 4815
rect 3100 4765 3115 4785
rect 3135 4765 3150 4785
rect 3100 4735 3150 4765
rect 3100 4715 3115 4735
rect 3135 4715 3150 4735
rect 2800 4665 2815 4685
rect 2835 4665 2850 4685
rect 2800 4650 2850 4665
rect 3100 4685 3150 4715
rect 3250 4985 3300 5015
rect 3550 5035 3600 5050
rect 3550 5015 3565 5035
rect 3585 5015 3600 5035
rect 3250 4965 3265 4985
rect 3285 4965 3300 4985
rect 3250 4935 3300 4965
rect 3250 4915 3265 4935
rect 3285 4915 3300 4935
rect 3250 4885 3300 4915
rect 3250 4865 3265 4885
rect 3285 4865 3300 4885
rect 3250 4835 3300 4865
rect 3250 4815 3265 4835
rect 3285 4815 3300 4835
rect 3250 4785 3300 4815
rect 3250 4765 3265 4785
rect 3285 4765 3300 4785
rect 3250 4735 3300 4765
rect 3250 4715 3265 4735
rect 3285 4715 3300 4735
rect 3250 4700 3300 4715
rect 3400 4985 3450 5000
rect 3400 4965 3415 4985
rect 3435 4965 3450 4985
rect 3400 4935 3450 4965
rect 3400 4915 3415 4935
rect 3435 4915 3450 4935
rect 3400 4885 3450 4915
rect 3400 4865 3415 4885
rect 3435 4865 3450 4885
rect 3400 4835 3450 4865
rect 3400 4815 3415 4835
rect 3435 4815 3450 4835
rect 3400 4785 3450 4815
rect 3400 4765 3415 4785
rect 3435 4765 3450 4785
rect 3400 4735 3450 4765
rect 3400 4715 3415 4735
rect 3435 4715 3450 4735
rect 3100 4665 3115 4685
rect 3135 4665 3150 4685
rect 3100 4650 3150 4665
rect 3400 4685 3450 4715
rect 3400 4665 3415 4685
rect 3435 4665 3450 4685
rect 3400 4650 3450 4665
rect 2500 4635 3450 4650
rect 2500 4615 3415 4635
rect 3435 4615 3450 4635
rect 2500 4600 3450 4615
rect 3550 4985 3600 5015
rect 3550 4965 3565 4985
rect 3585 4965 3600 4985
rect 3550 4935 3600 4965
rect 3550 4915 3565 4935
rect 3585 4915 3600 4935
rect 3550 4885 3600 4915
rect 3550 4865 3565 4885
rect 3585 4865 3600 4885
rect 3550 4835 3600 4865
rect 3550 4815 3565 4835
rect 3585 4815 3600 4835
rect 3550 4785 3600 4815
rect 3550 4765 3565 4785
rect 3585 4765 3600 4785
rect 3550 4735 3600 4765
rect 3550 4715 3565 4735
rect 3585 4715 3600 4735
rect 3550 4685 3600 4715
rect 3550 4665 3565 4685
rect 3585 4665 3600 4685
rect 3550 4635 3600 4665
rect 3550 4615 3565 4635
rect 3585 4615 3600 4635
rect 3550 4600 3600 4615
rect 4150 5085 4200 5160
rect 8350 5190 8400 5200
rect 8350 5160 8360 5190
rect 8390 5160 8400 5190
rect 4150 5065 4165 5085
rect 4185 5065 4200 5085
rect 4150 5035 4200 5065
rect 4150 5015 4165 5035
rect 4185 5015 4200 5035
rect 4150 4985 4200 5015
rect 4150 4965 4165 4985
rect 4185 4965 4200 4985
rect 4150 4935 4200 4965
rect 4150 4915 4165 4935
rect 4185 4915 4200 4935
rect 4150 4885 4200 4915
rect 4150 4865 4165 4885
rect 4185 4865 4200 4885
rect 4150 4835 4200 4865
rect 4150 4815 4165 4835
rect 4185 4815 4200 4835
rect 4150 4785 4200 4815
rect 4150 4765 4165 4785
rect 4185 4765 4200 4785
rect 4150 4735 4200 4765
rect 4150 4715 4165 4735
rect 4185 4715 4200 4735
rect 2500 4540 2550 4550
rect 2500 4510 2510 4540
rect 2540 4510 2550 4540
rect 2500 4500 2550 4510
rect 2800 4540 2850 4550
rect 2800 4510 2810 4540
rect 2840 4510 2850 4540
rect 2800 4500 2850 4510
rect 2950 4540 3000 4550
rect 2950 4510 2960 4540
rect 2990 4510 3000 4540
rect 2950 4500 3000 4510
rect 3100 4540 3150 4550
rect 3100 4510 3110 4540
rect 3140 4510 3150 4540
rect 3100 4500 3150 4510
rect 3400 4540 3450 4550
rect 3400 4510 3410 4540
rect 3440 4510 3450 4540
rect 3400 4500 3450 4510
rect 3700 4540 3750 4550
rect 3700 4510 3710 4540
rect 3740 4510 3750 4540
rect 3700 4500 3750 4510
rect 4000 4540 4050 4550
rect 4000 4510 4010 4540
rect 4040 4510 4050 4540
rect 4000 4500 4050 4510
rect 2350 4415 2365 4435
rect 2385 4415 2400 4435
rect 2350 4385 2400 4415
rect 2350 4365 2365 4385
rect 2385 4365 2400 4385
rect 2350 4335 2400 4365
rect 2350 4315 2365 4335
rect 2385 4315 2400 4335
rect 2350 4285 2400 4315
rect 2350 4265 2365 4285
rect 2385 4265 2400 4285
rect 2350 4235 2400 4265
rect 2350 4215 2365 4235
rect 2385 4215 2400 4235
rect 2350 4185 2400 4215
rect 2350 4165 2365 4185
rect 2385 4165 2400 4185
rect 2350 4135 2400 4165
rect 2350 4115 2365 4135
rect 2385 4115 2400 4135
rect 2350 4085 2400 4115
rect 2350 4065 2365 4085
rect 2385 4065 2400 4085
rect 2050 4015 2065 4035
rect 2085 4015 2100 4035
rect 2050 4000 2100 4015
rect 2350 4035 2400 4065
rect 2500 4435 3450 4450
rect 2500 4415 3415 4435
rect 3435 4415 3450 4435
rect 2500 4400 3450 4415
rect 2500 4385 2550 4400
rect 2500 4365 2515 4385
rect 2535 4365 2550 4385
rect 2500 4335 2550 4365
rect 2800 4385 2850 4400
rect 2800 4365 2815 4385
rect 2835 4365 2850 4385
rect 2500 4315 2515 4335
rect 2535 4315 2550 4335
rect 2500 4285 2550 4315
rect 2500 4265 2515 4285
rect 2535 4265 2550 4285
rect 2500 4235 2550 4265
rect 2500 4215 2515 4235
rect 2535 4215 2550 4235
rect 2500 4185 2550 4215
rect 2500 4165 2515 4185
rect 2535 4165 2550 4185
rect 2500 4135 2550 4165
rect 2500 4115 2515 4135
rect 2535 4115 2550 4135
rect 2500 4085 2550 4115
rect 2500 4065 2515 4085
rect 2535 4065 2550 4085
rect 2500 4050 2550 4065
rect 2650 4335 2700 4350
rect 2650 4315 2665 4335
rect 2685 4315 2700 4335
rect 2650 4285 2700 4315
rect 2650 4265 2665 4285
rect 2685 4265 2700 4285
rect 2650 4235 2700 4265
rect 2650 4215 2665 4235
rect 2685 4215 2700 4235
rect 2650 4185 2700 4215
rect 2650 4165 2665 4185
rect 2685 4165 2700 4185
rect 2650 4135 2700 4165
rect 2650 4115 2665 4135
rect 2685 4115 2700 4135
rect 2650 4085 2700 4115
rect 2650 4065 2665 4085
rect 2685 4065 2700 4085
rect 2350 4015 2365 4035
rect 2385 4015 2400 4035
rect 2350 4000 2400 4015
rect 2650 4035 2700 4065
rect 2800 4335 2850 4365
rect 3100 4385 3150 4400
rect 3100 4365 3115 4385
rect 3135 4365 3150 4385
rect 2800 4315 2815 4335
rect 2835 4315 2850 4335
rect 2800 4285 2850 4315
rect 2800 4265 2815 4285
rect 2835 4265 2850 4285
rect 2800 4235 2850 4265
rect 2800 4215 2815 4235
rect 2835 4215 2850 4235
rect 2800 4185 2850 4215
rect 2800 4165 2815 4185
rect 2835 4165 2850 4185
rect 2800 4135 2850 4165
rect 2800 4115 2815 4135
rect 2835 4115 2850 4135
rect 2800 4085 2850 4115
rect 2800 4065 2815 4085
rect 2835 4065 2850 4085
rect 2800 4050 2850 4065
rect 2950 4335 3000 4350
rect 2950 4315 2965 4335
rect 2985 4315 3000 4335
rect 2950 4285 3000 4315
rect 2950 4265 2965 4285
rect 2985 4265 3000 4285
rect 2950 4235 3000 4265
rect 2950 4215 2965 4235
rect 2985 4215 3000 4235
rect 2950 4185 3000 4215
rect 2950 4165 2965 4185
rect 2985 4165 3000 4185
rect 2950 4135 3000 4165
rect 2950 4115 2965 4135
rect 2985 4115 3000 4135
rect 2950 4085 3000 4115
rect 2950 4065 2965 4085
rect 2985 4065 3000 4085
rect 2650 4015 2665 4035
rect 2685 4015 2700 4035
rect 2650 4000 2700 4015
rect 2950 4035 3000 4065
rect 3100 4335 3150 4365
rect 3400 4385 3450 4400
rect 3400 4365 3415 4385
rect 3435 4365 3450 4385
rect 3100 4315 3115 4335
rect 3135 4315 3150 4335
rect 3100 4285 3150 4315
rect 3100 4265 3115 4285
rect 3135 4265 3150 4285
rect 3100 4235 3150 4265
rect 3100 4215 3115 4235
rect 3135 4215 3150 4235
rect 3100 4185 3150 4215
rect 3100 4165 3115 4185
rect 3135 4165 3150 4185
rect 3100 4135 3150 4165
rect 3100 4115 3115 4135
rect 3135 4115 3150 4135
rect 3100 4085 3150 4115
rect 3100 4065 3115 4085
rect 3135 4065 3150 4085
rect 3100 4050 3150 4065
rect 3250 4335 3300 4350
rect 3250 4315 3265 4335
rect 3285 4315 3300 4335
rect 3250 4285 3300 4315
rect 3250 4265 3265 4285
rect 3285 4265 3300 4285
rect 3250 4235 3300 4265
rect 3250 4215 3265 4235
rect 3285 4215 3300 4235
rect 3250 4185 3300 4215
rect 3250 4165 3265 4185
rect 3285 4165 3300 4185
rect 3250 4135 3300 4165
rect 3250 4115 3265 4135
rect 3285 4115 3300 4135
rect 3250 4085 3300 4115
rect 3250 4065 3265 4085
rect 3285 4065 3300 4085
rect 2950 4015 2965 4035
rect 2985 4015 3000 4035
rect 2950 4000 3000 4015
rect 3250 4035 3300 4065
rect 3400 4335 3450 4365
rect 3400 4315 3415 4335
rect 3435 4315 3450 4335
rect 3400 4285 3450 4315
rect 3400 4265 3415 4285
rect 3435 4265 3450 4285
rect 3400 4235 3450 4265
rect 3400 4215 3415 4235
rect 3435 4215 3450 4235
rect 3400 4185 3450 4215
rect 3400 4165 3415 4185
rect 3435 4165 3450 4185
rect 3400 4135 3450 4165
rect 3400 4115 3415 4135
rect 3435 4115 3450 4135
rect 3400 4085 3450 4115
rect 3400 4065 3415 4085
rect 3435 4065 3450 4085
rect 3400 4050 3450 4065
rect 3550 4435 3600 4450
rect 3550 4415 3565 4435
rect 3585 4415 3600 4435
rect 3550 4385 3600 4415
rect 3550 4365 3565 4385
rect 3585 4365 3600 4385
rect 3550 4335 3600 4365
rect 3550 4315 3565 4335
rect 3585 4315 3600 4335
rect 3550 4285 3600 4315
rect 3550 4265 3565 4285
rect 3585 4265 3600 4285
rect 3550 4235 3600 4265
rect 3550 4215 3565 4235
rect 3585 4215 3600 4235
rect 3550 4185 3600 4215
rect 3550 4165 3565 4185
rect 3585 4165 3600 4185
rect 3550 4135 3600 4165
rect 3550 4115 3565 4135
rect 3585 4115 3600 4135
rect 3550 4085 3600 4115
rect 3550 4065 3565 4085
rect 3585 4065 3600 4085
rect 3250 4015 3265 4035
rect 3285 4015 3300 4035
rect 3250 4000 3300 4015
rect 3550 4035 3600 4065
rect 3550 4015 3565 4035
rect 3585 4015 3600 4035
rect 3550 4000 3600 4015
rect 550 3985 3600 4000
rect 550 3965 565 3985
rect 585 3965 865 3985
rect 885 3965 1165 3985
rect 1185 3965 1465 3985
rect 1485 3965 1765 3985
rect 1785 3965 2065 3985
rect 2085 3965 2365 3985
rect 2385 3965 2665 3985
rect 2685 3965 2965 3985
rect 2985 3965 3265 3985
rect 3285 3965 3565 3985
rect 3585 3965 3600 3985
rect 550 3950 3600 3965
rect 4150 4440 4200 4715
rect 4750 5085 7800 5100
rect 4750 5065 4765 5085
rect 4785 5065 5065 5085
rect 5085 5065 5365 5085
rect 5385 5065 5665 5085
rect 5685 5065 5965 5085
rect 5985 5065 6265 5085
rect 6285 5065 6565 5085
rect 6585 5065 6865 5085
rect 6885 5065 7165 5085
rect 7185 5065 7465 5085
rect 7485 5065 7765 5085
rect 7785 5065 7800 5085
rect 4750 5050 7800 5065
rect 4750 5035 4800 5050
rect 4750 5015 4765 5035
rect 4785 5015 4800 5035
rect 4750 4985 4800 5015
rect 5050 5035 5100 5050
rect 5050 5015 5065 5035
rect 5085 5015 5100 5035
rect 4750 4965 4765 4985
rect 4785 4965 4800 4985
rect 4750 4935 4800 4965
rect 4750 4915 4765 4935
rect 4785 4915 4800 4935
rect 4750 4885 4800 4915
rect 4750 4865 4765 4885
rect 4785 4865 4800 4885
rect 4750 4835 4800 4865
rect 4750 4815 4765 4835
rect 4785 4815 4800 4835
rect 4750 4785 4800 4815
rect 4750 4765 4765 4785
rect 4785 4765 4800 4785
rect 4750 4735 4800 4765
rect 4750 4715 4765 4735
rect 4785 4715 4800 4735
rect 4750 4685 4800 4715
rect 4750 4665 4765 4685
rect 4785 4665 4800 4685
rect 4750 4635 4800 4665
rect 4750 4615 4765 4635
rect 4785 4615 4800 4635
rect 4750 4600 4800 4615
rect 4900 4985 4950 5000
rect 4900 4965 4915 4985
rect 4935 4965 4950 4985
rect 4900 4935 4950 4965
rect 4900 4915 4915 4935
rect 4935 4915 4950 4935
rect 4900 4885 4950 4915
rect 4900 4865 4915 4885
rect 4935 4865 4950 4885
rect 4900 4835 4950 4865
rect 4900 4815 4915 4835
rect 4935 4815 4950 4835
rect 4900 4785 4950 4815
rect 4900 4765 4915 4785
rect 4935 4765 4950 4785
rect 4900 4735 4950 4765
rect 4900 4715 4915 4735
rect 4935 4715 4950 4735
rect 4900 4685 4950 4715
rect 5050 4985 5100 5015
rect 5350 5035 5400 5050
rect 5350 5015 5365 5035
rect 5385 5015 5400 5035
rect 5050 4965 5065 4985
rect 5085 4965 5100 4985
rect 5050 4935 5100 4965
rect 5050 4915 5065 4935
rect 5085 4915 5100 4935
rect 5050 4885 5100 4915
rect 5050 4865 5065 4885
rect 5085 4865 5100 4885
rect 5050 4835 5100 4865
rect 5050 4815 5065 4835
rect 5085 4815 5100 4835
rect 5050 4785 5100 4815
rect 5050 4765 5065 4785
rect 5085 4765 5100 4785
rect 5050 4735 5100 4765
rect 5050 4715 5065 4735
rect 5085 4715 5100 4735
rect 5050 4700 5100 4715
rect 5200 4985 5250 5000
rect 5200 4965 5215 4985
rect 5235 4965 5250 4985
rect 5200 4935 5250 4965
rect 5200 4915 5215 4935
rect 5235 4915 5250 4935
rect 5200 4885 5250 4915
rect 5200 4865 5215 4885
rect 5235 4865 5250 4885
rect 5200 4835 5250 4865
rect 5200 4815 5215 4835
rect 5235 4815 5250 4835
rect 5200 4785 5250 4815
rect 5200 4765 5215 4785
rect 5235 4765 5250 4785
rect 5200 4735 5250 4765
rect 5200 4715 5215 4735
rect 5235 4715 5250 4735
rect 4900 4665 4915 4685
rect 4935 4665 4950 4685
rect 4900 4650 4950 4665
rect 5200 4685 5250 4715
rect 5350 4985 5400 5015
rect 5650 5035 5700 5050
rect 5650 5015 5665 5035
rect 5685 5015 5700 5035
rect 5350 4965 5365 4985
rect 5385 4965 5400 4985
rect 5350 4935 5400 4965
rect 5350 4915 5365 4935
rect 5385 4915 5400 4935
rect 5350 4885 5400 4915
rect 5350 4865 5365 4885
rect 5385 4865 5400 4885
rect 5350 4835 5400 4865
rect 5350 4815 5365 4835
rect 5385 4815 5400 4835
rect 5350 4785 5400 4815
rect 5350 4765 5365 4785
rect 5385 4765 5400 4785
rect 5350 4735 5400 4765
rect 5350 4715 5365 4735
rect 5385 4715 5400 4735
rect 5350 4700 5400 4715
rect 5500 4985 5550 5000
rect 5500 4965 5515 4985
rect 5535 4965 5550 4985
rect 5500 4935 5550 4965
rect 5500 4915 5515 4935
rect 5535 4915 5550 4935
rect 5500 4885 5550 4915
rect 5500 4865 5515 4885
rect 5535 4865 5550 4885
rect 5500 4835 5550 4865
rect 5500 4815 5515 4835
rect 5535 4815 5550 4835
rect 5500 4785 5550 4815
rect 5500 4765 5515 4785
rect 5535 4765 5550 4785
rect 5500 4735 5550 4765
rect 5500 4715 5515 4735
rect 5535 4715 5550 4735
rect 5200 4665 5215 4685
rect 5235 4665 5250 4685
rect 5200 4650 5250 4665
rect 5500 4685 5550 4715
rect 5650 4985 5700 5015
rect 5950 5035 6000 5050
rect 5950 5015 5965 5035
rect 5985 5015 6000 5035
rect 5650 4965 5665 4985
rect 5685 4965 5700 4985
rect 5650 4935 5700 4965
rect 5650 4915 5665 4935
rect 5685 4915 5700 4935
rect 5650 4885 5700 4915
rect 5650 4865 5665 4885
rect 5685 4865 5700 4885
rect 5650 4835 5700 4865
rect 5650 4815 5665 4835
rect 5685 4815 5700 4835
rect 5650 4785 5700 4815
rect 5650 4765 5665 4785
rect 5685 4765 5700 4785
rect 5650 4735 5700 4765
rect 5650 4715 5665 4735
rect 5685 4715 5700 4735
rect 5650 4700 5700 4715
rect 5800 4985 5850 5000
rect 5800 4965 5815 4985
rect 5835 4965 5850 4985
rect 5800 4935 5850 4965
rect 5800 4915 5815 4935
rect 5835 4915 5850 4935
rect 5800 4885 5850 4915
rect 5800 4865 5815 4885
rect 5835 4865 5850 4885
rect 5800 4835 5850 4865
rect 5800 4815 5815 4835
rect 5835 4815 5850 4835
rect 5800 4785 5850 4815
rect 5800 4765 5815 4785
rect 5835 4765 5850 4785
rect 5800 4735 5850 4765
rect 5800 4715 5815 4735
rect 5835 4715 5850 4735
rect 5500 4665 5515 4685
rect 5535 4665 5550 4685
rect 5500 4650 5550 4665
rect 5800 4685 5850 4715
rect 5800 4665 5815 4685
rect 5835 4665 5850 4685
rect 5800 4650 5850 4665
rect 4900 4635 5850 4650
rect 4900 4615 4915 4635
rect 4935 4615 5850 4635
rect 4900 4600 5850 4615
rect 5950 4985 6000 5015
rect 6250 5035 6300 5050
rect 6250 5015 6265 5035
rect 6285 5015 6300 5035
rect 5950 4965 5965 4985
rect 5985 4965 6000 4985
rect 5950 4935 6000 4965
rect 5950 4915 5965 4935
rect 5985 4915 6000 4935
rect 5950 4885 6000 4915
rect 5950 4865 5965 4885
rect 5985 4865 6000 4885
rect 5950 4835 6000 4865
rect 5950 4815 5965 4835
rect 5985 4815 6000 4835
rect 5950 4785 6000 4815
rect 5950 4765 5965 4785
rect 5985 4765 6000 4785
rect 5950 4735 6000 4765
rect 5950 4715 5965 4735
rect 5985 4715 6000 4735
rect 5950 4685 6000 4715
rect 5950 4665 5965 4685
rect 5985 4665 6000 4685
rect 5950 4635 6000 4665
rect 5950 4615 5965 4635
rect 5985 4615 6000 4635
rect 4300 4540 4350 4550
rect 4300 4510 4310 4540
rect 4340 4510 4350 4540
rect 4300 4500 4350 4510
rect 4600 4540 4650 4550
rect 4600 4510 4610 4540
rect 4640 4510 4650 4540
rect 4600 4500 4650 4510
rect 4900 4540 4950 4550
rect 4900 4510 4910 4540
rect 4940 4510 4950 4540
rect 4900 4500 4950 4510
rect 5200 4540 5250 4550
rect 5200 4510 5210 4540
rect 5240 4510 5250 4540
rect 5200 4500 5250 4510
rect 5350 4540 5400 4550
rect 5350 4510 5360 4540
rect 5390 4510 5400 4540
rect 5350 4500 5400 4510
rect 5500 4540 5550 4550
rect 5500 4510 5510 4540
rect 5540 4510 5550 4540
rect 5500 4500 5550 4510
rect 5800 4540 5850 4550
rect 5800 4510 5810 4540
rect 5840 4510 5850 4540
rect 5800 4500 5850 4510
rect 4150 4410 4160 4440
rect 4190 4410 4200 4440
rect 4150 4340 4200 4410
rect 4150 4310 4160 4340
rect 4190 4310 4200 4340
rect 4150 4285 4200 4310
rect 4150 4265 4165 4285
rect 4185 4265 4200 4285
rect 4150 4240 4200 4265
rect 4150 4210 4160 4240
rect 4190 4210 4200 4240
rect 4150 4185 4200 4210
rect 4150 4165 4165 4185
rect 4185 4165 4200 4185
rect 4150 4140 4200 4165
rect 4150 4110 4160 4140
rect 4190 4110 4200 4140
rect 4150 4085 4200 4110
rect 4150 4065 4165 4085
rect 4185 4065 4200 4085
rect 4150 4040 4200 4065
rect 4150 4010 4160 4040
rect 4190 4010 4200 4040
rect 4150 3985 4200 4010
rect 4150 3965 4165 3985
rect 4185 3965 4200 3985
rect -50 3860 -40 3890
rect -10 3860 0 3890
rect -650 3765 -635 3785
rect -615 3765 -600 3785
rect -650 3740 -600 3765
rect -650 3710 -640 3740
rect -610 3710 -600 3740
rect -650 3685 -600 3710
rect -650 3665 -635 3685
rect -615 3665 -600 3685
rect -650 3640 -600 3665
rect -650 3610 -640 3640
rect -610 3610 -600 3640
rect -650 3585 -600 3610
rect -650 3565 -635 3585
rect -615 3565 -600 3585
rect -650 3540 -600 3565
rect -650 3510 -640 3540
rect -610 3510 -600 3540
rect -650 3485 -600 3510
rect -650 3465 -635 3485
rect -615 3465 -600 3485
rect -650 3440 -600 3465
rect -650 3410 -640 3440
rect -610 3410 -600 3440
rect -650 3385 -600 3410
rect -650 3365 -635 3385
rect -615 3365 -600 3385
rect -650 3340 -600 3365
rect -650 3310 -640 3340
rect -610 3310 -600 3340
rect -650 3140 -600 3310
rect -500 3785 -450 3800
rect -500 3765 -485 3785
rect -465 3765 -450 3785
rect -500 3735 -450 3765
rect -500 3715 -485 3735
rect -465 3715 -450 3735
rect -500 3685 -450 3715
rect -500 3665 -485 3685
rect -465 3665 -450 3685
rect -500 3635 -450 3665
rect -500 3615 -485 3635
rect -465 3615 -450 3635
rect -500 3585 -450 3615
rect -500 3565 -485 3585
rect -465 3565 -450 3585
rect -500 3535 -450 3565
rect -500 3515 -485 3535
rect -465 3515 -450 3535
rect -500 3485 -450 3515
rect -500 3465 -485 3485
rect -465 3465 -450 3485
rect -500 3435 -450 3465
rect -500 3415 -485 3435
rect -465 3415 -450 3435
rect -500 3385 -450 3415
rect -350 3785 -300 3800
rect -350 3765 -335 3785
rect -315 3765 -300 3785
rect -350 3735 -300 3765
rect -350 3715 -335 3735
rect -315 3715 -300 3735
rect -350 3685 -300 3715
rect -350 3665 -335 3685
rect -315 3665 -300 3685
rect -350 3635 -300 3665
rect -350 3615 -335 3635
rect -315 3615 -300 3635
rect -350 3585 -300 3615
rect -350 3565 -335 3585
rect -315 3565 -300 3585
rect -350 3535 -300 3565
rect -350 3515 -335 3535
rect -315 3515 -300 3535
rect -350 3485 -300 3515
rect -350 3465 -335 3485
rect -315 3465 -300 3485
rect -350 3435 -300 3465
rect -350 3415 -335 3435
rect -315 3415 -300 3435
rect -350 3400 -300 3415
rect -200 3785 -150 3800
rect -200 3765 -185 3785
rect -165 3765 -150 3785
rect -200 3735 -150 3765
rect -200 3715 -185 3735
rect -165 3715 -150 3735
rect -200 3685 -150 3715
rect -200 3665 -185 3685
rect -165 3665 -150 3685
rect -200 3635 -150 3665
rect -200 3615 -185 3635
rect -165 3615 -150 3635
rect -200 3585 -150 3615
rect -200 3565 -185 3585
rect -165 3565 -150 3585
rect -200 3535 -150 3565
rect -200 3515 -185 3535
rect -165 3515 -150 3535
rect -200 3485 -150 3515
rect -200 3465 -185 3485
rect -165 3465 -150 3485
rect -200 3435 -150 3465
rect -200 3415 -185 3435
rect -165 3415 -150 3435
rect -500 3365 -485 3385
rect -465 3365 -450 3385
rect -500 3350 -450 3365
rect -200 3385 -150 3415
rect -200 3365 -185 3385
rect -165 3365 -150 3385
rect -200 3350 -150 3365
rect -500 3335 -150 3350
rect -500 3315 -485 3335
rect -465 3315 -185 3335
rect -165 3315 -150 3335
rect -500 3300 -150 3315
rect -50 3785 0 3860
rect 4150 3890 4200 3965
rect 4750 4435 4800 4450
rect 4750 4415 4765 4435
rect 4785 4415 4800 4435
rect 4750 4385 4800 4415
rect 4750 4365 4765 4385
rect 4785 4365 4800 4385
rect 4750 4335 4800 4365
rect 4750 4315 4765 4335
rect 4785 4315 4800 4335
rect 4750 4285 4800 4315
rect 4750 4265 4765 4285
rect 4785 4265 4800 4285
rect 4750 4235 4800 4265
rect 4750 4215 4765 4235
rect 4785 4215 4800 4235
rect 4750 4185 4800 4215
rect 4750 4165 4765 4185
rect 4785 4165 4800 4185
rect 4750 4135 4800 4165
rect 4750 4115 4765 4135
rect 4785 4115 4800 4135
rect 4750 4085 4800 4115
rect 4750 4065 4765 4085
rect 4785 4065 4800 4085
rect 4750 4035 4800 4065
rect 4900 4435 5850 4450
rect 4900 4415 4915 4435
rect 4935 4415 5850 4435
rect 4900 4400 5850 4415
rect 4900 4385 4950 4400
rect 4900 4365 4915 4385
rect 4935 4365 4950 4385
rect 4900 4335 4950 4365
rect 5200 4385 5250 4400
rect 5200 4365 5215 4385
rect 5235 4365 5250 4385
rect 4900 4315 4915 4335
rect 4935 4315 4950 4335
rect 4900 4285 4950 4315
rect 4900 4265 4915 4285
rect 4935 4265 4950 4285
rect 4900 4235 4950 4265
rect 4900 4215 4915 4235
rect 4935 4215 4950 4235
rect 4900 4185 4950 4215
rect 4900 4165 4915 4185
rect 4935 4165 4950 4185
rect 4900 4135 4950 4165
rect 4900 4115 4915 4135
rect 4935 4115 4950 4135
rect 4900 4085 4950 4115
rect 4900 4065 4915 4085
rect 4935 4065 4950 4085
rect 4900 4050 4950 4065
rect 5050 4335 5100 4350
rect 5050 4315 5065 4335
rect 5085 4315 5100 4335
rect 5050 4285 5100 4315
rect 5050 4265 5065 4285
rect 5085 4265 5100 4285
rect 5050 4235 5100 4265
rect 5050 4215 5065 4235
rect 5085 4215 5100 4235
rect 5050 4185 5100 4215
rect 5050 4165 5065 4185
rect 5085 4165 5100 4185
rect 5050 4135 5100 4165
rect 5050 4115 5065 4135
rect 5085 4115 5100 4135
rect 5050 4085 5100 4115
rect 5050 4065 5065 4085
rect 5085 4065 5100 4085
rect 4750 4015 4765 4035
rect 4785 4015 4800 4035
rect 4750 4000 4800 4015
rect 5050 4035 5100 4065
rect 5200 4335 5250 4365
rect 5500 4385 5550 4400
rect 5500 4365 5515 4385
rect 5535 4365 5550 4385
rect 5200 4315 5215 4335
rect 5235 4315 5250 4335
rect 5200 4285 5250 4315
rect 5200 4265 5215 4285
rect 5235 4265 5250 4285
rect 5200 4235 5250 4265
rect 5200 4215 5215 4235
rect 5235 4215 5250 4235
rect 5200 4185 5250 4215
rect 5200 4165 5215 4185
rect 5235 4165 5250 4185
rect 5200 4135 5250 4165
rect 5200 4115 5215 4135
rect 5235 4115 5250 4135
rect 5200 4085 5250 4115
rect 5200 4065 5215 4085
rect 5235 4065 5250 4085
rect 5200 4050 5250 4065
rect 5350 4335 5400 4350
rect 5350 4315 5365 4335
rect 5385 4315 5400 4335
rect 5350 4285 5400 4315
rect 5350 4265 5365 4285
rect 5385 4265 5400 4285
rect 5350 4235 5400 4265
rect 5350 4215 5365 4235
rect 5385 4215 5400 4235
rect 5350 4185 5400 4215
rect 5350 4165 5365 4185
rect 5385 4165 5400 4185
rect 5350 4135 5400 4165
rect 5350 4115 5365 4135
rect 5385 4115 5400 4135
rect 5350 4085 5400 4115
rect 5350 4065 5365 4085
rect 5385 4065 5400 4085
rect 5050 4015 5065 4035
rect 5085 4015 5100 4035
rect 5050 4000 5100 4015
rect 5350 4035 5400 4065
rect 5500 4335 5550 4365
rect 5800 4385 5850 4400
rect 5800 4365 5815 4385
rect 5835 4365 5850 4385
rect 5500 4315 5515 4335
rect 5535 4315 5550 4335
rect 5500 4285 5550 4315
rect 5500 4265 5515 4285
rect 5535 4265 5550 4285
rect 5500 4235 5550 4265
rect 5500 4215 5515 4235
rect 5535 4215 5550 4235
rect 5500 4185 5550 4215
rect 5500 4165 5515 4185
rect 5535 4165 5550 4185
rect 5500 4135 5550 4165
rect 5500 4115 5515 4135
rect 5535 4115 5550 4135
rect 5500 4085 5550 4115
rect 5500 4065 5515 4085
rect 5535 4065 5550 4085
rect 5500 4050 5550 4065
rect 5650 4335 5700 4350
rect 5650 4315 5665 4335
rect 5685 4315 5700 4335
rect 5650 4285 5700 4315
rect 5650 4265 5665 4285
rect 5685 4265 5700 4285
rect 5650 4235 5700 4265
rect 5650 4215 5665 4235
rect 5685 4215 5700 4235
rect 5650 4185 5700 4215
rect 5650 4165 5665 4185
rect 5685 4165 5700 4185
rect 5650 4135 5700 4165
rect 5650 4115 5665 4135
rect 5685 4115 5700 4135
rect 5650 4085 5700 4115
rect 5650 4065 5665 4085
rect 5685 4065 5700 4085
rect 5350 4015 5365 4035
rect 5385 4015 5400 4035
rect 5350 4000 5400 4015
rect 5650 4035 5700 4065
rect 5800 4335 5850 4365
rect 5800 4315 5815 4335
rect 5835 4315 5850 4335
rect 5800 4285 5850 4315
rect 5800 4265 5815 4285
rect 5835 4265 5850 4285
rect 5800 4235 5850 4265
rect 5800 4215 5815 4235
rect 5835 4215 5850 4235
rect 5800 4185 5850 4215
rect 5800 4165 5815 4185
rect 5835 4165 5850 4185
rect 5800 4135 5850 4165
rect 5800 4115 5815 4135
rect 5835 4115 5850 4135
rect 5800 4085 5850 4115
rect 5800 4065 5815 4085
rect 5835 4065 5850 4085
rect 5800 4050 5850 4065
rect 5950 4435 6000 4615
rect 6100 4985 6150 5000
rect 6100 4965 6115 4985
rect 6135 4965 6150 4985
rect 6100 4935 6150 4965
rect 6100 4915 6115 4935
rect 6135 4915 6150 4935
rect 6100 4885 6150 4915
rect 6100 4865 6115 4885
rect 6135 4865 6150 4885
rect 6100 4835 6150 4865
rect 6100 4815 6115 4835
rect 6135 4815 6150 4835
rect 6100 4785 6150 4815
rect 6100 4765 6115 4785
rect 6135 4765 6150 4785
rect 6100 4735 6150 4765
rect 6100 4715 6115 4735
rect 6135 4715 6150 4735
rect 6100 4685 6150 4715
rect 6250 4985 6300 5015
rect 6550 5035 6600 5050
rect 6550 5015 6565 5035
rect 6585 5015 6600 5035
rect 6250 4965 6265 4985
rect 6285 4965 6300 4985
rect 6250 4935 6300 4965
rect 6250 4915 6265 4935
rect 6285 4915 6300 4935
rect 6250 4885 6300 4915
rect 6250 4865 6265 4885
rect 6285 4865 6300 4885
rect 6250 4835 6300 4865
rect 6250 4815 6265 4835
rect 6285 4815 6300 4835
rect 6250 4785 6300 4815
rect 6250 4765 6265 4785
rect 6285 4765 6300 4785
rect 6250 4735 6300 4765
rect 6250 4715 6265 4735
rect 6285 4715 6300 4735
rect 6250 4700 6300 4715
rect 6400 4985 6450 5000
rect 6400 4965 6415 4985
rect 6435 4965 6450 4985
rect 6400 4935 6450 4965
rect 6400 4915 6415 4935
rect 6435 4915 6450 4935
rect 6400 4885 6450 4915
rect 6400 4865 6415 4885
rect 6435 4865 6450 4885
rect 6400 4835 6450 4865
rect 6400 4815 6415 4835
rect 6435 4815 6450 4835
rect 6400 4785 6450 4815
rect 6400 4765 6415 4785
rect 6435 4765 6450 4785
rect 6400 4735 6450 4765
rect 6400 4715 6415 4735
rect 6435 4715 6450 4735
rect 6100 4665 6115 4685
rect 6135 4665 6150 4685
rect 6100 4650 6150 4665
rect 6400 4685 6450 4715
rect 6400 4665 6415 4685
rect 6435 4665 6450 4685
rect 6400 4650 6450 4665
rect 6100 4635 6450 4650
rect 6100 4615 6115 4635
rect 6135 4615 6415 4635
rect 6435 4615 6450 4635
rect 6100 4600 6450 4615
rect 6550 4985 6600 5015
rect 6850 5035 6900 5050
rect 6850 5015 6865 5035
rect 6885 5015 6900 5035
rect 6550 4965 6565 4985
rect 6585 4965 6600 4985
rect 6550 4935 6600 4965
rect 6550 4915 6565 4935
rect 6585 4915 6600 4935
rect 6550 4885 6600 4915
rect 6550 4865 6565 4885
rect 6585 4865 6600 4885
rect 6550 4835 6600 4865
rect 6550 4815 6565 4835
rect 6585 4815 6600 4835
rect 6550 4785 6600 4815
rect 6550 4765 6565 4785
rect 6585 4765 6600 4785
rect 6550 4735 6600 4765
rect 6550 4715 6565 4735
rect 6585 4715 6600 4735
rect 6550 4685 6600 4715
rect 6550 4665 6565 4685
rect 6585 4665 6600 4685
rect 6550 4635 6600 4665
rect 6550 4615 6565 4635
rect 6585 4615 6600 4635
rect 6100 4540 6150 4550
rect 6100 4510 6110 4540
rect 6140 4510 6150 4540
rect 6100 4500 6150 4510
rect 6250 4540 6300 4600
rect 6250 4510 6260 4540
rect 6290 4510 6300 4540
rect 6250 4450 6300 4510
rect 6400 4540 6450 4550
rect 6400 4510 6410 4540
rect 6440 4510 6450 4540
rect 6400 4500 6450 4510
rect 5950 4415 5965 4435
rect 5985 4415 6000 4435
rect 5950 4385 6000 4415
rect 5950 4365 5965 4385
rect 5985 4365 6000 4385
rect 5950 4335 6000 4365
rect 5950 4315 5965 4335
rect 5985 4315 6000 4335
rect 5950 4285 6000 4315
rect 5950 4265 5965 4285
rect 5985 4265 6000 4285
rect 5950 4235 6000 4265
rect 5950 4215 5965 4235
rect 5985 4215 6000 4235
rect 5950 4185 6000 4215
rect 5950 4165 5965 4185
rect 5985 4165 6000 4185
rect 5950 4135 6000 4165
rect 5950 4115 5965 4135
rect 5985 4115 6000 4135
rect 5950 4085 6000 4115
rect 5950 4065 5965 4085
rect 5985 4065 6000 4085
rect 5650 4015 5665 4035
rect 5685 4015 5700 4035
rect 5650 4000 5700 4015
rect 5950 4035 6000 4065
rect 6100 4435 6450 4450
rect 6100 4415 6115 4435
rect 6135 4415 6415 4435
rect 6435 4415 6450 4435
rect 6100 4400 6450 4415
rect 6100 4385 6150 4400
rect 6100 4365 6115 4385
rect 6135 4365 6150 4385
rect 6100 4335 6150 4365
rect 6400 4385 6450 4400
rect 6400 4365 6415 4385
rect 6435 4365 6450 4385
rect 6100 4315 6115 4335
rect 6135 4315 6150 4335
rect 6100 4285 6150 4315
rect 6100 4265 6115 4285
rect 6135 4265 6150 4285
rect 6100 4235 6150 4265
rect 6100 4215 6115 4235
rect 6135 4215 6150 4235
rect 6100 4185 6150 4215
rect 6100 4165 6115 4185
rect 6135 4165 6150 4185
rect 6100 4135 6150 4165
rect 6100 4115 6115 4135
rect 6135 4115 6150 4135
rect 6100 4085 6150 4115
rect 6100 4065 6115 4085
rect 6135 4065 6150 4085
rect 6100 4050 6150 4065
rect 6250 4335 6300 4350
rect 6250 4315 6265 4335
rect 6285 4315 6300 4335
rect 6250 4285 6300 4315
rect 6250 4265 6265 4285
rect 6285 4265 6300 4285
rect 6250 4235 6300 4265
rect 6250 4215 6265 4235
rect 6285 4215 6300 4235
rect 6250 4185 6300 4215
rect 6250 4165 6265 4185
rect 6285 4165 6300 4185
rect 6250 4135 6300 4165
rect 6250 4115 6265 4135
rect 6285 4115 6300 4135
rect 6250 4085 6300 4115
rect 6250 4065 6265 4085
rect 6285 4065 6300 4085
rect 5950 4015 5965 4035
rect 5985 4015 6000 4035
rect 5950 4000 6000 4015
rect 6250 4035 6300 4065
rect 6400 4335 6450 4365
rect 6400 4315 6415 4335
rect 6435 4315 6450 4335
rect 6400 4285 6450 4315
rect 6400 4265 6415 4285
rect 6435 4265 6450 4285
rect 6400 4235 6450 4265
rect 6400 4215 6415 4235
rect 6435 4215 6450 4235
rect 6400 4185 6450 4215
rect 6400 4165 6415 4185
rect 6435 4165 6450 4185
rect 6400 4135 6450 4165
rect 6400 4115 6415 4135
rect 6435 4115 6450 4135
rect 6400 4085 6450 4115
rect 6400 4065 6415 4085
rect 6435 4065 6450 4085
rect 6400 4050 6450 4065
rect 6550 4435 6600 4615
rect 6700 4985 6750 5000
rect 6700 4965 6715 4985
rect 6735 4965 6750 4985
rect 6700 4935 6750 4965
rect 6700 4915 6715 4935
rect 6735 4915 6750 4935
rect 6700 4885 6750 4915
rect 6700 4865 6715 4885
rect 6735 4865 6750 4885
rect 6700 4835 6750 4865
rect 6700 4815 6715 4835
rect 6735 4815 6750 4835
rect 6700 4785 6750 4815
rect 6700 4765 6715 4785
rect 6735 4765 6750 4785
rect 6700 4735 6750 4765
rect 6700 4715 6715 4735
rect 6735 4715 6750 4735
rect 6700 4685 6750 4715
rect 6850 4985 6900 5015
rect 7150 5035 7200 5050
rect 7150 5015 7165 5035
rect 7185 5015 7200 5035
rect 6850 4965 6865 4985
rect 6885 4965 6900 4985
rect 6850 4935 6900 4965
rect 6850 4915 6865 4935
rect 6885 4915 6900 4935
rect 6850 4885 6900 4915
rect 6850 4865 6865 4885
rect 6885 4865 6900 4885
rect 6850 4835 6900 4865
rect 6850 4815 6865 4835
rect 6885 4815 6900 4835
rect 6850 4785 6900 4815
rect 6850 4765 6865 4785
rect 6885 4765 6900 4785
rect 6850 4735 6900 4765
rect 6850 4715 6865 4735
rect 6885 4715 6900 4735
rect 6850 4700 6900 4715
rect 7000 4985 7050 5000
rect 7000 4965 7015 4985
rect 7035 4965 7050 4985
rect 7000 4935 7050 4965
rect 7000 4915 7015 4935
rect 7035 4915 7050 4935
rect 7000 4885 7050 4915
rect 7000 4865 7015 4885
rect 7035 4865 7050 4885
rect 7000 4835 7050 4865
rect 7000 4815 7015 4835
rect 7035 4815 7050 4835
rect 7000 4785 7050 4815
rect 7000 4765 7015 4785
rect 7035 4765 7050 4785
rect 7000 4735 7050 4765
rect 7000 4715 7015 4735
rect 7035 4715 7050 4735
rect 6700 4665 6715 4685
rect 6735 4665 6750 4685
rect 6700 4650 6750 4665
rect 7000 4685 7050 4715
rect 7150 4985 7200 5015
rect 7450 5035 7500 5050
rect 7450 5015 7465 5035
rect 7485 5015 7500 5035
rect 7150 4965 7165 4985
rect 7185 4965 7200 4985
rect 7150 4935 7200 4965
rect 7150 4915 7165 4935
rect 7185 4915 7200 4935
rect 7150 4885 7200 4915
rect 7150 4865 7165 4885
rect 7185 4865 7200 4885
rect 7150 4835 7200 4865
rect 7150 4815 7165 4835
rect 7185 4815 7200 4835
rect 7150 4785 7200 4815
rect 7150 4765 7165 4785
rect 7185 4765 7200 4785
rect 7150 4735 7200 4765
rect 7150 4715 7165 4735
rect 7185 4715 7200 4735
rect 7150 4700 7200 4715
rect 7300 4985 7350 5000
rect 7300 4965 7315 4985
rect 7335 4965 7350 4985
rect 7300 4935 7350 4965
rect 7300 4915 7315 4935
rect 7335 4915 7350 4935
rect 7300 4885 7350 4915
rect 7300 4865 7315 4885
rect 7335 4865 7350 4885
rect 7300 4835 7350 4865
rect 7300 4815 7315 4835
rect 7335 4815 7350 4835
rect 7300 4785 7350 4815
rect 7300 4765 7315 4785
rect 7335 4765 7350 4785
rect 7300 4735 7350 4765
rect 7300 4715 7315 4735
rect 7335 4715 7350 4735
rect 7000 4665 7015 4685
rect 7035 4665 7050 4685
rect 7000 4650 7050 4665
rect 7300 4685 7350 4715
rect 7450 4985 7500 5015
rect 7750 5035 7800 5050
rect 7750 5015 7765 5035
rect 7785 5015 7800 5035
rect 7450 4965 7465 4985
rect 7485 4965 7500 4985
rect 7450 4935 7500 4965
rect 7450 4915 7465 4935
rect 7485 4915 7500 4935
rect 7450 4885 7500 4915
rect 7450 4865 7465 4885
rect 7485 4865 7500 4885
rect 7450 4835 7500 4865
rect 7450 4815 7465 4835
rect 7485 4815 7500 4835
rect 7450 4785 7500 4815
rect 7450 4765 7465 4785
rect 7485 4765 7500 4785
rect 7450 4735 7500 4765
rect 7450 4715 7465 4735
rect 7485 4715 7500 4735
rect 7450 4700 7500 4715
rect 7600 4985 7650 5000
rect 7600 4965 7615 4985
rect 7635 4965 7650 4985
rect 7600 4935 7650 4965
rect 7600 4915 7615 4935
rect 7635 4915 7650 4935
rect 7600 4885 7650 4915
rect 7600 4865 7615 4885
rect 7635 4865 7650 4885
rect 7600 4835 7650 4865
rect 7600 4815 7615 4835
rect 7635 4815 7650 4835
rect 7600 4785 7650 4815
rect 7600 4765 7615 4785
rect 7635 4765 7650 4785
rect 7600 4735 7650 4765
rect 7600 4715 7615 4735
rect 7635 4715 7650 4735
rect 7300 4665 7315 4685
rect 7335 4665 7350 4685
rect 7300 4650 7350 4665
rect 7600 4685 7650 4715
rect 7600 4665 7615 4685
rect 7635 4665 7650 4685
rect 7600 4650 7650 4665
rect 6700 4635 7650 4650
rect 6700 4615 7615 4635
rect 7635 4615 7650 4635
rect 6700 4600 7650 4615
rect 7750 4985 7800 5015
rect 7750 4965 7765 4985
rect 7785 4965 7800 4985
rect 7750 4935 7800 4965
rect 7750 4915 7765 4935
rect 7785 4915 7800 4935
rect 7750 4885 7800 4915
rect 7750 4865 7765 4885
rect 7785 4865 7800 4885
rect 7750 4835 7800 4865
rect 7750 4815 7765 4835
rect 7785 4815 7800 4835
rect 7750 4785 7800 4815
rect 7750 4765 7765 4785
rect 7785 4765 7800 4785
rect 7750 4735 7800 4765
rect 7750 4715 7765 4735
rect 7785 4715 7800 4735
rect 7750 4685 7800 4715
rect 7750 4665 7765 4685
rect 7785 4665 7800 4685
rect 7750 4635 7800 4665
rect 7750 4615 7765 4635
rect 7785 4615 7800 4635
rect 7750 4600 7800 4615
rect 8350 5085 8400 5160
rect 8650 5190 8700 5200
rect 8650 5160 8660 5190
rect 8690 5160 8700 5190
rect 8350 5065 8365 5085
rect 8385 5065 8400 5085
rect 8350 5040 8400 5065
rect 8350 5010 8360 5040
rect 8390 5010 8400 5040
rect 8350 4985 8400 5010
rect 8350 4965 8365 4985
rect 8385 4965 8400 4985
rect 8350 4940 8400 4965
rect 8350 4910 8360 4940
rect 8390 4910 8400 4940
rect 8350 4885 8400 4910
rect 8350 4865 8365 4885
rect 8385 4865 8400 4885
rect 8350 4840 8400 4865
rect 8350 4810 8360 4840
rect 8390 4810 8400 4840
rect 8350 4785 8400 4810
rect 8350 4765 8365 4785
rect 8385 4765 8400 4785
rect 8350 4740 8400 4765
rect 8350 4710 8360 4740
rect 8390 4710 8400 4740
rect 8350 4685 8400 4710
rect 8350 4665 8365 4685
rect 8385 4665 8400 4685
rect 8350 4640 8400 4665
rect 8350 4610 8360 4640
rect 8390 4610 8400 4640
rect 6700 4540 6750 4550
rect 6700 4510 6710 4540
rect 6740 4510 6750 4540
rect 6700 4500 6750 4510
rect 7000 4540 7050 4550
rect 7000 4510 7010 4540
rect 7040 4510 7050 4540
rect 7000 4500 7050 4510
rect 7150 4540 7200 4550
rect 7150 4510 7160 4540
rect 7190 4510 7200 4540
rect 7150 4500 7200 4510
rect 7300 4540 7350 4550
rect 7300 4510 7310 4540
rect 7340 4510 7350 4540
rect 7300 4500 7350 4510
rect 7600 4540 7650 4550
rect 7600 4510 7610 4540
rect 7640 4510 7650 4540
rect 7600 4500 7650 4510
rect 7900 4540 7950 4550
rect 7900 4510 7910 4540
rect 7940 4510 7950 4540
rect 7900 4500 7950 4510
rect 8200 4540 8250 4550
rect 8200 4510 8210 4540
rect 8240 4510 8250 4540
rect 8200 4500 8250 4510
rect 6550 4415 6565 4435
rect 6585 4415 6600 4435
rect 6550 4385 6600 4415
rect 6550 4365 6565 4385
rect 6585 4365 6600 4385
rect 6550 4335 6600 4365
rect 6550 4315 6565 4335
rect 6585 4315 6600 4335
rect 6550 4285 6600 4315
rect 6550 4265 6565 4285
rect 6585 4265 6600 4285
rect 6550 4235 6600 4265
rect 6550 4215 6565 4235
rect 6585 4215 6600 4235
rect 6550 4185 6600 4215
rect 6550 4165 6565 4185
rect 6585 4165 6600 4185
rect 6550 4135 6600 4165
rect 6550 4115 6565 4135
rect 6585 4115 6600 4135
rect 6550 4085 6600 4115
rect 6550 4065 6565 4085
rect 6585 4065 6600 4085
rect 6250 4015 6265 4035
rect 6285 4015 6300 4035
rect 6250 4000 6300 4015
rect 6550 4035 6600 4065
rect 6700 4435 7650 4450
rect 6700 4415 7615 4435
rect 7635 4415 7650 4435
rect 6700 4400 7650 4415
rect 6700 4385 6750 4400
rect 6700 4365 6715 4385
rect 6735 4365 6750 4385
rect 6700 4335 6750 4365
rect 7000 4385 7050 4400
rect 7000 4365 7015 4385
rect 7035 4365 7050 4385
rect 6700 4315 6715 4335
rect 6735 4315 6750 4335
rect 6700 4285 6750 4315
rect 6700 4265 6715 4285
rect 6735 4265 6750 4285
rect 6700 4235 6750 4265
rect 6700 4215 6715 4235
rect 6735 4215 6750 4235
rect 6700 4185 6750 4215
rect 6700 4165 6715 4185
rect 6735 4165 6750 4185
rect 6700 4135 6750 4165
rect 6700 4115 6715 4135
rect 6735 4115 6750 4135
rect 6700 4085 6750 4115
rect 6700 4065 6715 4085
rect 6735 4065 6750 4085
rect 6700 4050 6750 4065
rect 6850 4335 6900 4350
rect 6850 4315 6865 4335
rect 6885 4315 6900 4335
rect 6850 4285 6900 4315
rect 6850 4265 6865 4285
rect 6885 4265 6900 4285
rect 6850 4235 6900 4265
rect 6850 4215 6865 4235
rect 6885 4215 6900 4235
rect 6850 4185 6900 4215
rect 6850 4165 6865 4185
rect 6885 4165 6900 4185
rect 6850 4135 6900 4165
rect 6850 4115 6865 4135
rect 6885 4115 6900 4135
rect 6850 4085 6900 4115
rect 6850 4065 6865 4085
rect 6885 4065 6900 4085
rect 6550 4015 6565 4035
rect 6585 4015 6600 4035
rect 6550 4000 6600 4015
rect 6850 4035 6900 4065
rect 7000 4335 7050 4365
rect 7300 4385 7350 4400
rect 7300 4365 7315 4385
rect 7335 4365 7350 4385
rect 7000 4315 7015 4335
rect 7035 4315 7050 4335
rect 7000 4285 7050 4315
rect 7000 4265 7015 4285
rect 7035 4265 7050 4285
rect 7000 4235 7050 4265
rect 7000 4215 7015 4235
rect 7035 4215 7050 4235
rect 7000 4185 7050 4215
rect 7000 4165 7015 4185
rect 7035 4165 7050 4185
rect 7000 4135 7050 4165
rect 7000 4115 7015 4135
rect 7035 4115 7050 4135
rect 7000 4085 7050 4115
rect 7000 4065 7015 4085
rect 7035 4065 7050 4085
rect 7000 4050 7050 4065
rect 7150 4335 7200 4350
rect 7150 4315 7165 4335
rect 7185 4315 7200 4335
rect 7150 4285 7200 4315
rect 7150 4265 7165 4285
rect 7185 4265 7200 4285
rect 7150 4235 7200 4265
rect 7150 4215 7165 4235
rect 7185 4215 7200 4235
rect 7150 4185 7200 4215
rect 7150 4165 7165 4185
rect 7185 4165 7200 4185
rect 7150 4135 7200 4165
rect 7150 4115 7165 4135
rect 7185 4115 7200 4135
rect 7150 4085 7200 4115
rect 7150 4065 7165 4085
rect 7185 4065 7200 4085
rect 6850 4015 6865 4035
rect 6885 4015 6900 4035
rect 6850 4000 6900 4015
rect 7150 4035 7200 4065
rect 7300 4335 7350 4365
rect 7600 4385 7650 4400
rect 7600 4365 7615 4385
rect 7635 4365 7650 4385
rect 7300 4315 7315 4335
rect 7335 4315 7350 4335
rect 7300 4285 7350 4315
rect 7300 4265 7315 4285
rect 7335 4265 7350 4285
rect 7300 4235 7350 4265
rect 7300 4215 7315 4235
rect 7335 4215 7350 4235
rect 7300 4185 7350 4215
rect 7300 4165 7315 4185
rect 7335 4165 7350 4185
rect 7300 4135 7350 4165
rect 7300 4115 7315 4135
rect 7335 4115 7350 4135
rect 7300 4085 7350 4115
rect 7300 4065 7315 4085
rect 7335 4065 7350 4085
rect 7300 4050 7350 4065
rect 7450 4335 7500 4350
rect 7450 4315 7465 4335
rect 7485 4315 7500 4335
rect 7450 4285 7500 4315
rect 7450 4265 7465 4285
rect 7485 4265 7500 4285
rect 7450 4235 7500 4265
rect 7450 4215 7465 4235
rect 7485 4215 7500 4235
rect 7450 4185 7500 4215
rect 7450 4165 7465 4185
rect 7485 4165 7500 4185
rect 7450 4135 7500 4165
rect 7450 4115 7465 4135
rect 7485 4115 7500 4135
rect 7450 4085 7500 4115
rect 7450 4065 7465 4085
rect 7485 4065 7500 4085
rect 7150 4015 7165 4035
rect 7185 4015 7200 4035
rect 7150 4000 7200 4015
rect 7450 4035 7500 4065
rect 7600 4335 7650 4365
rect 7600 4315 7615 4335
rect 7635 4315 7650 4335
rect 7600 4285 7650 4315
rect 7600 4265 7615 4285
rect 7635 4265 7650 4285
rect 7600 4235 7650 4265
rect 7600 4215 7615 4235
rect 7635 4215 7650 4235
rect 7600 4185 7650 4215
rect 7600 4165 7615 4185
rect 7635 4165 7650 4185
rect 7600 4135 7650 4165
rect 7600 4115 7615 4135
rect 7635 4115 7650 4135
rect 7600 4085 7650 4115
rect 7600 4065 7615 4085
rect 7635 4065 7650 4085
rect 7600 4050 7650 4065
rect 7750 4435 7800 4450
rect 7750 4415 7765 4435
rect 7785 4415 7800 4435
rect 7750 4385 7800 4415
rect 7750 4365 7765 4385
rect 7785 4365 7800 4385
rect 7750 4335 7800 4365
rect 7750 4315 7765 4335
rect 7785 4315 7800 4335
rect 7750 4285 7800 4315
rect 7750 4265 7765 4285
rect 7785 4265 7800 4285
rect 7750 4235 7800 4265
rect 7750 4215 7765 4235
rect 7785 4215 7800 4235
rect 7750 4185 7800 4215
rect 7750 4165 7765 4185
rect 7785 4165 7800 4185
rect 7750 4135 7800 4165
rect 7750 4115 7765 4135
rect 7785 4115 7800 4135
rect 7750 4085 7800 4115
rect 7750 4065 7765 4085
rect 7785 4065 7800 4085
rect 7450 4015 7465 4035
rect 7485 4015 7500 4035
rect 7450 4000 7500 4015
rect 7750 4035 7800 4065
rect 7750 4015 7765 4035
rect 7785 4015 7800 4035
rect 7750 4000 7800 4015
rect 4750 3985 7800 4000
rect 4750 3965 4765 3985
rect 4785 3965 5065 3985
rect 5085 3965 5365 3985
rect 5385 3965 5665 3985
rect 5685 3965 5965 3985
rect 5985 3965 6265 3985
rect 6285 3965 6565 3985
rect 6585 3965 6865 3985
rect 6885 3965 7165 3985
rect 7185 3965 7465 3985
rect 7485 3965 7765 3985
rect 7785 3965 7800 3985
rect 4750 3950 7800 3965
rect 8350 4440 8400 4610
rect 8500 5085 8550 5100
rect 8500 5065 8515 5085
rect 8535 5065 8550 5085
rect 8500 5035 8550 5065
rect 8500 5015 8515 5035
rect 8535 5015 8550 5035
rect 8500 4985 8550 5015
rect 8500 4965 8515 4985
rect 8535 4965 8550 4985
rect 8500 4935 8550 4965
rect 8500 4915 8515 4935
rect 8535 4915 8550 4935
rect 8500 4885 8550 4915
rect 8500 4865 8515 4885
rect 8535 4865 8550 4885
rect 8500 4835 8550 4865
rect 8500 4815 8515 4835
rect 8535 4815 8550 4835
rect 8500 4785 8550 4815
rect 8500 4765 8515 4785
rect 8535 4765 8550 4785
rect 8500 4735 8550 4765
rect 8500 4715 8515 4735
rect 8535 4715 8550 4735
rect 8500 4685 8550 4715
rect 8500 4665 8515 4685
rect 8535 4665 8550 4685
rect 8500 4635 8550 4665
rect 8500 4615 8515 4635
rect 8535 4615 8550 4635
rect 8500 4600 8550 4615
rect 8650 5085 8700 5160
rect 8950 5190 9000 5200
rect 8950 5160 8960 5190
rect 8990 5160 9000 5190
rect 8650 5065 8665 5085
rect 8685 5065 8700 5085
rect 8650 5040 8700 5065
rect 8650 5010 8660 5040
rect 8690 5010 8700 5040
rect 8650 4985 8700 5010
rect 8650 4965 8665 4985
rect 8685 4965 8700 4985
rect 8650 4940 8700 4965
rect 8650 4910 8660 4940
rect 8690 4910 8700 4940
rect 8650 4885 8700 4910
rect 8650 4865 8665 4885
rect 8685 4865 8700 4885
rect 8650 4840 8700 4865
rect 8650 4810 8660 4840
rect 8690 4810 8700 4840
rect 8650 4785 8700 4810
rect 8650 4765 8665 4785
rect 8685 4765 8700 4785
rect 8650 4740 8700 4765
rect 8650 4710 8660 4740
rect 8690 4710 8700 4740
rect 8650 4685 8700 4710
rect 8650 4665 8665 4685
rect 8685 4665 8700 4685
rect 8650 4640 8700 4665
rect 8650 4610 8660 4640
rect 8690 4610 8700 4640
rect 8500 4540 8550 4550
rect 8500 4510 8510 4540
rect 8540 4510 8550 4540
rect 8500 4500 8550 4510
rect 8350 4410 8360 4440
rect 8390 4410 8400 4440
rect 8350 4385 8400 4410
rect 8350 4365 8365 4385
rect 8385 4365 8400 4385
rect 8350 4340 8400 4365
rect 8350 4310 8360 4340
rect 8390 4310 8400 4340
rect 8350 4285 8400 4310
rect 8350 4265 8365 4285
rect 8385 4265 8400 4285
rect 8350 4240 8400 4265
rect 8350 4210 8360 4240
rect 8390 4210 8400 4240
rect 8350 4185 8400 4210
rect 8350 4165 8365 4185
rect 8385 4165 8400 4185
rect 8350 4140 8400 4165
rect 8350 4110 8360 4140
rect 8390 4110 8400 4140
rect 8350 4085 8400 4110
rect 8350 4065 8365 4085
rect 8385 4065 8400 4085
rect 8350 4040 8400 4065
rect 8350 4010 8360 4040
rect 8390 4010 8400 4040
rect 8350 3985 8400 4010
rect 8350 3965 8365 3985
rect 8385 3965 8400 3985
rect 4150 3860 4160 3890
rect 4190 3860 4200 3890
rect -50 3765 -35 3785
rect -15 3765 0 3785
rect -50 3735 0 3765
rect -50 3715 -35 3735
rect -15 3715 0 3735
rect -50 3685 0 3715
rect -50 3665 -35 3685
rect -15 3665 0 3685
rect -50 3635 0 3665
rect -50 3615 -35 3635
rect -15 3615 0 3635
rect -50 3585 0 3615
rect -50 3565 -35 3585
rect -15 3565 0 3585
rect -50 3535 0 3565
rect -50 3515 -35 3535
rect -15 3515 0 3535
rect -50 3485 0 3515
rect -50 3465 -35 3485
rect -15 3465 0 3485
rect -50 3435 0 3465
rect -50 3415 -35 3435
rect -15 3415 0 3435
rect -500 3240 -450 3250
rect -500 3210 -490 3240
rect -460 3210 -450 3240
rect -500 3200 -450 3210
rect -350 3240 -300 3300
rect -350 3210 -340 3240
rect -310 3210 -300 3240
rect -350 3150 -300 3210
rect -200 3240 -150 3250
rect -200 3210 -190 3240
rect -160 3210 -150 3240
rect -200 3200 -150 3210
rect -650 3110 -640 3140
rect -610 3110 -600 3140
rect -650 3085 -600 3110
rect -650 3065 -635 3085
rect -615 3065 -600 3085
rect -650 3040 -600 3065
rect -650 3010 -640 3040
rect -610 3010 -600 3040
rect -650 2985 -600 3010
rect -650 2965 -635 2985
rect -615 2965 -600 2985
rect -650 2940 -600 2965
rect -650 2910 -640 2940
rect -610 2910 -600 2940
rect -650 2885 -600 2910
rect -650 2865 -635 2885
rect -615 2865 -600 2885
rect -650 2840 -600 2865
rect -650 2810 -640 2840
rect -610 2810 -600 2840
rect -650 2785 -600 2810
rect -650 2765 -635 2785
rect -615 2765 -600 2785
rect -650 2740 -600 2765
rect -650 2710 -640 2740
rect -610 2710 -600 2740
rect -650 2685 -600 2710
rect -650 2665 -635 2685
rect -615 2665 -600 2685
rect -650 2590 -600 2665
rect -500 3135 -150 3150
rect -500 3115 -485 3135
rect -465 3115 -185 3135
rect -165 3115 -150 3135
rect -500 3100 -150 3115
rect -500 3085 -450 3100
rect -500 3065 -485 3085
rect -465 3065 -450 3085
rect -500 3035 -450 3065
rect -200 3085 -150 3100
rect -200 3065 -185 3085
rect -165 3065 -150 3085
rect -500 3015 -485 3035
rect -465 3015 -450 3035
rect -500 2985 -450 3015
rect -500 2965 -485 2985
rect -465 2965 -450 2985
rect -500 2935 -450 2965
rect -500 2915 -485 2935
rect -465 2915 -450 2935
rect -500 2885 -450 2915
rect -500 2865 -485 2885
rect -465 2865 -450 2885
rect -500 2835 -450 2865
rect -500 2815 -485 2835
rect -465 2815 -450 2835
rect -500 2785 -450 2815
rect -500 2765 -485 2785
rect -465 2765 -450 2785
rect -500 2735 -450 2765
rect -500 2715 -485 2735
rect -465 2715 -450 2735
rect -500 2685 -450 2715
rect -500 2665 -485 2685
rect -465 2665 -450 2685
rect -500 2650 -450 2665
rect -350 3035 -300 3050
rect -350 3015 -335 3035
rect -315 3015 -300 3035
rect -350 2985 -300 3015
rect -350 2965 -335 2985
rect -315 2965 -300 2985
rect -350 2935 -300 2965
rect -350 2915 -335 2935
rect -315 2915 -300 2935
rect -350 2885 -300 2915
rect -350 2865 -335 2885
rect -315 2865 -300 2885
rect -350 2835 -300 2865
rect -350 2815 -335 2835
rect -315 2815 -300 2835
rect -350 2785 -300 2815
rect -350 2765 -335 2785
rect -315 2765 -300 2785
rect -350 2735 -300 2765
rect -350 2715 -335 2735
rect -315 2715 -300 2735
rect -350 2685 -300 2715
rect -350 2665 -335 2685
rect -315 2665 -300 2685
rect -350 2650 -300 2665
rect -200 3035 -150 3065
rect -200 3015 -185 3035
rect -165 3015 -150 3035
rect -200 2985 -150 3015
rect -200 2965 -185 2985
rect -165 2965 -150 2985
rect -200 2935 -150 2965
rect -200 2915 -185 2935
rect -165 2915 -150 2935
rect -200 2885 -150 2915
rect -200 2865 -185 2885
rect -165 2865 -150 2885
rect -200 2835 -150 2865
rect -200 2815 -185 2835
rect -165 2815 -150 2835
rect -200 2785 -150 2815
rect -200 2765 -185 2785
rect -165 2765 -150 2785
rect -200 2735 -150 2765
rect -200 2715 -185 2735
rect -165 2715 -150 2735
rect -200 2685 -150 2715
rect -200 2665 -185 2685
rect -165 2665 -150 2685
rect -200 2650 -150 2665
rect -50 3140 0 3415
rect 550 3785 3600 3800
rect 550 3765 565 3785
rect 585 3765 865 3785
rect 885 3765 1165 3785
rect 1185 3765 1465 3785
rect 1485 3765 1765 3785
rect 1785 3765 2065 3785
rect 2085 3765 2365 3785
rect 2385 3765 2665 3785
rect 2685 3765 2965 3785
rect 2985 3765 3265 3785
rect 3285 3765 3565 3785
rect 3585 3765 3600 3785
rect 550 3750 3600 3765
rect 550 3735 600 3750
rect 550 3715 565 3735
rect 585 3715 600 3735
rect 550 3685 600 3715
rect 850 3735 900 3750
rect 850 3715 865 3735
rect 885 3715 900 3735
rect 550 3665 565 3685
rect 585 3665 600 3685
rect 550 3635 600 3665
rect 550 3615 565 3635
rect 585 3615 600 3635
rect 550 3585 600 3615
rect 550 3565 565 3585
rect 585 3565 600 3585
rect 550 3535 600 3565
rect 550 3515 565 3535
rect 585 3515 600 3535
rect 550 3485 600 3515
rect 550 3465 565 3485
rect 585 3465 600 3485
rect 550 3435 600 3465
rect 550 3415 565 3435
rect 585 3415 600 3435
rect 550 3385 600 3415
rect 550 3365 565 3385
rect 585 3365 600 3385
rect 550 3335 600 3365
rect 550 3315 565 3335
rect 585 3315 600 3335
rect 100 3240 150 3250
rect 100 3210 110 3240
rect 140 3210 150 3240
rect 100 3200 150 3210
rect 400 3240 450 3250
rect 400 3210 410 3240
rect 440 3210 450 3240
rect 400 3200 450 3210
rect -50 3110 -40 3140
rect -10 3110 0 3140
rect -50 3040 0 3110
rect -50 3010 -40 3040
rect -10 3010 0 3040
rect -50 2985 0 3010
rect -50 2965 -35 2985
rect -15 2965 0 2985
rect -50 2940 0 2965
rect -50 2910 -40 2940
rect -10 2910 0 2940
rect -50 2885 0 2910
rect -50 2865 -35 2885
rect -15 2865 0 2885
rect -50 2840 0 2865
rect -50 2810 -40 2840
rect -10 2810 0 2840
rect -50 2785 0 2810
rect -50 2765 -35 2785
rect -15 2765 0 2785
rect -50 2740 0 2765
rect -50 2710 -40 2740
rect -10 2710 0 2740
rect -50 2685 0 2710
rect -50 2665 -35 2685
rect -15 2665 0 2685
rect -650 2560 -640 2590
rect -610 2560 -600 2590
rect -650 2550 -600 2560
rect -50 2590 0 2665
rect 550 3135 600 3315
rect 700 3685 750 3700
rect 700 3665 715 3685
rect 735 3665 750 3685
rect 700 3635 750 3665
rect 700 3615 715 3635
rect 735 3615 750 3635
rect 700 3585 750 3615
rect 700 3565 715 3585
rect 735 3565 750 3585
rect 700 3535 750 3565
rect 700 3515 715 3535
rect 735 3515 750 3535
rect 700 3485 750 3515
rect 700 3465 715 3485
rect 735 3465 750 3485
rect 700 3435 750 3465
rect 700 3415 715 3435
rect 735 3415 750 3435
rect 700 3385 750 3415
rect 850 3685 900 3715
rect 1150 3735 1200 3750
rect 1150 3715 1165 3735
rect 1185 3715 1200 3735
rect 850 3665 865 3685
rect 885 3665 900 3685
rect 850 3635 900 3665
rect 850 3615 865 3635
rect 885 3615 900 3635
rect 850 3585 900 3615
rect 850 3565 865 3585
rect 885 3565 900 3585
rect 850 3535 900 3565
rect 850 3515 865 3535
rect 885 3515 900 3535
rect 850 3485 900 3515
rect 850 3465 865 3485
rect 885 3465 900 3485
rect 850 3435 900 3465
rect 850 3415 865 3435
rect 885 3415 900 3435
rect 850 3400 900 3415
rect 1000 3685 1050 3700
rect 1000 3665 1015 3685
rect 1035 3665 1050 3685
rect 1000 3635 1050 3665
rect 1000 3615 1015 3635
rect 1035 3615 1050 3635
rect 1000 3585 1050 3615
rect 1000 3565 1015 3585
rect 1035 3565 1050 3585
rect 1000 3535 1050 3565
rect 1000 3515 1015 3535
rect 1035 3515 1050 3535
rect 1000 3485 1050 3515
rect 1000 3465 1015 3485
rect 1035 3465 1050 3485
rect 1000 3435 1050 3465
rect 1000 3415 1015 3435
rect 1035 3415 1050 3435
rect 700 3365 715 3385
rect 735 3365 750 3385
rect 700 3350 750 3365
rect 1000 3385 1050 3415
rect 1150 3685 1200 3715
rect 1450 3735 1500 3750
rect 1450 3715 1465 3735
rect 1485 3715 1500 3735
rect 1150 3665 1165 3685
rect 1185 3665 1200 3685
rect 1150 3635 1200 3665
rect 1150 3615 1165 3635
rect 1185 3615 1200 3635
rect 1150 3585 1200 3615
rect 1150 3565 1165 3585
rect 1185 3565 1200 3585
rect 1150 3535 1200 3565
rect 1150 3515 1165 3535
rect 1185 3515 1200 3535
rect 1150 3485 1200 3515
rect 1150 3465 1165 3485
rect 1185 3465 1200 3485
rect 1150 3435 1200 3465
rect 1150 3415 1165 3435
rect 1185 3415 1200 3435
rect 1150 3400 1200 3415
rect 1300 3685 1350 3700
rect 1300 3665 1315 3685
rect 1335 3665 1350 3685
rect 1300 3635 1350 3665
rect 1300 3615 1315 3635
rect 1335 3615 1350 3635
rect 1300 3585 1350 3615
rect 1300 3565 1315 3585
rect 1335 3565 1350 3585
rect 1300 3535 1350 3565
rect 1300 3515 1315 3535
rect 1335 3515 1350 3535
rect 1300 3485 1350 3515
rect 1300 3465 1315 3485
rect 1335 3465 1350 3485
rect 1300 3435 1350 3465
rect 1300 3415 1315 3435
rect 1335 3415 1350 3435
rect 1000 3365 1015 3385
rect 1035 3365 1050 3385
rect 1000 3350 1050 3365
rect 1300 3385 1350 3415
rect 1450 3685 1500 3715
rect 1750 3735 1800 3750
rect 1750 3715 1765 3735
rect 1785 3715 1800 3735
rect 1450 3665 1465 3685
rect 1485 3665 1500 3685
rect 1450 3635 1500 3665
rect 1450 3615 1465 3635
rect 1485 3615 1500 3635
rect 1450 3585 1500 3615
rect 1450 3565 1465 3585
rect 1485 3565 1500 3585
rect 1450 3535 1500 3565
rect 1450 3515 1465 3535
rect 1485 3515 1500 3535
rect 1450 3485 1500 3515
rect 1450 3465 1465 3485
rect 1485 3465 1500 3485
rect 1450 3435 1500 3465
rect 1450 3415 1465 3435
rect 1485 3415 1500 3435
rect 1450 3400 1500 3415
rect 1600 3685 1650 3700
rect 1600 3665 1615 3685
rect 1635 3665 1650 3685
rect 1600 3635 1650 3665
rect 1600 3615 1615 3635
rect 1635 3615 1650 3635
rect 1600 3585 1650 3615
rect 1600 3565 1615 3585
rect 1635 3565 1650 3585
rect 1600 3535 1650 3565
rect 1600 3515 1615 3535
rect 1635 3515 1650 3535
rect 1600 3485 1650 3515
rect 1600 3465 1615 3485
rect 1635 3465 1650 3485
rect 1600 3435 1650 3465
rect 1600 3415 1615 3435
rect 1635 3415 1650 3435
rect 1300 3365 1315 3385
rect 1335 3365 1350 3385
rect 1300 3350 1350 3365
rect 1600 3385 1650 3415
rect 1600 3365 1615 3385
rect 1635 3365 1650 3385
rect 1600 3350 1650 3365
rect 700 3335 1650 3350
rect 700 3315 715 3335
rect 735 3315 1650 3335
rect 700 3300 1650 3315
rect 1750 3685 1800 3715
rect 2050 3735 2100 3750
rect 2050 3715 2065 3735
rect 2085 3715 2100 3735
rect 1750 3665 1765 3685
rect 1785 3665 1800 3685
rect 1750 3635 1800 3665
rect 1750 3615 1765 3635
rect 1785 3615 1800 3635
rect 1750 3585 1800 3615
rect 1750 3565 1765 3585
rect 1785 3565 1800 3585
rect 1750 3535 1800 3565
rect 1750 3515 1765 3535
rect 1785 3515 1800 3535
rect 1750 3485 1800 3515
rect 1750 3465 1765 3485
rect 1785 3465 1800 3485
rect 1750 3435 1800 3465
rect 1750 3415 1765 3435
rect 1785 3415 1800 3435
rect 1750 3385 1800 3415
rect 1750 3365 1765 3385
rect 1785 3365 1800 3385
rect 1750 3335 1800 3365
rect 1750 3315 1765 3335
rect 1785 3315 1800 3335
rect 700 3240 750 3250
rect 700 3210 710 3240
rect 740 3210 750 3240
rect 700 3200 750 3210
rect 1000 3240 1050 3250
rect 1000 3210 1010 3240
rect 1040 3210 1050 3240
rect 1000 3200 1050 3210
rect 1150 3240 1200 3300
rect 1150 3210 1160 3240
rect 1190 3210 1200 3240
rect 1150 3150 1200 3210
rect 1300 3240 1350 3250
rect 1300 3210 1310 3240
rect 1340 3210 1350 3240
rect 1300 3200 1350 3210
rect 1600 3240 1650 3250
rect 1600 3210 1610 3240
rect 1640 3210 1650 3240
rect 1600 3200 1650 3210
rect 550 3115 565 3135
rect 585 3115 600 3135
rect 550 3085 600 3115
rect 550 3065 565 3085
rect 585 3065 600 3085
rect 550 3035 600 3065
rect 550 3015 565 3035
rect 585 3015 600 3035
rect 550 2985 600 3015
rect 550 2965 565 2985
rect 585 2965 600 2985
rect 550 2935 600 2965
rect 550 2915 565 2935
rect 585 2915 600 2935
rect 550 2885 600 2915
rect 550 2865 565 2885
rect 585 2865 600 2885
rect 550 2835 600 2865
rect 550 2815 565 2835
rect 585 2815 600 2835
rect 550 2785 600 2815
rect 550 2765 565 2785
rect 585 2765 600 2785
rect 550 2735 600 2765
rect 700 3135 1650 3150
rect 700 3115 715 3135
rect 735 3115 1015 3135
rect 1035 3115 1315 3135
rect 1335 3115 1615 3135
rect 1635 3115 1650 3135
rect 700 3100 1650 3115
rect 700 3085 750 3100
rect 700 3065 715 3085
rect 735 3065 750 3085
rect 700 3035 750 3065
rect 1000 3085 1050 3100
rect 1000 3065 1015 3085
rect 1035 3065 1050 3085
rect 700 3015 715 3035
rect 735 3015 750 3035
rect 700 2985 750 3015
rect 700 2965 715 2985
rect 735 2965 750 2985
rect 700 2935 750 2965
rect 700 2915 715 2935
rect 735 2915 750 2935
rect 700 2885 750 2915
rect 700 2865 715 2885
rect 735 2865 750 2885
rect 700 2835 750 2865
rect 700 2815 715 2835
rect 735 2815 750 2835
rect 700 2785 750 2815
rect 700 2765 715 2785
rect 735 2765 750 2785
rect 700 2750 750 2765
rect 850 3035 900 3050
rect 850 3015 865 3035
rect 885 3015 900 3035
rect 850 2985 900 3015
rect 850 2965 865 2985
rect 885 2965 900 2985
rect 850 2935 900 2965
rect 850 2915 865 2935
rect 885 2915 900 2935
rect 850 2885 900 2915
rect 850 2865 865 2885
rect 885 2865 900 2885
rect 850 2835 900 2865
rect 850 2815 865 2835
rect 885 2815 900 2835
rect 850 2785 900 2815
rect 850 2765 865 2785
rect 885 2765 900 2785
rect 550 2715 565 2735
rect 585 2715 600 2735
rect 550 2700 600 2715
rect 850 2735 900 2765
rect 1000 3035 1050 3065
rect 1300 3085 1350 3100
rect 1300 3065 1315 3085
rect 1335 3065 1350 3085
rect 1000 3015 1015 3035
rect 1035 3015 1050 3035
rect 1000 2985 1050 3015
rect 1000 2965 1015 2985
rect 1035 2965 1050 2985
rect 1000 2935 1050 2965
rect 1000 2915 1015 2935
rect 1035 2915 1050 2935
rect 1000 2885 1050 2915
rect 1000 2865 1015 2885
rect 1035 2865 1050 2885
rect 1000 2835 1050 2865
rect 1000 2815 1015 2835
rect 1035 2815 1050 2835
rect 1000 2785 1050 2815
rect 1000 2765 1015 2785
rect 1035 2765 1050 2785
rect 1000 2750 1050 2765
rect 1150 3035 1200 3050
rect 1150 3015 1165 3035
rect 1185 3015 1200 3035
rect 1150 2985 1200 3015
rect 1150 2965 1165 2985
rect 1185 2965 1200 2985
rect 1150 2935 1200 2965
rect 1150 2915 1165 2935
rect 1185 2915 1200 2935
rect 1150 2885 1200 2915
rect 1150 2865 1165 2885
rect 1185 2865 1200 2885
rect 1150 2835 1200 2865
rect 1150 2815 1165 2835
rect 1185 2815 1200 2835
rect 1150 2785 1200 2815
rect 1150 2765 1165 2785
rect 1185 2765 1200 2785
rect 850 2715 865 2735
rect 885 2715 900 2735
rect 850 2700 900 2715
rect 1150 2735 1200 2765
rect 1300 3035 1350 3065
rect 1600 3085 1650 3100
rect 1600 3065 1615 3085
rect 1635 3065 1650 3085
rect 1300 3015 1315 3035
rect 1335 3015 1350 3035
rect 1300 2985 1350 3015
rect 1300 2965 1315 2985
rect 1335 2965 1350 2985
rect 1300 2935 1350 2965
rect 1300 2915 1315 2935
rect 1335 2915 1350 2935
rect 1300 2885 1350 2915
rect 1300 2865 1315 2885
rect 1335 2865 1350 2885
rect 1300 2835 1350 2865
rect 1300 2815 1315 2835
rect 1335 2815 1350 2835
rect 1300 2785 1350 2815
rect 1300 2765 1315 2785
rect 1335 2765 1350 2785
rect 1300 2750 1350 2765
rect 1450 3035 1500 3050
rect 1450 3015 1465 3035
rect 1485 3015 1500 3035
rect 1450 2985 1500 3015
rect 1450 2965 1465 2985
rect 1485 2965 1500 2985
rect 1450 2935 1500 2965
rect 1450 2915 1465 2935
rect 1485 2915 1500 2935
rect 1450 2885 1500 2915
rect 1450 2865 1465 2885
rect 1485 2865 1500 2885
rect 1450 2835 1500 2865
rect 1450 2815 1465 2835
rect 1485 2815 1500 2835
rect 1450 2785 1500 2815
rect 1450 2765 1465 2785
rect 1485 2765 1500 2785
rect 1150 2715 1165 2735
rect 1185 2715 1200 2735
rect 1150 2700 1200 2715
rect 1450 2735 1500 2765
rect 1600 3035 1650 3065
rect 1600 3015 1615 3035
rect 1635 3015 1650 3035
rect 1600 2985 1650 3015
rect 1600 2965 1615 2985
rect 1635 2965 1650 2985
rect 1600 2935 1650 2965
rect 1600 2915 1615 2935
rect 1635 2915 1650 2935
rect 1600 2885 1650 2915
rect 1600 2865 1615 2885
rect 1635 2865 1650 2885
rect 1600 2835 1650 2865
rect 1600 2815 1615 2835
rect 1635 2815 1650 2835
rect 1600 2785 1650 2815
rect 1600 2765 1615 2785
rect 1635 2765 1650 2785
rect 1600 2750 1650 2765
rect 1750 3135 1800 3315
rect 1900 3685 1950 3700
rect 1900 3665 1915 3685
rect 1935 3665 1950 3685
rect 1900 3635 1950 3665
rect 1900 3615 1915 3635
rect 1935 3615 1950 3635
rect 1900 3585 1950 3615
rect 1900 3565 1915 3585
rect 1935 3565 1950 3585
rect 1900 3535 1950 3565
rect 1900 3515 1915 3535
rect 1935 3515 1950 3535
rect 1900 3485 1950 3515
rect 1900 3465 1915 3485
rect 1935 3465 1950 3485
rect 1900 3435 1950 3465
rect 1900 3415 1915 3435
rect 1935 3415 1950 3435
rect 1900 3385 1950 3415
rect 2050 3685 2100 3715
rect 2350 3735 2400 3750
rect 2350 3715 2365 3735
rect 2385 3715 2400 3735
rect 2050 3665 2065 3685
rect 2085 3665 2100 3685
rect 2050 3635 2100 3665
rect 2050 3615 2065 3635
rect 2085 3615 2100 3635
rect 2050 3585 2100 3615
rect 2050 3565 2065 3585
rect 2085 3565 2100 3585
rect 2050 3535 2100 3565
rect 2050 3515 2065 3535
rect 2085 3515 2100 3535
rect 2050 3485 2100 3515
rect 2050 3465 2065 3485
rect 2085 3465 2100 3485
rect 2050 3435 2100 3465
rect 2050 3415 2065 3435
rect 2085 3415 2100 3435
rect 2050 3400 2100 3415
rect 2200 3685 2250 3700
rect 2200 3665 2215 3685
rect 2235 3665 2250 3685
rect 2200 3635 2250 3665
rect 2200 3615 2215 3635
rect 2235 3615 2250 3635
rect 2200 3585 2250 3615
rect 2200 3565 2215 3585
rect 2235 3565 2250 3585
rect 2200 3535 2250 3565
rect 2200 3515 2215 3535
rect 2235 3515 2250 3535
rect 2200 3485 2250 3515
rect 2200 3465 2215 3485
rect 2235 3465 2250 3485
rect 2200 3435 2250 3465
rect 2200 3415 2215 3435
rect 2235 3415 2250 3435
rect 1900 3365 1915 3385
rect 1935 3365 1950 3385
rect 1900 3350 1950 3365
rect 2200 3385 2250 3415
rect 2200 3365 2215 3385
rect 2235 3365 2250 3385
rect 2200 3350 2250 3365
rect 1900 3335 2250 3350
rect 1900 3315 1915 3335
rect 1935 3315 2215 3335
rect 2235 3315 2250 3335
rect 1900 3300 2250 3315
rect 2350 3685 2400 3715
rect 2650 3735 2700 3750
rect 2650 3715 2665 3735
rect 2685 3715 2700 3735
rect 2350 3665 2365 3685
rect 2385 3665 2400 3685
rect 2350 3635 2400 3665
rect 2350 3615 2365 3635
rect 2385 3615 2400 3635
rect 2350 3585 2400 3615
rect 2350 3565 2365 3585
rect 2385 3565 2400 3585
rect 2350 3535 2400 3565
rect 2350 3515 2365 3535
rect 2385 3515 2400 3535
rect 2350 3485 2400 3515
rect 2350 3465 2365 3485
rect 2385 3465 2400 3485
rect 2350 3435 2400 3465
rect 2350 3415 2365 3435
rect 2385 3415 2400 3435
rect 2350 3385 2400 3415
rect 2350 3365 2365 3385
rect 2385 3365 2400 3385
rect 2350 3335 2400 3365
rect 2350 3315 2365 3335
rect 2385 3315 2400 3335
rect 1900 3240 1950 3250
rect 1900 3210 1910 3240
rect 1940 3210 1950 3240
rect 1900 3200 1950 3210
rect 2050 3240 2100 3300
rect 2050 3210 2060 3240
rect 2090 3210 2100 3240
rect 2050 3150 2100 3210
rect 2200 3240 2250 3250
rect 2200 3210 2210 3240
rect 2240 3210 2250 3240
rect 2200 3200 2250 3210
rect 1750 3115 1765 3135
rect 1785 3115 1800 3135
rect 1750 3085 1800 3115
rect 1750 3065 1765 3085
rect 1785 3065 1800 3085
rect 1750 3035 1800 3065
rect 1750 3015 1765 3035
rect 1785 3015 1800 3035
rect 1750 2985 1800 3015
rect 1750 2965 1765 2985
rect 1785 2965 1800 2985
rect 1750 2935 1800 2965
rect 1750 2915 1765 2935
rect 1785 2915 1800 2935
rect 1750 2885 1800 2915
rect 1750 2865 1765 2885
rect 1785 2865 1800 2885
rect 1750 2835 1800 2865
rect 1750 2815 1765 2835
rect 1785 2815 1800 2835
rect 1750 2785 1800 2815
rect 1750 2765 1765 2785
rect 1785 2765 1800 2785
rect 1450 2715 1465 2735
rect 1485 2715 1500 2735
rect 1450 2700 1500 2715
rect 1750 2735 1800 2765
rect 1900 3135 2250 3150
rect 1900 3115 1915 3135
rect 1935 3115 2215 3135
rect 2235 3115 2250 3135
rect 1900 3100 2250 3115
rect 1900 3085 1950 3100
rect 1900 3065 1915 3085
rect 1935 3065 1950 3085
rect 1900 3035 1950 3065
rect 2200 3085 2250 3100
rect 2200 3065 2215 3085
rect 2235 3065 2250 3085
rect 1900 3015 1915 3035
rect 1935 3015 1950 3035
rect 1900 2985 1950 3015
rect 1900 2965 1915 2985
rect 1935 2965 1950 2985
rect 1900 2935 1950 2965
rect 1900 2915 1915 2935
rect 1935 2915 1950 2935
rect 1900 2885 1950 2915
rect 1900 2865 1915 2885
rect 1935 2865 1950 2885
rect 1900 2835 1950 2865
rect 1900 2815 1915 2835
rect 1935 2815 1950 2835
rect 1900 2785 1950 2815
rect 1900 2765 1915 2785
rect 1935 2765 1950 2785
rect 1900 2750 1950 2765
rect 2050 3035 2100 3050
rect 2050 3015 2065 3035
rect 2085 3015 2100 3035
rect 2050 2985 2100 3015
rect 2050 2965 2065 2985
rect 2085 2965 2100 2985
rect 2050 2935 2100 2965
rect 2050 2915 2065 2935
rect 2085 2915 2100 2935
rect 2050 2885 2100 2915
rect 2050 2865 2065 2885
rect 2085 2865 2100 2885
rect 2050 2835 2100 2865
rect 2050 2815 2065 2835
rect 2085 2815 2100 2835
rect 2050 2785 2100 2815
rect 2050 2765 2065 2785
rect 2085 2765 2100 2785
rect 1750 2715 1765 2735
rect 1785 2715 1800 2735
rect 1750 2700 1800 2715
rect 2050 2735 2100 2765
rect 2200 3035 2250 3065
rect 2200 3015 2215 3035
rect 2235 3015 2250 3035
rect 2200 2985 2250 3015
rect 2200 2965 2215 2985
rect 2235 2965 2250 2985
rect 2200 2935 2250 2965
rect 2200 2915 2215 2935
rect 2235 2915 2250 2935
rect 2200 2885 2250 2915
rect 2200 2865 2215 2885
rect 2235 2865 2250 2885
rect 2200 2835 2250 2865
rect 2200 2815 2215 2835
rect 2235 2815 2250 2835
rect 2200 2785 2250 2815
rect 2200 2765 2215 2785
rect 2235 2765 2250 2785
rect 2200 2750 2250 2765
rect 2350 3135 2400 3315
rect 2500 3685 2550 3700
rect 2500 3665 2515 3685
rect 2535 3665 2550 3685
rect 2500 3635 2550 3665
rect 2500 3615 2515 3635
rect 2535 3615 2550 3635
rect 2500 3585 2550 3615
rect 2500 3565 2515 3585
rect 2535 3565 2550 3585
rect 2500 3535 2550 3565
rect 2500 3515 2515 3535
rect 2535 3515 2550 3535
rect 2500 3485 2550 3515
rect 2500 3465 2515 3485
rect 2535 3465 2550 3485
rect 2500 3435 2550 3465
rect 2500 3415 2515 3435
rect 2535 3415 2550 3435
rect 2500 3385 2550 3415
rect 2650 3685 2700 3715
rect 2950 3735 3000 3750
rect 2950 3715 2965 3735
rect 2985 3715 3000 3735
rect 2650 3665 2665 3685
rect 2685 3665 2700 3685
rect 2650 3635 2700 3665
rect 2650 3615 2665 3635
rect 2685 3615 2700 3635
rect 2650 3585 2700 3615
rect 2650 3565 2665 3585
rect 2685 3565 2700 3585
rect 2650 3535 2700 3565
rect 2650 3515 2665 3535
rect 2685 3515 2700 3535
rect 2650 3485 2700 3515
rect 2650 3465 2665 3485
rect 2685 3465 2700 3485
rect 2650 3435 2700 3465
rect 2650 3415 2665 3435
rect 2685 3415 2700 3435
rect 2650 3400 2700 3415
rect 2800 3685 2850 3700
rect 2800 3665 2815 3685
rect 2835 3665 2850 3685
rect 2800 3635 2850 3665
rect 2800 3615 2815 3635
rect 2835 3615 2850 3635
rect 2800 3585 2850 3615
rect 2800 3565 2815 3585
rect 2835 3565 2850 3585
rect 2800 3535 2850 3565
rect 2800 3515 2815 3535
rect 2835 3515 2850 3535
rect 2800 3485 2850 3515
rect 2800 3465 2815 3485
rect 2835 3465 2850 3485
rect 2800 3435 2850 3465
rect 2800 3415 2815 3435
rect 2835 3415 2850 3435
rect 2500 3365 2515 3385
rect 2535 3365 2550 3385
rect 2500 3350 2550 3365
rect 2800 3385 2850 3415
rect 2950 3685 3000 3715
rect 3250 3735 3300 3750
rect 3250 3715 3265 3735
rect 3285 3715 3300 3735
rect 2950 3665 2965 3685
rect 2985 3665 3000 3685
rect 2950 3635 3000 3665
rect 2950 3615 2965 3635
rect 2985 3615 3000 3635
rect 2950 3585 3000 3615
rect 2950 3565 2965 3585
rect 2985 3565 3000 3585
rect 2950 3535 3000 3565
rect 2950 3515 2965 3535
rect 2985 3515 3000 3535
rect 2950 3485 3000 3515
rect 2950 3465 2965 3485
rect 2985 3465 3000 3485
rect 2950 3435 3000 3465
rect 2950 3415 2965 3435
rect 2985 3415 3000 3435
rect 2950 3400 3000 3415
rect 3100 3685 3150 3700
rect 3100 3665 3115 3685
rect 3135 3665 3150 3685
rect 3100 3635 3150 3665
rect 3100 3615 3115 3635
rect 3135 3615 3150 3635
rect 3100 3585 3150 3615
rect 3100 3565 3115 3585
rect 3135 3565 3150 3585
rect 3100 3535 3150 3565
rect 3100 3515 3115 3535
rect 3135 3515 3150 3535
rect 3100 3485 3150 3515
rect 3100 3465 3115 3485
rect 3135 3465 3150 3485
rect 3100 3435 3150 3465
rect 3100 3415 3115 3435
rect 3135 3415 3150 3435
rect 2800 3365 2815 3385
rect 2835 3365 2850 3385
rect 2800 3350 2850 3365
rect 3100 3385 3150 3415
rect 3250 3685 3300 3715
rect 3550 3735 3600 3750
rect 3550 3715 3565 3735
rect 3585 3715 3600 3735
rect 3250 3665 3265 3685
rect 3285 3665 3300 3685
rect 3250 3635 3300 3665
rect 3250 3615 3265 3635
rect 3285 3615 3300 3635
rect 3250 3585 3300 3615
rect 3250 3565 3265 3585
rect 3285 3565 3300 3585
rect 3250 3535 3300 3565
rect 3250 3515 3265 3535
rect 3285 3515 3300 3535
rect 3250 3485 3300 3515
rect 3250 3465 3265 3485
rect 3285 3465 3300 3485
rect 3250 3435 3300 3465
rect 3250 3415 3265 3435
rect 3285 3415 3300 3435
rect 3250 3400 3300 3415
rect 3400 3685 3450 3700
rect 3400 3665 3415 3685
rect 3435 3665 3450 3685
rect 3400 3635 3450 3665
rect 3400 3615 3415 3635
rect 3435 3615 3450 3635
rect 3400 3585 3450 3615
rect 3400 3565 3415 3585
rect 3435 3565 3450 3585
rect 3400 3535 3450 3565
rect 3400 3515 3415 3535
rect 3435 3515 3450 3535
rect 3400 3485 3450 3515
rect 3400 3465 3415 3485
rect 3435 3465 3450 3485
rect 3400 3435 3450 3465
rect 3400 3415 3415 3435
rect 3435 3415 3450 3435
rect 3100 3365 3115 3385
rect 3135 3365 3150 3385
rect 3100 3350 3150 3365
rect 3400 3385 3450 3415
rect 3400 3365 3415 3385
rect 3435 3365 3450 3385
rect 3400 3350 3450 3365
rect 2500 3335 3450 3350
rect 2500 3315 3415 3335
rect 3435 3315 3450 3335
rect 2500 3300 3450 3315
rect 3550 3685 3600 3715
rect 3550 3665 3565 3685
rect 3585 3665 3600 3685
rect 3550 3635 3600 3665
rect 3550 3615 3565 3635
rect 3585 3615 3600 3635
rect 3550 3585 3600 3615
rect 3550 3565 3565 3585
rect 3585 3565 3600 3585
rect 3550 3535 3600 3565
rect 3550 3515 3565 3535
rect 3585 3515 3600 3535
rect 3550 3485 3600 3515
rect 3550 3465 3565 3485
rect 3585 3465 3600 3485
rect 3550 3435 3600 3465
rect 3550 3415 3565 3435
rect 3585 3415 3600 3435
rect 3550 3385 3600 3415
rect 3550 3365 3565 3385
rect 3585 3365 3600 3385
rect 3550 3335 3600 3365
rect 3550 3315 3565 3335
rect 3585 3315 3600 3335
rect 2500 3240 2550 3250
rect 2500 3210 2510 3240
rect 2540 3210 2550 3240
rect 2500 3200 2550 3210
rect 2800 3240 2850 3250
rect 2800 3210 2810 3240
rect 2840 3210 2850 3240
rect 2800 3200 2850 3210
rect 2950 3240 3000 3300
rect 2950 3210 2960 3240
rect 2990 3210 3000 3240
rect 2950 3150 3000 3210
rect 3100 3240 3150 3250
rect 3100 3210 3110 3240
rect 3140 3210 3150 3240
rect 3100 3200 3150 3210
rect 3400 3240 3450 3250
rect 3400 3210 3410 3240
rect 3440 3210 3450 3240
rect 3400 3200 3450 3210
rect 2350 3115 2365 3135
rect 2385 3115 2400 3135
rect 2350 3085 2400 3115
rect 2350 3065 2365 3085
rect 2385 3065 2400 3085
rect 2350 3035 2400 3065
rect 2350 3015 2365 3035
rect 2385 3015 2400 3035
rect 2350 2985 2400 3015
rect 2350 2965 2365 2985
rect 2385 2965 2400 2985
rect 2350 2935 2400 2965
rect 2350 2915 2365 2935
rect 2385 2915 2400 2935
rect 2350 2885 2400 2915
rect 2350 2865 2365 2885
rect 2385 2865 2400 2885
rect 2350 2835 2400 2865
rect 2350 2815 2365 2835
rect 2385 2815 2400 2835
rect 2350 2785 2400 2815
rect 2350 2765 2365 2785
rect 2385 2765 2400 2785
rect 2050 2715 2065 2735
rect 2085 2715 2100 2735
rect 2050 2700 2100 2715
rect 2350 2735 2400 2765
rect 2500 3135 3450 3150
rect 2500 3115 2515 3135
rect 2535 3115 2815 3135
rect 2835 3115 3115 3135
rect 3135 3115 3415 3135
rect 3435 3115 3450 3135
rect 2500 3100 3450 3115
rect 2500 3085 2550 3100
rect 2500 3065 2515 3085
rect 2535 3065 2550 3085
rect 2500 3035 2550 3065
rect 2800 3085 2850 3100
rect 2800 3065 2815 3085
rect 2835 3065 2850 3085
rect 2500 3015 2515 3035
rect 2535 3015 2550 3035
rect 2500 2985 2550 3015
rect 2500 2965 2515 2985
rect 2535 2965 2550 2985
rect 2500 2935 2550 2965
rect 2500 2915 2515 2935
rect 2535 2915 2550 2935
rect 2500 2885 2550 2915
rect 2500 2865 2515 2885
rect 2535 2865 2550 2885
rect 2500 2835 2550 2865
rect 2500 2815 2515 2835
rect 2535 2815 2550 2835
rect 2500 2785 2550 2815
rect 2500 2765 2515 2785
rect 2535 2765 2550 2785
rect 2500 2750 2550 2765
rect 2650 3035 2700 3050
rect 2650 3015 2665 3035
rect 2685 3015 2700 3035
rect 2650 2985 2700 3015
rect 2650 2965 2665 2985
rect 2685 2965 2700 2985
rect 2650 2935 2700 2965
rect 2650 2915 2665 2935
rect 2685 2915 2700 2935
rect 2650 2885 2700 2915
rect 2650 2865 2665 2885
rect 2685 2865 2700 2885
rect 2650 2835 2700 2865
rect 2650 2815 2665 2835
rect 2685 2815 2700 2835
rect 2650 2785 2700 2815
rect 2650 2765 2665 2785
rect 2685 2765 2700 2785
rect 2350 2715 2365 2735
rect 2385 2715 2400 2735
rect 2350 2700 2400 2715
rect 2650 2735 2700 2765
rect 2800 3035 2850 3065
rect 3100 3085 3150 3100
rect 3100 3065 3115 3085
rect 3135 3065 3150 3085
rect 2800 3015 2815 3035
rect 2835 3015 2850 3035
rect 2800 2985 2850 3015
rect 2800 2965 2815 2985
rect 2835 2965 2850 2985
rect 2800 2935 2850 2965
rect 2800 2915 2815 2935
rect 2835 2915 2850 2935
rect 2800 2885 2850 2915
rect 2800 2865 2815 2885
rect 2835 2865 2850 2885
rect 2800 2835 2850 2865
rect 2800 2815 2815 2835
rect 2835 2815 2850 2835
rect 2800 2785 2850 2815
rect 2800 2765 2815 2785
rect 2835 2765 2850 2785
rect 2800 2750 2850 2765
rect 2950 3035 3000 3050
rect 2950 3015 2965 3035
rect 2985 3015 3000 3035
rect 2950 2985 3000 3015
rect 2950 2965 2965 2985
rect 2985 2965 3000 2985
rect 2950 2935 3000 2965
rect 2950 2915 2965 2935
rect 2985 2915 3000 2935
rect 2950 2885 3000 2915
rect 2950 2865 2965 2885
rect 2985 2865 3000 2885
rect 2950 2835 3000 2865
rect 2950 2815 2965 2835
rect 2985 2815 3000 2835
rect 2950 2785 3000 2815
rect 2950 2765 2965 2785
rect 2985 2765 3000 2785
rect 2650 2715 2665 2735
rect 2685 2715 2700 2735
rect 2650 2700 2700 2715
rect 2950 2735 3000 2765
rect 3100 3035 3150 3065
rect 3400 3085 3450 3100
rect 3400 3065 3415 3085
rect 3435 3065 3450 3085
rect 3100 3015 3115 3035
rect 3135 3015 3150 3035
rect 3100 2985 3150 3015
rect 3100 2965 3115 2985
rect 3135 2965 3150 2985
rect 3100 2935 3150 2965
rect 3100 2915 3115 2935
rect 3135 2915 3150 2935
rect 3100 2885 3150 2915
rect 3100 2865 3115 2885
rect 3135 2865 3150 2885
rect 3100 2835 3150 2865
rect 3100 2815 3115 2835
rect 3135 2815 3150 2835
rect 3100 2785 3150 2815
rect 3100 2765 3115 2785
rect 3135 2765 3150 2785
rect 3100 2750 3150 2765
rect 3250 3035 3300 3050
rect 3250 3015 3265 3035
rect 3285 3015 3300 3035
rect 3250 2985 3300 3015
rect 3250 2965 3265 2985
rect 3285 2965 3300 2985
rect 3250 2935 3300 2965
rect 3250 2915 3265 2935
rect 3285 2915 3300 2935
rect 3250 2885 3300 2915
rect 3250 2865 3265 2885
rect 3285 2865 3300 2885
rect 3250 2835 3300 2865
rect 3250 2815 3265 2835
rect 3285 2815 3300 2835
rect 3250 2785 3300 2815
rect 3250 2765 3265 2785
rect 3285 2765 3300 2785
rect 2950 2715 2965 2735
rect 2985 2715 3000 2735
rect 2950 2700 3000 2715
rect 3250 2735 3300 2765
rect 3400 3035 3450 3065
rect 3400 3015 3415 3035
rect 3435 3015 3450 3035
rect 3400 2985 3450 3015
rect 3400 2965 3415 2985
rect 3435 2965 3450 2985
rect 3400 2935 3450 2965
rect 3400 2915 3415 2935
rect 3435 2915 3450 2935
rect 3400 2885 3450 2915
rect 3400 2865 3415 2885
rect 3435 2865 3450 2885
rect 3400 2835 3450 2865
rect 3400 2815 3415 2835
rect 3435 2815 3450 2835
rect 3400 2785 3450 2815
rect 3400 2765 3415 2785
rect 3435 2765 3450 2785
rect 3400 2750 3450 2765
rect 3550 3135 3600 3315
rect 4150 3785 4200 3860
rect 8350 3890 8400 3965
rect 8500 4435 8550 4450
rect 8500 4415 8515 4435
rect 8535 4415 8550 4435
rect 8500 4385 8550 4415
rect 8500 4365 8515 4385
rect 8535 4365 8550 4385
rect 8500 4335 8550 4365
rect 8500 4315 8515 4335
rect 8535 4315 8550 4335
rect 8500 4285 8550 4315
rect 8500 4265 8515 4285
rect 8535 4265 8550 4285
rect 8500 4235 8550 4265
rect 8500 4215 8515 4235
rect 8535 4215 8550 4235
rect 8500 4185 8550 4215
rect 8500 4165 8515 4185
rect 8535 4165 8550 4185
rect 8500 4135 8550 4165
rect 8500 4115 8515 4135
rect 8535 4115 8550 4135
rect 8500 4085 8550 4115
rect 8500 4065 8515 4085
rect 8535 4065 8550 4085
rect 8500 4035 8550 4065
rect 8500 4015 8515 4035
rect 8535 4015 8550 4035
rect 8500 3985 8550 4015
rect 8500 3965 8515 3985
rect 8535 3965 8550 3985
rect 8500 3950 8550 3965
rect 8650 4440 8700 4610
rect 8800 5085 8850 5100
rect 8800 5065 8815 5085
rect 8835 5065 8850 5085
rect 8800 5035 8850 5065
rect 8800 5015 8815 5035
rect 8835 5015 8850 5035
rect 8800 4985 8850 5015
rect 8800 4965 8815 4985
rect 8835 4965 8850 4985
rect 8800 4935 8850 4965
rect 8800 4915 8815 4935
rect 8835 4915 8850 4935
rect 8800 4885 8850 4915
rect 8800 4865 8815 4885
rect 8835 4865 8850 4885
rect 8800 4835 8850 4865
rect 8800 4815 8815 4835
rect 8835 4815 8850 4835
rect 8800 4785 8850 4815
rect 8800 4765 8815 4785
rect 8835 4765 8850 4785
rect 8800 4735 8850 4765
rect 8800 4715 8815 4735
rect 8835 4715 8850 4735
rect 8800 4685 8850 4715
rect 8800 4665 8815 4685
rect 8835 4665 8850 4685
rect 8800 4635 8850 4665
rect 8800 4615 8815 4635
rect 8835 4615 8850 4635
rect 8800 4600 8850 4615
rect 8950 5085 9000 5160
rect 9250 5190 9300 5200
rect 9250 5160 9260 5190
rect 9290 5160 9300 5190
rect 8950 5065 8965 5085
rect 8985 5065 9000 5085
rect 8950 5040 9000 5065
rect 8950 5010 8960 5040
rect 8990 5010 9000 5040
rect 8950 4985 9000 5010
rect 8950 4965 8965 4985
rect 8985 4965 9000 4985
rect 8950 4940 9000 4965
rect 8950 4910 8960 4940
rect 8990 4910 9000 4940
rect 8950 4885 9000 4910
rect 8950 4865 8965 4885
rect 8985 4865 9000 4885
rect 8950 4840 9000 4865
rect 8950 4810 8960 4840
rect 8990 4810 9000 4840
rect 8950 4785 9000 4810
rect 8950 4765 8965 4785
rect 8985 4765 9000 4785
rect 8950 4740 9000 4765
rect 8950 4710 8960 4740
rect 8990 4710 9000 4740
rect 8950 4685 9000 4710
rect 8950 4665 8965 4685
rect 8985 4665 9000 4685
rect 8950 4640 9000 4665
rect 8950 4610 8960 4640
rect 8990 4610 9000 4640
rect 8800 4540 8850 4550
rect 8800 4510 8810 4540
rect 8840 4510 8850 4540
rect 8800 4500 8850 4510
rect 8650 4410 8660 4440
rect 8690 4410 8700 4440
rect 8650 4385 8700 4410
rect 8650 4365 8665 4385
rect 8685 4365 8700 4385
rect 8650 4340 8700 4365
rect 8650 4310 8660 4340
rect 8690 4310 8700 4340
rect 8650 4285 8700 4310
rect 8650 4265 8665 4285
rect 8685 4265 8700 4285
rect 8650 4240 8700 4265
rect 8650 4210 8660 4240
rect 8690 4210 8700 4240
rect 8650 4185 8700 4210
rect 8650 4165 8665 4185
rect 8685 4165 8700 4185
rect 8650 4140 8700 4165
rect 8650 4110 8660 4140
rect 8690 4110 8700 4140
rect 8650 4085 8700 4110
rect 8650 4065 8665 4085
rect 8685 4065 8700 4085
rect 8650 4040 8700 4065
rect 8650 4010 8660 4040
rect 8690 4010 8700 4040
rect 8650 3985 8700 4010
rect 8650 3965 8665 3985
rect 8685 3965 8700 3985
rect 8350 3860 8360 3890
rect 8390 3860 8400 3890
rect 4150 3765 4165 3785
rect 4185 3765 4200 3785
rect 4150 3735 4200 3765
rect 4150 3715 4165 3735
rect 4185 3715 4200 3735
rect 4150 3685 4200 3715
rect 4150 3665 4165 3685
rect 4185 3665 4200 3685
rect 4150 3635 4200 3665
rect 4150 3615 4165 3635
rect 4185 3615 4200 3635
rect 4150 3585 4200 3615
rect 4150 3565 4165 3585
rect 4185 3565 4200 3585
rect 4150 3535 4200 3565
rect 4150 3515 4165 3535
rect 4185 3515 4200 3535
rect 4150 3485 4200 3515
rect 4150 3465 4165 3485
rect 4185 3465 4200 3485
rect 4150 3435 4200 3465
rect 4150 3415 4165 3435
rect 4185 3415 4200 3435
rect 3700 3240 3750 3250
rect 3700 3210 3710 3240
rect 3740 3210 3750 3240
rect 3700 3200 3750 3210
rect 4000 3240 4050 3250
rect 4000 3210 4010 3240
rect 4040 3210 4050 3240
rect 4000 3200 4050 3210
rect 3550 3115 3565 3135
rect 3585 3115 3600 3135
rect 3550 3085 3600 3115
rect 3550 3065 3565 3085
rect 3585 3065 3600 3085
rect 3550 3035 3600 3065
rect 3550 3015 3565 3035
rect 3585 3015 3600 3035
rect 3550 2985 3600 3015
rect 3550 2965 3565 2985
rect 3585 2965 3600 2985
rect 3550 2935 3600 2965
rect 3550 2915 3565 2935
rect 3585 2915 3600 2935
rect 3550 2885 3600 2915
rect 3550 2865 3565 2885
rect 3585 2865 3600 2885
rect 3550 2835 3600 2865
rect 3550 2815 3565 2835
rect 3585 2815 3600 2835
rect 3550 2785 3600 2815
rect 3550 2765 3565 2785
rect 3585 2765 3600 2785
rect 3250 2715 3265 2735
rect 3285 2715 3300 2735
rect 3250 2700 3300 2715
rect 3550 2735 3600 2765
rect 3550 2715 3565 2735
rect 3585 2715 3600 2735
rect 3550 2700 3600 2715
rect 550 2685 3600 2700
rect 550 2665 565 2685
rect 585 2665 865 2685
rect 885 2665 1165 2685
rect 1185 2665 1465 2685
rect 1485 2665 1765 2685
rect 1785 2665 2065 2685
rect 2085 2665 2365 2685
rect 2385 2665 2665 2685
rect 2685 2665 2965 2685
rect 2985 2665 3265 2685
rect 3285 2665 3565 2685
rect 3585 2665 3600 2685
rect 550 2650 3600 2665
rect 4150 3140 4200 3415
rect 4750 3785 7800 3800
rect 4750 3765 4765 3785
rect 4785 3765 5065 3785
rect 5085 3765 5365 3785
rect 5385 3765 5665 3785
rect 5685 3765 5965 3785
rect 5985 3765 6265 3785
rect 6285 3765 6565 3785
rect 6585 3765 6865 3785
rect 6885 3765 7165 3785
rect 7185 3765 7465 3785
rect 7485 3765 7765 3785
rect 7785 3765 7800 3785
rect 4750 3750 7800 3765
rect 4750 3735 4800 3750
rect 4750 3715 4765 3735
rect 4785 3715 4800 3735
rect 4750 3685 4800 3715
rect 5050 3735 5100 3750
rect 5050 3715 5065 3735
rect 5085 3715 5100 3735
rect 4750 3665 4765 3685
rect 4785 3665 4800 3685
rect 4750 3635 4800 3665
rect 4750 3615 4765 3635
rect 4785 3615 4800 3635
rect 4750 3585 4800 3615
rect 4750 3565 4765 3585
rect 4785 3565 4800 3585
rect 4750 3535 4800 3565
rect 4750 3515 4765 3535
rect 4785 3515 4800 3535
rect 4750 3485 4800 3515
rect 4750 3465 4765 3485
rect 4785 3465 4800 3485
rect 4750 3435 4800 3465
rect 4750 3415 4765 3435
rect 4785 3415 4800 3435
rect 4750 3385 4800 3415
rect 4750 3365 4765 3385
rect 4785 3365 4800 3385
rect 4750 3335 4800 3365
rect 4750 3315 4765 3335
rect 4785 3315 4800 3335
rect 4300 3240 4350 3250
rect 4300 3210 4310 3240
rect 4340 3210 4350 3240
rect 4300 3200 4350 3210
rect 4600 3240 4650 3250
rect 4600 3210 4610 3240
rect 4640 3210 4650 3240
rect 4600 3200 4650 3210
rect 4150 3110 4160 3140
rect 4190 3110 4200 3140
rect 4150 3040 4200 3110
rect 4150 3010 4160 3040
rect 4190 3010 4200 3040
rect 4150 2985 4200 3010
rect 4150 2965 4165 2985
rect 4185 2965 4200 2985
rect 4150 2940 4200 2965
rect 4150 2910 4160 2940
rect 4190 2910 4200 2940
rect 4150 2885 4200 2910
rect 4150 2865 4165 2885
rect 4185 2865 4200 2885
rect 4150 2840 4200 2865
rect 4150 2810 4160 2840
rect 4190 2810 4200 2840
rect 4150 2785 4200 2810
rect 4150 2765 4165 2785
rect 4185 2765 4200 2785
rect 4150 2740 4200 2765
rect 4150 2710 4160 2740
rect 4190 2710 4200 2740
rect 4150 2685 4200 2710
rect 4150 2665 4165 2685
rect 4185 2665 4200 2685
rect -50 2560 -40 2590
rect -10 2560 0 2590
rect -50 2550 0 2560
rect 4150 2590 4200 2665
rect 4750 3135 4800 3315
rect 4900 3685 4950 3700
rect 4900 3665 4915 3685
rect 4935 3665 4950 3685
rect 4900 3635 4950 3665
rect 4900 3615 4915 3635
rect 4935 3615 4950 3635
rect 4900 3585 4950 3615
rect 4900 3565 4915 3585
rect 4935 3565 4950 3585
rect 4900 3535 4950 3565
rect 4900 3515 4915 3535
rect 4935 3515 4950 3535
rect 4900 3485 4950 3515
rect 4900 3465 4915 3485
rect 4935 3465 4950 3485
rect 4900 3435 4950 3465
rect 4900 3415 4915 3435
rect 4935 3415 4950 3435
rect 4900 3385 4950 3415
rect 5050 3685 5100 3715
rect 5350 3735 5400 3750
rect 5350 3715 5365 3735
rect 5385 3715 5400 3735
rect 5050 3665 5065 3685
rect 5085 3665 5100 3685
rect 5050 3635 5100 3665
rect 5050 3615 5065 3635
rect 5085 3615 5100 3635
rect 5050 3585 5100 3615
rect 5050 3565 5065 3585
rect 5085 3565 5100 3585
rect 5050 3535 5100 3565
rect 5050 3515 5065 3535
rect 5085 3515 5100 3535
rect 5050 3485 5100 3515
rect 5050 3465 5065 3485
rect 5085 3465 5100 3485
rect 5050 3435 5100 3465
rect 5050 3415 5065 3435
rect 5085 3415 5100 3435
rect 5050 3400 5100 3415
rect 5200 3685 5250 3700
rect 5200 3665 5215 3685
rect 5235 3665 5250 3685
rect 5200 3635 5250 3665
rect 5200 3615 5215 3635
rect 5235 3615 5250 3635
rect 5200 3585 5250 3615
rect 5200 3565 5215 3585
rect 5235 3565 5250 3585
rect 5200 3535 5250 3565
rect 5200 3515 5215 3535
rect 5235 3515 5250 3535
rect 5200 3485 5250 3515
rect 5200 3465 5215 3485
rect 5235 3465 5250 3485
rect 5200 3435 5250 3465
rect 5200 3415 5215 3435
rect 5235 3415 5250 3435
rect 4900 3365 4915 3385
rect 4935 3365 4950 3385
rect 4900 3350 4950 3365
rect 5200 3385 5250 3415
rect 5350 3685 5400 3715
rect 5650 3735 5700 3750
rect 5650 3715 5665 3735
rect 5685 3715 5700 3735
rect 5350 3665 5365 3685
rect 5385 3665 5400 3685
rect 5350 3635 5400 3665
rect 5350 3615 5365 3635
rect 5385 3615 5400 3635
rect 5350 3585 5400 3615
rect 5350 3565 5365 3585
rect 5385 3565 5400 3585
rect 5350 3535 5400 3565
rect 5350 3515 5365 3535
rect 5385 3515 5400 3535
rect 5350 3485 5400 3515
rect 5350 3465 5365 3485
rect 5385 3465 5400 3485
rect 5350 3435 5400 3465
rect 5350 3415 5365 3435
rect 5385 3415 5400 3435
rect 5350 3400 5400 3415
rect 5500 3685 5550 3700
rect 5500 3665 5515 3685
rect 5535 3665 5550 3685
rect 5500 3635 5550 3665
rect 5500 3615 5515 3635
rect 5535 3615 5550 3635
rect 5500 3585 5550 3615
rect 5500 3565 5515 3585
rect 5535 3565 5550 3585
rect 5500 3535 5550 3565
rect 5500 3515 5515 3535
rect 5535 3515 5550 3535
rect 5500 3485 5550 3515
rect 5500 3465 5515 3485
rect 5535 3465 5550 3485
rect 5500 3435 5550 3465
rect 5500 3415 5515 3435
rect 5535 3415 5550 3435
rect 5200 3365 5215 3385
rect 5235 3365 5250 3385
rect 5200 3350 5250 3365
rect 5500 3385 5550 3415
rect 5650 3685 5700 3715
rect 5950 3735 6000 3750
rect 5950 3715 5965 3735
rect 5985 3715 6000 3735
rect 5650 3665 5665 3685
rect 5685 3665 5700 3685
rect 5650 3635 5700 3665
rect 5650 3615 5665 3635
rect 5685 3615 5700 3635
rect 5650 3585 5700 3615
rect 5650 3565 5665 3585
rect 5685 3565 5700 3585
rect 5650 3535 5700 3565
rect 5650 3515 5665 3535
rect 5685 3515 5700 3535
rect 5650 3485 5700 3515
rect 5650 3465 5665 3485
rect 5685 3465 5700 3485
rect 5650 3435 5700 3465
rect 5650 3415 5665 3435
rect 5685 3415 5700 3435
rect 5650 3400 5700 3415
rect 5800 3685 5850 3700
rect 5800 3665 5815 3685
rect 5835 3665 5850 3685
rect 5800 3635 5850 3665
rect 5800 3615 5815 3635
rect 5835 3615 5850 3635
rect 5800 3585 5850 3615
rect 5800 3565 5815 3585
rect 5835 3565 5850 3585
rect 5800 3535 5850 3565
rect 5800 3515 5815 3535
rect 5835 3515 5850 3535
rect 5800 3485 5850 3515
rect 5800 3465 5815 3485
rect 5835 3465 5850 3485
rect 5800 3435 5850 3465
rect 5800 3415 5815 3435
rect 5835 3415 5850 3435
rect 5500 3365 5515 3385
rect 5535 3365 5550 3385
rect 5500 3350 5550 3365
rect 5800 3385 5850 3415
rect 5800 3365 5815 3385
rect 5835 3365 5850 3385
rect 5800 3350 5850 3365
rect 4900 3335 5850 3350
rect 4900 3315 4915 3335
rect 4935 3315 5850 3335
rect 4900 3300 5850 3315
rect 5950 3685 6000 3715
rect 6250 3735 6300 3750
rect 6250 3715 6265 3735
rect 6285 3715 6300 3735
rect 5950 3665 5965 3685
rect 5985 3665 6000 3685
rect 5950 3635 6000 3665
rect 5950 3615 5965 3635
rect 5985 3615 6000 3635
rect 5950 3585 6000 3615
rect 5950 3565 5965 3585
rect 5985 3565 6000 3585
rect 5950 3535 6000 3565
rect 5950 3515 5965 3535
rect 5985 3515 6000 3535
rect 5950 3485 6000 3515
rect 5950 3465 5965 3485
rect 5985 3465 6000 3485
rect 5950 3435 6000 3465
rect 5950 3415 5965 3435
rect 5985 3415 6000 3435
rect 5950 3385 6000 3415
rect 5950 3365 5965 3385
rect 5985 3365 6000 3385
rect 5950 3335 6000 3365
rect 5950 3315 5965 3335
rect 5985 3315 6000 3335
rect 4900 3240 4950 3250
rect 4900 3210 4910 3240
rect 4940 3210 4950 3240
rect 4900 3200 4950 3210
rect 5200 3240 5250 3250
rect 5200 3210 5210 3240
rect 5240 3210 5250 3240
rect 5200 3200 5250 3210
rect 5350 3240 5400 3300
rect 5350 3210 5360 3240
rect 5390 3210 5400 3240
rect 5350 3150 5400 3210
rect 5500 3240 5550 3250
rect 5500 3210 5510 3240
rect 5540 3210 5550 3240
rect 5500 3200 5550 3210
rect 5800 3240 5850 3250
rect 5800 3210 5810 3240
rect 5840 3210 5850 3240
rect 5800 3200 5850 3210
rect 4750 3115 4765 3135
rect 4785 3115 4800 3135
rect 4750 3085 4800 3115
rect 4750 3065 4765 3085
rect 4785 3065 4800 3085
rect 4750 3035 4800 3065
rect 4750 3015 4765 3035
rect 4785 3015 4800 3035
rect 4750 2985 4800 3015
rect 4750 2965 4765 2985
rect 4785 2965 4800 2985
rect 4750 2935 4800 2965
rect 4750 2915 4765 2935
rect 4785 2915 4800 2935
rect 4750 2885 4800 2915
rect 4750 2865 4765 2885
rect 4785 2865 4800 2885
rect 4750 2835 4800 2865
rect 4750 2815 4765 2835
rect 4785 2815 4800 2835
rect 4750 2785 4800 2815
rect 4750 2765 4765 2785
rect 4785 2765 4800 2785
rect 4750 2735 4800 2765
rect 4900 3135 5850 3150
rect 4900 3115 4915 3135
rect 4935 3115 5215 3135
rect 5235 3115 5515 3135
rect 5535 3115 5815 3135
rect 5835 3115 5850 3135
rect 4900 3100 5850 3115
rect 4900 3085 4950 3100
rect 4900 3065 4915 3085
rect 4935 3065 4950 3085
rect 4900 3035 4950 3065
rect 5200 3085 5250 3100
rect 5200 3065 5215 3085
rect 5235 3065 5250 3085
rect 4900 3015 4915 3035
rect 4935 3015 4950 3035
rect 4900 2985 4950 3015
rect 4900 2965 4915 2985
rect 4935 2965 4950 2985
rect 4900 2935 4950 2965
rect 4900 2915 4915 2935
rect 4935 2915 4950 2935
rect 4900 2885 4950 2915
rect 4900 2865 4915 2885
rect 4935 2865 4950 2885
rect 4900 2835 4950 2865
rect 4900 2815 4915 2835
rect 4935 2815 4950 2835
rect 4900 2785 4950 2815
rect 4900 2765 4915 2785
rect 4935 2765 4950 2785
rect 4900 2750 4950 2765
rect 5050 3035 5100 3050
rect 5050 3015 5065 3035
rect 5085 3015 5100 3035
rect 5050 2985 5100 3015
rect 5050 2965 5065 2985
rect 5085 2965 5100 2985
rect 5050 2935 5100 2965
rect 5050 2915 5065 2935
rect 5085 2915 5100 2935
rect 5050 2885 5100 2915
rect 5050 2865 5065 2885
rect 5085 2865 5100 2885
rect 5050 2835 5100 2865
rect 5050 2815 5065 2835
rect 5085 2815 5100 2835
rect 5050 2785 5100 2815
rect 5050 2765 5065 2785
rect 5085 2765 5100 2785
rect 4750 2715 4765 2735
rect 4785 2715 4800 2735
rect 4750 2700 4800 2715
rect 5050 2735 5100 2765
rect 5200 3035 5250 3065
rect 5500 3085 5550 3100
rect 5500 3065 5515 3085
rect 5535 3065 5550 3085
rect 5200 3015 5215 3035
rect 5235 3015 5250 3035
rect 5200 2985 5250 3015
rect 5200 2965 5215 2985
rect 5235 2965 5250 2985
rect 5200 2935 5250 2965
rect 5200 2915 5215 2935
rect 5235 2915 5250 2935
rect 5200 2885 5250 2915
rect 5200 2865 5215 2885
rect 5235 2865 5250 2885
rect 5200 2835 5250 2865
rect 5200 2815 5215 2835
rect 5235 2815 5250 2835
rect 5200 2785 5250 2815
rect 5200 2765 5215 2785
rect 5235 2765 5250 2785
rect 5200 2750 5250 2765
rect 5350 3035 5400 3050
rect 5350 3015 5365 3035
rect 5385 3015 5400 3035
rect 5350 2985 5400 3015
rect 5350 2965 5365 2985
rect 5385 2965 5400 2985
rect 5350 2935 5400 2965
rect 5350 2915 5365 2935
rect 5385 2915 5400 2935
rect 5350 2885 5400 2915
rect 5350 2865 5365 2885
rect 5385 2865 5400 2885
rect 5350 2835 5400 2865
rect 5350 2815 5365 2835
rect 5385 2815 5400 2835
rect 5350 2785 5400 2815
rect 5350 2765 5365 2785
rect 5385 2765 5400 2785
rect 5050 2715 5065 2735
rect 5085 2715 5100 2735
rect 5050 2700 5100 2715
rect 5350 2735 5400 2765
rect 5500 3035 5550 3065
rect 5800 3085 5850 3100
rect 5800 3065 5815 3085
rect 5835 3065 5850 3085
rect 5500 3015 5515 3035
rect 5535 3015 5550 3035
rect 5500 2985 5550 3015
rect 5500 2965 5515 2985
rect 5535 2965 5550 2985
rect 5500 2935 5550 2965
rect 5500 2915 5515 2935
rect 5535 2915 5550 2935
rect 5500 2885 5550 2915
rect 5500 2865 5515 2885
rect 5535 2865 5550 2885
rect 5500 2835 5550 2865
rect 5500 2815 5515 2835
rect 5535 2815 5550 2835
rect 5500 2785 5550 2815
rect 5500 2765 5515 2785
rect 5535 2765 5550 2785
rect 5500 2750 5550 2765
rect 5650 3035 5700 3050
rect 5650 3015 5665 3035
rect 5685 3015 5700 3035
rect 5650 2985 5700 3015
rect 5650 2965 5665 2985
rect 5685 2965 5700 2985
rect 5650 2935 5700 2965
rect 5650 2915 5665 2935
rect 5685 2915 5700 2935
rect 5650 2885 5700 2915
rect 5650 2865 5665 2885
rect 5685 2865 5700 2885
rect 5650 2835 5700 2865
rect 5650 2815 5665 2835
rect 5685 2815 5700 2835
rect 5650 2785 5700 2815
rect 5650 2765 5665 2785
rect 5685 2765 5700 2785
rect 5350 2715 5365 2735
rect 5385 2715 5400 2735
rect 5350 2700 5400 2715
rect 5650 2735 5700 2765
rect 5800 3035 5850 3065
rect 5800 3015 5815 3035
rect 5835 3015 5850 3035
rect 5800 2985 5850 3015
rect 5800 2965 5815 2985
rect 5835 2965 5850 2985
rect 5800 2935 5850 2965
rect 5800 2915 5815 2935
rect 5835 2915 5850 2935
rect 5800 2885 5850 2915
rect 5800 2865 5815 2885
rect 5835 2865 5850 2885
rect 5800 2835 5850 2865
rect 5800 2815 5815 2835
rect 5835 2815 5850 2835
rect 5800 2785 5850 2815
rect 5800 2765 5815 2785
rect 5835 2765 5850 2785
rect 5800 2750 5850 2765
rect 5950 3135 6000 3315
rect 6100 3685 6150 3700
rect 6100 3665 6115 3685
rect 6135 3665 6150 3685
rect 6100 3635 6150 3665
rect 6100 3615 6115 3635
rect 6135 3615 6150 3635
rect 6100 3585 6150 3615
rect 6100 3565 6115 3585
rect 6135 3565 6150 3585
rect 6100 3535 6150 3565
rect 6100 3515 6115 3535
rect 6135 3515 6150 3535
rect 6100 3485 6150 3515
rect 6100 3465 6115 3485
rect 6135 3465 6150 3485
rect 6100 3435 6150 3465
rect 6100 3415 6115 3435
rect 6135 3415 6150 3435
rect 6100 3385 6150 3415
rect 6250 3685 6300 3715
rect 6550 3735 6600 3750
rect 6550 3715 6565 3735
rect 6585 3715 6600 3735
rect 6250 3665 6265 3685
rect 6285 3665 6300 3685
rect 6250 3635 6300 3665
rect 6250 3615 6265 3635
rect 6285 3615 6300 3635
rect 6250 3585 6300 3615
rect 6250 3565 6265 3585
rect 6285 3565 6300 3585
rect 6250 3535 6300 3565
rect 6250 3515 6265 3535
rect 6285 3515 6300 3535
rect 6250 3485 6300 3515
rect 6250 3465 6265 3485
rect 6285 3465 6300 3485
rect 6250 3435 6300 3465
rect 6250 3415 6265 3435
rect 6285 3415 6300 3435
rect 6250 3400 6300 3415
rect 6400 3685 6450 3700
rect 6400 3665 6415 3685
rect 6435 3665 6450 3685
rect 6400 3635 6450 3665
rect 6400 3615 6415 3635
rect 6435 3615 6450 3635
rect 6400 3585 6450 3615
rect 6400 3565 6415 3585
rect 6435 3565 6450 3585
rect 6400 3535 6450 3565
rect 6400 3515 6415 3535
rect 6435 3515 6450 3535
rect 6400 3485 6450 3515
rect 6400 3465 6415 3485
rect 6435 3465 6450 3485
rect 6400 3435 6450 3465
rect 6400 3415 6415 3435
rect 6435 3415 6450 3435
rect 6100 3365 6115 3385
rect 6135 3365 6150 3385
rect 6100 3350 6150 3365
rect 6400 3385 6450 3415
rect 6400 3365 6415 3385
rect 6435 3365 6450 3385
rect 6400 3350 6450 3365
rect 6100 3335 6450 3350
rect 6100 3315 6115 3335
rect 6135 3315 6415 3335
rect 6435 3315 6450 3335
rect 6100 3300 6450 3315
rect 6550 3685 6600 3715
rect 6850 3735 6900 3750
rect 6850 3715 6865 3735
rect 6885 3715 6900 3735
rect 6550 3665 6565 3685
rect 6585 3665 6600 3685
rect 6550 3635 6600 3665
rect 6550 3615 6565 3635
rect 6585 3615 6600 3635
rect 6550 3585 6600 3615
rect 6550 3565 6565 3585
rect 6585 3565 6600 3585
rect 6550 3535 6600 3565
rect 6550 3515 6565 3535
rect 6585 3515 6600 3535
rect 6550 3485 6600 3515
rect 6550 3465 6565 3485
rect 6585 3465 6600 3485
rect 6550 3435 6600 3465
rect 6550 3415 6565 3435
rect 6585 3415 6600 3435
rect 6550 3385 6600 3415
rect 6550 3365 6565 3385
rect 6585 3365 6600 3385
rect 6550 3335 6600 3365
rect 6550 3315 6565 3335
rect 6585 3315 6600 3335
rect 6100 3240 6150 3250
rect 6100 3210 6110 3240
rect 6140 3210 6150 3240
rect 6100 3200 6150 3210
rect 6250 3240 6300 3300
rect 6250 3210 6260 3240
rect 6290 3210 6300 3240
rect 6250 3150 6300 3210
rect 6400 3240 6450 3250
rect 6400 3210 6410 3240
rect 6440 3210 6450 3240
rect 6400 3200 6450 3210
rect 5950 3115 5965 3135
rect 5985 3115 6000 3135
rect 5950 3085 6000 3115
rect 5950 3065 5965 3085
rect 5985 3065 6000 3085
rect 5950 3035 6000 3065
rect 5950 3015 5965 3035
rect 5985 3015 6000 3035
rect 5950 2985 6000 3015
rect 5950 2965 5965 2985
rect 5985 2965 6000 2985
rect 5950 2935 6000 2965
rect 5950 2915 5965 2935
rect 5985 2915 6000 2935
rect 5950 2885 6000 2915
rect 5950 2865 5965 2885
rect 5985 2865 6000 2885
rect 5950 2835 6000 2865
rect 5950 2815 5965 2835
rect 5985 2815 6000 2835
rect 5950 2785 6000 2815
rect 5950 2765 5965 2785
rect 5985 2765 6000 2785
rect 5650 2715 5665 2735
rect 5685 2715 5700 2735
rect 5650 2700 5700 2715
rect 5950 2735 6000 2765
rect 6100 3135 6450 3150
rect 6100 3115 6115 3135
rect 6135 3115 6415 3135
rect 6435 3115 6450 3135
rect 6100 3100 6450 3115
rect 6100 3085 6150 3100
rect 6100 3065 6115 3085
rect 6135 3065 6150 3085
rect 6100 3035 6150 3065
rect 6400 3085 6450 3100
rect 6400 3065 6415 3085
rect 6435 3065 6450 3085
rect 6100 3015 6115 3035
rect 6135 3015 6150 3035
rect 6100 2985 6150 3015
rect 6100 2965 6115 2985
rect 6135 2965 6150 2985
rect 6100 2935 6150 2965
rect 6100 2915 6115 2935
rect 6135 2915 6150 2935
rect 6100 2885 6150 2915
rect 6100 2865 6115 2885
rect 6135 2865 6150 2885
rect 6100 2835 6150 2865
rect 6100 2815 6115 2835
rect 6135 2815 6150 2835
rect 6100 2785 6150 2815
rect 6100 2765 6115 2785
rect 6135 2765 6150 2785
rect 6100 2750 6150 2765
rect 6250 3035 6300 3050
rect 6250 3015 6265 3035
rect 6285 3015 6300 3035
rect 6250 2985 6300 3015
rect 6250 2965 6265 2985
rect 6285 2965 6300 2985
rect 6250 2935 6300 2965
rect 6250 2915 6265 2935
rect 6285 2915 6300 2935
rect 6250 2885 6300 2915
rect 6250 2865 6265 2885
rect 6285 2865 6300 2885
rect 6250 2835 6300 2865
rect 6250 2815 6265 2835
rect 6285 2815 6300 2835
rect 6250 2785 6300 2815
rect 6250 2765 6265 2785
rect 6285 2765 6300 2785
rect 5950 2715 5965 2735
rect 5985 2715 6000 2735
rect 5950 2700 6000 2715
rect 6250 2735 6300 2765
rect 6400 3035 6450 3065
rect 6400 3015 6415 3035
rect 6435 3015 6450 3035
rect 6400 2985 6450 3015
rect 6400 2965 6415 2985
rect 6435 2965 6450 2985
rect 6400 2935 6450 2965
rect 6400 2915 6415 2935
rect 6435 2915 6450 2935
rect 6400 2885 6450 2915
rect 6400 2865 6415 2885
rect 6435 2865 6450 2885
rect 6400 2835 6450 2865
rect 6400 2815 6415 2835
rect 6435 2815 6450 2835
rect 6400 2785 6450 2815
rect 6400 2765 6415 2785
rect 6435 2765 6450 2785
rect 6400 2750 6450 2765
rect 6550 3135 6600 3315
rect 6700 3685 6750 3700
rect 6700 3665 6715 3685
rect 6735 3665 6750 3685
rect 6700 3635 6750 3665
rect 6700 3615 6715 3635
rect 6735 3615 6750 3635
rect 6700 3585 6750 3615
rect 6700 3565 6715 3585
rect 6735 3565 6750 3585
rect 6700 3535 6750 3565
rect 6700 3515 6715 3535
rect 6735 3515 6750 3535
rect 6700 3485 6750 3515
rect 6700 3465 6715 3485
rect 6735 3465 6750 3485
rect 6700 3435 6750 3465
rect 6700 3415 6715 3435
rect 6735 3415 6750 3435
rect 6700 3385 6750 3415
rect 6850 3685 6900 3715
rect 7150 3735 7200 3750
rect 7150 3715 7165 3735
rect 7185 3715 7200 3735
rect 6850 3665 6865 3685
rect 6885 3665 6900 3685
rect 6850 3635 6900 3665
rect 6850 3615 6865 3635
rect 6885 3615 6900 3635
rect 6850 3585 6900 3615
rect 6850 3565 6865 3585
rect 6885 3565 6900 3585
rect 6850 3535 6900 3565
rect 6850 3515 6865 3535
rect 6885 3515 6900 3535
rect 6850 3485 6900 3515
rect 6850 3465 6865 3485
rect 6885 3465 6900 3485
rect 6850 3435 6900 3465
rect 6850 3415 6865 3435
rect 6885 3415 6900 3435
rect 6850 3400 6900 3415
rect 7000 3685 7050 3700
rect 7000 3665 7015 3685
rect 7035 3665 7050 3685
rect 7000 3635 7050 3665
rect 7000 3615 7015 3635
rect 7035 3615 7050 3635
rect 7000 3585 7050 3615
rect 7000 3565 7015 3585
rect 7035 3565 7050 3585
rect 7000 3535 7050 3565
rect 7000 3515 7015 3535
rect 7035 3515 7050 3535
rect 7000 3485 7050 3515
rect 7000 3465 7015 3485
rect 7035 3465 7050 3485
rect 7000 3435 7050 3465
rect 7000 3415 7015 3435
rect 7035 3415 7050 3435
rect 6700 3365 6715 3385
rect 6735 3365 6750 3385
rect 6700 3350 6750 3365
rect 7000 3385 7050 3415
rect 7150 3685 7200 3715
rect 7450 3735 7500 3750
rect 7450 3715 7465 3735
rect 7485 3715 7500 3735
rect 7150 3665 7165 3685
rect 7185 3665 7200 3685
rect 7150 3635 7200 3665
rect 7150 3615 7165 3635
rect 7185 3615 7200 3635
rect 7150 3585 7200 3615
rect 7150 3565 7165 3585
rect 7185 3565 7200 3585
rect 7150 3535 7200 3565
rect 7150 3515 7165 3535
rect 7185 3515 7200 3535
rect 7150 3485 7200 3515
rect 7150 3465 7165 3485
rect 7185 3465 7200 3485
rect 7150 3435 7200 3465
rect 7150 3415 7165 3435
rect 7185 3415 7200 3435
rect 7150 3400 7200 3415
rect 7300 3685 7350 3700
rect 7300 3665 7315 3685
rect 7335 3665 7350 3685
rect 7300 3635 7350 3665
rect 7300 3615 7315 3635
rect 7335 3615 7350 3635
rect 7300 3585 7350 3615
rect 7300 3565 7315 3585
rect 7335 3565 7350 3585
rect 7300 3535 7350 3565
rect 7300 3515 7315 3535
rect 7335 3515 7350 3535
rect 7300 3485 7350 3515
rect 7300 3465 7315 3485
rect 7335 3465 7350 3485
rect 7300 3435 7350 3465
rect 7300 3415 7315 3435
rect 7335 3415 7350 3435
rect 7000 3365 7015 3385
rect 7035 3365 7050 3385
rect 7000 3350 7050 3365
rect 7300 3385 7350 3415
rect 7450 3685 7500 3715
rect 7750 3735 7800 3750
rect 7750 3715 7765 3735
rect 7785 3715 7800 3735
rect 7450 3665 7465 3685
rect 7485 3665 7500 3685
rect 7450 3635 7500 3665
rect 7450 3615 7465 3635
rect 7485 3615 7500 3635
rect 7450 3585 7500 3615
rect 7450 3565 7465 3585
rect 7485 3565 7500 3585
rect 7450 3535 7500 3565
rect 7450 3515 7465 3535
rect 7485 3515 7500 3535
rect 7450 3485 7500 3515
rect 7450 3465 7465 3485
rect 7485 3465 7500 3485
rect 7450 3435 7500 3465
rect 7450 3415 7465 3435
rect 7485 3415 7500 3435
rect 7450 3400 7500 3415
rect 7600 3685 7650 3700
rect 7600 3665 7615 3685
rect 7635 3665 7650 3685
rect 7600 3635 7650 3665
rect 7600 3615 7615 3635
rect 7635 3615 7650 3635
rect 7600 3585 7650 3615
rect 7600 3565 7615 3585
rect 7635 3565 7650 3585
rect 7600 3535 7650 3565
rect 7600 3515 7615 3535
rect 7635 3515 7650 3535
rect 7600 3485 7650 3515
rect 7600 3465 7615 3485
rect 7635 3465 7650 3485
rect 7600 3435 7650 3465
rect 7600 3415 7615 3435
rect 7635 3415 7650 3435
rect 7300 3365 7315 3385
rect 7335 3365 7350 3385
rect 7300 3350 7350 3365
rect 7600 3385 7650 3415
rect 7600 3365 7615 3385
rect 7635 3365 7650 3385
rect 7600 3350 7650 3365
rect 6700 3335 7650 3350
rect 6700 3315 7615 3335
rect 7635 3315 7650 3335
rect 6700 3300 7650 3315
rect 7750 3685 7800 3715
rect 7750 3665 7765 3685
rect 7785 3665 7800 3685
rect 7750 3635 7800 3665
rect 7750 3615 7765 3635
rect 7785 3615 7800 3635
rect 7750 3585 7800 3615
rect 7750 3565 7765 3585
rect 7785 3565 7800 3585
rect 7750 3535 7800 3565
rect 7750 3515 7765 3535
rect 7785 3515 7800 3535
rect 7750 3485 7800 3515
rect 7750 3465 7765 3485
rect 7785 3465 7800 3485
rect 7750 3435 7800 3465
rect 7750 3415 7765 3435
rect 7785 3415 7800 3435
rect 7750 3385 7800 3415
rect 7750 3365 7765 3385
rect 7785 3365 7800 3385
rect 7750 3335 7800 3365
rect 7750 3315 7765 3335
rect 7785 3315 7800 3335
rect 6700 3240 6750 3250
rect 6700 3210 6710 3240
rect 6740 3210 6750 3240
rect 6700 3200 6750 3210
rect 7000 3240 7050 3250
rect 7000 3210 7010 3240
rect 7040 3210 7050 3240
rect 7000 3200 7050 3210
rect 7150 3240 7200 3300
rect 7150 3210 7160 3240
rect 7190 3210 7200 3240
rect 7150 3150 7200 3210
rect 7300 3240 7350 3250
rect 7300 3210 7310 3240
rect 7340 3210 7350 3240
rect 7300 3200 7350 3210
rect 7600 3240 7650 3250
rect 7600 3210 7610 3240
rect 7640 3210 7650 3240
rect 7600 3200 7650 3210
rect 6550 3115 6565 3135
rect 6585 3115 6600 3135
rect 6550 3085 6600 3115
rect 6550 3065 6565 3085
rect 6585 3065 6600 3085
rect 6550 3035 6600 3065
rect 6550 3015 6565 3035
rect 6585 3015 6600 3035
rect 6550 2985 6600 3015
rect 6550 2965 6565 2985
rect 6585 2965 6600 2985
rect 6550 2935 6600 2965
rect 6550 2915 6565 2935
rect 6585 2915 6600 2935
rect 6550 2885 6600 2915
rect 6550 2865 6565 2885
rect 6585 2865 6600 2885
rect 6550 2835 6600 2865
rect 6550 2815 6565 2835
rect 6585 2815 6600 2835
rect 6550 2785 6600 2815
rect 6550 2765 6565 2785
rect 6585 2765 6600 2785
rect 6250 2715 6265 2735
rect 6285 2715 6300 2735
rect 6250 2700 6300 2715
rect 6550 2735 6600 2765
rect 6700 3135 7650 3150
rect 6700 3115 6715 3135
rect 6735 3115 7015 3135
rect 7035 3115 7315 3135
rect 7335 3115 7615 3135
rect 7635 3115 7650 3135
rect 6700 3100 7650 3115
rect 6700 3085 6750 3100
rect 6700 3065 6715 3085
rect 6735 3065 6750 3085
rect 6700 3035 6750 3065
rect 7000 3085 7050 3100
rect 7000 3065 7015 3085
rect 7035 3065 7050 3085
rect 6700 3015 6715 3035
rect 6735 3015 6750 3035
rect 6700 2985 6750 3015
rect 6700 2965 6715 2985
rect 6735 2965 6750 2985
rect 6700 2935 6750 2965
rect 6700 2915 6715 2935
rect 6735 2915 6750 2935
rect 6700 2885 6750 2915
rect 6700 2865 6715 2885
rect 6735 2865 6750 2885
rect 6700 2835 6750 2865
rect 6700 2815 6715 2835
rect 6735 2815 6750 2835
rect 6700 2785 6750 2815
rect 6700 2765 6715 2785
rect 6735 2765 6750 2785
rect 6700 2750 6750 2765
rect 6850 3035 6900 3050
rect 6850 3015 6865 3035
rect 6885 3015 6900 3035
rect 6850 2985 6900 3015
rect 6850 2965 6865 2985
rect 6885 2965 6900 2985
rect 6850 2935 6900 2965
rect 6850 2915 6865 2935
rect 6885 2915 6900 2935
rect 6850 2885 6900 2915
rect 6850 2865 6865 2885
rect 6885 2865 6900 2885
rect 6850 2835 6900 2865
rect 6850 2815 6865 2835
rect 6885 2815 6900 2835
rect 6850 2785 6900 2815
rect 6850 2765 6865 2785
rect 6885 2765 6900 2785
rect 6550 2715 6565 2735
rect 6585 2715 6600 2735
rect 6550 2700 6600 2715
rect 6850 2735 6900 2765
rect 7000 3035 7050 3065
rect 7300 3085 7350 3100
rect 7300 3065 7315 3085
rect 7335 3065 7350 3085
rect 7000 3015 7015 3035
rect 7035 3015 7050 3035
rect 7000 2985 7050 3015
rect 7000 2965 7015 2985
rect 7035 2965 7050 2985
rect 7000 2935 7050 2965
rect 7000 2915 7015 2935
rect 7035 2915 7050 2935
rect 7000 2885 7050 2915
rect 7000 2865 7015 2885
rect 7035 2865 7050 2885
rect 7000 2835 7050 2865
rect 7000 2815 7015 2835
rect 7035 2815 7050 2835
rect 7000 2785 7050 2815
rect 7000 2765 7015 2785
rect 7035 2765 7050 2785
rect 7000 2750 7050 2765
rect 7150 3035 7200 3050
rect 7150 3015 7165 3035
rect 7185 3015 7200 3035
rect 7150 2985 7200 3015
rect 7150 2965 7165 2985
rect 7185 2965 7200 2985
rect 7150 2935 7200 2965
rect 7150 2915 7165 2935
rect 7185 2915 7200 2935
rect 7150 2885 7200 2915
rect 7150 2865 7165 2885
rect 7185 2865 7200 2885
rect 7150 2835 7200 2865
rect 7150 2815 7165 2835
rect 7185 2815 7200 2835
rect 7150 2785 7200 2815
rect 7150 2765 7165 2785
rect 7185 2765 7200 2785
rect 6850 2715 6865 2735
rect 6885 2715 6900 2735
rect 6850 2700 6900 2715
rect 7150 2735 7200 2765
rect 7300 3035 7350 3065
rect 7600 3085 7650 3100
rect 7600 3065 7615 3085
rect 7635 3065 7650 3085
rect 7300 3015 7315 3035
rect 7335 3015 7350 3035
rect 7300 2985 7350 3015
rect 7300 2965 7315 2985
rect 7335 2965 7350 2985
rect 7300 2935 7350 2965
rect 7300 2915 7315 2935
rect 7335 2915 7350 2935
rect 7300 2885 7350 2915
rect 7300 2865 7315 2885
rect 7335 2865 7350 2885
rect 7300 2835 7350 2865
rect 7300 2815 7315 2835
rect 7335 2815 7350 2835
rect 7300 2785 7350 2815
rect 7300 2765 7315 2785
rect 7335 2765 7350 2785
rect 7300 2750 7350 2765
rect 7450 3035 7500 3050
rect 7450 3015 7465 3035
rect 7485 3015 7500 3035
rect 7450 2985 7500 3015
rect 7450 2965 7465 2985
rect 7485 2965 7500 2985
rect 7450 2935 7500 2965
rect 7450 2915 7465 2935
rect 7485 2915 7500 2935
rect 7450 2885 7500 2915
rect 7450 2865 7465 2885
rect 7485 2865 7500 2885
rect 7450 2835 7500 2865
rect 7450 2815 7465 2835
rect 7485 2815 7500 2835
rect 7450 2785 7500 2815
rect 7450 2765 7465 2785
rect 7485 2765 7500 2785
rect 7150 2715 7165 2735
rect 7185 2715 7200 2735
rect 7150 2700 7200 2715
rect 7450 2735 7500 2765
rect 7600 3035 7650 3065
rect 7600 3015 7615 3035
rect 7635 3015 7650 3035
rect 7600 2985 7650 3015
rect 7600 2965 7615 2985
rect 7635 2965 7650 2985
rect 7600 2935 7650 2965
rect 7600 2915 7615 2935
rect 7635 2915 7650 2935
rect 7600 2885 7650 2915
rect 7600 2865 7615 2885
rect 7635 2865 7650 2885
rect 7600 2835 7650 2865
rect 7600 2815 7615 2835
rect 7635 2815 7650 2835
rect 7600 2785 7650 2815
rect 7600 2765 7615 2785
rect 7635 2765 7650 2785
rect 7600 2750 7650 2765
rect 7750 3135 7800 3315
rect 8350 3785 8400 3860
rect 8650 3890 8700 3965
rect 8800 4435 8850 4450
rect 8800 4415 8815 4435
rect 8835 4415 8850 4435
rect 8800 4385 8850 4415
rect 8800 4365 8815 4385
rect 8835 4365 8850 4385
rect 8800 4335 8850 4365
rect 8800 4315 8815 4335
rect 8835 4315 8850 4335
rect 8800 4285 8850 4315
rect 8800 4265 8815 4285
rect 8835 4265 8850 4285
rect 8800 4235 8850 4265
rect 8800 4215 8815 4235
rect 8835 4215 8850 4235
rect 8800 4185 8850 4215
rect 8800 4165 8815 4185
rect 8835 4165 8850 4185
rect 8800 4135 8850 4165
rect 8800 4115 8815 4135
rect 8835 4115 8850 4135
rect 8800 4085 8850 4115
rect 8800 4065 8815 4085
rect 8835 4065 8850 4085
rect 8800 4035 8850 4065
rect 8800 4015 8815 4035
rect 8835 4015 8850 4035
rect 8800 3985 8850 4015
rect 8800 3965 8815 3985
rect 8835 3965 8850 3985
rect 8800 3950 8850 3965
rect 8950 4440 9000 4610
rect 9100 5085 9150 5100
rect 9100 5065 9115 5085
rect 9135 5065 9150 5085
rect 9100 5035 9150 5065
rect 9100 5015 9115 5035
rect 9135 5015 9150 5035
rect 9100 4985 9150 5015
rect 9100 4965 9115 4985
rect 9135 4965 9150 4985
rect 9100 4935 9150 4965
rect 9100 4915 9115 4935
rect 9135 4915 9150 4935
rect 9100 4885 9150 4915
rect 9100 4865 9115 4885
rect 9135 4865 9150 4885
rect 9100 4835 9150 4865
rect 9100 4815 9115 4835
rect 9135 4815 9150 4835
rect 9100 4785 9150 4815
rect 9100 4765 9115 4785
rect 9135 4765 9150 4785
rect 9100 4735 9150 4765
rect 9100 4715 9115 4735
rect 9135 4715 9150 4735
rect 9100 4685 9150 4715
rect 9100 4665 9115 4685
rect 9135 4665 9150 4685
rect 9100 4635 9150 4665
rect 9100 4615 9115 4635
rect 9135 4615 9150 4635
rect 9100 4600 9150 4615
rect 9250 5085 9300 5160
rect 9550 5190 9600 5200
rect 9550 5160 9560 5190
rect 9590 5160 9600 5190
rect 9250 5065 9265 5085
rect 9285 5065 9300 5085
rect 9250 5040 9300 5065
rect 9250 5010 9260 5040
rect 9290 5010 9300 5040
rect 9250 4985 9300 5010
rect 9250 4965 9265 4985
rect 9285 4965 9300 4985
rect 9250 4940 9300 4965
rect 9250 4910 9260 4940
rect 9290 4910 9300 4940
rect 9250 4885 9300 4910
rect 9250 4865 9265 4885
rect 9285 4865 9300 4885
rect 9250 4840 9300 4865
rect 9250 4810 9260 4840
rect 9290 4810 9300 4840
rect 9250 4785 9300 4810
rect 9250 4765 9265 4785
rect 9285 4765 9300 4785
rect 9250 4740 9300 4765
rect 9250 4710 9260 4740
rect 9290 4710 9300 4740
rect 9250 4685 9300 4710
rect 9250 4665 9265 4685
rect 9285 4665 9300 4685
rect 9250 4640 9300 4665
rect 9250 4610 9260 4640
rect 9290 4610 9300 4640
rect 9100 4540 9150 4550
rect 9100 4510 9110 4540
rect 9140 4510 9150 4540
rect 9100 4500 9150 4510
rect 8950 4410 8960 4440
rect 8990 4410 9000 4440
rect 8950 4385 9000 4410
rect 8950 4365 8965 4385
rect 8985 4365 9000 4385
rect 8950 4340 9000 4365
rect 8950 4310 8960 4340
rect 8990 4310 9000 4340
rect 8950 4285 9000 4310
rect 8950 4265 8965 4285
rect 8985 4265 9000 4285
rect 8950 4240 9000 4265
rect 8950 4210 8960 4240
rect 8990 4210 9000 4240
rect 8950 4185 9000 4210
rect 8950 4165 8965 4185
rect 8985 4165 9000 4185
rect 8950 4140 9000 4165
rect 8950 4110 8960 4140
rect 8990 4110 9000 4140
rect 8950 4085 9000 4110
rect 8950 4065 8965 4085
rect 8985 4065 9000 4085
rect 8950 4040 9000 4065
rect 8950 4010 8960 4040
rect 8990 4010 9000 4040
rect 8950 3985 9000 4010
rect 8950 3965 8965 3985
rect 8985 3965 9000 3985
rect 8650 3860 8660 3890
rect 8690 3860 8700 3890
rect 8350 3765 8365 3785
rect 8385 3765 8400 3785
rect 8350 3740 8400 3765
rect 8350 3710 8360 3740
rect 8390 3710 8400 3740
rect 8350 3685 8400 3710
rect 8350 3665 8365 3685
rect 8385 3665 8400 3685
rect 8350 3640 8400 3665
rect 8350 3610 8360 3640
rect 8390 3610 8400 3640
rect 8350 3585 8400 3610
rect 8350 3565 8365 3585
rect 8385 3565 8400 3585
rect 8350 3540 8400 3565
rect 8350 3510 8360 3540
rect 8390 3510 8400 3540
rect 8350 3485 8400 3510
rect 8350 3465 8365 3485
rect 8385 3465 8400 3485
rect 8350 3440 8400 3465
rect 8350 3410 8360 3440
rect 8390 3410 8400 3440
rect 8350 3385 8400 3410
rect 8350 3365 8365 3385
rect 8385 3365 8400 3385
rect 8350 3340 8400 3365
rect 8350 3310 8360 3340
rect 8390 3310 8400 3340
rect 7900 3240 7950 3250
rect 7900 3210 7910 3240
rect 7940 3210 7950 3240
rect 7900 3200 7950 3210
rect 8200 3240 8250 3250
rect 8200 3210 8210 3240
rect 8240 3210 8250 3240
rect 8200 3200 8250 3210
rect 7750 3115 7765 3135
rect 7785 3115 7800 3135
rect 7750 3085 7800 3115
rect 7750 3065 7765 3085
rect 7785 3065 7800 3085
rect 7750 3035 7800 3065
rect 7750 3015 7765 3035
rect 7785 3015 7800 3035
rect 7750 2985 7800 3015
rect 7750 2965 7765 2985
rect 7785 2965 7800 2985
rect 7750 2935 7800 2965
rect 7750 2915 7765 2935
rect 7785 2915 7800 2935
rect 7750 2885 7800 2915
rect 7750 2865 7765 2885
rect 7785 2865 7800 2885
rect 7750 2835 7800 2865
rect 7750 2815 7765 2835
rect 7785 2815 7800 2835
rect 7750 2785 7800 2815
rect 7750 2765 7765 2785
rect 7785 2765 7800 2785
rect 7450 2715 7465 2735
rect 7485 2715 7500 2735
rect 7450 2700 7500 2715
rect 7750 2735 7800 2765
rect 7750 2715 7765 2735
rect 7785 2715 7800 2735
rect 7750 2700 7800 2715
rect 4750 2685 7800 2700
rect 4750 2665 4765 2685
rect 4785 2665 5065 2685
rect 5085 2665 5365 2685
rect 5385 2665 5665 2685
rect 5685 2665 5965 2685
rect 5985 2665 6265 2685
rect 6285 2665 6565 2685
rect 6585 2665 6865 2685
rect 6885 2665 7165 2685
rect 7185 2665 7465 2685
rect 7485 2665 7765 2685
rect 7785 2665 7800 2685
rect 4750 2650 7800 2665
rect 8350 3140 8400 3310
rect 8500 3785 8550 3800
rect 8500 3765 8515 3785
rect 8535 3765 8550 3785
rect 8500 3735 8550 3765
rect 8500 3715 8515 3735
rect 8535 3715 8550 3735
rect 8500 3685 8550 3715
rect 8500 3665 8515 3685
rect 8535 3665 8550 3685
rect 8500 3635 8550 3665
rect 8500 3615 8515 3635
rect 8535 3615 8550 3635
rect 8500 3585 8550 3615
rect 8500 3565 8515 3585
rect 8535 3565 8550 3585
rect 8500 3535 8550 3565
rect 8500 3515 8515 3535
rect 8535 3515 8550 3535
rect 8500 3485 8550 3515
rect 8500 3465 8515 3485
rect 8535 3465 8550 3485
rect 8500 3435 8550 3465
rect 8500 3415 8515 3435
rect 8535 3415 8550 3435
rect 8500 3385 8550 3415
rect 8500 3365 8515 3385
rect 8535 3365 8550 3385
rect 8500 3335 8550 3365
rect 8500 3315 8515 3335
rect 8535 3315 8550 3335
rect 8500 3300 8550 3315
rect 8650 3785 8700 3860
rect 8950 3890 9000 3965
rect 9100 4435 9150 4450
rect 9100 4415 9115 4435
rect 9135 4415 9150 4435
rect 9100 4385 9150 4415
rect 9100 4365 9115 4385
rect 9135 4365 9150 4385
rect 9100 4335 9150 4365
rect 9100 4315 9115 4335
rect 9135 4315 9150 4335
rect 9100 4285 9150 4315
rect 9100 4265 9115 4285
rect 9135 4265 9150 4285
rect 9100 4235 9150 4265
rect 9100 4215 9115 4235
rect 9135 4215 9150 4235
rect 9100 4185 9150 4215
rect 9100 4165 9115 4185
rect 9135 4165 9150 4185
rect 9100 4135 9150 4165
rect 9100 4115 9115 4135
rect 9135 4115 9150 4135
rect 9100 4085 9150 4115
rect 9100 4065 9115 4085
rect 9135 4065 9150 4085
rect 9100 4035 9150 4065
rect 9100 4015 9115 4035
rect 9135 4015 9150 4035
rect 9100 3985 9150 4015
rect 9100 3965 9115 3985
rect 9135 3965 9150 3985
rect 9100 3950 9150 3965
rect 9250 4440 9300 4610
rect 9400 5085 9450 5100
rect 9400 5065 9415 5085
rect 9435 5065 9450 5085
rect 9400 5035 9450 5065
rect 9400 5015 9415 5035
rect 9435 5015 9450 5035
rect 9400 4985 9450 5015
rect 9400 4965 9415 4985
rect 9435 4965 9450 4985
rect 9400 4935 9450 4965
rect 9400 4915 9415 4935
rect 9435 4915 9450 4935
rect 9400 4885 9450 4915
rect 9400 4865 9415 4885
rect 9435 4865 9450 4885
rect 9400 4835 9450 4865
rect 9400 4815 9415 4835
rect 9435 4815 9450 4835
rect 9400 4785 9450 4815
rect 9400 4765 9415 4785
rect 9435 4765 9450 4785
rect 9400 4735 9450 4765
rect 9400 4715 9415 4735
rect 9435 4715 9450 4735
rect 9400 4685 9450 4715
rect 9400 4665 9415 4685
rect 9435 4665 9450 4685
rect 9400 4635 9450 4665
rect 9400 4615 9415 4635
rect 9435 4615 9450 4635
rect 9400 4600 9450 4615
rect 9550 5085 9600 5160
rect 9850 5190 9900 5200
rect 9850 5160 9860 5190
rect 9890 5160 9900 5190
rect 9550 5065 9565 5085
rect 9585 5065 9600 5085
rect 9550 5040 9600 5065
rect 9550 5010 9560 5040
rect 9590 5010 9600 5040
rect 9550 4985 9600 5010
rect 9550 4965 9565 4985
rect 9585 4965 9600 4985
rect 9550 4940 9600 4965
rect 9550 4910 9560 4940
rect 9590 4910 9600 4940
rect 9550 4885 9600 4910
rect 9550 4865 9565 4885
rect 9585 4865 9600 4885
rect 9550 4840 9600 4865
rect 9550 4810 9560 4840
rect 9590 4810 9600 4840
rect 9550 4785 9600 4810
rect 9550 4765 9565 4785
rect 9585 4765 9600 4785
rect 9550 4740 9600 4765
rect 9550 4710 9560 4740
rect 9590 4710 9600 4740
rect 9550 4685 9600 4710
rect 9550 4665 9565 4685
rect 9585 4665 9600 4685
rect 9550 4640 9600 4665
rect 9550 4610 9560 4640
rect 9590 4610 9600 4640
rect 9400 4540 9450 4550
rect 9400 4510 9410 4540
rect 9440 4510 9450 4540
rect 9400 4500 9450 4510
rect 9250 4410 9260 4440
rect 9290 4410 9300 4440
rect 9250 4385 9300 4410
rect 9250 4365 9265 4385
rect 9285 4365 9300 4385
rect 9250 4340 9300 4365
rect 9250 4310 9260 4340
rect 9290 4310 9300 4340
rect 9250 4285 9300 4310
rect 9250 4265 9265 4285
rect 9285 4265 9300 4285
rect 9250 4240 9300 4265
rect 9250 4210 9260 4240
rect 9290 4210 9300 4240
rect 9250 4185 9300 4210
rect 9250 4165 9265 4185
rect 9285 4165 9300 4185
rect 9250 4140 9300 4165
rect 9250 4110 9260 4140
rect 9290 4110 9300 4140
rect 9250 4085 9300 4110
rect 9250 4065 9265 4085
rect 9285 4065 9300 4085
rect 9250 4040 9300 4065
rect 9250 4010 9260 4040
rect 9290 4010 9300 4040
rect 9250 3985 9300 4010
rect 9250 3965 9265 3985
rect 9285 3965 9300 3985
rect 8950 3860 8960 3890
rect 8990 3860 9000 3890
rect 8650 3765 8665 3785
rect 8685 3765 8700 3785
rect 8650 3740 8700 3765
rect 8650 3710 8660 3740
rect 8690 3710 8700 3740
rect 8650 3685 8700 3710
rect 8650 3665 8665 3685
rect 8685 3665 8700 3685
rect 8650 3640 8700 3665
rect 8650 3610 8660 3640
rect 8690 3610 8700 3640
rect 8650 3585 8700 3610
rect 8650 3565 8665 3585
rect 8685 3565 8700 3585
rect 8650 3540 8700 3565
rect 8650 3510 8660 3540
rect 8690 3510 8700 3540
rect 8650 3485 8700 3510
rect 8650 3465 8665 3485
rect 8685 3465 8700 3485
rect 8650 3440 8700 3465
rect 8650 3410 8660 3440
rect 8690 3410 8700 3440
rect 8650 3385 8700 3410
rect 8650 3365 8665 3385
rect 8685 3365 8700 3385
rect 8650 3340 8700 3365
rect 8650 3310 8660 3340
rect 8690 3310 8700 3340
rect 8500 3240 8550 3250
rect 8500 3210 8510 3240
rect 8540 3210 8550 3240
rect 8500 3200 8550 3210
rect 8350 3110 8360 3140
rect 8390 3110 8400 3140
rect 8350 3085 8400 3110
rect 8350 3065 8365 3085
rect 8385 3065 8400 3085
rect 8350 3040 8400 3065
rect 8350 3010 8360 3040
rect 8390 3010 8400 3040
rect 8350 2985 8400 3010
rect 8350 2965 8365 2985
rect 8385 2965 8400 2985
rect 8350 2940 8400 2965
rect 8350 2910 8360 2940
rect 8390 2910 8400 2940
rect 8350 2885 8400 2910
rect 8350 2865 8365 2885
rect 8385 2865 8400 2885
rect 8350 2840 8400 2865
rect 8350 2810 8360 2840
rect 8390 2810 8400 2840
rect 8350 2785 8400 2810
rect 8350 2765 8365 2785
rect 8385 2765 8400 2785
rect 8350 2740 8400 2765
rect 8350 2710 8360 2740
rect 8390 2710 8400 2740
rect 8350 2685 8400 2710
rect 8350 2665 8365 2685
rect 8385 2665 8400 2685
rect 4150 2560 4160 2590
rect 4190 2560 4200 2590
rect 4150 2550 4200 2560
rect 8350 2590 8400 2665
rect 8500 3135 8550 3150
rect 8500 3115 8515 3135
rect 8535 3115 8550 3135
rect 8500 3085 8550 3115
rect 8500 3065 8515 3085
rect 8535 3065 8550 3085
rect 8500 3035 8550 3065
rect 8500 3015 8515 3035
rect 8535 3015 8550 3035
rect 8500 2985 8550 3015
rect 8500 2965 8515 2985
rect 8535 2965 8550 2985
rect 8500 2935 8550 2965
rect 8500 2915 8515 2935
rect 8535 2915 8550 2935
rect 8500 2885 8550 2915
rect 8500 2865 8515 2885
rect 8535 2865 8550 2885
rect 8500 2835 8550 2865
rect 8500 2815 8515 2835
rect 8535 2815 8550 2835
rect 8500 2785 8550 2815
rect 8500 2765 8515 2785
rect 8535 2765 8550 2785
rect 8500 2735 8550 2765
rect 8500 2715 8515 2735
rect 8535 2715 8550 2735
rect 8500 2685 8550 2715
rect 8500 2665 8515 2685
rect 8535 2665 8550 2685
rect 8500 2650 8550 2665
rect 8650 3140 8700 3310
rect 8800 3785 8850 3800
rect 8800 3765 8815 3785
rect 8835 3765 8850 3785
rect 8800 3735 8850 3765
rect 8800 3715 8815 3735
rect 8835 3715 8850 3735
rect 8800 3685 8850 3715
rect 8800 3665 8815 3685
rect 8835 3665 8850 3685
rect 8800 3635 8850 3665
rect 8800 3615 8815 3635
rect 8835 3615 8850 3635
rect 8800 3585 8850 3615
rect 8800 3565 8815 3585
rect 8835 3565 8850 3585
rect 8800 3535 8850 3565
rect 8800 3515 8815 3535
rect 8835 3515 8850 3535
rect 8800 3485 8850 3515
rect 8800 3465 8815 3485
rect 8835 3465 8850 3485
rect 8800 3435 8850 3465
rect 8800 3415 8815 3435
rect 8835 3415 8850 3435
rect 8800 3385 8850 3415
rect 8800 3365 8815 3385
rect 8835 3365 8850 3385
rect 8800 3335 8850 3365
rect 8800 3315 8815 3335
rect 8835 3315 8850 3335
rect 8800 3300 8850 3315
rect 8950 3785 9000 3860
rect 9250 3890 9300 3965
rect 9400 4435 9450 4450
rect 9400 4415 9415 4435
rect 9435 4415 9450 4435
rect 9400 4385 9450 4415
rect 9400 4365 9415 4385
rect 9435 4365 9450 4385
rect 9400 4335 9450 4365
rect 9400 4315 9415 4335
rect 9435 4315 9450 4335
rect 9400 4285 9450 4315
rect 9400 4265 9415 4285
rect 9435 4265 9450 4285
rect 9400 4235 9450 4265
rect 9400 4215 9415 4235
rect 9435 4215 9450 4235
rect 9400 4185 9450 4215
rect 9400 4165 9415 4185
rect 9435 4165 9450 4185
rect 9400 4135 9450 4165
rect 9400 4115 9415 4135
rect 9435 4115 9450 4135
rect 9400 4085 9450 4115
rect 9400 4065 9415 4085
rect 9435 4065 9450 4085
rect 9400 4035 9450 4065
rect 9400 4015 9415 4035
rect 9435 4015 9450 4035
rect 9400 3985 9450 4015
rect 9400 3965 9415 3985
rect 9435 3965 9450 3985
rect 9400 3950 9450 3965
rect 9550 4440 9600 4610
rect 9700 5085 9750 5100
rect 9700 5065 9715 5085
rect 9735 5065 9750 5085
rect 9700 5035 9750 5065
rect 9700 5015 9715 5035
rect 9735 5015 9750 5035
rect 9700 4985 9750 5015
rect 9700 4965 9715 4985
rect 9735 4965 9750 4985
rect 9700 4935 9750 4965
rect 9700 4915 9715 4935
rect 9735 4915 9750 4935
rect 9700 4885 9750 4915
rect 9700 4865 9715 4885
rect 9735 4865 9750 4885
rect 9700 4835 9750 4865
rect 9700 4815 9715 4835
rect 9735 4815 9750 4835
rect 9700 4785 9750 4815
rect 9700 4765 9715 4785
rect 9735 4765 9750 4785
rect 9700 4735 9750 4765
rect 9700 4715 9715 4735
rect 9735 4715 9750 4735
rect 9700 4685 9750 4715
rect 9700 4665 9715 4685
rect 9735 4665 9750 4685
rect 9700 4635 9750 4665
rect 9700 4615 9715 4635
rect 9735 4615 9750 4635
rect 9700 4600 9750 4615
rect 9850 5085 9900 5160
rect 10150 5190 10200 5200
rect 10150 5160 10160 5190
rect 10190 5160 10200 5190
rect 9850 5065 9865 5085
rect 9885 5065 9900 5085
rect 9850 5040 9900 5065
rect 9850 5010 9860 5040
rect 9890 5010 9900 5040
rect 9850 4985 9900 5010
rect 9850 4965 9865 4985
rect 9885 4965 9900 4985
rect 9850 4940 9900 4965
rect 9850 4910 9860 4940
rect 9890 4910 9900 4940
rect 9850 4885 9900 4910
rect 9850 4865 9865 4885
rect 9885 4865 9900 4885
rect 9850 4840 9900 4865
rect 9850 4810 9860 4840
rect 9890 4810 9900 4840
rect 9850 4785 9900 4810
rect 9850 4765 9865 4785
rect 9885 4765 9900 4785
rect 9850 4740 9900 4765
rect 9850 4710 9860 4740
rect 9890 4710 9900 4740
rect 9850 4685 9900 4710
rect 9850 4665 9865 4685
rect 9885 4665 9900 4685
rect 9850 4640 9900 4665
rect 9850 4610 9860 4640
rect 9890 4610 9900 4640
rect 9700 4540 9750 4550
rect 9700 4510 9710 4540
rect 9740 4510 9750 4540
rect 9700 4500 9750 4510
rect 9550 4410 9560 4440
rect 9590 4410 9600 4440
rect 9550 4385 9600 4410
rect 9550 4365 9565 4385
rect 9585 4365 9600 4385
rect 9550 4340 9600 4365
rect 9550 4310 9560 4340
rect 9590 4310 9600 4340
rect 9550 4285 9600 4310
rect 9550 4265 9565 4285
rect 9585 4265 9600 4285
rect 9550 4240 9600 4265
rect 9550 4210 9560 4240
rect 9590 4210 9600 4240
rect 9550 4185 9600 4210
rect 9550 4165 9565 4185
rect 9585 4165 9600 4185
rect 9550 4140 9600 4165
rect 9550 4110 9560 4140
rect 9590 4110 9600 4140
rect 9550 4085 9600 4110
rect 9550 4065 9565 4085
rect 9585 4065 9600 4085
rect 9550 4040 9600 4065
rect 9550 4010 9560 4040
rect 9590 4010 9600 4040
rect 9550 3985 9600 4010
rect 9550 3965 9565 3985
rect 9585 3965 9600 3985
rect 9250 3860 9260 3890
rect 9290 3860 9300 3890
rect 8950 3765 8965 3785
rect 8985 3765 9000 3785
rect 8950 3740 9000 3765
rect 8950 3710 8960 3740
rect 8990 3710 9000 3740
rect 8950 3685 9000 3710
rect 8950 3665 8965 3685
rect 8985 3665 9000 3685
rect 8950 3640 9000 3665
rect 8950 3610 8960 3640
rect 8990 3610 9000 3640
rect 8950 3585 9000 3610
rect 8950 3565 8965 3585
rect 8985 3565 9000 3585
rect 8950 3540 9000 3565
rect 8950 3510 8960 3540
rect 8990 3510 9000 3540
rect 8950 3485 9000 3510
rect 8950 3465 8965 3485
rect 8985 3465 9000 3485
rect 8950 3440 9000 3465
rect 8950 3410 8960 3440
rect 8990 3410 9000 3440
rect 8950 3385 9000 3410
rect 8950 3365 8965 3385
rect 8985 3365 9000 3385
rect 8950 3340 9000 3365
rect 8950 3310 8960 3340
rect 8990 3310 9000 3340
rect 8800 3240 8850 3250
rect 8800 3210 8810 3240
rect 8840 3210 8850 3240
rect 8800 3200 8850 3210
rect 8650 3110 8660 3140
rect 8690 3110 8700 3140
rect 8650 3085 8700 3110
rect 8650 3065 8665 3085
rect 8685 3065 8700 3085
rect 8650 3040 8700 3065
rect 8650 3010 8660 3040
rect 8690 3010 8700 3040
rect 8650 2985 8700 3010
rect 8650 2965 8665 2985
rect 8685 2965 8700 2985
rect 8650 2940 8700 2965
rect 8650 2910 8660 2940
rect 8690 2910 8700 2940
rect 8650 2885 8700 2910
rect 8650 2865 8665 2885
rect 8685 2865 8700 2885
rect 8650 2840 8700 2865
rect 8650 2810 8660 2840
rect 8690 2810 8700 2840
rect 8650 2785 8700 2810
rect 8650 2765 8665 2785
rect 8685 2765 8700 2785
rect 8650 2740 8700 2765
rect 8650 2710 8660 2740
rect 8690 2710 8700 2740
rect 8650 2685 8700 2710
rect 8650 2665 8665 2685
rect 8685 2665 8700 2685
rect 8350 2560 8360 2590
rect 8390 2560 8400 2590
rect 8350 2550 8400 2560
rect 8650 2590 8700 2665
rect 8800 3135 8850 3150
rect 8800 3115 8815 3135
rect 8835 3115 8850 3135
rect 8800 3085 8850 3115
rect 8800 3065 8815 3085
rect 8835 3065 8850 3085
rect 8800 3035 8850 3065
rect 8800 3015 8815 3035
rect 8835 3015 8850 3035
rect 8800 2985 8850 3015
rect 8800 2965 8815 2985
rect 8835 2965 8850 2985
rect 8800 2935 8850 2965
rect 8800 2915 8815 2935
rect 8835 2915 8850 2935
rect 8800 2885 8850 2915
rect 8800 2865 8815 2885
rect 8835 2865 8850 2885
rect 8800 2835 8850 2865
rect 8800 2815 8815 2835
rect 8835 2815 8850 2835
rect 8800 2785 8850 2815
rect 8800 2765 8815 2785
rect 8835 2765 8850 2785
rect 8800 2735 8850 2765
rect 8800 2715 8815 2735
rect 8835 2715 8850 2735
rect 8800 2685 8850 2715
rect 8800 2665 8815 2685
rect 8835 2665 8850 2685
rect 8800 2650 8850 2665
rect 8950 3140 9000 3310
rect 9100 3785 9150 3800
rect 9100 3765 9115 3785
rect 9135 3765 9150 3785
rect 9100 3735 9150 3765
rect 9100 3715 9115 3735
rect 9135 3715 9150 3735
rect 9100 3685 9150 3715
rect 9100 3665 9115 3685
rect 9135 3665 9150 3685
rect 9100 3635 9150 3665
rect 9100 3615 9115 3635
rect 9135 3615 9150 3635
rect 9100 3585 9150 3615
rect 9100 3565 9115 3585
rect 9135 3565 9150 3585
rect 9100 3535 9150 3565
rect 9100 3515 9115 3535
rect 9135 3515 9150 3535
rect 9100 3485 9150 3515
rect 9100 3465 9115 3485
rect 9135 3465 9150 3485
rect 9100 3435 9150 3465
rect 9100 3415 9115 3435
rect 9135 3415 9150 3435
rect 9100 3385 9150 3415
rect 9100 3365 9115 3385
rect 9135 3365 9150 3385
rect 9100 3335 9150 3365
rect 9100 3315 9115 3335
rect 9135 3315 9150 3335
rect 9100 3300 9150 3315
rect 9250 3785 9300 3860
rect 9550 3890 9600 3965
rect 9700 4435 9750 4450
rect 9700 4415 9715 4435
rect 9735 4415 9750 4435
rect 9700 4385 9750 4415
rect 9700 4365 9715 4385
rect 9735 4365 9750 4385
rect 9700 4335 9750 4365
rect 9700 4315 9715 4335
rect 9735 4315 9750 4335
rect 9700 4285 9750 4315
rect 9700 4265 9715 4285
rect 9735 4265 9750 4285
rect 9700 4235 9750 4265
rect 9700 4215 9715 4235
rect 9735 4215 9750 4235
rect 9700 4185 9750 4215
rect 9700 4165 9715 4185
rect 9735 4165 9750 4185
rect 9700 4135 9750 4165
rect 9700 4115 9715 4135
rect 9735 4115 9750 4135
rect 9700 4085 9750 4115
rect 9700 4065 9715 4085
rect 9735 4065 9750 4085
rect 9700 4035 9750 4065
rect 9700 4015 9715 4035
rect 9735 4015 9750 4035
rect 9700 3985 9750 4015
rect 9700 3965 9715 3985
rect 9735 3965 9750 3985
rect 9700 3950 9750 3965
rect 9850 4440 9900 4610
rect 10000 5085 10050 5100
rect 10000 5065 10015 5085
rect 10035 5065 10050 5085
rect 10000 5035 10050 5065
rect 10000 5015 10015 5035
rect 10035 5015 10050 5035
rect 10000 4985 10050 5015
rect 10000 4965 10015 4985
rect 10035 4965 10050 4985
rect 10000 4935 10050 4965
rect 10000 4915 10015 4935
rect 10035 4915 10050 4935
rect 10000 4885 10050 4915
rect 10000 4865 10015 4885
rect 10035 4865 10050 4885
rect 10000 4835 10050 4865
rect 10000 4815 10015 4835
rect 10035 4815 10050 4835
rect 10000 4785 10050 4815
rect 10000 4765 10015 4785
rect 10035 4765 10050 4785
rect 10000 4735 10050 4765
rect 10000 4715 10015 4735
rect 10035 4715 10050 4735
rect 10000 4685 10050 4715
rect 10000 4665 10015 4685
rect 10035 4665 10050 4685
rect 10000 4635 10050 4665
rect 10000 4615 10015 4635
rect 10035 4615 10050 4635
rect 10000 4600 10050 4615
rect 10150 5085 10200 5160
rect 10450 5190 10500 5200
rect 10450 5160 10460 5190
rect 10490 5160 10500 5190
rect 10150 5065 10165 5085
rect 10185 5065 10200 5085
rect 10150 5040 10200 5065
rect 10150 5010 10160 5040
rect 10190 5010 10200 5040
rect 10150 4985 10200 5010
rect 10150 4965 10165 4985
rect 10185 4965 10200 4985
rect 10150 4940 10200 4965
rect 10150 4910 10160 4940
rect 10190 4910 10200 4940
rect 10150 4885 10200 4910
rect 10150 4865 10165 4885
rect 10185 4865 10200 4885
rect 10150 4840 10200 4865
rect 10150 4810 10160 4840
rect 10190 4810 10200 4840
rect 10150 4785 10200 4810
rect 10150 4765 10165 4785
rect 10185 4765 10200 4785
rect 10150 4740 10200 4765
rect 10150 4710 10160 4740
rect 10190 4710 10200 4740
rect 10150 4685 10200 4710
rect 10150 4665 10165 4685
rect 10185 4665 10200 4685
rect 10150 4640 10200 4665
rect 10150 4610 10160 4640
rect 10190 4610 10200 4640
rect 10000 4540 10050 4550
rect 10000 4510 10010 4540
rect 10040 4510 10050 4540
rect 10000 4500 10050 4510
rect 9850 4410 9860 4440
rect 9890 4410 9900 4440
rect 9850 4385 9900 4410
rect 9850 4365 9865 4385
rect 9885 4365 9900 4385
rect 9850 4340 9900 4365
rect 9850 4310 9860 4340
rect 9890 4310 9900 4340
rect 9850 4285 9900 4310
rect 9850 4265 9865 4285
rect 9885 4265 9900 4285
rect 9850 4240 9900 4265
rect 9850 4210 9860 4240
rect 9890 4210 9900 4240
rect 9850 4185 9900 4210
rect 9850 4165 9865 4185
rect 9885 4165 9900 4185
rect 9850 4140 9900 4165
rect 9850 4110 9860 4140
rect 9890 4110 9900 4140
rect 9850 4085 9900 4110
rect 9850 4065 9865 4085
rect 9885 4065 9900 4085
rect 9850 4040 9900 4065
rect 9850 4010 9860 4040
rect 9890 4010 9900 4040
rect 9850 3985 9900 4010
rect 9850 3965 9865 3985
rect 9885 3965 9900 3985
rect 9550 3860 9560 3890
rect 9590 3860 9600 3890
rect 9250 3765 9265 3785
rect 9285 3765 9300 3785
rect 9250 3740 9300 3765
rect 9250 3710 9260 3740
rect 9290 3710 9300 3740
rect 9250 3685 9300 3710
rect 9250 3665 9265 3685
rect 9285 3665 9300 3685
rect 9250 3640 9300 3665
rect 9250 3610 9260 3640
rect 9290 3610 9300 3640
rect 9250 3585 9300 3610
rect 9250 3565 9265 3585
rect 9285 3565 9300 3585
rect 9250 3540 9300 3565
rect 9250 3510 9260 3540
rect 9290 3510 9300 3540
rect 9250 3485 9300 3510
rect 9250 3465 9265 3485
rect 9285 3465 9300 3485
rect 9250 3440 9300 3465
rect 9250 3410 9260 3440
rect 9290 3410 9300 3440
rect 9250 3385 9300 3410
rect 9250 3365 9265 3385
rect 9285 3365 9300 3385
rect 9250 3340 9300 3365
rect 9250 3310 9260 3340
rect 9290 3310 9300 3340
rect 9100 3240 9150 3250
rect 9100 3210 9110 3240
rect 9140 3210 9150 3240
rect 9100 3200 9150 3210
rect 8950 3110 8960 3140
rect 8990 3110 9000 3140
rect 8950 3085 9000 3110
rect 8950 3065 8965 3085
rect 8985 3065 9000 3085
rect 8950 3040 9000 3065
rect 8950 3010 8960 3040
rect 8990 3010 9000 3040
rect 8950 2985 9000 3010
rect 8950 2965 8965 2985
rect 8985 2965 9000 2985
rect 8950 2940 9000 2965
rect 8950 2910 8960 2940
rect 8990 2910 9000 2940
rect 8950 2885 9000 2910
rect 8950 2865 8965 2885
rect 8985 2865 9000 2885
rect 8950 2840 9000 2865
rect 8950 2810 8960 2840
rect 8990 2810 9000 2840
rect 8950 2785 9000 2810
rect 8950 2765 8965 2785
rect 8985 2765 9000 2785
rect 8950 2740 9000 2765
rect 8950 2710 8960 2740
rect 8990 2710 9000 2740
rect 8950 2685 9000 2710
rect 8950 2665 8965 2685
rect 8985 2665 9000 2685
rect 8650 2560 8660 2590
rect 8690 2560 8700 2590
rect 8650 2550 8700 2560
rect 8950 2590 9000 2665
rect 9100 3135 9150 3150
rect 9100 3115 9115 3135
rect 9135 3115 9150 3135
rect 9100 3085 9150 3115
rect 9100 3065 9115 3085
rect 9135 3065 9150 3085
rect 9100 3035 9150 3065
rect 9100 3015 9115 3035
rect 9135 3015 9150 3035
rect 9100 2985 9150 3015
rect 9100 2965 9115 2985
rect 9135 2965 9150 2985
rect 9100 2935 9150 2965
rect 9100 2915 9115 2935
rect 9135 2915 9150 2935
rect 9100 2885 9150 2915
rect 9100 2865 9115 2885
rect 9135 2865 9150 2885
rect 9100 2835 9150 2865
rect 9100 2815 9115 2835
rect 9135 2815 9150 2835
rect 9100 2785 9150 2815
rect 9100 2765 9115 2785
rect 9135 2765 9150 2785
rect 9100 2735 9150 2765
rect 9100 2715 9115 2735
rect 9135 2715 9150 2735
rect 9100 2685 9150 2715
rect 9100 2665 9115 2685
rect 9135 2665 9150 2685
rect 9100 2650 9150 2665
rect 9250 3140 9300 3310
rect 9400 3785 9450 3800
rect 9400 3765 9415 3785
rect 9435 3765 9450 3785
rect 9400 3735 9450 3765
rect 9400 3715 9415 3735
rect 9435 3715 9450 3735
rect 9400 3685 9450 3715
rect 9400 3665 9415 3685
rect 9435 3665 9450 3685
rect 9400 3635 9450 3665
rect 9400 3615 9415 3635
rect 9435 3615 9450 3635
rect 9400 3585 9450 3615
rect 9400 3565 9415 3585
rect 9435 3565 9450 3585
rect 9400 3535 9450 3565
rect 9400 3515 9415 3535
rect 9435 3515 9450 3535
rect 9400 3485 9450 3515
rect 9400 3465 9415 3485
rect 9435 3465 9450 3485
rect 9400 3435 9450 3465
rect 9400 3415 9415 3435
rect 9435 3415 9450 3435
rect 9400 3385 9450 3415
rect 9400 3365 9415 3385
rect 9435 3365 9450 3385
rect 9400 3335 9450 3365
rect 9400 3315 9415 3335
rect 9435 3315 9450 3335
rect 9400 3300 9450 3315
rect 9550 3785 9600 3860
rect 9850 3890 9900 3965
rect 10000 4435 10050 4450
rect 10000 4415 10015 4435
rect 10035 4415 10050 4435
rect 10000 4385 10050 4415
rect 10000 4365 10015 4385
rect 10035 4365 10050 4385
rect 10000 4335 10050 4365
rect 10000 4315 10015 4335
rect 10035 4315 10050 4335
rect 10000 4285 10050 4315
rect 10000 4265 10015 4285
rect 10035 4265 10050 4285
rect 10000 4235 10050 4265
rect 10000 4215 10015 4235
rect 10035 4215 10050 4235
rect 10000 4185 10050 4215
rect 10000 4165 10015 4185
rect 10035 4165 10050 4185
rect 10000 4135 10050 4165
rect 10000 4115 10015 4135
rect 10035 4115 10050 4135
rect 10000 4085 10050 4115
rect 10000 4065 10015 4085
rect 10035 4065 10050 4085
rect 10000 4035 10050 4065
rect 10000 4015 10015 4035
rect 10035 4015 10050 4035
rect 10000 3985 10050 4015
rect 10000 3965 10015 3985
rect 10035 3965 10050 3985
rect 10000 3950 10050 3965
rect 10150 4440 10200 4610
rect 10300 5085 10350 5100
rect 10300 5065 10315 5085
rect 10335 5065 10350 5085
rect 10300 5035 10350 5065
rect 10300 5015 10315 5035
rect 10335 5015 10350 5035
rect 10300 4985 10350 5015
rect 10300 4965 10315 4985
rect 10335 4965 10350 4985
rect 10300 4935 10350 4965
rect 10300 4915 10315 4935
rect 10335 4915 10350 4935
rect 10300 4885 10350 4915
rect 10300 4865 10315 4885
rect 10335 4865 10350 4885
rect 10300 4835 10350 4865
rect 10300 4815 10315 4835
rect 10335 4815 10350 4835
rect 10300 4785 10350 4815
rect 10300 4765 10315 4785
rect 10335 4765 10350 4785
rect 10300 4735 10350 4765
rect 10300 4715 10315 4735
rect 10335 4715 10350 4735
rect 10300 4685 10350 4715
rect 10300 4665 10315 4685
rect 10335 4665 10350 4685
rect 10300 4635 10350 4665
rect 10300 4615 10315 4635
rect 10335 4615 10350 4635
rect 10300 4600 10350 4615
rect 10450 5085 10500 5160
rect 10750 5190 10800 5200
rect 10750 5160 10760 5190
rect 10790 5160 10800 5190
rect 10450 5065 10465 5085
rect 10485 5065 10500 5085
rect 10450 5040 10500 5065
rect 10450 5010 10460 5040
rect 10490 5010 10500 5040
rect 10450 4985 10500 5010
rect 10450 4965 10465 4985
rect 10485 4965 10500 4985
rect 10450 4940 10500 4965
rect 10450 4910 10460 4940
rect 10490 4910 10500 4940
rect 10450 4885 10500 4910
rect 10450 4865 10465 4885
rect 10485 4865 10500 4885
rect 10450 4840 10500 4865
rect 10450 4810 10460 4840
rect 10490 4810 10500 4840
rect 10450 4785 10500 4810
rect 10450 4765 10465 4785
rect 10485 4765 10500 4785
rect 10450 4740 10500 4765
rect 10450 4710 10460 4740
rect 10490 4710 10500 4740
rect 10450 4685 10500 4710
rect 10450 4665 10465 4685
rect 10485 4665 10500 4685
rect 10450 4640 10500 4665
rect 10450 4610 10460 4640
rect 10490 4610 10500 4640
rect 10300 4540 10350 4550
rect 10300 4510 10310 4540
rect 10340 4510 10350 4540
rect 10300 4500 10350 4510
rect 10150 4410 10160 4440
rect 10190 4410 10200 4440
rect 10150 4385 10200 4410
rect 10150 4365 10165 4385
rect 10185 4365 10200 4385
rect 10150 4340 10200 4365
rect 10150 4310 10160 4340
rect 10190 4310 10200 4340
rect 10150 4285 10200 4310
rect 10150 4265 10165 4285
rect 10185 4265 10200 4285
rect 10150 4240 10200 4265
rect 10150 4210 10160 4240
rect 10190 4210 10200 4240
rect 10150 4185 10200 4210
rect 10150 4165 10165 4185
rect 10185 4165 10200 4185
rect 10150 4140 10200 4165
rect 10150 4110 10160 4140
rect 10190 4110 10200 4140
rect 10150 4085 10200 4110
rect 10150 4065 10165 4085
rect 10185 4065 10200 4085
rect 10150 4040 10200 4065
rect 10150 4010 10160 4040
rect 10190 4010 10200 4040
rect 10150 3985 10200 4010
rect 10150 3965 10165 3985
rect 10185 3965 10200 3985
rect 9850 3860 9860 3890
rect 9890 3860 9900 3890
rect 9550 3765 9565 3785
rect 9585 3765 9600 3785
rect 9550 3740 9600 3765
rect 9550 3710 9560 3740
rect 9590 3710 9600 3740
rect 9550 3685 9600 3710
rect 9550 3665 9565 3685
rect 9585 3665 9600 3685
rect 9550 3640 9600 3665
rect 9550 3610 9560 3640
rect 9590 3610 9600 3640
rect 9550 3585 9600 3610
rect 9550 3565 9565 3585
rect 9585 3565 9600 3585
rect 9550 3540 9600 3565
rect 9550 3510 9560 3540
rect 9590 3510 9600 3540
rect 9550 3485 9600 3510
rect 9550 3465 9565 3485
rect 9585 3465 9600 3485
rect 9550 3440 9600 3465
rect 9550 3410 9560 3440
rect 9590 3410 9600 3440
rect 9550 3385 9600 3410
rect 9550 3365 9565 3385
rect 9585 3365 9600 3385
rect 9550 3340 9600 3365
rect 9550 3310 9560 3340
rect 9590 3310 9600 3340
rect 9400 3240 9450 3250
rect 9400 3210 9410 3240
rect 9440 3210 9450 3240
rect 9400 3200 9450 3210
rect 9250 3110 9260 3140
rect 9290 3110 9300 3140
rect 9250 3085 9300 3110
rect 9250 3065 9265 3085
rect 9285 3065 9300 3085
rect 9250 3040 9300 3065
rect 9250 3010 9260 3040
rect 9290 3010 9300 3040
rect 9250 2985 9300 3010
rect 9250 2965 9265 2985
rect 9285 2965 9300 2985
rect 9250 2940 9300 2965
rect 9250 2910 9260 2940
rect 9290 2910 9300 2940
rect 9250 2885 9300 2910
rect 9250 2865 9265 2885
rect 9285 2865 9300 2885
rect 9250 2840 9300 2865
rect 9250 2810 9260 2840
rect 9290 2810 9300 2840
rect 9250 2785 9300 2810
rect 9250 2765 9265 2785
rect 9285 2765 9300 2785
rect 9250 2740 9300 2765
rect 9250 2710 9260 2740
rect 9290 2710 9300 2740
rect 9250 2685 9300 2710
rect 9250 2665 9265 2685
rect 9285 2665 9300 2685
rect 8950 2560 8960 2590
rect 8990 2560 9000 2590
rect 8950 2550 9000 2560
rect 9250 2590 9300 2665
rect 9400 3135 9450 3150
rect 9400 3115 9415 3135
rect 9435 3115 9450 3135
rect 9400 3085 9450 3115
rect 9400 3065 9415 3085
rect 9435 3065 9450 3085
rect 9400 3035 9450 3065
rect 9400 3015 9415 3035
rect 9435 3015 9450 3035
rect 9400 2985 9450 3015
rect 9400 2965 9415 2985
rect 9435 2965 9450 2985
rect 9400 2935 9450 2965
rect 9400 2915 9415 2935
rect 9435 2915 9450 2935
rect 9400 2885 9450 2915
rect 9400 2865 9415 2885
rect 9435 2865 9450 2885
rect 9400 2835 9450 2865
rect 9400 2815 9415 2835
rect 9435 2815 9450 2835
rect 9400 2785 9450 2815
rect 9400 2765 9415 2785
rect 9435 2765 9450 2785
rect 9400 2735 9450 2765
rect 9400 2715 9415 2735
rect 9435 2715 9450 2735
rect 9400 2685 9450 2715
rect 9400 2665 9415 2685
rect 9435 2665 9450 2685
rect 9400 2650 9450 2665
rect 9550 3140 9600 3310
rect 9700 3785 9750 3800
rect 9700 3765 9715 3785
rect 9735 3765 9750 3785
rect 9700 3735 9750 3765
rect 9700 3715 9715 3735
rect 9735 3715 9750 3735
rect 9700 3685 9750 3715
rect 9700 3665 9715 3685
rect 9735 3665 9750 3685
rect 9700 3635 9750 3665
rect 9700 3615 9715 3635
rect 9735 3615 9750 3635
rect 9700 3585 9750 3615
rect 9700 3565 9715 3585
rect 9735 3565 9750 3585
rect 9700 3535 9750 3565
rect 9700 3515 9715 3535
rect 9735 3515 9750 3535
rect 9700 3485 9750 3515
rect 9700 3465 9715 3485
rect 9735 3465 9750 3485
rect 9700 3435 9750 3465
rect 9700 3415 9715 3435
rect 9735 3415 9750 3435
rect 9700 3385 9750 3415
rect 9700 3365 9715 3385
rect 9735 3365 9750 3385
rect 9700 3335 9750 3365
rect 9700 3315 9715 3335
rect 9735 3315 9750 3335
rect 9700 3300 9750 3315
rect 9850 3785 9900 3860
rect 10150 3890 10200 3965
rect 10300 4435 10350 4450
rect 10300 4415 10315 4435
rect 10335 4415 10350 4435
rect 10300 4385 10350 4415
rect 10300 4365 10315 4385
rect 10335 4365 10350 4385
rect 10300 4335 10350 4365
rect 10300 4315 10315 4335
rect 10335 4315 10350 4335
rect 10300 4285 10350 4315
rect 10300 4265 10315 4285
rect 10335 4265 10350 4285
rect 10300 4235 10350 4265
rect 10300 4215 10315 4235
rect 10335 4215 10350 4235
rect 10300 4185 10350 4215
rect 10300 4165 10315 4185
rect 10335 4165 10350 4185
rect 10300 4135 10350 4165
rect 10300 4115 10315 4135
rect 10335 4115 10350 4135
rect 10300 4085 10350 4115
rect 10300 4065 10315 4085
rect 10335 4065 10350 4085
rect 10300 4035 10350 4065
rect 10300 4015 10315 4035
rect 10335 4015 10350 4035
rect 10300 3985 10350 4015
rect 10300 3965 10315 3985
rect 10335 3965 10350 3985
rect 10300 3950 10350 3965
rect 10450 4440 10500 4610
rect 10600 5085 10650 5100
rect 10600 5065 10615 5085
rect 10635 5065 10650 5085
rect 10600 5035 10650 5065
rect 10600 5015 10615 5035
rect 10635 5015 10650 5035
rect 10600 4985 10650 5015
rect 10600 4965 10615 4985
rect 10635 4965 10650 4985
rect 10600 4935 10650 4965
rect 10600 4915 10615 4935
rect 10635 4915 10650 4935
rect 10600 4885 10650 4915
rect 10600 4865 10615 4885
rect 10635 4865 10650 4885
rect 10600 4835 10650 4865
rect 10600 4815 10615 4835
rect 10635 4815 10650 4835
rect 10600 4785 10650 4815
rect 10600 4765 10615 4785
rect 10635 4765 10650 4785
rect 10600 4735 10650 4765
rect 10600 4715 10615 4735
rect 10635 4715 10650 4735
rect 10600 4685 10650 4715
rect 10600 4665 10615 4685
rect 10635 4665 10650 4685
rect 10600 4635 10650 4665
rect 10600 4615 10615 4635
rect 10635 4615 10650 4635
rect 10600 4600 10650 4615
rect 10750 5085 10800 5160
rect 11950 5190 12000 5200
rect 11950 5160 11960 5190
rect 11990 5160 12000 5190
rect 10750 5065 10765 5085
rect 10785 5065 10800 5085
rect 10750 5040 10800 5065
rect 10750 5010 10760 5040
rect 10790 5010 10800 5040
rect 10750 4985 10800 5010
rect 10750 4965 10765 4985
rect 10785 4965 10800 4985
rect 10750 4940 10800 4965
rect 10750 4910 10760 4940
rect 10790 4910 10800 4940
rect 10750 4885 10800 4910
rect 10750 4865 10765 4885
rect 10785 4865 10800 4885
rect 10750 4840 10800 4865
rect 10750 4810 10760 4840
rect 10790 4810 10800 4840
rect 10750 4785 10800 4810
rect 10750 4765 10765 4785
rect 10785 4765 10800 4785
rect 10750 4740 10800 4765
rect 10750 4710 10760 4740
rect 10790 4710 10800 4740
rect 10750 4685 10800 4710
rect 10750 4665 10765 4685
rect 10785 4665 10800 4685
rect 10750 4640 10800 4665
rect 10750 4610 10760 4640
rect 10790 4610 10800 4640
rect 10600 4540 10650 4550
rect 10600 4510 10610 4540
rect 10640 4510 10650 4540
rect 10600 4500 10650 4510
rect 10450 4410 10460 4440
rect 10490 4410 10500 4440
rect 10450 4385 10500 4410
rect 10450 4365 10465 4385
rect 10485 4365 10500 4385
rect 10450 4340 10500 4365
rect 10450 4310 10460 4340
rect 10490 4310 10500 4340
rect 10450 4285 10500 4310
rect 10450 4265 10465 4285
rect 10485 4265 10500 4285
rect 10450 4240 10500 4265
rect 10450 4210 10460 4240
rect 10490 4210 10500 4240
rect 10450 4185 10500 4210
rect 10450 4165 10465 4185
rect 10485 4165 10500 4185
rect 10450 4140 10500 4165
rect 10450 4110 10460 4140
rect 10490 4110 10500 4140
rect 10450 4085 10500 4110
rect 10450 4065 10465 4085
rect 10485 4065 10500 4085
rect 10450 4040 10500 4065
rect 10450 4010 10460 4040
rect 10490 4010 10500 4040
rect 10450 3985 10500 4010
rect 10450 3965 10465 3985
rect 10485 3965 10500 3985
rect 10150 3860 10160 3890
rect 10190 3860 10200 3890
rect 9850 3765 9865 3785
rect 9885 3765 9900 3785
rect 9850 3740 9900 3765
rect 9850 3710 9860 3740
rect 9890 3710 9900 3740
rect 9850 3685 9900 3710
rect 9850 3665 9865 3685
rect 9885 3665 9900 3685
rect 9850 3640 9900 3665
rect 9850 3610 9860 3640
rect 9890 3610 9900 3640
rect 9850 3585 9900 3610
rect 9850 3565 9865 3585
rect 9885 3565 9900 3585
rect 9850 3540 9900 3565
rect 9850 3510 9860 3540
rect 9890 3510 9900 3540
rect 9850 3485 9900 3510
rect 9850 3465 9865 3485
rect 9885 3465 9900 3485
rect 9850 3440 9900 3465
rect 9850 3410 9860 3440
rect 9890 3410 9900 3440
rect 9850 3385 9900 3410
rect 9850 3365 9865 3385
rect 9885 3365 9900 3385
rect 9850 3340 9900 3365
rect 9850 3310 9860 3340
rect 9890 3310 9900 3340
rect 9700 3240 9750 3250
rect 9700 3210 9710 3240
rect 9740 3210 9750 3240
rect 9700 3200 9750 3210
rect 9550 3110 9560 3140
rect 9590 3110 9600 3140
rect 9550 3085 9600 3110
rect 9550 3065 9565 3085
rect 9585 3065 9600 3085
rect 9550 3040 9600 3065
rect 9550 3010 9560 3040
rect 9590 3010 9600 3040
rect 9550 2985 9600 3010
rect 9550 2965 9565 2985
rect 9585 2965 9600 2985
rect 9550 2940 9600 2965
rect 9550 2910 9560 2940
rect 9590 2910 9600 2940
rect 9550 2885 9600 2910
rect 9550 2865 9565 2885
rect 9585 2865 9600 2885
rect 9550 2840 9600 2865
rect 9550 2810 9560 2840
rect 9590 2810 9600 2840
rect 9550 2785 9600 2810
rect 9550 2765 9565 2785
rect 9585 2765 9600 2785
rect 9550 2740 9600 2765
rect 9550 2710 9560 2740
rect 9590 2710 9600 2740
rect 9550 2685 9600 2710
rect 9550 2665 9565 2685
rect 9585 2665 9600 2685
rect 9250 2560 9260 2590
rect 9290 2560 9300 2590
rect 9250 2550 9300 2560
rect 9550 2590 9600 2665
rect 9700 3135 9750 3150
rect 9700 3115 9715 3135
rect 9735 3115 9750 3135
rect 9700 3085 9750 3115
rect 9700 3065 9715 3085
rect 9735 3065 9750 3085
rect 9700 3035 9750 3065
rect 9700 3015 9715 3035
rect 9735 3015 9750 3035
rect 9700 2985 9750 3015
rect 9700 2965 9715 2985
rect 9735 2965 9750 2985
rect 9700 2935 9750 2965
rect 9700 2915 9715 2935
rect 9735 2915 9750 2935
rect 9700 2885 9750 2915
rect 9700 2865 9715 2885
rect 9735 2865 9750 2885
rect 9700 2835 9750 2865
rect 9700 2815 9715 2835
rect 9735 2815 9750 2835
rect 9700 2785 9750 2815
rect 9700 2765 9715 2785
rect 9735 2765 9750 2785
rect 9700 2735 9750 2765
rect 9700 2715 9715 2735
rect 9735 2715 9750 2735
rect 9700 2685 9750 2715
rect 9700 2665 9715 2685
rect 9735 2665 9750 2685
rect 9700 2650 9750 2665
rect 9850 3140 9900 3310
rect 10000 3785 10050 3800
rect 10000 3765 10015 3785
rect 10035 3765 10050 3785
rect 10000 3735 10050 3765
rect 10000 3715 10015 3735
rect 10035 3715 10050 3735
rect 10000 3685 10050 3715
rect 10000 3665 10015 3685
rect 10035 3665 10050 3685
rect 10000 3635 10050 3665
rect 10000 3615 10015 3635
rect 10035 3615 10050 3635
rect 10000 3585 10050 3615
rect 10000 3565 10015 3585
rect 10035 3565 10050 3585
rect 10000 3535 10050 3565
rect 10000 3515 10015 3535
rect 10035 3515 10050 3535
rect 10000 3485 10050 3515
rect 10000 3465 10015 3485
rect 10035 3465 10050 3485
rect 10000 3435 10050 3465
rect 10000 3415 10015 3435
rect 10035 3415 10050 3435
rect 10000 3385 10050 3415
rect 10000 3365 10015 3385
rect 10035 3365 10050 3385
rect 10000 3335 10050 3365
rect 10000 3315 10015 3335
rect 10035 3315 10050 3335
rect 10000 3300 10050 3315
rect 10150 3785 10200 3860
rect 10450 3890 10500 3965
rect 10600 4435 10650 4450
rect 10600 4415 10615 4435
rect 10635 4415 10650 4435
rect 10600 4385 10650 4415
rect 10600 4365 10615 4385
rect 10635 4365 10650 4385
rect 10600 4335 10650 4365
rect 10600 4315 10615 4335
rect 10635 4315 10650 4335
rect 10600 4285 10650 4315
rect 10600 4265 10615 4285
rect 10635 4265 10650 4285
rect 10600 4235 10650 4265
rect 10600 4215 10615 4235
rect 10635 4215 10650 4235
rect 10600 4185 10650 4215
rect 10600 4165 10615 4185
rect 10635 4165 10650 4185
rect 10600 4135 10650 4165
rect 10600 4115 10615 4135
rect 10635 4115 10650 4135
rect 10600 4085 10650 4115
rect 10600 4065 10615 4085
rect 10635 4065 10650 4085
rect 10600 4035 10650 4065
rect 10600 4015 10615 4035
rect 10635 4015 10650 4035
rect 10600 3985 10650 4015
rect 10600 3965 10615 3985
rect 10635 3965 10650 3985
rect 10600 3950 10650 3965
rect 10750 4440 10800 4610
rect 11350 5085 11400 5100
rect 11350 5065 11365 5085
rect 11385 5065 11400 5085
rect 11350 5035 11400 5065
rect 11350 5015 11365 5035
rect 11385 5015 11400 5035
rect 11350 4985 11400 5015
rect 11350 4965 11365 4985
rect 11385 4965 11400 4985
rect 11350 4935 11400 4965
rect 11350 4915 11365 4935
rect 11385 4915 11400 4935
rect 11350 4885 11400 4915
rect 11350 4865 11365 4885
rect 11385 4865 11400 4885
rect 11350 4835 11400 4865
rect 11350 4815 11365 4835
rect 11385 4815 11400 4835
rect 11350 4785 11400 4815
rect 11350 4765 11365 4785
rect 11385 4765 11400 4785
rect 11350 4735 11400 4765
rect 11350 4715 11365 4735
rect 11385 4715 11400 4735
rect 11350 4685 11400 4715
rect 11350 4665 11365 4685
rect 11385 4665 11400 4685
rect 11350 4635 11400 4665
rect 11350 4615 11365 4635
rect 11385 4615 11400 4635
rect 10900 4540 10950 4550
rect 10900 4510 10910 4540
rect 10940 4510 10950 4540
rect 10900 4500 10950 4510
rect 11200 4540 11250 4550
rect 11200 4510 11210 4540
rect 11240 4510 11250 4540
rect 11200 4500 11250 4510
rect 11350 4540 11400 4615
rect 11950 5085 12000 5160
rect 13150 5190 13200 5200
rect 13150 5160 13160 5190
rect 13190 5160 13200 5190
rect 11950 5065 11965 5085
rect 11985 5065 12000 5085
rect 11950 5040 12000 5065
rect 11950 5010 11960 5040
rect 11990 5010 12000 5040
rect 11950 4985 12000 5010
rect 11950 4965 11965 4985
rect 11985 4965 12000 4985
rect 11950 4940 12000 4965
rect 11950 4910 11960 4940
rect 11990 4910 12000 4940
rect 11950 4885 12000 4910
rect 11950 4865 11965 4885
rect 11985 4865 12000 4885
rect 11950 4840 12000 4865
rect 11950 4810 11960 4840
rect 11990 4810 12000 4840
rect 11950 4785 12000 4810
rect 11950 4765 11965 4785
rect 11985 4765 12000 4785
rect 11950 4740 12000 4765
rect 11950 4710 11960 4740
rect 11990 4710 12000 4740
rect 11950 4685 12000 4710
rect 11950 4665 11965 4685
rect 11985 4665 12000 4685
rect 11950 4640 12000 4665
rect 11950 4610 11960 4640
rect 11990 4610 12000 4640
rect 11350 4510 11360 4540
rect 11390 4510 11400 4540
rect 10750 4410 10760 4440
rect 10790 4410 10800 4440
rect 10750 4385 10800 4410
rect 10750 4365 10765 4385
rect 10785 4365 10800 4385
rect 10750 4340 10800 4365
rect 10750 4310 10760 4340
rect 10790 4310 10800 4340
rect 10750 4285 10800 4310
rect 10750 4265 10765 4285
rect 10785 4265 10800 4285
rect 10750 4240 10800 4265
rect 10750 4210 10760 4240
rect 10790 4210 10800 4240
rect 10750 4185 10800 4210
rect 10750 4165 10765 4185
rect 10785 4165 10800 4185
rect 10750 4140 10800 4165
rect 10750 4110 10760 4140
rect 10790 4110 10800 4140
rect 10750 4085 10800 4110
rect 10750 4065 10765 4085
rect 10785 4065 10800 4085
rect 10750 4040 10800 4065
rect 10750 4010 10760 4040
rect 10790 4010 10800 4040
rect 10750 3985 10800 4010
rect 10750 3965 10765 3985
rect 10785 3965 10800 3985
rect 10450 3860 10460 3890
rect 10490 3860 10500 3890
rect 10150 3765 10165 3785
rect 10185 3765 10200 3785
rect 10150 3740 10200 3765
rect 10150 3710 10160 3740
rect 10190 3710 10200 3740
rect 10150 3685 10200 3710
rect 10150 3665 10165 3685
rect 10185 3665 10200 3685
rect 10150 3640 10200 3665
rect 10150 3610 10160 3640
rect 10190 3610 10200 3640
rect 10150 3585 10200 3610
rect 10150 3565 10165 3585
rect 10185 3565 10200 3585
rect 10150 3540 10200 3565
rect 10150 3510 10160 3540
rect 10190 3510 10200 3540
rect 10150 3485 10200 3510
rect 10150 3465 10165 3485
rect 10185 3465 10200 3485
rect 10150 3440 10200 3465
rect 10150 3410 10160 3440
rect 10190 3410 10200 3440
rect 10150 3385 10200 3410
rect 10150 3365 10165 3385
rect 10185 3365 10200 3385
rect 10150 3340 10200 3365
rect 10150 3310 10160 3340
rect 10190 3310 10200 3340
rect 10000 3240 10050 3250
rect 10000 3210 10010 3240
rect 10040 3210 10050 3240
rect 10000 3200 10050 3210
rect 9850 3110 9860 3140
rect 9890 3110 9900 3140
rect 9850 3085 9900 3110
rect 9850 3065 9865 3085
rect 9885 3065 9900 3085
rect 9850 3040 9900 3065
rect 9850 3010 9860 3040
rect 9890 3010 9900 3040
rect 9850 2985 9900 3010
rect 9850 2965 9865 2985
rect 9885 2965 9900 2985
rect 9850 2940 9900 2965
rect 9850 2910 9860 2940
rect 9890 2910 9900 2940
rect 9850 2885 9900 2910
rect 9850 2865 9865 2885
rect 9885 2865 9900 2885
rect 9850 2840 9900 2865
rect 9850 2810 9860 2840
rect 9890 2810 9900 2840
rect 9850 2785 9900 2810
rect 9850 2765 9865 2785
rect 9885 2765 9900 2785
rect 9850 2740 9900 2765
rect 9850 2710 9860 2740
rect 9890 2710 9900 2740
rect 9850 2685 9900 2710
rect 9850 2665 9865 2685
rect 9885 2665 9900 2685
rect 9550 2560 9560 2590
rect 9590 2560 9600 2590
rect 9550 2550 9600 2560
rect 9850 2590 9900 2665
rect 10000 3135 10050 3150
rect 10000 3115 10015 3135
rect 10035 3115 10050 3135
rect 10000 3085 10050 3115
rect 10000 3065 10015 3085
rect 10035 3065 10050 3085
rect 10000 3035 10050 3065
rect 10000 3015 10015 3035
rect 10035 3015 10050 3035
rect 10000 2985 10050 3015
rect 10000 2965 10015 2985
rect 10035 2965 10050 2985
rect 10000 2935 10050 2965
rect 10000 2915 10015 2935
rect 10035 2915 10050 2935
rect 10000 2885 10050 2915
rect 10000 2865 10015 2885
rect 10035 2865 10050 2885
rect 10000 2835 10050 2865
rect 10000 2815 10015 2835
rect 10035 2815 10050 2835
rect 10000 2785 10050 2815
rect 10000 2765 10015 2785
rect 10035 2765 10050 2785
rect 10000 2735 10050 2765
rect 10000 2715 10015 2735
rect 10035 2715 10050 2735
rect 10000 2685 10050 2715
rect 10000 2665 10015 2685
rect 10035 2665 10050 2685
rect 10000 2650 10050 2665
rect 10150 3140 10200 3310
rect 10300 3785 10350 3800
rect 10300 3765 10315 3785
rect 10335 3765 10350 3785
rect 10300 3735 10350 3765
rect 10300 3715 10315 3735
rect 10335 3715 10350 3735
rect 10300 3685 10350 3715
rect 10300 3665 10315 3685
rect 10335 3665 10350 3685
rect 10300 3635 10350 3665
rect 10300 3615 10315 3635
rect 10335 3615 10350 3635
rect 10300 3585 10350 3615
rect 10300 3565 10315 3585
rect 10335 3565 10350 3585
rect 10300 3535 10350 3565
rect 10300 3515 10315 3535
rect 10335 3515 10350 3535
rect 10300 3485 10350 3515
rect 10300 3465 10315 3485
rect 10335 3465 10350 3485
rect 10300 3435 10350 3465
rect 10300 3415 10315 3435
rect 10335 3415 10350 3435
rect 10300 3385 10350 3415
rect 10300 3365 10315 3385
rect 10335 3365 10350 3385
rect 10300 3335 10350 3365
rect 10300 3315 10315 3335
rect 10335 3315 10350 3335
rect 10300 3300 10350 3315
rect 10450 3785 10500 3860
rect 10750 3890 10800 3965
rect 10750 3860 10760 3890
rect 10790 3860 10800 3890
rect 10450 3765 10465 3785
rect 10485 3765 10500 3785
rect 10450 3740 10500 3765
rect 10450 3710 10460 3740
rect 10490 3710 10500 3740
rect 10450 3685 10500 3710
rect 10450 3665 10465 3685
rect 10485 3665 10500 3685
rect 10450 3640 10500 3665
rect 10450 3610 10460 3640
rect 10490 3610 10500 3640
rect 10450 3585 10500 3610
rect 10450 3565 10465 3585
rect 10485 3565 10500 3585
rect 10450 3540 10500 3565
rect 10450 3510 10460 3540
rect 10490 3510 10500 3540
rect 10450 3485 10500 3510
rect 10450 3465 10465 3485
rect 10485 3465 10500 3485
rect 10450 3440 10500 3465
rect 10450 3410 10460 3440
rect 10490 3410 10500 3440
rect 10450 3385 10500 3410
rect 10450 3365 10465 3385
rect 10485 3365 10500 3385
rect 10450 3340 10500 3365
rect 10450 3310 10460 3340
rect 10490 3310 10500 3340
rect 10300 3240 10350 3250
rect 10300 3210 10310 3240
rect 10340 3210 10350 3240
rect 10300 3200 10350 3210
rect 10150 3110 10160 3140
rect 10190 3110 10200 3140
rect 10150 3085 10200 3110
rect 10150 3065 10165 3085
rect 10185 3065 10200 3085
rect 10150 3040 10200 3065
rect 10150 3010 10160 3040
rect 10190 3010 10200 3040
rect 10150 2985 10200 3010
rect 10150 2965 10165 2985
rect 10185 2965 10200 2985
rect 10150 2940 10200 2965
rect 10150 2910 10160 2940
rect 10190 2910 10200 2940
rect 10150 2885 10200 2910
rect 10150 2865 10165 2885
rect 10185 2865 10200 2885
rect 10150 2840 10200 2865
rect 10150 2810 10160 2840
rect 10190 2810 10200 2840
rect 10150 2785 10200 2810
rect 10150 2765 10165 2785
rect 10185 2765 10200 2785
rect 10150 2740 10200 2765
rect 10150 2710 10160 2740
rect 10190 2710 10200 2740
rect 10150 2685 10200 2710
rect 10150 2665 10165 2685
rect 10185 2665 10200 2685
rect 9850 2560 9860 2590
rect 9890 2560 9900 2590
rect 9850 2550 9900 2560
rect 10150 2590 10200 2665
rect 10300 3135 10350 3150
rect 10300 3115 10315 3135
rect 10335 3115 10350 3135
rect 10300 3085 10350 3115
rect 10300 3065 10315 3085
rect 10335 3065 10350 3085
rect 10300 3035 10350 3065
rect 10300 3015 10315 3035
rect 10335 3015 10350 3035
rect 10300 2985 10350 3015
rect 10300 2965 10315 2985
rect 10335 2965 10350 2985
rect 10300 2935 10350 2965
rect 10300 2915 10315 2935
rect 10335 2915 10350 2935
rect 10300 2885 10350 2915
rect 10300 2865 10315 2885
rect 10335 2865 10350 2885
rect 10300 2835 10350 2865
rect 10300 2815 10315 2835
rect 10335 2815 10350 2835
rect 10300 2785 10350 2815
rect 10300 2765 10315 2785
rect 10335 2765 10350 2785
rect 10300 2735 10350 2765
rect 10300 2715 10315 2735
rect 10335 2715 10350 2735
rect 10300 2685 10350 2715
rect 10300 2665 10315 2685
rect 10335 2665 10350 2685
rect 10300 2650 10350 2665
rect 10450 3140 10500 3310
rect 10600 3785 10650 3800
rect 10600 3765 10615 3785
rect 10635 3765 10650 3785
rect 10600 3735 10650 3765
rect 10600 3715 10615 3735
rect 10635 3715 10650 3735
rect 10600 3685 10650 3715
rect 10600 3665 10615 3685
rect 10635 3665 10650 3685
rect 10600 3635 10650 3665
rect 10600 3615 10615 3635
rect 10635 3615 10650 3635
rect 10600 3585 10650 3615
rect 10600 3565 10615 3585
rect 10635 3565 10650 3585
rect 10600 3535 10650 3565
rect 10600 3515 10615 3535
rect 10635 3515 10650 3535
rect 10600 3485 10650 3515
rect 10600 3465 10615 3485
rect 10635 3465 10650 3485
rect 10600 3435 10650 3465
rect 10600 3415 10615 3435
rect 10635 3415 10650 3435
rect 10600 3385 10650 3415
rect 10600 3365 10615 3385
rect 10635 3365 10650 3385
rect 10600 3335 10650 3365
rect 10600 3315 10615 3335
rect 10635 3315 10650 3335
rect 10600 3300 10650 3315
rect 10750 3785 10800 3860
rect 10750 3765 10765 3785
rect 10785 3765 10800 3785
rect 10750 3740 10800 3765
rect 10750 3710 10760 3740
rect 10790 3710 10800 3740
rect 10750 3685 10800 3710
rect 10750 3665 10765 3685
rect 10785 3665 10800 3685
rect 10750 3640 10800 3665
rect 10750 3610 10760 3640
rect 10790 3610 10800 3640
rect 10750 3585 10800 3610
rect 10750 3565 10765 3585
rect 10785 3565 10800 3585
rect 10750 3540 10800 3565
rect 10750 3510 10760 3540
rect 10790 3510 10800 3540
rect 10750 3485 10800 3510
rect 10750 3465 10765 3485
rect 10785 3465 10800 3485
rect 10750 3440 10800 3465
rect 10750 3410 10760 3440
rect 10790 3410 10800 3440
rect 10750 3385 10800 3410
rect 10750 3365 10765 3385
rect 10785 3365 10800 3385
rect 10750 3340 10800 3365
rect 10750 3310 10760 3340
rect 10790 3310 10800 3340
rect 10600 3240 10650 3250
rect 10600 3210 10610 3240
rect 10640 3210 10650 3240
rect 10600 3200 10650 3210
rect 10450 3110 10460 3140
rect 10490 3110 10500 3140
rect 10450 3085 10500 3110
rect 10450 3065 10465 3085
rect 10485 3065 10500 3085
rect 10450 3040 10500 3065
rect 10450 3010 10460 3040
rect 10490 3010 10500 3040
rect 10450 2985 10500 3010
rect 10450 2965 10465 2985
rect 10485 2965 10500 2985
rect 10450 2940 10500 2965
rect 10450 2910 10460 2940
rect 10490 2910 10500 2940
rect 10450 2885 10500 2910
rect 10450 2865 10465 2885
rect 10485 2865 10500 2885
rect 10450 2840 10500 2865
rect 10450 2810 10460 2840
rect 10490 2810 10500 2840
rect 10450 2785 10500 2810
rect 10450 2765 10465 2785
rect 10485 2765 10500 2785
rect 10450 2740 10500 2765
rect 10450 2710 10460 2740
rect 10490 2710 10500 2740
rect 10450 2685 10500 2710
rect 10450 2665 10465 2685
rect 10485 2665 10500 2685
rect 10150 2560 10160 2590
rect 10190 2560 10200 2590
rect 10150 2550 10200 2560
rect 10450 2590 10500 2665
rect 10600 3135 10650 3150
rect 10600 3115 10615 3135
rect 10635 3115 10650 3135
rect 10600 3085 10650 3115
rect 10600 3065 10615 3085
rect 10635 3065 10650 3085
rect 10600 3035 10650 3065
rect 10600 3015 10615 3035
rect 10635 3015 10650 3035
rect 10600 2985 10650 3015
rect 10600 2965 10615 2985
rect 10635 2965 10650 2985
rect 10600 2935 10650 2965
rect 10600 2915 10615 2935
rect 10635 2915 10650 2935
rect 10600 2885 10650 2915
rect 10600 2865 10615 2885
rect 10635 2865 10650 2885
rect 10600 2835 10650 2865
rect 10600 2815 10615 2835
rect 10635 2815 10650 2835
rect 10600 2785 10650 2815
rect 10600 2765 10615 2785
rect 10635 2765 10650 2785
rect 10600 2735 10650 2765
rect 10600 2715 10615 2735
rect 10635 2715 10650 2735
rect 10600 2685 10650 2715
rect 10600 2665 10615 2685
rect 10635 2665 10650 2685
rect 10600 2650 10650 2665
rect 10750 3140 10800 3310
rect 11350 4435 11400 4510
rect 11500 4540 11550 4550
rect 11500 4510 11510 4540
rect 11540 4510 11550 4540
rect 11500 4500 11550 4510
rect 11800 4540 11850 4550
rect 11800 4510 11810 4540
rect 11840 4510 11850 4540
rect 11800 4500 11850 4510
rect 11350 4415 11365 4435
rect 11385 4415 11400 4435
rect 11350 4385 11400 4415
rect 11350 4365 11365 4385
rect 11385 4365 11400 4385
rect 11350 4335 11400 4365
rect 11350 4315 11365 4335
rect 11385 4315 11400 4335
rect 11350 4285 11400 4315
rect 11350 4265 11365 4285
rect 11385 4265 11400 4285
rect 11350 4235 11400 4265
rect 11350 4215 11365 4235
rect 11385 4215 11400 4235
rect 11350 4185 11400 4215
rect 11350 4165 11365 4185
rect 11385 4165 11400 4185
rect 11350 4135 11400 4165
rect 11350 4115 11365 4135
rect 11385 4115 11400 4135
rect 11350 4085 11400 4115
rect 11350 4065 11365 4085
rect 11385 4065 11400 4085
rect 11350 4035 11400 4065
rect 11350 4015 11365 4035
rect 11385 4015 11400 4035
rect 11350 3985 11400 4015
rect 11350 3965 11365 3985
rect 11385 3965 11400 3985
rect 11350 3785 11400 3965
rect 11350 3765 11365 3785
rect 11385 3765 11400 3785
rect 11350 3735 11400 3765
rect 11350 3715 11365 3735
rect 11385 3715 11400 3735
rect 11350 3685 11400 3715
rect 11350 3665 11365 3685
rect 11385 3665 11400 3685
rect 11350 3635 11400 3665
rect 11350 3615 11365 3635
rect 11385 3615 11400 3635
rect 11350 3585 11400 3615
rect 11350 3565 11365 3585
rect 11385 3565 11400 3585
rect 11350 3535 11400 3565
rect 11350 3515 11365 3535
rect 11385 3515 11400 3535
rect 11350 3485 11400 3515
rect 11350 3465 11365 3485
rect 11385 3465 11400 3485
rect 11350 3435 11400 3465
rect 11350 3415 11365 3435
rect 11385 3415 11400 3435
rect 11350 3385 11400 3415
rect 11350 3365 11365 3385
rect 11385 3365 11400 3385
rect 11350 3335 11400 3365
rect 11350 3315 11365 3335
rect 11385 3315 11400 3335
rect 10900 3240 10950 3250
rect 10900 3210 10910 3240
rect 10940 3210 10950 3240
rect 10900 3200 10950 3210
rect 11200 3240 11250 3250
rect 11200 3210 11210 3240
rect 11240 3210 11250 3240
rect 11200 3200 11250 3210
rect 11350 3240 11400 3315
rect 11950 4440 12000 4610
rect 12550 5085 12600 5100
rect 12550 5065 12565 5085
rect 12585 5065 12600 5085
rect 12550 5035 12600 5065
rect 12550 5015 12565 5035
rect 12585 5015 12600 5035
rect 12550 4985 12600 5015
rect 12550 4965 12565 4985
rect 12585 4965 12600 4985
rect 12550 4935 12600 4965
rect 12550 4915 12565 4935
rect 12585 4915 12600 4935
rect 12550 4885 12600 4915
rect 12550 4865 12565 4885
rect 12585 4865 12600 4885
rect 12550 4835 12600 4865
rect 12550 4815 12565 4835
rect 12585 4815 12600 4835
rect 12550 4785 12600 4815
rect 12550 4765 12565 4785
rect 12585 4765 12600 4785
rect 12550 4735 12600 4765
rect 12550 4715 12565 4735
rect 12585 4715 12600 4735
rect 12550 4685 12600 4715
rect 12550 4665 12565 4685
rect 12585 4665 12600 4685
rect 12550 4635 12600 4665
rect 12550 4615 12565 4635
rect 12585 4615 12600 4635
rect 12100 4540 12150 4550
rect 12100 4510 12110 4540
rect 12140 4510 12150 4540
rect 12100 4500 12150 4510
rect 12400 4540 12450 4550
rect 12400 4510 12410 4540
rect 12440 4510 12450 4540
rect 12400 4500 12450 4510
rect 12550 4540 12600 4615
rect 13150 5085 13200 5160
rect 14350 5190 14400 5200
rect 14350 5160 14360 5190
rect 14390 5160 14400 5190
rect 13150 5065 13165 5085
rect 13185 5065 13200 5085
rect 13150 5040 13200 5065
rect 13150 5010 13160 5040
rect 13190 5010 13200 5040
rect 13150 4985 13200 5010
rect 13150 4965 13165 4985
rect 13185 4965 13200 4985
rect 13150 4940 13200 4965
rect 13150 4910 13160 4940
rect 13190 4910 13200 4940
rect 13150 4885 13200 4910
rect 13150 4865 13165 4885
rect 13185 4865 13200 4885
rect 13150 4840 13200 4865
rect 13150 4810 13160 4840
rect 13190 4810 13200 4840
rect 13150 4785 13200 4810
rect 13150 4765 13165 4785
rect 13185 4765 13200 4785
rect 13150 4740 13200 4765
rect 13150 4710 13160 4740
rect 13190 4710 13200 4740
rect 13150 4685 13200 4710
rect 13150 4665 13165 4685
rect 13185 4665 13200 4685
rect 13150 4640 13200 4665
rect 13150 4610 13160 4640
rect 13190 4610 13200 4640
rect 12550 4510 12560 4540
rect 12590 4510 12600 4540
rect 11950 4410 11960 4440
rect 11990 4410 12000 4440
rect 11950 4385 12000 4410
rect 11950 4365 11965 4385
rect 11985 4365 12000 4385
rect 11950 4340 12000 4365
rect 11950 4310 11960 4340
rect 11990 4310 12000 4340
rect 11950 4285 12000 4310
rect 11950 4265 11965 4285
rect 11985 4265 12000 4285
rect 11950 4240 12000 4265
rect 11950 4210 11960 4240
rect 11990 4210 12000 4240
rect 11950 4185 12000 4210
rect 11950 4165 11965 4185
rect 11985 4165 12000 4185
rect 11950 4140 12000 4165
rect 11950 4110 11960 4140
rect 11990 4110 12000 4140
rect 11950 4085 12000 4110
rect 11950 4065 11965 4085
rect 11985 4065 12000 4085
rect 11950 4040 12000 4065
rect 11950 4010 11960 4040
rect 11990 4010 12000 4040
rect 11950 3985 12000 4010
rect 11950 3965 11965 3985
rect 11985 3965 12000 3985
rect 11950 3890 12000 3965
rect 11950 3860 11960 3890
rect 11990 3860 12000 3890
rect 11950 3785 12000 3860
rect 11950 3765 11965 3785
rect 11985 3765 12000 3785
rect 11950 3740 12000 3765
rect 11950 3710 11960 3740
rect 11990 3710 12000 3740
rect 11950 3685 12000 3710
rect 11950 3665 11965 3685
rect 11985 3665 12000 3685
rect 11950 3640 12000 3665
rect 11950 3610 11960 3640
rect 11990 3610 12000 3640
rect 11950 3585 12000 3610
rect 11950 3565 11965 3585
rect 11985 3565 12000 3585
rect 11950 3540 12000 3565
rect 11950 3510 11960 3540
rect 11990 3510 12000 3540
rect 11950 3485 12000 3510
rect 11950 3465 11965 3485
rect 11985 3465 12000 3485
rect 11950 3440 12000 3465
rect 11950 3410 11960 3440
rect 11990 3410 12000 3440
rect 11950 3385 12000 3410
rect 11950 3365 11965 3385
rect 11985 3365 12000 3385
rect 11950 3340 12000 3365
rect 11950 3310 11960 3340
rect 11990 3310 12000 3340
rect 11350 3210 11360 3240
rect 11390 3210 11400 3240
rect 10750 3110 10760 3140
rect 10790 3110 10800 3140
rect 10750 3085 10800 3110
rect 10750 3065 10765 3085
rect 10785 3065 10800 3085
rect 10750 3040 10800 3065
rect 10750 3010 10760 3040
rect 10790 3010 10800 3040
rect 10750 2985 10800 3010
rect 10750 2965 10765 2985
rect 10785 2965 10800 2985
rect 10750 2940 10800 2965
rect 10750 2910 10760 2940
rect 10790 2910 10800 2940
rect 10750 2885 10800 2910
rect 10750 2865 10765 2885
rect 10785 2865 10800 2885
rect 10750 2840 10800 2865
rect 10750 2810 10760 2840
rect 10790 2810 10800 2840
rect 10750 2785 10800 2810
rect 10750 2765 10765 2785
rect 10785 2765 10800 2785
rect 10750 2740 10800 2765
rect 10750 2710 10760 2740
rect 10790 2710 10800 2740
rect 10750 2685 10800 2710
rect 10750 2665 10765 2685
rect 10785 2665 10800 2685
rect 10450 2560 10460 2590
rect 10490 2560 10500 2590
rect 10450 2550 10500 2560
rect 10750 2590 10800 2665
rect 11350 3135 11400 3210
rect 11500 3240 11550 3250
rect 11500 3210 11510 3240
rect 11540 3210 11550 3240
rect 11500 3200 11550 3210
rect 11800 3240 11850 3250
rect 11800 3210 11810 3240
rect 11840 3210 11850 3240
rect 11800 3200 11850 3210
rect 11350 3115 11365 3135
rect 11385 3115 11400 3135
rect 11350 3085 11400 3115
rect 11350 3065 11365 3085
rect 11385 3065 11400 3085
rect 11350 3035 11400 3065
rect 11350 3015 11365 3035
rect 11385 3015 11400 3035
rect 11350 2985 11400 3015
rect 11350 2965 11365 2985
rect 11385 2965 11400 2985
rect 11350 2935 11400 2965
rect 11350 2915 11365 2935
rect 11385 2915 11400 2935
rect 11350 2885 11400 2915
rect 11350 2865 11365 2885
rect 11385 2865 11400 2885
rect 11350 2835 11400 2865
rect 11350 2815 11365 2835
rect 11385 2815 11400 2835
rect 11350 2785 11400 2815
rect 11350 2765 11365 2785
rect 11385 2765 11400 2785
rect 11350 2735 11400 2765
rect 11350 2715 11365 2735
rect 11385 2715 11400 2735
rect 11350 2685 11400 2715
rect 11350 2665 11365 2685
rect 11385 2665 11400 2685
rect 11350 2650 11400 2665
rect 11950 3140 12000 3310
rect 12550 4435 12600 4510
rect 12700 4540 12750 4550
rect 12700 4510 12710 4540
rect 12740 4510 12750 4540
rect 12700 4500 12750 4510
rect 13000 4540 13050 4550
rect 13000 4510 13010 4540
rect 13040 4510 13050 4540
rect 13000 4500 13050 4510
rect 12550 4415 12565 4435
rect 12585 4415 12600 4435
rect 12550 4385 12600 4415
rect 12550 4365 12565 4385
rect 12585 4365 12600 4385
rect 12550 4335 12600 4365
rect 12550 4315 12565 4335
rect 12585 4315 12600 4335
rect 12550 4285 12600 4315
rect 12550 4265 12565 4285
rect 12585 4265 12600 4285
rect 12550 4235 12600 4265
rect 12550 4215 12565 4235
rect 12585 4215 12600 4235
rect 12550 4185 12600 4215
rect 12550 4165 12565 4185
rect 12585 4165 12600 4185
rect 12550 4135 12600 4165
rect 12550 4115 12565 4135
rect 12585 4115 12600 4135
rect 12550 4085 12600 4115
rect 12550 4065 12565 4085
rect 12585 4065 12600 4085
rect 12550 4035 12600 4065
rect 12550 4015 12565 4035
rect 12585 4015 12600 4035
rect 12550 3985 12600 4015
rect 12550 3965 12565 3985
rect 12585 3965 12600 3985
rect 12550 3785 12600 3965
rect 12550 3765 12565 3785
rect 12585 3765 12600 3785
rect 12550 3735 12600 3765
rect 12550 3715 12565 3735
rect 12585 3715 12600 3735
rect 12550 3685 12600 3715
rect 12550 3665 12565 3685
rect 12585 3665 12600 3685
rect 12550 3635 12600 3665
rect 12550 3615 12565 3635
rect 12585 3615 12600 3635
rect 12550 3585 12600 3615
rect 12550 3565 12565 3585
rect 12585 3565 12600 3585
rect 12550 3535 12600 3565
rect 12550 3515 12565 3535
rect 12585 3515 12600 3535
rect 12550 3485 12600 3515
rect 12550 3465 12565 3485
rect 12585 3465 12600 3485
rect 12550 3435 12600 3465
rect 12550 3415 12565 3435
rect 12585 3415 12600 3435
rect 12550 3385 12600 3415
rect 12550 3365 12565 3385
rect 12585 3365 12600 3385
rect 12550 3335 12600 3365
rect 12550 3315 12565 3335
rect 12585 3315 12600 3335
rect 12100 3240 12150 3250
rect 12100 3210 12110 3240
rect 12140 3210 12150 3240
rect 12100 3200 12150 3210
rect 12400 3240 12450 3250
rect 12400 3210 12410 3240
rect 12440 3210 12450 3240
rect 12400 3200 12450 3210
rect 12550 3240 12600 3315
rect 13150 4440 13200 4610
rect 13750 5085 13800 5100
rect 13750 5065 13765 5085
rect 13785 5065 13800 5085
rect 13750 5035 13800 5065
rect 13750 5015 13765 5035
rect 13785 5015 13800 5035
rect 13750 4985 13800 5015
rect 13750 4965 13765 4985
rect 13785 4965 13800 4985
rect 13750 4935 13800 4965
rect 13750 4915 13765 4935
rect 13785 4915 13800 4935
rect 13750 4885 13800 4915
rect 13750 4865 13765 4885
rect 13785 4865 13800 4885
rect 13750 4835 13800 4865
rect 13750 4815 13765 4835
rect 13785 4815 13800 4835
rect 13750 4785 13800 4815
rect 13750 4765 13765 4785
rect 13785 4765 13800 4785
rect 13750 4735 13800 4765
rect 13750 4715 13765 4735
rect 13785 4715 13800 4735
rect 13750 4685 13800 4715
rect 13750 4665 13765 4685
rect 13785 4665 13800 4685
rect 13750 4635 13800 4665
rect 13750 4615 13765 4635
rect 13785 4615 13800 4635
rect 13300 4540 13350 4550
rect 13300 4510 13310 4540
rect 13340 4510 13350 4540
rect 13300 4500 13350 4510
rect 13600 4540 13650 4550
rect 13600 4510 13610 4540
rect 13640 4510 13650 4540
rect 13600 4500 13650 4510
rect 13750 4540 13800 4615
rect 14350 5085 14400 5160
rect 15550 5190 15600 5200
rect 15550 5160 15560 5190
rect 15590 5160 15600 5190
rect 14350 5065 14365 5085
rect 14385 5065 14400 5085
rect 14350 5040 14400 5065
rect 14350 5010 14360 5040
rect 14390 5010 14400 5040
rect 14350 4985 14400 5010
rect 14350 4965 14365 4985
rect 14385 4965 14400 4985
rect 14350 4940 14400 4965
rect 14350 4910 14360 4940
rect 14390 4910 14400 4940
rect 14350 4885 14400 4910
rect 14350 4865 14365 4885
rect 14385 4865 14400 4885
rect 14350 4840 14400 4865
rect 14350 4810 14360 4840
rect 14390 4810 14400 4840
rect 14350 4785 14400 4810
rect 14350 4765 14365 4785
rect 14385 4765 14400 4785
rect 14350 4740 14400 4765
rect 14350 4710 14360 4740
rect 14390 4710 14400 4740
rect 14350 4685 14400 4710
rect 14350 4665 14365 4685
rect 14385 4665 14400 4685
rect 14350 4640 14400 4665
rect 14350 4610 14360 4640
rect 14390 4610 14400 4640
rect 13750 4510 13760 4540
rect 13790 4510 13800 4540
rect 13150 4410 13160 4440
rect 13190 4410 13200 4440
rect 13150 4385 13200 4410
rect 13150 4365 13165 4385
rect 13185 4365 13200 4385
rect 13150 4340 13200 4365
rect 13150 4310 13160 4340
rect 13190 4310 13200 4340
rect 13150 4285 13200 4310
rect 13150 4265 13165 4285
rect 13185 4265 13200 4285
rect 13150 4240 13200 4265
rect 13150 4210 13160 4240
rect 13190 4210 13200 4240
rect 13150 4185 13200 4210
rect 13150 4165 13165 4185
rect 13185 4165 13200 4185
rect 13150 4140 13200 4165
rect 13150 4110 13160 4140
rect 13190 4110 13200 4140
rect 13150 4085 13200 4110
rect 13150 4065 13165 4085
rect 13185 4065 13200 4085
rect 13150 4040 13200 4065
rect 13150 4010 13160 4040
rect 13190 4010 13200 4040
rect 13150 3985 13200 4010
rect 13150 3965 13165 3985
rect 13185 3965 13200 3985
rect 13150 3890 13200 3965
rect 13150 3860 13160 3890
rect 13190 3860 13200 3890
rect 13150 3785 13200 3860
rect 13150 3765 13165 3785
rect 13185 3765 13200 3785
rect 13150 3740 13200 3765
rect 13150 3710 13160 3740
rect 13190 3710 13200 3740
rect 13150 3685 13200 3710
rect 13150 3665 13165 3685
rect 13185 3665 13200 3685
rect 13150 3640 13200 3665
rect 13150 3610 13160 3640
rect 13190 3610 13200 3640
rect 13150 3585 13200 3610
rect 13150 3565 13165 3585
rect 13185 3565 13200 3585
rect 13150 3540 13200 3565
rect 13150 3510 13160 3540
rect 13190 3510 13200 3540
rect 13150 3485 13200 3510
rect 13150 3465 13165 3485
rect 13185 3465 13200 3485
rect 13150 3440 13200 3465
rect 13150 3410 13160 3440
rect 13190 3410 13200 3440
rect 13150 3385 13200 3410
rect 13150 3365 13165 3385
rect 13185 3365 13200 3385
rect 13150 3340 13200 3365
rect 13150 3310 13160 3340
rect 13190 3310 13200 3340
rect 12550 3210 12560 3240
rect 12590 3210 12600 3240
rect 11950 3110 11960 3140
rect 11990 3110 12000 3140
rect 11950 3085 12000 3110
rect 11950 3065 11965 3085
rect 11985 3065 12000 3085
rect 11950 3040 12000 3065
rect 11950 3010 11960 3040
rect 11990 3010 12000 3040
rect 11950 2985 12000 3010
rect 11950 2965 11965 2985
rect 11985 2965 12000 2985
rect 11950 2940 12000 2965
rect 11950 2910 11960 2940
rect 11990 2910 12000 2940
rect 11950 2885 12000 2910
rect 11950 2865 11965 2885
rect 11985 2865 12000 2885
rect 11950 2840 12000 2865
rect 11950 2810 11960 2840
rect 11990 2810 12000 2840
rect 11950 2785 12000 2810
rect 11950 2765 11965 2785
rect 11985 2765 12000 2785
rect 11950 2740 12000 2765
rect 11950 2710 11960 2740
rect 11990 2710 12000 2740
rect 11950 2685 12000 2710
rect 11950 2665 11965 2685
rect 11985 2665 12000 2685
rect 10750 2560 10760 2590
rect 10790 2560 10800 2590
rect 10750 2550 10800 2560
rect 11950 2590 12000 2665
rect 12550 3135 12600 3210
rect 12700 3240 12750 3250
rect 12700 3210 12710 3240
rect 12740 3210 12750 3240
rect 12700 3200 12750 3210
rect 13000 3240 13050 3250
rect 13000 3210 13010 3240
rect 13040 3210 13050 3240
rect 13000 3200 13050 3210
rect 12550 3115 12565 3135
rect 12585 3115 12600 3135
rect 12550 3085 12600 3115
rect 12550 3065 12565 3085
rect 12585 3065 12600 3085
rect 12550 3035 12600 3065
rect 12550 3015 12565 3035
rect 12585 3015 12600 3035
rect 12550 2985 12600 3015
rect 12550 2965 12565 2985
rect 12585 2965 12600 2985
rect 12550 2935 12600 2965
rect 12550 2915 12565 2935
rect 12585 2915 12600 2935
rect 12550 2885 12600 2915
rect 12550 2865 12565 2885
rect 12585 2865 12600 2885
rect 12550 2835 12600 2865
rect 12550 2815 12565 2835
rect 12585 2815 12600 2835
rect 12550 2785 12600 2815
rect 12550 2765 12565 2785
rect 12585 2765 12600 2785
rect 12550 2735 12600 2765
rect 12550 2715 12565 2735
rect 12585 2715 12600 2735
rect 12550 2685 12600 2715
rect 12550 2665 12565 2685
rect 12585 2665 12600 2685
rect 12550 2650 12600 2665
rect 13150 3140 13200 3310
rect 13750 4435 13800 4510
rect 13900 4540 13950 4550
rect 13900 4510 13910 4540
rect 13940 4510 13950 4540
rect 13900 4500 13950 4510
rect 14200 4540 14250 4550
rect 14200 4510 14210 4540
rect 14240 4510 14250 4540
rect 14200 4500 14250 4510
rect 13750 4415 13765 4435
rect 13785 4415 13800 4435
rect 13750 4385 13800 4415
rect 13750 4365 13765 4385
rect 13785 4365 13800 4385
rect 13750 4335 13800 4365
rect 13750 4315 13765 4335
rect 13785 4315 13800 4335
rect 13750 4285 13800 4315
rect 13750 4265 13765 4285
rect 13785 4265 13800 4285
rect 13750 4235 13800 4265
rect 13750 4215 13765 4235
rect 13785 4215 13800 4235
rect 13750 4185 13800 4215
rect 13750 4165 13765 4185
rect 13785 4165 13800 4185
rect 13750 4135 13800 4165
rect 13750 4115 13765 4135
rect 13785 4115 13800 4135
rect 13750 4085 13800 4115
rect 13750 4065 13765 4085
rect 13785 4065 13800 4085
rect 13750 4035 13800 4065
rect 13750 4015 13765 4035
rect 13785 4015 13800 4035
rect 13750 3985 13800 4015
rect 13750 3965 13765 3985
rect 13785 3965 13800 3985
rect 13750 3785 13800 3965
rect 13750 3765 13765 3785
rect 13785 3765 13800 3785
rect 13750 3735 13800 3765
rect 13750 3715 13765 3735
rect 13785 3715 13800 3735
rect 13750 3685 13800 3715
rect 13750 3665 13765 3685
rect 13785 3665 13800 3685
rect 13750 3635 13800 3665
rect 13750 3615 13765 3635
rect 13785 3615 13800 3635
rect 13750 3585 13800 3615
rect 13750 3565 13765 3585
rect 13785 3565 13800 3585
rect 13750 3535 13800 3565
rect 13750 3515 13765 3535
rect 13785 3515 13800 3535
rect 13750 3485 13800 3515
rect 13750 3465 13765 3485
rect 13785 3465 13800 3485
rect 13750 3435 13800 3465
rect 13750 3415 13765 3435
rect 13785 3415 13800 3435
rect 13750 3385 13800 3415
rect 13750 3365 13765 3385
rect 13785 3365 13800 3385
rect 13750 3335 13800 3365
rect 13750 3315 13765 3335
rect 13785 3315 13800 3335
rect 13300 3240 13350 3250
rect 13300 3210 13310 3240
rect 13340 3210 13350 3240
rect 13300 3200 13350 3210
rect 13600 3240 13650 3250
rect 13600 3210 13610 3240
rect 13640 3210 13650 3240
rect 13600 3200 13650 3210
rect 13750 3240 13800 3315
rect 14350 4440 14400 4610
rect 14950 5085 15000 5100
rect 14950 5065 14965 5085
rect 14985 5065 15000 5085
rect 14950 5035 15000 5065
rect 14950 5015 14965 5035
rect 14985 5015 15000 5035
rect 14950 4985 15000 5015
rect 14950 4965 14965 4985
rect 14985 4965 15000 4985
rect 14950 4935 15000 4965
rect 14950 4915 14965 4935
rect 14985 4915 15000 4935
rect 14950 4885 15000 4915
rect 14950 4865 14965 4885
rect 14985 4865 15000 4885
rect 14950 4835 15000 4865
rect 14950 4815 14965 4835
rect 14985 4815 15000 4835
rect 14950 4785 15000 4815
rect 14950 4765 14965 4785
rect 14985 4765 15000 4785
rect 14950 4735 15000 4765
rect 14950 4715 14965 4735
rect 14985 4715 15000 4735
rect 14950 4685 15000 4715
rect 14950 4665 14965 4685
rect 14985 4665 15000 4685
rect 14950 4635 15000 4665
rect 14950 4615 14965 4635
rect 14985 4615 15000 4635
rect 14500 4540 14550 4550
rect 14500 4510 14510 4540
rect 14540 4510 14550 4540
rect 14500 4500 14550 4510
rect 14800 4540 14850 4550
rect 14800 4510 14810 4540
rect 14840 4510 14850 4540
rect 14800 4500 14850 4510
rect 14950 4540 15000 4615
rect 15550 5085 15600 5160
rect 17950 5190 18000 5200
rect 17950 5160 17960 5190
rect 17990 5160 18000 5190
rect 17950 5100 18000 5160
rect 20350 5190 20400 5200
rect 20350 5160 20360 5190
rect 20390 5160 20400 5190
rect 15550 5065 15565 5085
rect 15585 5065 15600 5085
rect 15550 5040 15600 5065
rect 15550 5010 15560 5040
rect 15590 5010 15600 5040
rect 15550 4985 15600 5010
rect 15550 4965 15565 4985
rect 15585 4965 15600 4985
rect 15550 4940 15600 4965
rect 15550 4910 15560 4940
rect 15590 4910 15600 4940
rect 15550 4885 15600 4910
rect 15550 4865 15565 4885
rect 15585 4865 15600 4885
rect 15550 4840 15600 4865
rect 15550 4810 15560 4840
rect 15590 4810 15600 4840
rect 15550 4785 15600 4810
rect 15550 4765 15565 4785
rect 15585 4765 15600 4785
rect 15550 4740 15600 4765
rect 15550 4710 15560 4740
rect 15590 4710 15600 4740
rect 15550 4685 15600 4710
rect 15550 4665 15565 4685
rect 15585 4665 15600 4685
rect 15550 4640 15600 4665
rect 15550 4610 15560 4640
rect 15590 4610 15600 4640
rect 14950 4510 14960 4540
rect 14990 4510 15000 4540
rect 14350 4410 14360 4440
rect 14390 4410 14400 4440
rect 14350 4385 14400 4410
rect 14350 4365 14365 4385
rect 14385 4365 14400 4385
rect 14350 4340 14400 4365
rect 14350 4310 14360 4340
rect 14390 4310 14400 4340
rect 14350 4285 14400 4310
rect 14350 4265 14365 4285
rect 14385 4265 14400 4285
rect 14350 4240 14400 4265
rect 14350 4210 14360 4240
rect 14390 4210 14400 4240
rect 14350 4185 14400 4210
rect 14350 4165 14365 4185
rect 14385 4165 14400 4185
rect 14350 4140 14400 4165
rect 14350 4110 14360 4140
rect 14390 4110 14400 4140
rect 14350 4085 14400 4110
rect 14350 4065 14365 4085
rect 14385 4065 14400 4085
rect 14350 4040 14400 4065
rect 14350 4010 14360 4040
rect 14390 4010 14400 4040
rect 14350 3985 14400 4010
rect 14350 3965 14365 3985
rect 14385 3965 14400 3985
rect 14350 3890 14400 3965
rect 14350 3860 14360 3890
rect 14390 3860 14400 3890
rect 14350 3785 14400 3860
rect 14350 3765 14365 3785
rect 14385 3765 14400 3785
rect 14350 3740 14400 3765
rect 14350 3710 14360 3740
rect 14390 3710 14400 3740
rect 14350 3685 14400 3710
rect 14350 3665 14365 3685
rect 14385 3665 14400 3685
rect 14350 3640 14400 3665
rect 14350 3610 14360 3640
rect 14390 3610 14400 3640
rect 14350 3585 14400 3610
rect 14350 3565 14365 3585
rect 14385 3565 14400 3585
rect 14350 3540 14400 3565
rect 14350 3510 14360 3540
rect 14390 3510 14400 3540
rect 14350 3485 14400 3510
rect 14350 3465 14365 3485
rect 14385 3465 14400 3485
rect 14350 3440 14400 3465
rect 14350 3410 14360 3440
rect 14390 3410 14400 3440
rect 14350 3385 14400 3410
rect 14350 3365 14365 3385
rect 14385 3365 14400 3385
rect 14350 3340 14400 3365
rect 14350 3310 14360 3340
rect 14390 3310 14400 3340
rect 13750 3210 13760 3240
rect 13790 3210 13800 3240
rect 13150 3110 13160 3140
rect 13190 3110 13200 3140
rect 13150 3085 13200 3110
rect 13150 3065 13165 3085
rect 13185 3065 13200 3085
rect 13150 3040 13200 3065
rect 13150 3010 13160 3040
rect 13190 3010 13200 3040
rect 13150 2985 13200 3010
rect 13150 2965 13165 2985
rect 13185 2965 13200 2985
rect 13150 2940 13200 2965
rect 13150 2910 13160 2940
rect 13190 2910 13200 2940
rect 13150 2885 13200 2910
rect 13150 2865 13165 2885
rect 13185 2865 13200 2885
rect 13150 2840 13200 2865
rect 13150 2810 13160 2840
rect 13190 2810 13200 2840
rect 13150 2785 13200 2810
rect 13150 2765 13165 2785
rect 13185 2765 13200 2785
rect 13150 2740 13200 2765
rect 13150 2710 13160 2740
rect 13190 2710 13200 2740
rect 13150 2685 13200 2710
rect 13150 2665 13165 2685
rect 13185 2665 13200 2685
rect 11950 2560 11960 2590
rect 11990 2560 12000 2590
rect 11950 2550 12000 2560
rect 13150 2590 13200 2665
rect 13750 3135 13800 3210
rect 13900 3240 13950 3250
rect 13900 3210 13910 3240
rect 13940 3210 13950 3240
rect 13900 3200 13950 3210
rect 14200 3240 14250 3250
rect 14200 3210 14210 3240
rect 14240 3210 14250 3240
rect 14200 3200 14250 3210
rect 13750 3115 13765 3135
rect 13785 3115 13800 3135
rect 13750 3085 13800 3115
rect 13750 3065 13765 3085
rect 13785 3065 13800 3085
rect 13750 3035 13800 3065
rect 13750 3015 13765 3035
rect 13785 3015 13800 3035
rect 13750 2985 13800 3015
rect 13750 2965 13765 2985
rect 13785 2965 13800 2985
rect 13750 2935 13800 2965
rect 13750 2915 13765 2935
rect 13785 2915 13800 2935
rect 13750 2885 13800 2915
rect 13750 2865 13765 2885
rect 13785 2865 13800 2885
rect 13750 2835 13800 2865
rect 13750 2815 13765 2835
rect 13785 2815 13800 2835
rect 13750 2785 13800 2815
rect 13750 2765 13765 2785
rect 13785 2765 13800 2785
rect 13750 2735 13800 2765
rect 13750 2715 13765 2735
rect 13785 2715 13800 2735
rect 13750 2685 13800 2715
rect 13750 2665 13765 2685
rect 13785 2665 13800 2685
rect 13750 2650 13800 2665
rect 14350 3140 14400 3310
rect 14950 4435 15000 4510
rect 15100 4540 15150 4550
rect 15100 4510 15110 4540
rect 15140 4510 15150 4540
rect 15100 4500 15150 4510
rect 15400 4540 15450 4550
rect 15400 4510 15410 4540
rect 15440 4510 15450 4540
rect 15400 4500 15450 4510
rect 14950 4415 14965 4435
rect 14985 4415 15000 4435
rect 14950 4385 15000 4415
rect 14950 4365 14965 4385
rect 14985 4365 15000 4385
rect 14950 4335 15000 4365
rect 14950 4315 14965 4335
rect 14985 4315 15000 4335
rect 14950 4285 15000 4315
rect 14950 4265 14965 4285
rect 14985 4265 15000 4285
rect 14950 4235 15000 4265
rect 14950 4215 14965 4235
rect 14985 4215 15000 4235
rect 14950 4185 15000 4215
rect 14950 4165 14965 4185
rect 14985 4165 15000 4185
rect 14950 4135 15000 4165
rect 14950 4115 14965 4135
rect 14985 4115 15000 4135
rect 14950 4085 15000 4115
rect 14950 4065 14965 4085
rect 14985 4065 15000 4085
rect 14950 4035 15000 4065
rect 14950 4015 14965 4035
rect 14985 4015 15000 4035
rect 14950 3985 15000 4015
rect 14950 3965 14965 3985
rect 14985 3965 15000 3985
rect 14950 3785 15000 3965
rect 14950 3765 14965 3785
rect 14985 3765 15000 3785
rect 14950 3735 15000 3765
rect 14950 3715 14965 3735
rect 14985 3715 15000 3735
rect 14950 3685 15000 3715
rect 14950 3665 14965 3685
rect 14985 3665 15000 3685
rect 14950 3635 15000 3665
rect 14950 3615 14965 3635
rect 14985 3615 15000 3635
rect 14950 3585 15000 3615
rect 14950 3565 14965 3585
rect 14985 3565 15000 3585
rect 14950 3535 15000 3565
rect 14950 3515 14965 3535
rect 14985 3515 15000 3535
rect 14950 3485 15000 3515
rect 14950 3465 14965 3485
rect 14985 3465 15000 3485
rect 14950 3435 15000 3465
rect 14950 3415 14965 3435
rect 14985 3415 15000 3435
rect 14950 3385 15000 3415
rect 14950 3365 14965 3385
rect 14985 3365 15000 3385
rect 14950 3335 15000 3365
rect 14950 3315 14965 3335
rect 14985 3315 15000 3335
rect 14500 3240 14550 3250
rect 14500 3210 14510 3240
rect 14540 3210 14550 3240
rect 14500 3200 14550 3210
rect 14800 3240 14850 3250
rect 14800 3210 14810 3240
rect 14840 3210 14850 3240
rect 14800 3200 14850 3210
rect 14950 3240 15000 3315
rect 15550 4440 15600 4610
rect 16150 5085 19800 5100
rect 16150 5065 16165 5085
rect 16185 5065 16465 5085
rect 16485 5065 16765 5085
rect 16785 5065 17065 5085
rect 17085 5065 17365 5085
rect 17385 5065 18565 5085
rect 18585 5065 18865 5085
rect 18885 5065 19165 5085
rect 19185 5065 19465 5085
rect 19485 5065 19765 5085
rect 19785 5065 19800 5085
rect 16150 5050 19800 5065
rect 16150 5035 16200 5050
rect 16150 5015 16165 5035
rect 16185 5015 16200 5035
rect 16150 4985 16200 5015
rect 16450 5035 16500 5050
rect 16450 5015 16465 5035
rect 16485 5015 16500 5035
rect 16150 4965 16165 4985
rect 16185 4965 16200 4985
rect 16150 4935 16200 4965
rect 16150 4915 16165 4935
rect 16185 4915 16200 4935
rect 16150 4885 16200 4915
rect 16150 4865 16165 4885
rect 16185 4865 16200 4885
rect 16150 4835 16200 4865
rect 16150 4815 16165 4835
rect 16185 4815 16200 4835
rect 16150 4785 16200 4815
rect 16150 4765 16165 4785
rect 16185 4765 16200 4785
rect 16150 4735 16200 4765
rect 16150 4715 16165 4735
rect 16185 4715 16200 4735
rect 16150 4685 16200 4715
rect 16150 4665 16165 4685
rect 16185 4665 16200 4685
rect 16150 4635 16200 4665
rect 16150 4615 16165 4635
rect 16185 4615 16200 4635
rect 15700 4540 15750 4550
rect 15700 4510 15710 4540
rect 15740 4510 15750 4540
rect 15700 4500 15750 4510
rect 16000 4540 16050 4550
rect 16000 4510 16010 4540
rect 16040 4510 16050 4540
rect 16000 4500 16050 4510
rect 15550 4410 15560 4440
rect 15590 4410 15600 4440
rect 15550 4385 15600 4410
rect 15550 4365 15565 4385
rect 15585 4365 15600 4385
rect 15550 4340 15600 4365
rect 15550 4310 15560 4340
rect 15590 4310 15600 4340
rect 15550 4285 15600 4310
rect 15550 4265 15565 4285
rect 15585 4265 15600 4285
rect 15550 4240 15600 4265
rect 15550 4210 15560 4240
rect 15590 4210 15600 4240
rect 15550 4185 15600 4210
rect 15550 4165 15565 4185
rect 15585 4165 15600 4185
rect 15550 4140 15600 4165
rect 15550 4110 15560 4140
rect 15590 4110 15600 4140
rect 15550 4085 15600 4110
rect 15550 4065 15565 4085
rect 15585 4065 15600 4085
rect 15550 4040 15600 4065
rect 15550 4010 15560 4040
rect 15590 4010 15600 4040
rect 15550 3985 15600 4010
rect 15550 3965 15565 3985
rect 15585 3965 15600 3985
rect 15550 3890 15600 3965
rect 16150 4435 16200 4615
rect 16300 4985 16350 5000
rect 16300 4965 16315 4985
rect 16335 4965 16350 4985
rect 16300 4935 16350 4965
rect 16300 4915 16315 4935
rect 16335 4915 16350 4935
rect 16300 4885 16350 4915
rect 16300 4865 16315 4885
rect 16335 4865 16350 4885
rect 16300 4835 16350 4865
rect 16300 4815 16315 4835
rect 16335 4815 16350 4835
rect 16300 4785 16350 4815
rect 16300 4765 16315 4785
rect 16335 4765 16350 4785
rect 16300 4735 16350 4765
rect 16300 4715 16315 4735
rect 16335 4715 16350 4735
rect 16300 4685 16350 4715
rect 16450 4985 16500 5015
rect 16750 5035 16800 5050
rect 16750 5015 16765 5035
rect 16785 5015 16800 5035
rect 16450 4965 16465 4985
rect 16485 4965 16500 4985
rect 16450 4935 16500 4965
rect 16450 4915 16465 4935
rect 16485 4915 16500 4935
rect 16450 4885 16500 4915
rect 16450 4865 16465 4885
rect 16485 4865 16500 4885
rect 16450 4835 16500 4865
rect 16450 4815 16465 4835
rect 16485 4815 16500 4835
rect 16450 4785 16500 4815
rect 16450 4765 16465 4785
rect 16485 4765 16500 4785
rect 16450 4735 16500 4765
rect 16450 4715 16465 4735
rect 16485 4715 16500 4735
rect 16450 4700 16500 4715
rect 16600 4985 16650 5000
rect 16600 4965 16615 4985
rect 16635 4965 16650 4985
rect 16600 4935 16650 4965
rect 16600 4915 16615 4935
rect 16635 4915 16650 4935
rect 16600 4885 16650 4915
rect 16600 4865 16615 4885
rect 16635 4865 16650 4885
rect 16600 4835 16650 4865
rect 16600 4815 16615 4835
rect 16635 4815 16650 4835
rect 16600 4785 16650 4815
rect 16600 4765 16615 4785
rect 16635 4765 16650 4785
rect 16600 4735 16650 4765
rect 16600 4715 16615 4735
rect 16635 4715 16650 4735
rect 16300 4665 16315 4685
rect 16335 4665 16350 4685
rect 16300 4650 16350 4665
rect 16600 4685 16650 4715
rect 16750 4985 16800 5015
rect 17050 5035 17100 5050
rect 17050 5015 17065 5035
rect 17085 5015 17100 5035
rect 16750 4965 16765 4985
rect 16785 4965 16800 4985
rect 16750 4935 16800 4965
rect 16750 4915 16765 4935
rect 16785 4915 16800 4935
rect 16750 4885 16800 4915
rect 16750 4865 16765 4885
rect 16785 4865 16800 4885
rect 16750 4835 16800 4865
rect 16750 4815 16765 4835
rect 16785 4815 16800 4835
rect 16750 4785 16800 4815
rect 16750 4765 16765 4785
rect 16785 4765 16800 4785
rect 16750 4735 16800 4765
rect 16750 4715 16765 4735
rect 16785 4715 16800 4735
rect 16750 4700 16800 4715
rect 16900 4985 16950 5000
rect 16900 4965 16915 4985
rect 16935 4965 16950 4985
rect 16900 4935 16950 4965
rect 16900 4915 16915 4935
rect 16935 4915 16950 4935
rect 16900 4885 16950 4915
rect 16900 4865 16915 4885
rect 16935 4865 16950 4885
rect 16900 4835 16950 4865
rect 16900 4815 16915 4835
rect 16935 4815 16950 4835
rect 16900 4785 16950 4815
rect 16900 4765 16915 4785
rect 16935 4765 16950 4785
rect 16900 4735 16950 4765
rect 16900 4715 16915 4735
rect 16935 4715 16950 4735
rect 16600 4665 16615 4685
rect 16635 4665 16650 4685
rect 16600 4650 16650 4665
rect 16900 4685 16950 4715
rect 17050 4985 17100 5015
rect 17350 5035 17400 5050
rect 17350 5015 17365 5035
rect 17385 5015 17400 5035
rect 17050 4965 17065 4985
rect 17085 4965 17100 4985
rect 17050 4935 17100 4965
rect 17050 4915 17065 4935
rect 17085 4915 17100 4935
rect 17050 4885 17100 4915
rect 17050 4865 17065 4885
rect 17085 4865 17100 4885
rect 17050 4835 17100 4865
rect 17050 4815 17065 4835
rect 17085 4815 17100 4835
rect 17050 4785 17100 4815
rect 17050 4765 17065 4785
rect 17085 4765 17100 4785
rect 17050 4735 17100 4765
rect 17050 4715 17065 4735
rect 17085 4715 17100 4735
rect 17050 4700 17100 4715
rect 17200 4985 17250 5000
rect 17200 4965 17215 4985
rect 17235 4965 17250 4985
rect 17200 4935 17250 4965
rect 17200 4915 17215 4935
rect 17235 4915 17250 4935
rect 17200 4885 17250 4915
rect 17200 4865 17215 4885
rect 17235 4865 17250 4885
rect 17200 4835 17250 4865
rect 17200 4815 17215 4835
rect 17235 4815 17250 4835
rect 17200 4785 17250 4815
rect 17200 4765 17215 4785
rect 17235 4765 17250 4785
rect 17200 4735 17250 4765
rect 17200 4715 17215 4735
rect 17235 4715 17250 4735
rect 16900 4665 16915 4685
rect 16935 4665 16950 4685
rect 16900 4650 16950 4665
rect 17200 4685 17250 4715
rect 17200 4665 17215 4685
rect 17235 4665 17250 4685
rect 17200 4650 17250 4665
rect 16300 4635 17250 4650
rect 16300 4615 16315 4635
rect 16335 4615 16615 4635
rect 16635 4615 16915 4635
rect 16935 4615 17215 4635
rect 17235 4615 17250 4635
rect 16300 4600 17250 4615
rect 17350 4985 17400 5015
rect 18550 5035 18600 5050
rect 18550 5015 18565 5035
rect 18585 5015 18600 5035
rect 17350 4965 17365 4985
rect 17385 4965 17400 4985
rect 17350 4935 17400 4965
rect 17350 4915 17365 4935
rect 17385 4915 17400 4935
rect 17350 4885 17400 4915
rect 17350 4865 17365 4885
rect 17385 4865 17400 4885
rect 17350 4835 17400 4865
rect 17350 4815 17365 4835
rect 17385 4815 17400 4835
rect 17350 4785 17400 4815
rect 17350 4765 17365 4785
rect 17385 4765 17400 4785
rect 17350 4735 17400 4765
rect 17350 4715 17365 4735
rect 17385 4715 17400 4735
rect 17350 4685 17400 4715
rect 17350 4665 17365 4685
rect 17385 4665 17400 4685
rect 17350 4635 17400 4665
rect 17350 4615 17365 4635
rect 17385 4615 17400 4635
rect 16300 4540 16350 4550
rect 16300 4510 16310 4540
rect 16340 4510 16350 4540
rect 16300 4500 16350 4510
rect 16450 4450 16500 4600
rect 16600 4540 16650 4550
rect 16600 4510 16610 4540
rect 16640 4510 16650 4540
rect 16600 4500 16650 4510
rect 16750 4540 16800 4600
rect 16750 4510 16760 4540
rect 16790 4510 16800 4540
rect 16750 4450 16800 4510
rect 16900 4540 16950 4550
rect 16900 4510 16910 4540
rect 16940 4510 16950 4540
rect 16900 4500 16950 4510
rect 17050 4450 17100 4600
rect 17200 4540 17250 4550
rect 17200 4510 17210 4540
rect 17240 4510 17250 4540
rect 17200 4500 17250 4510
rect 16150 4415 16165 4435
rect 16185 4415 16200 4435
rect 16150 4385 16200 4415
rect 16150 4365 16165 4385
rect 16185 4365 16200 4385
rect 16150 4335 16200 4365
rect 16150 4315 16165 4335
rect 16185 4315 16200 4335
rect 16150 4285 16200 4315
rect 16150 4265 16165 4285
rect 16185 4265 16200 4285
rect 16150 4235 16200 4265
rect 16150 4215 16165 4235
rect 16185 4215 16200 4235
rect 16150 4185 16200 4215
rect 16150 4165 16165 4185
rect 16185 4165 16200 4185
rect 16150 4135 16200 4165
rect 16150 4115 16165 4135
rect 16185 4115 16200 4135
rect 16150 4085 16200 4115
rect 16150 4065 16165 4085
rect 16185 4065 16200 4085
rect 16150 4035 16200 4065
rect 16300 4435 17250 4450
rect 16300 4415 16315 4435
rect 16335 4415 16615 4435
rect 16635 4415 16915 4435
rect 16935 4415 17215 4435
rect 17235 4415 17250 4435
rect 16300 4400 17250 4415
rect 16300 4385 16350 4400
rect 16300 4365 16315 4385
rect 16335 4365 16350 4385
rect 16300 4335 16350 4365
rect 16600 4385 16650 4400
rect 16600 4365 16615 4385
rect 16635 4365 16650 4385
rect 16300 4315 16315 4335
rect 16335 4315 16350 4335
rect 16300 4285 16350 4315
rect 16300 4265 16315 4285
rect 16335 4265 16350 4285
rect 16300 4235 16350 4265
rect 16300 4215 16315 4235
rect 16335 4215 16350 4235
rect 16300 4185 16350 4215
rect 16300 4165 16315 4185
rect 16335 4165 16350 4185
rect 16300 4135 16350 4165
rect 16300 4115 16315 4135
rect 16335 4115 16350 4135
rect 16300 4085 16350 4115
rect 16300 4065 16315 4085
rect 16335 4065 16350 4085
rect 16300 4050 16350 4065
rect 16450 4335 16500 4350
rect 16450 4315 16465 4335
rect 16485 4315 16500 4335
rect 16450 4285 16500 4315
rect 16450 4265 16465 4285
rect 16485 4265 16500 4285
rect 16450 4235 16500 4265
rect 16450 4215 16465 4235
rect 16485 4215 16500 4235
rect 16450 4185 16500 4215
rect 16450 4165 16465 4185
rect 16485 4165 16500 4185
rect 16450 4135 16500 4165
rect 16450 4115 16465 4135
rect 16485 4115 16500 4135
rect 16450 4085 16500 4115
rect 16450 4065 16465 4085
rect 16485 4065 16500 4085
rect 16150 4015 16165 4035
rect 16185 4015 16200 4035
rect 16150 4000 16200 4015
rect 16450 4035 16500 4065
rect 16600 4335 16650 4365
rect 16900 4385 16950 4400
rect 16900 4365 16915 4385
rect 16935 4365 16950 4385
rect 16600 4315 16615 4335
rect 16635 4315 16650 4335
rect 16600 4285 16650 4315
rect 16600 4265 16615 4285
rect 16635 4265 16650 4285
rect 16600 4235 16650 4265
rect 16600 4215 16615 4235
rect 16635 4215 16650 4235
rect 16600 4185 16650 4215
rect 16600 4165 16615 4185
rect 16635 4165 16650 4185
rect 16600 4135 16650 4165
rect 16600 4115 16615 4135
rect 16635 4115 16650 4135
rect 16600 4085 16650 4115
rect 16600 4065 16615 4085
rect 16635 4065 16650 4085
rect 16600 4050 16650 4065
rect 16750 4335 16800 4350
rect 16750 4315 16765 4335
rect 16785 4315 16800 4335
rect 16750 4285 16800 4315
rect 16750 4265 16765 4285
rect 16785 4265 16800 4285
rect 16750 4235 16800 4265
rect 16750 4215 16765 4235
rect 16785 4215 16800 4235
rect 16750 4185 16800 4215
rect 16750 4165 16765 4185
rect 16785 4165 16800 4185
rect 16750 4135 16800 4165
rect 16750 4115 16765 4135
rect 16785 4115 16800 4135
rect 16750 4085 16800 4115
rect 16750 4065 16765 4085
rect 16785 4065 16800 4085
rect 16450 4015 16465 4035
rect 16485 4015 16500 4035
rect 16450 4000 16500 4015
rect 16750 4035 16800 4065
rect 16900 4335 16950 4365
rect 17200 4385 17250 4400
rect 17200 4365 17215 4385
rect 17235 4365 17250 4385
rect 16900 4315 16915 4335
rect 16935 4315 16950 4335
rect 16900 4285 16950 4315
rect 16900 4265 16915 4285
rect 16935 4265 16950 4285
rect 16900 4235 16950 4265
rect 16900 4215 16915 4235
rect 16935 4215 16950 4235
rect 16900 4185 16950 4215
rect 16900 4165 16915 4185
rect 16935 4165 16950 4185
rect 16900 4135 16950 4165
rect 16900 4115 16915 4135
rect 16935 4115 16950 4135
rect 16900 4085 16950 4115
rect 16900 4065 16915 4085
rect 16935 4065 16950 4085
rect 16900 4050 16950 4065
rect 17050 4335 17100 4350
rect 17050 4315 17065 4335
rect 17085 4315 17100 4335
rect 17050 4285 17100 4315
rect 17050 4265 17065 4285
rect 17085 4265 17100 4285
rect 17050 4235 17100 4265
rect 17050 4215 17065 4235
rect 17085 4215 17100 4235
rect 17050 4185 17100 4215
rect 17050 4165 17065 4185
rect 17085 4165 17100 4185
rect 17050 4135 17100 4165
rect 17050 4115 17065 4135
rect 17085 4115 17100 4135
rect 17050 4085 17100 4115
rect 17050 4065 17065 4085
rect 17085 4065 17100 4085
rect 16750 4015 16765 4035
rect 16785 4015 16800 4035
rect 16750 4000 16800 4015
rect 17050 4035 17100 4065
rect 17200 4335 17250 4365
rect 17200 4315 17215 4335
rect 17235 4315 17250 4335
rect 17200 4285 17250 4315
rect 17200 4265 17215 4285
rect 17235 4265 17250 4285
rect 17200 4235 17250 4265
rect 17200 4215 17215 4235
rect 17235 4215 17250 4235
rect 17200 4185 17250 4215
rect 17200 4165 17215 4185
rect 17235 4165 17250 4185
rect 17200 4135 17250 4165
rect 17200 4115 17215 4135
rect 17235 4115 17250 4135
rect 17200 4085 17250 4115
rect 17200 4065 17215 4085
rect 17235 4065 17250 4085
rect 17200 4050 17250 4065
rect 17350 4435 17400 4615
rect 17950 4985 18000 5000
rect 17950 4965 17965 4985
rect 17985 4965 18000 4985
rect 17950 4940 18000 4965
rect 17950 4910 17960 4940
rect 17990 4910 18000 4940
rect 17950 4885 18000 4910
rect 17950 4865 17965 4885
rect 17985 4865 18000 4885
rect 17950 4840 18000 4865
rect 17950 4810 17960 4840
rect 17990 4810 18000 4840
rect 17950 4785 18000 4810
rect 17950 4765 17965 4785
rect 17985 4765 18000 4785
rect 17950 4740 18000 4765
rect 17950 4710 17960 4740
rect 17990 4710 18000 4740
rect 17950 4685 18000 4710
rect 17950 4665 17965 4685
rect 17985 4665 18000 4685
rect 17950 4640 18000 4665
rect 17950 4610 17960 4640
rect 17990 4610 18000 4640
rect 17500 4540 17550 4550
rect 17500 4510 17510 4540
rect 17540 4510 17550 4540
rect 17500 4500 17550 4510
rect 17800 4540 17850 4550
rect 17800 4510 17810 4540
rect 17840 4510 17850 4540
rect 17800 4500 17850 4510
rect 17350 4415 17365 4435
rect 17385 4415 17400 4435
rect 17350 4385 17400 4415
rect 17350 4365 17365 4385
rect 17385 4365 17400 4385
rect 17350 4335 17400 4365
rect 17350 4315 17365 4335
rect 17385 4315 17400 4335
rect 17350 4285 17400 4315
rect 17350 4265 17365 4285
rect 17385 4265 17400 4285
rect 17350 4235 17400 4265
rect 17350 4215 17365 4235
rect 17385 4215 17400 4235
rect 17350 4185 17400 4215
rect 17350 4165 17365 4185
rect 17385 4165 17400 4185
rect 17350 4135 17400 4165
rect 17350 4115 17365 4135
rect 17385 4115 17400 4135
rect 17350 4085 17400 4115
rect 17350 4065 17365 4085
rect 17385 4065 17400 4085
rect 17050 4015 17065 4035
rect 17085 4015 17100 4035
rect 17050 4000 17100 4015
rect 17350 4035 17400 4065
rect 17950 4440 18000 4610
rect 18550 4985 18600 5015
rect 18850 5035 18900 5050
rect 18850 5015 18865 5035
rect 18885 5015 18900 5035
rect 18550 4965 18565 4985
rect 18585 4965 18600 4985
rect 18550 4935 18600 4965
rect 18550 4915 18565 4935
rect 18585 4915 18600 4935
rect 18550 4885 18600 4915
rect 18550 4865 18565 4885
rect 18585 4865 18600 4885
rect 18550 4835 18600 4865
rect 18550 4815 18565 4835
rect 18585 4815 18600 4835
rect 18550 4785 18600 4815
rect 18550 4765 18565 4785
rect 18585 4765 18600 4785
rect 18550 4735 18600 4765
rect 18550 4715 18565 4735
rect 18585 4715 18600 4735
rect 18550 4685 18600 4715
rect 18550 4665 18565 4685
rect 18585 4665 18600 4685
rect 18550 4635 18600 4665
rect 18550 4615 18565 4635
rect 18585 4615 18600 4635
rect 18100 4540 18150 4550
rect 18100 4510 18110 4540
rect 18140 4510 18150 4540
rect 18100 4500 18150 4510
rect 18400 4540 18450 4550
rect 18400 4510 18410 4540
rect 18440 4510 18450 4540
rect 18400 4500 18450 4510
rect 17950 4410 17960 4440
rect 17990 4410 18000 4440
rect 17950 4385 18000 4410
rect 17950 4365 17965 4385
rect 17985 4365 18000 4385
rect 17950 4340 18000 4365
rect 17950 4310 17960 4340
rect 17990 4310 18000 4340
rect 17950 4285 18000 4310
rect 17950 4265 17965 4285
rect 17985 4265 18000 4285
rect 17950 4240 18000 4265
rect 17950 4210 17960 4240
rect 17990 4210 18000 4240
rect 17950 4185 18000 4210
rect 17950 4165 17965 4185
rect 17985 4165 18000 4185
rect 17950 4140 18000 4165
rect 17950 4110 17960 4140
rect 17990 4110 18000 4140
rect 17950 4085 18000 4110
rect 17950 4065 17965 4085
rect 17985 4065 18000 4085
rect 17950 4050 18000 4065
rect 18550 4435 18600 4615
rect 18700 4985 18750 5000
rect 18700 4965 18715 4985
rect 18735 4965 18750 4985
rect 18700 4935 18750 4965
rect 18700 4915 18715 4935
rect 18735 4915 18750 4935
rect 18700 4885 18750 4915
rect 18700 4865 18715 4885
rect 18735 4865 18750 4885
rect 18700 4835 18750 4865
rect 18700 4815 18715 4835
rect 18735 4815 18750 4835
rect 18700 4785 18750 4815
rect 18700 4765 18715 4785
rect 18735 4765 18750 4785
rect 18700 4735 18750 4765
rect 18700 4715 18715 4735
rect 18735 4715 18750 4735
rect 18700 4685 18750 4715
rect 18850 4985 18900 5015
rect 19150 5035 19200 5050
rect 19150 5015 19165 5035
rect 19185 5015 19200 5035
rect 18850 4965 18865 4985
rect 18885 4965 18900 4985
rect 18850 4935 18900 4965
rect 18850 4915 18865 4935
rect 18885 4915 18900 4935
rect 18850 4885 18900 4915
rect 18850 4865 18865 4885
rect 18885 4865 18900 4885
rect 18850 4835 18900 4865
rect 18850 4815 18865 4835
rect 18885 4815 18900 4835
rect 18850 4785 18900 4815
rect 18850 4765 18865 4785
rect 18885 4765 18900 4785
rect 18850 4735 18900 4765
rect 18850 4715 18865 4735
rect 18885 4715 18900 4735
rect 18850 4700 18900 4715
rect 19000 4985 19050 5000
rect 19000 4965 19015 4985
rect 19035 4965 19050 4985
rect 19000 4935 19050 4965
rect 19000 4915 19015 4935
rect 19035 4915 19050 4935
rect 19000 4885 19050 4915
rect 19000 4865 19015 4885
rect 19035 4865 19050 4885
rect 19000 4835 19050 4865
rect 19000 4815 19015 4835
rect 19035 4815 19050 4835
rect 19000 4785 19050 4815
rect 19000 4765 19015 4785
rect 19035 4765 19050 4785
rect 19000 4735 19050 4765
rect 19000 4715 19015 4735
rect 19035 4715 19050 4735
rect 18700 4665 18715 4685
rect 18735 4665 18750 4685
rect 18700 4650 18750 4665
rect 19000 4685 19050 4715
rect 19150 4985 19200 5015
rect 19450 5035 19500 5050
rect 19450 5015 19465 5035
rect 19485 5015 19500 5035
rect 19150 4965 19165 4985
rect 19185 4965 19200 4985
rect 19150 4935 19200 4965
rect 19150 4915 19165 4935
rect 19185 4915 19200 4935
rect 19150 4885 19200 4915
rect 19150 4865 19165 4885
rect 19185 4865 19200 4885
rect 19150 4835 19200 4865
rect 19150 4815 19165 4835
rect 19185 4815 19200 4835
rect 19150 4785 19200 4815
rect 19150 4765 19165 4785
rect 19185 4765 19200 4785
rect 19150 4735 19200 4765
rect 19150 4715 19165 4735
rect 19185 4715 19200 4735
rect 19150 4700 19200 4715
rect 19300 4985 19350 5000
rect 19300 4965 19315 4985
rect 19335 4965 19350 4985
rect 19300 4935 19350 4965
rect 19300 4915 19315 4935
rect 19335 4915 19350 4935
rect 19300 4885 19350 4915
rect 19300 4865 19315 4885
rect 19335 4865 19350 4885
rect 19300 4835 19350 4865
rect 19300 4815 19315 4835
rect 19335 4815 19350 4835
rect 19300 4785 19350 4815
rect 19300 4765 19315 4785
rect 19335 4765 19350 4785
rect 19300 4735 19350 4765
rect 19300 4715 19315 4735
rect 19335 4715 19350 4735
rect 19000 4665 19015 4685
rect 19035 4665 19050 4685
rect 19000 4650 19050 4665
rect 19300 4685 19350 4715
rect 19450 4985 19500 5015
rect 19750 5035 19800 5050
rect 19750 5015 19765 5035
rect 19785 5015 19800 5035
rect 19450 4965 19465 4985
rect 19485 4965 19500 4985
rect 19450 4935 19500 4965
rect 19450 4915 19465 4935
rect 19485 4915 19500 4935
rect 19450 4885 19500 4915
rect 19450 4865 19465 4885
rect 19485 4865 19500 4885
rect 19450 4835 19500 4865
rect 19450 4815 19465 4835
rect 19485 4815 19500 4835
rect 19450 4785 19500 4815
rect 19450 4765 19465 4785
rect 19485 4765 19500 4785
rect 19450 4735 19500 4765
rect 19450 4715 19465 4735
rect 19485 4715 19500 4735
rect 19450 4700 19500 4715
rect 19600 4985 19650 5000
rect 19600 4965 19615 4985
rect 19635 4965 19650 4985
rect 19600 4935 19650 4965
rect 19600 4915 19615 4935
rect 19635 4915 19650 4935
rect 19600 4885 19650 4915
rect 19600 4865 19615 4885
rect 19635 4865 19650 4885
rect 19600 4835 19650 4865
rect 19600 4815 19615 4835
rect 19635 4815 19650 4835
rect 19600 4785 19650 4815
rect 19600 4765 19615 4785
rect 19635 4765 19650 4785
rect 19600 4735 19650 4765
rect 19600 4715 19615 4735
rect 19635 4715 19650 4735
rect 19300 4665 19315 4685
rect 19335 4665 19350 4685
rect 19300 4650 19350 4665
rect 19600 4685 19650 4715
rect 19600 4665 19615 4685
rect 19635 4665 19650 4685
rect 19600 4650 19650 4665
rect 18700 4635 19650 4650
rect 18700 4615 18715 4635
rect 18735 4615 19015 4635
rect 19035 4615 19315 4635
rect 19335 4615 19615 4635
rect 19635 4615 19650 4635
rect 18700 4600 19650 4615
rect 19750 4985 19800 5015
rect 19750 4965 19765 4985
rect 19785 4965 19800 4985
rect 19750 4935 19800 4965
rect 19750 4915 19765 4935
rect 19785 4915 19800 4935
rect 19750 4885 19800 4915
rect 19750 4865 19765 4885
rect 19785 4865 19800 4885
rect 19750 4835 19800 4865
rect 19750 4815 19765 4835
rect 19785 4815 19800 4835
rect 19750 4785 19800 4815
rect 19750 4765 19765 4785
rect 19785 4765 19800 4785
rect 19750 4735 19800 4765
rect 19750 4715 19765 4735
rect 19785 4715 19800 4735
rect 19750 4685 19800 4715
rect 19750 4665 19765 4685
rect 19785 4665 19800 4685
rect 19750 4635 19800 4665
rect 19750 4615 19765 4635
rect 19785 4615 19800 4635
rect 18700 4540 18750 4550
rect 18700 4510 18710 4540
rect 18740 4510 18750 4540
rect 18700 4500 18750 4510
rect 19000 4540 19050 4550
rect 19000 4510 19010 4540
rect 19040 4510 19050 4540
rect 19000 4500 19050 4510
rect 19150 4540 19200 4600
rect 19150 4510 19160 4540
rect 19190 4510 19200 4540
rect 19150 4450 19200 4510
rect 19300 4540 19350 4550
rect 19300 4510 19310 4540
rect 19340 4510 19350 4540
rect 19300 4500 19350 4510
rect 19600 4540 19650 4550
rect 19600 4510 19610 4540
rect 19640 4510 19650 4540
rect 19600 4500 19650 4510
rect 18550 4415 18565 4435
rect 18585 4415 18600 4435
rect 18550 4385 18600 4415
rect 18550 4365 18565 4385
rect 18585 4365 18600 4385
rect 18550 4335 18600 4365
rect 18550 4315 18565 4335
rect 18585 4315 18600 4335
rect 18550 4285 18600 4315
rect 18550 4265 18565 4285
rect 18585 4265 18600 4285
rect 18550 4235 18600 4265
rect 18550 4215 18565 4235
rect 18585 4215 18600 4235
rect 18550 4185 18600 4215
rect 18550 4165 18565 4185
rect 18585 4165 18600 4185
rect 18550 4135 18600 4165
rect 18550 4115 18565 4135
rect 18585 4115 18600 4135
rect 18550 4085 18600 4115
rect 18550 4065 18565 4085
rect 18585 4065 18600 4085
rect 17350 4015 17365 4035
rect 17385 4015 17400 4035
rect 17350 4000 17400 4015
rect 18550 4035 18600 4065
rect 18700 4435 19650 4450
rect 18700 4415 18715 4435
rect 18735 4415 19015 4435
rect 19035 4415 19315 4435
rect 19335 4415 19615 4435
rect 19635 4415 19650 4435
rect 18700 4400 19650 4415
rect 18700 4385 18750 4400
rect 18700 4365 18715 4385
rect 18735 4365 18750 4385
rect 18700 4335 18750 4365
rect 19000 4385 19050 4400
rect 19000 4365 19015 4385
rect 19035 4365 19050 4385
rect 18700 4315 18715 4335
rect 18735 4315 18750 4335
rect 18700 4285 18750 4315
rect 18700 4265 18715 4285
rect 18735 4265 18750 4285
rect 18700 4235 18750 4265
rect 18700 4215 18715 4235
rect 18735 4215 18750 4235
rect 18700 4185 18750 4215
rect 18700 4165 18715 4185
rect 18735 4165 18750 4185
rect 18700 4135 18750 4165
rect 18700 4115 18715 4135
rect 18735 4115 18750 4135
rect 18700 4085 18750 4115
rect 18700 4065 18715 4085
rect 18735 4065 18750 4085
rect 18700 4050 18750 4065
rect 18850 4335 18900 4350
rect 18850 4315 18865 4335
rect 18885 4315 18900 4335
rect 18850 4285 18900 4315
rect 18850 4265 18865 4285
rect 18885 4265 18900 4285
rect 18850 4235 18900 4265
rect 18850 4215 18865 4235
rect 18885 4215 18900 4235
rect 18850 4185 18900 4215
rect 18850 4165 18865 4185
rect 18885 4165 18900 4185
rect 18850 4135 18900 4165
rect 18850 4115 18865 4135
rect 18885 4115 18900 4135
rect 18850 4085 18900 4115
rect 18850 4065 18865 4085
rect 18885 4065 18900 4085
rect 18550 4015 18565 4035
rect 18585 4015 18600 4035
rect 18550 4000 18600 4015
rect 18850 4035 18900 4065
rect 19000 4335 19050 4365
rect 19300 4385 19350 4400
rect 19300 4365 19315 4385
rect 19335 4365 19350 4385
rect 19000 4315 19015 4335
rect 19035 4315 19050 4335
rect 19000 4285 19050 4315
rect 19000 4265 19015 4285
rect 19035 4265 19050 4285
rect 19000 4235 19050 4265
rect 19000 4215 19015 4235
rect 19035 4215 19050 4235
rect 19000 4185 19050 4215
rect 19000 4165 19015 4185
rect 19035 4165 19050 4185
rect 19000 4135 19050 4165
rect 19000 4115 19015 4135
rect 19035 4115 19050 4135
rect 19000 4085 19050 4115
rect 19000 4065 19015 4085
rect 19035 4065 19050 4085
rect 19000 4050 19050 4065
rect 19150 4335 19200 4350
rect 19150 4315 19165 4335
rect 19185 4315 19200 4335
rect 19150 4285 19200 4315
rect 19150 4265 19165 4285
rect 19185 4265 19200 4285
rect 19150 4235 19200 4265
rect 19150 4215 19165 4235
rect 19185 4215 19200 4235
rect 19150 4185 19200 4215
rect 19150 4165 19165 4185
rect 19185 4165 19200 4185
rect 19150 4135 19200 4165
rect 19150 4115 19165 4135
rect 19185 4115 19200 4135
rect 19150 4085 19200 4115
rect 19150 4065 19165 4085
rect 19185 4065 19200 4085
rect 18850 4015 18865 4035
rect 18885 4015 18900 4035
rect 18850 4000 18900 4015
rect 19150 4035 19200 4065
rect 19300 4335 19350 4365
rect 19600 4385 19650 4400
rect 19600 4365 19615 4385
rect 19635 4365 19650 4385
rect 19300 4315 19315 4335
rect 19335 4315 19350 4335
rect 19300 4285 19350 4315
rect 19300 4265 19315 4285
rect 19335 4265 19350 4285
rect 19300 4235 19350 4265
rect 19300 4215 19315 4235
rect 19335 4215 19350 4235
rect 19300 4185 19350 4215
rect 19300 4165 19315 4185
rect 19335 4165 19350 4185
rect 19300 4135 19350 4165
rect 19300 4115 19315 4135
rect 19335 4115 19350 4135
rect 19300 4085 19350 4115
rect 19300 4065 19315 4085
rect 19335 4065 19350 4085
rect 19300 4050 19350 4065
rect 19450 4335 19500 4350
rect 19450 4315 19465 4335
rect 19485 4315 19500 4335
rect 19450 4285 19500 4315
rect 19450 4265 19465 4285
rect 19485 4265 19500 4285
rect 19450 4235 19500 4265
rect 19450 4215 19465 4235
rect 19485 4215 19500 4235
rect 19450 4185 19500 4215
rect 19450 4165 19465 4185
rect 19485 4165 19500 4185
rect 19450 4135 19500 4165
rect 19450 4115 19465 4135
rect 19485 4115 19500 4135
rect 19450 4085 19500 4115
rect 19450 4065 19465 4085
rect 19485 4065 19500 4085
rect 19150 4015 19165 4035
rect 19185 4015 19200 4035
rect 19150 4000 19200 4015
rect 19450 4035 19500 4065
rect 19600 4335 19650 4365
rect 19600 4315 19615 4335
rect 19635 4315 19650 4335
rect 19600 4285 19650 4315
rect 19600 4265 19615 4285
rect 19635 4265 19650 4285
rect 19600 4235 19650 4265
rect 19600 4215 19615 4235
rect 19635 4215 19650 4235
rect 19600 4185 19650 4215
rect 19600 4165 19615 4185
rect 19635 4165 19650 4185
rect 19600 4135 19650 4165
rect 19600 4115 19615 4135
rect 19635 4115 19650 4135
rect 19600 4085 19650 4115
rect 19600 4065 19615 4085
rect 19635 4065 19650 4085
rect 19600 4050 19650 4065
rect 19750 4435 19800 4615
rect 20350 5085 20400 5160
rect 20350 5065 20365 5085
rect 20385 5065 20400 5085
rect 20350 5040 20400 5065
rect 20350 5010 20360 5040
rect 20390 5010 20400 5040
rect 20350 4985 20400 5010
rect 20350 4965 20365 4985
rect 20385 4965 20400 4985
rect 20350 4940 20400 4965
rect 20350 4910 20360 4940
rect 20390 4910 20400 4940
rect 20350 4885 20400 4910
rect 20350 4865 20365 4885
rect 20385 4865 20400 4885
rect 20350 4840 20400 4865
rect 20350 4810 20360 4840
rect 20390 4810 20400 4840
rect 20350 4785 20400 4810
rect 20350 4765 20365 4785
rect 20385 4765 20400 4785
rect 20350 4740 20400 4765
rect 20350 4710 20360 4740
rect 20390 4710 20400 4740
rect 20350 4685 20400 4710
rect 20350 4665 20365 4685
rect 20385 4665 20400 4685
rect 20350 4640 20400 4665
rect 20350 4610 20360 4640
rect 20390 4610 20400 4640
rect 19900 4540 19950 4550
rect 19900 4510 19910 4540
rect 19940 4510 19950 4540
rect 19900 4500 19950 4510
rect 20200 4540 20250 4550
rect 20200 4510 20210 4540
rect 20240 4510 20250 4540
rect 20200 4500 20250 4510
rect 19750 4415 19765 4435
rect 19785 4415 19800 4435
rect 19750 4385 19800 4415
rect 19750 4365 19765 4385
rect 19785 4365 19800 4385
rect 19750 4335 19800 4365
rect 19750 4315 19765 4335
rect 19785 4315 19800 4335
rect 19750 4285 19800 4315
rect 19750 4265 19765 4285
rect 19785 4265 19800 4285
rect 19750 4235 19800 4265
rect 19750 4215 19765 4235
rect 19785 4215 19800 4235
rect 19750 4185 19800 4215
rect 19750 4165 19765 4185
rect 19785 4165 19800 4185
rect 19750 4135 19800 4165
rect 19750 4115 19765 4135
rect 19785 4115 19800 4135
rect 19750 4085 19800 4115
rect 19750 4065 19765 4085
rect 19785 4065 19800 4085
rect 19450 4015 19465 4035
rect 19485 4015 19500 4035
rect 19450 4000 19500 4015
rect 19750 4035 19800 4065
rect 19750 4015 19765 4035
rect 19785 4015 19800 4035
rect 19750 4000 19800 4015
rect 16150 3985 19800 4000
rect 16150 3965 16165 3985
rect 16185 3965 16465 3985
rect 16485 3965 16765 3985
rect 16785 3965 17065 3985
rect 17085 3965 17365 3985
rect 17385 3965 18565 3985
rect 18585 3965 18865 3985
rect 18885 3965 19165 3985
rect 19185 3965 19465 3985
rect 19485 3965 19765 3985
rect 19785 3965 19800 3985
rect 16150 3950 19800 3965
rect 20350 4440 20400 4610
rect 20350 4410 20360 4440
rect 20390 4410 20400 4440
rect 20350 4385 20400 4410
rect 20350 4365 20365 4385
rect 20385 4365 20400 4385
rect 20350 4340 20400 4365
rect 20350 4310 20360 4340
rect 20390 4310 20400 4340
rect 20350 4285 20400 4310
rect 20350 4265 20365 4285
rect 20385 4265 20400 4285
rect 20350 4240 20400 4265
rect 20350 4210 20360 4240
rect 20390 4210 20400 4240
rect 20350 4185 20400 4210
rect 20350 4165 20365 4185
rect 20385 4165 20400 4185
rect 20350 4140 20400 4165
rect 20350 4110 20360 4140
rect 20390 4110 20400 4140
rect 20350 4085 20400 4110
rect 20350 4065 20365 4085
rect 20385 4065 20400 4085
rect 20350 4040 20400 4065
rect 20350 4010 20360 4040
rect 20390 4010 20400 4040
rect 20350 3985 20400 4010
rect 20350 3965 20365 3985
rect 20385 3965 20400 3985
rect 15550 3860 15560 3890
rect 15590 3860 15600 3890
rect 15550 3785 15600 3860
rect 17950 3800 18000 3950
rect 20350 3890 20400 3965
rect 20350 3860 20360 3890
rect 20390 3860 20400 3890
rect 15550 3765 15565 3785
rect 15585 3765 15600 3785
rect 15550 3740 15600 3765
rect 15550 3710 15560 3740
rect 15590 3710 15600 3740
rect 15550 3685 15600 3710
rect 15550 3665 15565 3685
rect 15585 3665 15600 3685
rect 15550 3640 15600 3665
rect 15550 3610 15560 3640
rect 15590 3610 15600 3640
rect 15550 3585 15600 3610
rect 15550 3565 15565 3585
rect 15585 3565 15600 3585
rect 15550 3540 15600 3565
rect 15550 3510 15560 3540
rect 15590 3510 15600 3540
rect 15550 3485 15600 3510
rect 15550 3465 15565 3485
rect 15585 3465 15600 3485
rect 15550 3440 15600 3465
rect 15550 3410 15560 3440
rect 15590 3410 15600 3440
rect 15550 3385 15600 3410
rect 15550 3365 15565 3385
rect 15585 3365 15600 3385
rect 15550 3340 15600 3365
rect 15550 3310 15560 3340
rect 15590 3310 15600 3340
rect 14950 3210 14960 3240
rect 14990 3210 15000 3240
rect 14350 3110 14360 3140
rect 14390 3110 14400 3140
rect 14350 3085 14400 3110
rect 14350 3065 14365 3085
rect 14385 3065 14400 3085
rect 14350 3040 14400 3065
rect 14350 3010 14360 3040
rect 14390 3010 14400 3040
rect 14350 2985 14400 3010
rect 14350 2965 14365 2985
rect 14385 2965 14400 2985
rect 14350 2940 14400 2965
rect 14350 2910 14360 2940
rect 14390 2910 14400 2940
rect 14350 2885 14400 2910
rect 14350 2865 14365 2885
rect 14385 2865 14400 2885
rect 14350 2840 14400 2865
rect 14350 2810 14360 2840
rect 14390 2810 14400 2840
rect 14350 2785 14400 2810
rect 14350 2765 14365 2785
rect 14385 2765 14400 2785
rect 14350 2740 14400 2765
rect 14350 2710 14360 2740
rect 14390 2710 14400 2740
rect 14350 2685 14400 2710
rect 14350 2665 14365 2685
rect 14385 2665 14400 2685
rect 13150 2560 13160 2590
rect 13190 2560 13200 2590
rect 13150 2550 13200 2560
rect 14350 2590 14400 2665
rect 14950 3135 15000 3210
rect 15100 3240 15150 3250
rect 15100 3210 15110 3240
rect 15140 3210 15150 3240
rect 15100 3200 15150 3210
rect 15400 3240 15450 3250
rect 15400 3210 15410 3240
rect 15440 3210 15450 3240
rect 15400 3200 15450 3210
rect 14950 3115 14965 3135
rect 14985 3115 15000 3135
rect 14950 3085 15000 3115
rect 14950 3065 14965 3085
rect 14985 3065 15000 3085
rect 14950 3035 15000 3065
rect 14950 3015 14965 3035
rect 14985 3015 15000 3035
rect 14950 2985 15000 3015
rect 14950 2965 14965 2985
rect 14985 2965 15000 2985
rect 14950 2935 15000 2965
rect 14950 2915 14965 2935
rect 14985 2915 15000 2935
rect 14950 2885 15000 2915
rect 14950 2865 14965 2885
rect 14985 2865 15000 2885
rect 14950 2835 15000 2865
rect 14950 2815 14965 2835
rect 14985 2815 15000 2835
rect 14950 2785 15000 2815
rect 14950 2765 14965 2785
rect 14985 2765 15000 2785
rect 14950 2735 15000 2765
rect 14950 2715 14965 2735
rect 14985 2715 15000 2735
rect 14950 2685 15000 2715
rect 14950 2665 14965 2685
rect 14985 2665 15000 2685
rect 14950 2650 15000 2665
rect 15550 3140 15600 3310
rect 16150 3785 19800 3800
rect 16150 3765 16165 3785
rect 16185 3765 16465 3785
rect 16485 3765 16765 3785
rect 16785 3765 17065 3785
rect 17085 3765 17365 3785
rect 17385 3765 18565 3785
rect 18585 3765 18865 3785
rect 18885 3765 19165 3785
rect 19185 3765 19465 3785
rect 19485 3765 19765 3785
rect 19785 3765 19800 3785
rect 16150 3750 19800 3765
rect 16150 3735 16200 3750
rect 16150 3715 16165 3735
rect 16185 3715 16200 3735
rect 16150 3685 16200 3715
rect 16450 3735 16500 3750
rect 16450 3715 16465 3735
rect 16485 3715 16500 3735
rect 16150 3665 16165 3685
rect 16185 3665 16200 3685
rect 16150 3635 16200 3665
rect 16150 3615 16165 3635
rect 16185 3615 16200 3635
rect 16150 3585 16200 3615
rect 16150 3565 16165 3585
rect 16185 3565 16200 3585
rect 16150 3535 16200 3565
rect 16150 3515 16165 3535
rect 16185 3515 16200 3535
rect 16150 3485 16200 3515
rect 16150 3465 16165 3485
rect 16185 3465 16200 3485
rect 16150 3435 16200 3465
rect 16150 3415 16165 3435
rect 16185 3415 16200 3435
rect 16150 3385 16200 3415
rect 16150 3365 16165 3385
rect 16185 3365 16200 3385
rect 16150 3335 16200 3365
rect 16150 3315 16165 3335
rect 16185 3315 16200 3335
rect 15700 3240 15750 3250
rect 15700 3210 15710 3240
rect 15740 3210 15750 3240
rect 15700 3200 15750 3210
rect 16000 3240 16050 3250
rect 16000 3210 16010 3240
rect 16040 3210 16050 3240
rect 16000 3200 16050 3210
rect 15550 3110 15560 3140
rect 15590 3110 15600 3140
rect 15550 3085 15600 3110
rect 15550 3065 15565 3085
rect 15585 3065 15600 3085
rect 15550 3040 15600 3065
rect 15550 3010 15560 3040
rect 15590 3010 15600 3040
rect 15550 2985 15600 3010
rect 15550 2965 15565 2985
rect 15585 2965 15600 2985
rect 15550 2940 15600 2965
rect 15550 2910 15560 2940
rect 15590 2910 15600 2940
rect 15550 2885 15600 2910
rect 15550 2865 15565 2885
rect 15585 2865 15600 2885
rect 15550 2840 15600 2865
rect 15550 2810 15560 2840
rect 15590 2810 15600 2840
rect 15550 2785 15600 2810
rect 15550 2765 15565 2785
rect 15585 2765 15600 2785
rect 15550 2740 15600 2765
rect 15550 2710 15560 2740
rect 15590 2710 15600 2740
rect 15550 2685 15600 2710
rect 15550 2665 15565 2685
rect 15585 2665 15600 2685
rect 14350 2560 14360 2590
rect 14390 2560 14400 2590
rect 14350 2550 14400 2560
rect 15550 2590 15600 2665
rect 16150 3135 16200 3315
rect 16300 3685 16350 3700
rect 16300 3665 16315 3685
rect 16335 3665 16350 3685
rect 16300 3635 16350 3665
rect 16300 3615 16315 3635
rect 16335 3615 16350 3635
rect 16300 3585 16350 3615
rect 16300 3565 16315 3585
rect 16335 3565 16350 3585
rect 16300 3535 16350 3565
rect 16300 3515 16315 3535
rect 16335 3515 16350 3535
rect 16300 3485 16350 3515
rect 16300 3465 16315 3485
rect 16335 3465 16350 3485
rect 16300 3435 16350 3465
rect 16300 3415 16315 3435
rect 16335 3415 16350 3435
rect 16300 3385 16350 3415
rect 16450 3685 16500 3715
rect 16750 3735 16800 3750
rect 16750 3715 16765 3735
rect 16785 3715 16800 3735
rect 16450 3665 16465 3685
rect 16485 3665 16500 3685
rect 16450 3635 16500 3665
rect 16450 3615 16465 3635
rect 16485 3615 16500 3635
rect 16450 3585 16500 3615
rect 16450 3565 16465 3585
rect 16485 3565 16500 3585
rect 16450 3535 16500 3565
rect 16450 3515 16465 3535
rect 16485 3515 16500 3535
rect 16450 3485 16500 3515
rect 16450 3465 16465 3485
rect 16485 3465 16500 3485
rect 16450 3435 16500 3465
rect 16450 3415 16465 3435
rect 16485 3415 16500 3435
rect 16450 3400 16500 3415
rect 16600 3685 16650 3700
rect 16600 3665 16615 3685
rect 16635 3665 16650 3685
rect 16600 3635 16650 3665
rect 16600 3615 16615 3635
rect 16635 3615 16650 3635
rect 16600 3585 16650 3615
rect 16600 3565 16615 3585
rect 16635 3565 16650 3585
rect 16600 3535 16650 3565
rect 16600 3515 16615 3535
rect 16635 3515 16650 3535
rect 16600 3485 16650 3515
rect 16600 3465 16615 3485
rect 16635 3465 16650 3485
rect 16600 3435 16650 3465
rect 16600 3415 16615 3435
rect 16635 3415 16650 3435
rect 16300 3365 16315 3385
rect 16335 3365 16350 3385
rect 16300 3350 16350 3365
rect 16600 3385 16650 3415
rect 16750 3685 16800 3715
rect 17050 3735 17100 3750
rect 17050 3715 17065 3735
rect 17085 3715 17100 3735
rect 16750 3665 16765 3685
rect 16785 3665 16800 3685
rect 16750 3635 16800 3665
rect 16750 3615 16765 3635
rect 16785 3615 16800 3635
rect 16750 3585 16800 3615
rect 16750 3565 16765 3585
rect 16785 3565 16800 3585
rect 16750 3535 16800 3565
rect 16750 3515 16765 3535
rect 16785 3515 16800 3535
rect 16750 3485 16800 3515
rect 16750 3465 16765 3485
rect 16785 3465 16800 3485
rect 16750 3435 16800 3465
rect 16750 3415 16765 3435
rect 16785 3415 16800 3435
rect 16750 3400 16800 3415
rect 16900 3685 16950 3700
rect 16900 3665 16915 3685
rect 16935 3665 16950 3685
rect 16900 3635 16950 3665
rect 16900 3615 16915 3635
rect 16935 3615 16950 3635
rect 16900 3585 16950 3615
rect 16900 3565 16915 3585
rect 16935 3565 16950 3585
rect 16900 3535 16950 3565
rect 16900 3515 16915 3535
rect 16935 3515 16950 3535
rect 16900 3485 16950 3515
rect 16900 3465 16915 3485
rect 16935 3465 16950 3485
rect 16900 3435 16950 3465
rect 16900 3415 16915 3435
rect 16935 3415 16950 3435
rect 16600 3365 16615 3385
rect 16635 3365 16650 3385
rect 16600 3350 16650 3365
rect 16900 3385 16950 3415
rect 17050 3685 17100 3715
rect 17350 3735 17400 3750
rect 17350 3715 17365 3735
rect 17385 3715 17400 3735
rect 17050 3665 17065 3685
rect 17085 3665 17100 3685
rect 17050 3635 17100 3665
rect 17050 3615 17065 3635
rect 17085 3615 17100 3635
rect 17050 3585 17100 3615
rect 17050 3565 17065 3585
rect 17085 3565 17100 3585
rect 17050 3535 17100 3565
rect 17050 3515 17065 3535
rect 17085 3515 17100 3535
rect 17050 3485 17100 3515
rect 17050 3465 17065 3485
rect 17085 3465 17100 3485
rect 17050 3435 17100 3465
rect 17050 3415 17065 3435
rect 17085 3415 17100 3435
rect 17050 3400 17100 3415
rect 17200 3685 17250 3700
rect 17200 3665 17215 3685
rect 17235 3665 17250 3685
rect 17200 3635 17250 3665
rect 17200 3615 17215 3635
rect 17235 3615 17250 3635
rect 17200 3585 17250 3615
rect 17200 3565 17215 3585
rect 17235 3565 17250 3585
rect 17200 3535 17250 3565
rect 17200 3515 17215 3535
rect 17235 3515 17250 3535
rect 17200 3485 17250 3515
rect 17200 3465 17215 3485
rect 17235 3465 17250 3485
rect 17200 3435 17250 3465
rect 17200 3415 17215 3435
rect 17235 3415 17250 3435
rect 16900 3365 16915 3385
rect 16935 3365 16950 3385
rect 16900 3350 16950 3365
rect 17200 3385 17250 3415
rect 17200 3365 17215 3385
rect 17235 3365 17250 3385
rect 17200 3350 17250 3365
rect 16300 3335 17250 3350
rect 16300 3315 16315 3335
rect 16335 3315 16615 3335
rect 16635 3315 16915 3335
rect 16935 3315 17215 3335
rect 17235 3315 17250 3335
rect 16300 3300 17250 3315
rect 17350 3685 17400 3715
rect 18550 3735 18600 3750
rect 18550 3715 18565 3735
rect 18585 3715 18600 3735
rect 17350 3665 17365 3685
rect 17385 3665 17400 3685
rect 17350 3635 17400 3665
rect 17350 3615 17365 3635
rect 17385 3615 17400 3635
rect 17350 3585 17400 3615
rect 17350 3565 17365 3585
rect 17385 3565 17400 3585
rect 17350 3535 17400 3565
rect 17350 3515 17365 3535
rect 17385 3515 17400 3535
rect 17350 3485 17400 3515
rect 17350 3465 17365 3485
rect 17385 3465 17400 3485
rect 17350 3435 17400 3465
rect 17350 3415 17365 3435
rect 17385 3415 17400 3435
rect 17350 3385 17400 3415
rect 17350 3365 17365 3385
rect 17385 3365 17400 3385
rect 17350 3335 17400 3365
rect 17350 3315 17365 3335
rect 17385 3315 17400 3335
rect 16300 3240 16350 3250
rect 16300 3210 16310 3240
rect 16340 3210 16350 3240
rect 16300 3200 16350 3210
rect 16600 3240 16650 3250
rect 16600 3210 16610 3240
rect 16640 3210 16650 3240
rect 16600 3200 16650 3210
rect 16750 3240 16800 3300
rect 16750 3210 16760 3240
rect 16790 3210 16800 3240
rect 16750 3150 16800 3210
rect 16900 3240 16950 3250
rect 16900 3210 16910 3240
rect 16940 3210 16950 3240
rect 16900 3200 16950 3210
rect 17200 3240 17250 3250
rect 17200 3210 17210 3240
rect 17240 3210 17250 3240
rect 17200 3200 17250 3210
rect 16150 3115 16165 3135
rect 16185 3115 16200 3135
rect 16150 3085 16200 3115
rect 16150 3065 16165 3085
rect 16185 3065 16200 3085
rect 16150 3035 16200 3065
rect 16150 3015 16165 3035
rect 16185 3015 16200 3035
rect 16150 2985 16200 3015
rect 16150 2965 16165 2985
rect 16185 2965 16200 2985
rect 16150 2935 16200 2965
rect 16150 2915 16165 2935
rect 16185 2915 16200 2935
rect 16150 2885 16200 2915
rect 16150 2865 16165 2885
rect 16185 2865 16200 2885
rect 16150 2835 16200 2865
rect 16150 2815 16165 2835
rect 16185 2815 16200 2835
rect 16150 2785 16200 2815
rect 16150 2765 16165 2785
rect 16185 2765 16200 2785
rect 16150 2735 16200 2765
rect 16300 3135 17250 3150
rect 16300 3115 16315 3135
rect 16335 3115 16615 3135
rect 16635 3115 16915 3135
rect 16935 3115 17215 3135
rect 17235 3115 17250 3135
rect 16300 3100 17250 3115
rect 16300 3085 16350 3100
rect 16300 3065 16315 3085
rect 16335 3065 16350 3085
rect 16300 3035 16350 3065
rect 16600 3085 16650 3100
rect 16600 3065 16615 3085
rect 16635 3065 16650 3085
rect 16300 3015 16315 3035
rect 16335 3015 16350 3035
rect 16300 2985 16350 3015
rect 16300 2965 16315 2985
rect 16335 2965 16350 2985
rect 16300 2935 16350 2965
rect 16300 2915 16315 2935
rect 16335 2915 16350 2935
rect 16300 2885 16350 2915
rect 16300 2865 16315 2885
rect 16335 2865 16350 2885
rect 16300 2835 16350 2865
rect 16300 2815 16315 2835
rect 16335 2815 16350 2835
rect 16300 2785 16350 2815
rect 16300 2765 16315 2785
rect 16335 2765 16350 2785
rect 16300 2750 16350 2765
rect 16450 3035 16500 3050
rect 16450 3015 16465 3035
rect 16485 3015 16500 3035
rect 16450 2985 16500 3015
rect 16450 2965 16465 2985
rect 16485 2965 16500 2985
rect 16450 2935 16500 2965
rect 16450 2915 16465 2935
rect 16485 2915 16500 2935
rect 16450 2885 16500 2915
rect 16450 2865 16465 2885
rect 16485 2865 16500 2885
rect 16450 2835 16500 2865
rect 16450 2815 16465 2835
rect 16485 2815 16500 2835
rect 16450 2785 16500 2815
rect 16450 2765 16465 2785
rect 16485 2765 16500 2785
rect 16150 2715 16165 2735
rect 16185 2715 16200 2735
rect 16150 2700 16200 2715
rect 16450 2735 16500 2765
rect 16600 3035 16650 3065
rect 16900 3085 16950 3100
rect 16900 3065 16915 3085
rect 16935 3065 16950 3085
rect 16600 3015 16615 3035
rect 16635 3015 16650 3035
rect 16600 2985 16650 3015
rect 16600 2965 16615 2985
rect 16635 2965 16650 2985
rect 16600 2935 16650 2965
rect 16600 2915 16615 2935
rect 16635 2915 16650 2935
rect 16600 2885 16650 2915
rect 16600 2865 16615 2885
rect 16635 2865 16650 2885
rect 16600 2835 16650 2865
rect 16600 2815 16615 2835
rect 16635 2815 16650 2835
rect 16600 2785 16650 2815
rect 16600 2765 16615 2785
rect 16635 2765 16650 2785
rect 16600 2750 16650 2765
rect 16750 3035 16800 3050
rect 16750 3015 16765 3035
rect 16785 3015 16800 3035
rect 16750 2985 16800 3015
rect 16750 2965 16765 2985
rect 16785 2965 16800 2985
rect 16750 2935 16800 2965
rect 16750 2915 16765 2935
rect 16785 2915 16800 2935
rect 16750 2885 16800 2915
rect 16750 2865 16765 2885
rect 16785 2865 16800 2885
rect 16750 2835 16800 2865
rect 16750 2815 16765 2835
rect 16785 2815 16800 2835
rect 16750 2785 16800 2815
rect 16750 2765 16765 2785
rect 16785 2765 16800 2785
rect 16450 2715 16465 2735
rect 16485 2715 16500 2735
rect 16450 2700 16500 2715
rect 16750 2735 16800 2765
rect 16900 3035 16950 3065
rect 17200 3085 17250 3100
rect 17200 3065 17215 3085
rect 17235 3065 17250 3085
rect 16900 3015 16915 3035
rect 16935 3015 16950 3035
rect 16900 2985 16950 3015
rect 16900 2965 16915 2985
rect 16935 2965 16950 2985
rect 16900 2935 16950 2965
rect 16900 2915 16915 2935
rect 16935 2915 16950 2935
rect 16900 2885 16950 2915
rect 16900 2865 16915 2885
rect 16935 2865 16950 2885
rect 16900 2835 16950 2865
rect 16900 2815 16915 2835
rect 16935 2815 16950 2835
rect 16900 2785 16950 2815
rect 16900 2765 16915 2785
rect 16935 2765 16950 2785
rect 16900 2750 16950 2765
rect 17050 3035 17100 3050
rect 17050 3015 17065 3035
rect 17085 3015 17100 3035
rect 17050 2985 17100 3015
rect 17050 2965 17065 2985
rect 17085 2965 17100 2985
rect 17050 2935 17100 2965
rect 17050 2915 17065 2935
rect 17085 2915 17100 2935
rect 17050 2885 17100 2915
rect 17050 2865 17065 2885
rect 17085 2865 17100 2885
rect 17050 2835 17100 2865
rect 17050 2815 17065 2835
rect 17085 2815 17100 2835
rect 17050 2785 17100 2815
rect 17050 2765 17065 2785
rect 17085 2765 17100 2785
rect 16750 2715 16765 2735
rect 16785 2715 16800 2735
rect 16750 2700 16800 2715
rect 17050 2735 17100 2765
rect 17200 3035 17250 3065
rect 17200 3015 17215 3035
rect 17235 3015 17250 3035
rect 17200 2985 17250 3015
rect 17200 2965 17215 2985
rect 17235 2965 17250 2985
rect 17200 2935 17250 2965
rect 17200 2915 17215 2935
rect 17235 2915 17250 2935
rect 17200 2885 17250 2915
rect 17200 2865 17215 2885
rect 17235 2865 17250 2885
rect 17200 2835 17250 2865
rect 17200 2815 17215 2835
rect 17235 2815 17250 2835
rect 17200 2785 17250 2815
rect 17200 2765 17215 2785
rect 17235 2765 17250 2785
rect 17200 2750 17250 2765
rect 17350 3135 17400 3315
rect 17950 3685 18000 3700
rect 17950 3665 17965 3685
rect 17985 3665 18000 3685
rect 17950 3640 18000 3665
rect 17950 3610 17960 3640
rect 17990 3610 18000 3640
rect 17950 3585 18000 3610
rect 17950 3565 17965 3585
rect 17985 3565 18000 3585
rect 17950 3540 18000 3565
rect 17950 3510 17960 3540
rect 17990 3510 18000 3540
rect 17950 3485 18000 3510
rect 17950 3465 17965 3485
rect 17985 3465 18000 3485
rect 17950 3440 18000 3465
rect 17950 3410 17960 3440
rect 17990 3410 18000 3440
rect 17950 3385 18000 3410
rect 17950 3365 17965 3385
rect 17985 3365 18000 3385
rect 17950 3340 18000 3365
rect 17950 3310 17960 3340
rect 17990 3310 18000 3340
rect 17500 3240 17550 3250
rect 17500 3210 17510 3240
rect 17540 3210 17550 3240
rect 17500 3200 17550 3210
rect 17800 3240 17850 3250
rect 17800 3210 17810 3240
rect 17840 3210 17850 3240
rect 17800 3200 17850 3210
rect 17350 3115 17365 3135
rect 17385 3115 17400 3135
rect 17350 3085 17400 3115
rect 17350 3065 17365 3085
rect 17385 3065 17400 3085
rect 17350 3035 17400 3065
rect 17350 3015 17365 3035
rect 17385 3015 17400 3035
rect 17350 2985 17400 3015
rect 17350 2965 17365 2985
rect 17385 2965 17400 2985
rect 17350 2935 17400 2965
rect 17350 2915 17365 2935
rect 17385 2915 17400 2935
rect 17350 2885 17400 2915
rect 17350 2865 17365 2885
rect 17385 2865 17400 2885
rect 17350 2835 17400 2865
rect 17350 2815 17365 2835
rect 17385 2815 17400 2835
rect 17350 2785 17400 2815
rect 17350 2765 17365 2785
rect 17385 2765 17400 2785
rect 17050 2715 17065 2735
rect 17085 2715 17100 2735
rect 17050 2700 17100 2715
rect 17350 2735 17400 2765
rect 17950 3140 18000 3310
rect 18550 3685 18600 3715
rect 18850 3735 18900 3750
rect 18850 3715 18865 3735
rect 18885 3715 18900 3735
rect 18550 3665 18565 3685
rect 18585 3665 18600 3685
rect 18550 3635 18600 3665
rect 18550 3615 18565 3635
rect 18585 3615 18600 3635
rect 18550 3585 18600 3615
rect 18550 3565 18565 3585
rect 18585 3565 18600 3585
rect 18550 3535 18600 3565
rect 18550 3515 18565 3535
rect 18585 3515 18600 3535
rect 18550 3485 18600 3515
rect 18550 3465 18565 3485
rect 18585 3465 18600 3485
rect 18550 3435 18600 3465
rect 18550 3415 18565 3435
rect 18585 3415 18600 3435
rect 18550 3385 18600 3415
rect 18550 3365 18565 3385
rect 18585 3365 18600 3385
rect 18550 3335 18600 3365
rect 18550 3315 18565 3335
rect 18585 3315 18600 3335
rect 18100 3240 18150 3250
rect 18100 3210 18110 3240
rect 18140 3210 18150 3240
rect 18100 3200 18150 3210
rect 18400 3240 18450 3250
rect 18400 3210 18410 3240
rect 18440 3210 18450 3240
rect 18400 3200 18450 3210
rect 17950 3110 17960 3140
rect 17990 3110 18000 3140
rect 17950 3085 18000 3110
rect 17950 3065 17965 3085
rect 17985 3065 18000 3085
rect 17950 3040 18000 3065
rect 17950 3010 17960 3040
rect 17990 3010 18000 3040
rect 17950 2985 18000 3010
rect 17950 2965 17965 2985
rect 17985 2965 18000 2985
rect 17950 2940 18000 2965
rect 17950 2910 17960 2940
rect 17990 2910 18000 2940
rect 17950 2885 18000 2910
rect 17950 2865 17965 2885
rect 17985 2865 18000 2885
rect 17950 2840 18000 2865
rect 17950 2810 17960 2840
rect 17990 2810 18000 2840
rect 17950 2785 18000 2810
rect 17950 2765 17965 2785
rect 17985 2765 18000 2785
rect 17950 2750 18000 2765
rect 18550 3135 18600 3315
rect 18700 3685 18750 3700
rect 18700 3665 18715 3685
rect 18735 3665 18750 3685
rect 18700 3635 18750 3665
rect 18700 3615 18715 3635
rect 18735 3615 18750 3635
rect 18700 3585 18750 3615
rect 18700 3565 18715 3585
rect 18735 3565 18750 3585
rect 18700 3535 18750 3565
rect 18700 3515 18715 3535
rect 18735 3515 18750 3535
rect 18700 3485 18750 3515
rect 18700 3465 18715 3485
rect 18735 3465 18750 3485
rect 18700 3435 18750 3465
rect 18700 3415 18715 3435
rect 18735 3415 18750 3435
rect 18700 3385 18750 3415
rect 18850 3685 18900 3715
rect 19150 3735 19200 3750
rect 19150 3715 19165 3735
rect 19185 3715 19200 3735
rect 18850 3665 18865 3685
rect 18885 3665 18900 3685
rect 18850 3635 18900 3665
rect 18850 3615 18865 3635
rect 18885 3615 18900 3635
rect 18850 3585 18900 3615
rect 18850 3565 18865 3585
rect 18885 3565 18900 3585
rect 18850 3535 18900 3565
rect 18850 3515 18865 3535
rect 18885 3515 18900 3535
rect 18850 3485 18900 3515
rect 18850 3465 18865 3485
rect 18885 3465 18900 3485
rect 18850 3435 18900 3465
rect 18850 3415 18865 3435
rect 18885 3415 18900 3435
rect 18850 3400 18900 3415
rect 19000 3685 19050 3700
rect 19000 3665 19015 3685
rect 19035 3665 19050 3685
rect 19000 3635 19050 3665
rect 19000 3615 19015 3635
rect 19035 3615 19050 3635
rect 19000 3585 19050 3615
rect 19000 3565 19015 3585
rect 19035 3565 19050 3585
rect 19000 3535 19050 3565
rect 19000 3515 19015 3535
rect 19035 3515 19050 3535
rect 19000 3485 19050 3515
rect 19000 3465 19015 3485
rect 19035 3465 19050 3485
rect 19000 3435 19050 3465
rect 19000 3415 19015 3435
rect 19035 3415 19050 3435
rect 18700 3365 18715 3385
rect 18735 3365 18750 3385
rect 18700 3350 18750 3365
rect 19000 3385 19050 3415
rect 19150 3685 19200 3715
rect 19450 3735 19500 3750
rect 19450 3715 19465 3735
rect 19485 3715 19500 3735
rect 19150 3665 19165 3685
rect 19185 3665 19200 3685
rect 19150 3635 19200 3665
rect 19150 3615 19165 3635
rect 19185 3615 19200 3635
rect 19150 3585 19200 3615
rect 19150 3565 19165 3585
rect 19185 3565 19200 3585
rect 19150 3535 19200 3565
rect 19150 3515 19165 3535
rect 19185 3515 19200 3535
rect 19150 3485 19200 3515
rect 19150 3465 19165 3485
rect 19185 3465 19200 3485
rect 19150 3435 19200 3465
rect 19150 3415 19165 3435
rect 19185 3415 19200 3435
rect 19150 3400 19200 3415
rect 19300 3685 19350 3700
rect 19300 3665 19315 3685
rect 19335 3665 19350 3685
rect 19300 3635 19350 3665
rect 19300 3615 19315 3635
rect 19335 3615 19350 3635
rect 19300 3585 19350 3615
rect 19300 3565 19315 3585
rect 19335 3565 19350 3585
rect 19300 3535 19350 3565
rect 19300 3515 19315 3535
rect 19335 3515 19350 3535
rect 19300 3485 19350 3515
rect 19300 3465 19315 3485
rect 19335 3465 19350 3485
rect 19300 3435 19350 3465
rect 19300 3415 19315 3435
rect 19335 3415 19350 3435
rect 19000 3365 19015 3385
rect 19035 3365 19050 3385
rect 19000 3350 19050 3365
rect 19300 3385 19350 3415
rect 19450 3685 19500 3715
rect 19750 3735 19800 3750
rect 19750 3715 19765 3735
rect 19785 3715 19800 3735
rect 19450 3665 19465 3685
rect 19485 3665 19500 3685
rect 19450 3635 19500 3665
rect 19450 3615 19465 3635
rect 19485 3615 19500 3635
rect 19450 3585 19500 3615
rect 19450 3565 19465 3585
rect 19485 3565 19500 3585
rect 19450 3535 19500 3565
rect 19450 3515 19465 3535
rect 19485 3515 19500 3535
rect 19450 3485 19500 3515
rect 19450 3465 19465 3485
rect 19485 3465 19500 3485
rect 19450 3435 19500 3465
rect 19450 3415 19465 3435
rect 19485 3415 19500 3435
rect 19450 3400 19500 3415
rect 19600 3685 19650 3700
rect 19600 3665 19615 3685
rect 19635 3665 19650 3685
rect 19600 3635 19650 3665
rect 19600 3615 19615 3635
rect 19635 3615 19650 3635
rect 19600 3585 19650 3615
rect 19600 3565 19615 3585
rect 19635 3565 19650 3585
rect 19600 3535 19650 3565
rect 19600 3515 19615 3535
rect 19635 3515 19650 3535
rect 19600 3485 19650 3515
rect 19600 3465 19615 3485
rect 19635 3465 19650 3485
rect 19600 3435 19650 3465
rect 19600 3415 19615 3435
rect 19635 3415 19650 3435
rect 19300 3365 19315 3385
rect 19335 3365 19350 3385
rect 19300 3350 19350 3365
rect 19600 3385 19650 3415
rect 19600 3365 19615 3385
rect 19635 3365 19650 3385
rect 19600 3350 19650 3365
rect 18700 3335 19650 3350
rect 18700 3315 18715 3335
rect 18735 3315 19015 3335
rect 19035 3315 19315 3335
rect 19335 3315 19615 3335
rect 19635 3315 19650 3335
rect 18700 3300 19650 3315
rect 19750 3685 19800 3715
rect 19750 3665 19765 3685
rect 19785 3665 19800 3685
rect 19750 3635 19800 3665
rect 19750 3615 19765 3635
rect 19785 3615 19800 3635
rect 19750 3585 19800 3615
rect 19750 3565 19765 3585
rect 19785 3565 19800 3585
rect 19750 3535 19800 3565
rect 19750 3515 19765 3535
rect 19785 3515 19800 3535
rect 19750 3485 19800 3515
rect 19750 3465 19765 3485
rect 19785 3465 19800 3485
rect 19750 3435 19800 3465
rect 19750 3415 19765 3435
rect 19785 3415 19800 3435
rect 19750 3385 19800 3415
rect 19750 3365 19765 3385
rect 19785 3365 19800 3385
rect 19750 3335 19800 3365
rect 19750 3315 19765 3335
rect 19785 3315 19800 3335
rect 18700 3240 18750 3250
rect 18700 3210 18710 3240
rect 18740 3210 18750 3240
rect 18700 3200 18750 3210
rect 19000 3240 19050 3250
rect 19000 3210 19010 3240
rect 19040 3210 19050 3240
rect 19000 3200 19050 3210
rect 19150 3240 19200 3300
rect 19150 3210 19160 3240
rect 19190 3210 19200 3240
rect 19150 3150 19200 3210
rect 19300 3240 19350 3250
rect 19300 3210 19310 3240
rect 19340 3210 19350 3240
rect 19300 3200 19350 3210
rect 19600 3240 19650 3250
rect 19600 3210 19610 3240
rect 19640 3210 19650 3240
rect 19600 3200 19650 3210
rect 18550 3115 18565 3135
rect 18585 3115 18600 3135
rect 18550 3085 18600 3115
rect 18550 3065 18565 3085
rect 18585 3065 18600 3085
rect 18550 3035 18600 3065
rect 18550 3015 18565 3035
rect 18585 3015 18600 3035
rect 18550 2985 18600 3015
rect 18550 2965 18565 2985
rect 18585 2965 18600 2985
rect 18550 2935 18600 2965
rect 18550 2915 18565 2935
rect 18585 2915 18600 2935
rect 18550 2885 18600 2915
rect 18550 2865 18565 2885
rect 18585 2865 18600 2885
rect 18550 2835 18600 2865
rect 18550 2815 18565 2835
rect 18585 2815 18600 2835
rect 18550 2785 18600 2815
rect 18550 2765 18565 2785
rect 18585 2765 18600 2785
rect 17350 2715 17365 2735
rect 17385 2715 17400 2735
rect 17350 2700 17400 2715
rect 18550 2735 18600 2765
rect 18700 3135 19650 3150
rect 18700 3115 18715 3135
rect 18735 3115 19015 3135
rect 19035 3115 19315 3135
rect 19335 3115 19615 3135
rect 19635 3115 19650 3135
rect 18700 3100 19650 3115
rect 18700 3085 18750 3100
rect 18700 3065 18715 3085
rect 18735 3065 18750 3085
rect 18700 3035 18750 3065
rect 19000 3085 19050 3100
rect 19000 3065 19015 3085
rect 19035 3065 19050 3085
rect 18700 3015 18715 3035
rect 18735 3015 18750 3035
rect 18700 2985 18750 3015
rect 18700 2965 18715 2985
rect 18735 2965 18750 2985
rect 18700 2935 18750 2965
rect 18700 2915 18715 2935
rect 18735 2915 18750 2935
rect 18700 2885 18750 2915
rect 18700 2865 18715 2885
rect 18735 2865 18750 2885
rect 18700 2835 18750 2865
rect 18700 2815 18715 2835
rect 18735 2815 18750 2835
rect 18700 2785 18750 2815
rect 18700 2765 18715 2785
rect 18735 2765 18750 2785
rect 18700 2750 18750 2765
rect 18850 3035 18900 3050
rect 18850 3015 18865 3035
rect 18885 3015 18900 3035
rect 18850 2985 18900 3015
rect 18850 2965 18865 2985
rect 18885 2965 18900 2985
rect 18850 2935 18900 2965
rect 18850 2915 18865 2935
rect 18885 2915 18900 2935
rect 18850 2885 18900 2915
rect 18850 2865 18865 2885
rect 18885 2865 18900 2885
rect 18850 2835 18900 2865
rect 18850 2815 18865 2835
rect 18885 2815 18900 2835
rect 18850 2785 18900 2815
rect 18850 2765 18865 2785
rect 18885 2765 18900 2785
rect 18550 2715 18565 2735
rect 18585 2715 18600 2735
rect 18550 2700 18600 2715
rect 18850 2735 18900 2765
rect 19000 3035 19050 3065
rect 19300 3085 19350 3100
rect 19300 3065 19315 3085
rect 19335 3065 19350 3085
rect 19000 3015 19015 3035
rect 19035 3015 19050 3035
rect 19000 2985 19050 3015
rect 19000 2965 19015 2985
rect 19035 2965 19050 2985
rect 19000 2935 19050 2965
rect 19000 2915 19015 2935
rect 19035 2915 19050 2935
rect 19000 2885 19050 2915
rect 19000 2865 19015 2885
rect 19035 2865 19050 2885
rect 19000 2835 19050 2865
rect 19000 2815 19015 2835
rect 19035 2815 19050 2835
rect 19000 2785 19050 2815
rect 19000 2765 19015 2785
rect 19035 2765 19050 2785
rect 19000 2750 19050 2765
rect 19150 3035 19200 3050
rect 19150 3015 19165 3035
rect 19185 3015 19200 3035
rect 19150 2985 19200 3015
rect 19150 2965 19165 2985
rect 19185 2965 19200 2985
rect 19150 2935 19200 2965
rect 19150 2915 19165 2935
rect 19185 2915 19200 2935
rect 19150 2885 19200 2915
rect 19150 2865 19165 2885
rect 19185 2865 19200 2885
rect 19150 2835 19200 2865
rect 19150 2815 19165 2835
rect 19185 2815 19200 2835
rect 19150 2785 19200 2815
rect 19150 2765 19165 2785
rect 19185 2765 19200 2785
rect 18850 2715 18865 2735
rect 18885 2715 18900 2735
rect 18850 2700 18900 2715
rect 19150 2735 19200 2765
rect 19300 3035 19350 3065
rect 19600 3085 19650 3100
rect 19600 3065 19615 3085
rect 19635 3065 19650 3085
rect 19300 3015 19315 3035
rect 19335 3015 19350 3035
rect 19300 2985 19350 3015
rect 19300 2965 19315 2985
rect 19335 2965 19350 2985
rect 19300 2935 19350 2965
rect 19300 2915 19315 2935
rect 19335 2915 19350 2935
rect 19300 2885 19350 2915
rect 19300 2865 19315 2885
rect 19335 2865 19350 2885
rect 19300 2835 19350 2865
rect 19300 2815 19315 2835
rect 19335 2815 19350 2835
rect 19300 2785 19350 2815
rect 19300 2765 19315 2785
rect 19335 2765 19350 2785
rect 19300 2750 19350 2765
rect 19450 3035 19500 3050
rect 19450 3015 19465 3035
rect 19485 3015 19500 3035
rect 19450 2985 19500 3015
rect 19450 2965 19465 2985
rect 19485 2965 19500 2985
rect 19450 2935 19500 2965
rect 19450 2915 19465 2935
rect 19485 2915 19500 2935
rect 19450 2885 19500 2915
rect 19450 2865 19465 2885
rect 19485 2865 19500 2885
rect 19450 2835 19500 2865
rect 19450 2815 19465 2835
rect 19485 2815 19500 2835
rect 19450 2785 19500 2815
rect 19450 2765 19465 2785
rect 19485 2765 19500 2785
rect 19150 2715 19165 2735
rect 19185 2715 19200 2735
rect 19150 2700 19200 2715
rect 19450 2735 19500 2765
rect 19600 3035 19650 3065
rect 19600 3015 19615 3035
rect 19635 3015 19650 3035
rect 19600 2985 19650 3015
rect 19600 2965 19615 2985
rect 19635 2965 19650 2985
rect 19600 2935 19650 2965
rect 19600 2915 19615 2935
rect 19635 2915 19650 2935
rect 19600 2885 19650 2915
rect 19600 2865 19615 2885
rect 19635 2865 19650 2885
rect 19600 2835 19650 2865
rect 19600 2815 19615 2835
rect 19635 2815 19650 2835
rect 19600 2785 19650 2815
rect 19600 2765 19615 2785
rect 19635 2765 19650 2785
rect 19600 2750 19650 2765
rect 19750 3135 19800 3315
rect 20350 3785 20400 3860
rect 20350 3765 20365 3785
rect 20385 3765 20400 3785
rect 20350 3740 20400 3765
rect 20350 3710 20360 3740
rect 20390 3710 20400 3740
rect 20350 3685 20400 3710
rect 20350 3665 20365 3685
rect 20385 3665 20400 3685
rect 20350 3640 20400 3665
rect 20350 3610 20360 3640
rect 20390 3610 20400 3640
rect 20350 3585 20400 3610
rect 20350 3565 20365 3585
rect 20385 3565 20400 3585
rect 20350 3540 20400 3565
rect 20350 3510 20360 3540
rect 20390 3510 20400 3540
rect 20350 3485 20400 3510
rect 20350 3465 20365 3485
rect 20385 3465 20400 3485
rect 20350 3440 20400 3465
rect 20350 3410 20360 3440
rect 20390 3410 20400 3440
rect 20350 3385 20400 3410
rect 20350 3365 20365 3385
rect 20385 3365 20400 3385
rect 20350 3340 20400 3365
rect 20350 3310 20360 3340
rect 20390 3310 20400 3340
rect 19900 3240 19950 3250
rect 19900 3210 19910 3240
rect 19940 3210 19950 3240
rect 19900 3200 19950 3210
rect 20200 3240 20250 3250
rect 20200 3210 20210 3240
rect 20240 3210 20250 3240
rect 20200 3200 20250 3210
rect 19750 3115 19765 3135
rect 19785 3115 19800 3135
rect 19750 3085 19800 3115
rect 19750 3065 19765 3085
rect 19785 3065 19800 3085
rect 19750 3035 19800 3065
rect 19750 3015 19765 3035
rect 19785 3015 19800 3035
rect 19750 2985 19800 3015
rect 19750 2965 19765 2985
rect 19785 2965 19800 2985
rect 19750 2935 19800 2965
rect 19750 2915 19765 2935
rect 19785 2915 19800 2935
rect 19750 2885 19800 2915
rect 19750 2865 19765 2885
rect 19785 2865 19800 2885
rect 19750 2835 19800 2865
rect 19750 2815 19765 2835
rect 19785 2815 19800 2835
rect 19750 2785 19800 2815
rect 19750 2765 19765 2785
rect 19785 2765 19800 2785
rect 19450 2715 19465 2735
rect 19485 2715 19500 2735
rect 19450 2700 19500 2715
rect 19750 2735 19800 2765
rect 19750 2715 19765 2735
rect 19785 2715 19800 2735
rect 19750 2700 19800 2715
rect 16150 2685 19800 2700
rect 16150 2665 16165 2685
rect 16185 2665 16465 2685
rect 16485 2665 16765 2685
rect 16785 2665 17065 2685
rect 17085 2665 17365 2685
rect 17385 2665 18565 2685
rect 18585 2665 18865 2685
rect 18885 2665 19165 2685
rect 19185 2665 19465 2685
rect 19485 2665 19765 2685
rect 19785 2665 19800 2685
rect 16150 2650 19800 2665
rect 20350 3140 20400 3310
rect 20350 3110 20360 3140
rect 20390 3110 20400 3140
rect 20350 3085 20400 3110
rect 20350 3065 20365 3085
rect 20385 3065 20400 3085
rect 20350 3040 20400 3065
rect 20350 3010 20360 3040
rect 20390 3010 20400 3040
rect 20350 2985 20400 3010
rect 20350 2965 20365 2985
rect 20385 2965 20400 2985
rect 20350 2940 20400 2965
rect 20350 2910 20360 2940
rect 20390 2910 20400 2940
rect 20350 2885 20400 2910
rect 20350 2865 20365 2885
rect 20385 2865 20400 2885
rect 20350 2840 20400 2865
rect 20350 2810 20360 2840
rect 20390 2810 20400 2840
rect 20350 2785 20400 2810
rect 20350 2765 20365 2785
rect 20385 2765 20400 2785
rect 20350 2740 20400 2765
rect 20350 2710 20360 2740
rect 20390 2710 20400 2740
rect 20350 2685 20400 2710
rect 20350 2665 20365 2685
rect 20385 2665 20400 2685
rect 15550 2560 15560 2590
rect 15590 2560 15600 2590
rect 15550 2550 15600 2560
rect 17950 2590 18000 2650
rect 17950 2560 17960 2590
rect 17990 2560 18000 2590
rect 17950 2550 18000 2560
rect 20350 2590 20400 2665
rect 20350 2560 20360 2590
rect 20390 2560 20400 2590
rect 20350 2550 20400 2560
rect -650 1690 -600 1700
rect -650 1660 -640 1690
rect -610 1660 -600 1690
rect -650 1585 -600 1660
rect -50 1690 0 1700
rect -50 1660 -40 1690
rect -10 1660 0 1690
rect -650 1565 -635 1585
rect -615 1565 -600 1585
rect -650 1540 -600 1565
rect -650 1510 -640 1540
rect -610 1510 -600 1540
rect -650 1485 -600 1510
rect -650 1465 -635 1485
rect -615 1465 -600 1485
rect -650 1440 -600 1465
rect -650 1410 -640 1440
rect -610 1410 -600 1440
rect -650 1385 -600 1410
rect -650 1365 -635 1385
rect -615 1365 -600 1385
rect -650 1340 -600 1365
rect -650 1310 -640 1340
rect -610 1310 -600 1340
rect -650 1285 -600 1310
rect -650 1265 -635 1285
rect -615 1265 -600 1285
rect -650 1240 -600 1265
rect -650 1210 -640 1240
rect -610 1210 -600 1240
rect -650 1185 -600 1210
rect -650 1165 -635 1185
rect -615 1165 -600 1185
rect -650 1140 -600 1165
rect -650 1110 -640 1140
rect -610 1110 -600 1140
rect -650 1085 -600 1110
rect -650 1065 -635 1085
rect -615 1065 -600 1085
rect -650 1040 -600 1065
rect -650 1010 -640 1040
rect -610 1010 -600 1040
rect -650 985 -600 1010
rect -650 965 -635 985
rect -615 965 -600 985
rect -650 940 -600 965
rect -650 910 -640 940
rect -610 910 -600 940
rect -650 740 -600 910
rect -500 1585 -450 1600
rect -500 1565 -485 1585
rect -465 1565 -450 1585
rect -500 1535 -450 1565
rect -500 1515 -485 1535
rect -465 1515 -450 1535
rect -500 1485 -450 1515
rect -500 1465 -485 1485
rect -465 1465 -450 1485
rect -500 1435 -450 1465
rect -500 1415 -485 1435
rect -465 1415 -450 1435
rect -500 1385 -450 1415
rect -500 1365 -485 1385
rect -465 1365 -450 1385
rect -500 1335 -450 1365
rect -500 1315 -485 1335
rect -465 1315 -450 1335
rect -500 1285 -450 1315
rect -500 1265 -485 1285
rect -465 1265 -450 1285
rect -500 1235 -450 1265
rect -500 1215 -485 1235
rect -465 1215 -450 1235
rect -500 1185 -450 1215
rect -500 1165 -485 1185
rect -465 1165 -450 1185
rect -500 1135 -450 1165
rect -500 1115 -485 1135
rect -465 1115 -450 1135
rect -500 1085 -450 1115
rect -500 1065 -485 1085
rect -465 1065 -450 1085
rect -500 1035 -450 1065
rect -500 1015 -485 1035
rect -465 1015 -450 1035
rect -500 985 -450 1015
rect -500 965 -485 985
rect -465 965 -450 985
rect -500 935 -450 965
rect -500 915 -485 935
rect -465 915 -450 935
rect -500 900 -450 915
rect -350 1585 -300 1600
rect -350 1565 -335 1585
rect -315 1565 -300 1585
rect -350 1535 -300 1565
rect -350 1515 -335 1535
rect -315 1515 -300 1535
rect -350 1485 -300 1515
rect -350 1465 -335 1485
rect -315 1465 -300 1485
rect -350 1435 -300 1465
rect -350 1415 -335 1435
rect -315 1415 -300 1435
rect -350 1385 -300 1415
rect -350 1365 -335 1385
rect -315 1365 -300 1385
rect -350 1335 -300 1365
rect -350 1315 -335 1335
rect -315 1315 -300 1335
rect -350 1285 -300 1315
rect -350 1265 -335 1285
rect -315 1265 -300 1285
rect -350 1235 -300 1265
rect -350 1215 -335 1235
rect -315 1215 -300 1235
rect -350 1185 -300 1215
rect -350 1165 -335 1185
rect -315 1165 -300 1185
rect -350 1135 -300 1165
rect -350 1115 -335 1135
rect -315 1115 -300 1135
rect -350 1085 -300 1115
rect -350 1065 -335 1085
rect -315 1065 -300 1085
rect -350 1035 -300 1065
rect -350 1015 -335 1035
rect -315 1015 -300 1035
rect -350 985 -300 1015
rect -350 965 -335 985
rect -315 965 -300 985
rect -350 935 -300 965
rect -350 915 -335 935
rect -315 915 -300 935
rect -500 840 -450 850
rect -500 810 -490 840
rect -460 810 -450 840
rect -500 800 -450 810
rect -350 840 -300 915
rect -200 1585 -150 1600
rect -200 1565 -185 1585
rect -165 1565 -150 1585
rect -200 1535 -150 1565
rect -200 1515 -185 1535
rect -165 1515 -150 1535
rect -200 1485 -150 1515
rect -200 1465 -185 1485
rect -165 1465 -150 1485
rect -200 1435 -150 1465
rect -200 1415 -185 1435
rect -165 1415 -150 1435
rect -200 1385 -150 1415
rect -200 1365 -185 1385
rect -165 1365 -150 1385
rect -200 1335 -150 1365
rect -200 1315 -185 1335
rect -165 1315 -150 1335
rect -200 1285 -150 1315
rect -200 1265 -185 1285
rect -165 1265 -150 1285
rect -200 1235 -150 1265
rect -200 1215 -185 1235
rect -165 1215 -150 1235
rect -200 1185 -150 1215
rect -200 1165 -185 1185
rect -165 1165 -150 1185
rect -200 1135 -150 1165
rect -200 1115 -185 1135
rect -165 1115 -150 1135
rect -200 1085 -150 1115
rect -200 1065 -185 1085
rect -165 1065 -150 1085
rect -200 1035 -150 1065
rect -200 1015 -185 1035
rect -165 1015 -150 1035
rect -200 985 -150 1015
rect -200 965 -185 985
rect -165 965 -150 985
rect -200 935 -150 965
rect -200 915 -185 935
rect -165 915 -150 935
rect -200 900 -150 915
rect -50 1585 0 1660
rect 8350 1690 8400 1700
rect 8350 1660 8360 1690
rect 8390 1660 8400 1690
rect -50 1565 -35 1585
rect -15 1565 0 1585
rect -50 1540 0 1565
rect -50 1510 -40 1540
rect -10 1510 0 1540
rect -50 1485 0 1510
rect -50 1465 -35 1485
rect -15 1465 0 1485
rect -50 1440 0 1465
rect -50 1410 -40 1440
rect -10 1410 0 1440
rect -50 1385 0 1410
rect -50 1365 -35 1385
rect -15 1365 0 1385
rect -50 1340 0 1365
rect -50 1310 -40 1340
rect -10 1310 0 1340
rect -50 1285 0 1310
rect -50 1265 -35 1285
rect -15 1265 0 1285
rect -50 1240 0 1265
rect -50 1210 -40 1240
rect -10 1210 0 1240
rect -50 1185 0 1210
rect -50 1165 -35 1185
rect -15 1165 0 1185
rect -50 1140 0 1165
rect -50 1110 -40 1140
rect -10 1110 0 1140
rect -50 1085 0 1110
rect -50 1065 -35 1085
rect -15 1065 0 1085
rect -50 1040 0 1065
rect -50 1010 -40 1040
rect -10 1010 0 1040
rect -50 985 0 1010
rect -50 965 -35 985
rect -15 965 0 985
rect -50 940 0 965
rect -50 910 -40 940
rect -10 910 0 940
rect -350 810 -340 840
rect -310 810 -300 840
rect -650 710 -640 740
rect -610 710 -600 740
rect -650 685 -600 710
rect -650 665 -635 685
rect -615 665 -600 685
rect -650 640 -600 665
rect -650 610 -640 640
rect -610 610 -600 640
rect -650 585 -600 610
rect -650 565 -635 585
rect -615 565 -600 585
rect -650 540 -600 565
rect -650 510 -640 540
rect -610 510 -600 540
rect -650 485 -600 510
rect -650 465 -635 485
rect -615 465 -600 485
rect -650 440 -600 465
rect -650 410 -640 440
rect -610 410 -600 440
rect -650 385 -600 410
rect -650 365 -635 385
rect -615 365 -600 385
rect -650 340 -600 365
rect -650 310 -640 340
rect -610 310 -600 340
rect -650 285 -600 310
rect -650 265 -635 285
rect -615 265 -600 285
rect -650 240 -600 265
rect -650 210 -640 240
rect -610 210 -600 240
rect -650 185 -600 210
rect -650 165 -635 185
rect -615 165 -600 185
rect -650 140 -600 165
rect -650 110 -640 140
rect -610 110 -600 140
rect -650 85 -600 110
rect -650 65 -635 85
rect -615 65 -600 85
rect -650 -10 -600 65
rect -500 735 -450 750
rect -500 715 -485 735
rect -465 715 -450 735
rect -500 685 -450 715
rect -500 665 -485 685
rect -465 665 -450 685
rect -500 635 -450 665
rect -500 615 -485 635
rect -465 615 -450 635
rect -500 585 -450 615
rect -500 565 -485 585
rect -465 565 -450 585
rect -500 535 -450 565
rect -500 515 -485 535
rect -465 515 -450 535
rect -500 485 -450 515
rect -500 465 -485 485
rect -465 465 -450 485
rect -500 435 -450 465
rect -500 415 -485 435
rect -465 415 -450 435
rect -500 385 -450 415
rect -500 365 -485 385
rect -465 365 -450 385
rect -500 335 -450 365
rect -500 315 -485 335
rect -465 315 -450 335
rect -500 285 -450 315
rect -500 265 -485 285
rect -465 265 -450 285
rect -500 235 -450 265
rect -500 215 -485 235
rect -465 215 -450 235
rect -500 185 -450 215
rect -500 165 -485 185
rect -465 165 -450 185
rect -500 135 -450 165
rect -500 115 -485 135
rect -465 115 -450 135
rect -500 85 -450 115
rect -500 65 -485 85
rect -465 65 -450 85
rect -500 50 -450 65
rect -350 735 -300 810
rect -200 840 -150 850
rect -200 810 -190 840
rect -160 810 -150 840
rect -200 800 -150 810
rect -350 715 -335 735
rect -315 715 -300 735
rect -350 685 -300 715
rect -350 665 -335 685
rect -315 665 -300 685
rect -350 635 -300 665
rect -350 615 -335 635
rect -315 615 -300 635
rect -350 585 -300 615
rect -350 565 -335 585
rect -315 565 -300 585
rect -350 535 -300 565
rect -350 515 -335 535
rect -315 515 -300 535
rect -350 485 -300 515
rect -350 465 -335 485
rect -315 465 -300 485
rect -350 435 -300 465
rect -350 415 -335 435
rect -315 415 -300 435
rect -350 385 -300 415
rect -350 365 -335 385
rect -315 365 -300 385
rect -350 335 -300 365
rect -350 315 -335 335
rect -315 315 -300 335
rect -350 285 -300 315
rect -350 265 -335 285
rect -315 265 -300 285
rect -350 235 -300 265
rect -350 215 -335 235
rect -315 215 -300 235
rect -350 185 -300 215
rect -350 165 -335 185
rect -315 165 -300 185
rect -350 135 -300 165
rect -350 115 -335 135
rect -315 115 -300 135
rect -350 85 -300 115
rect -350 65 -335 85
rect -315 65 -300 85
rect -350 50 -300 65
rect -200 735 -150 750
rect -200 715 -185 735
rect -165 715 -150 735
rect -200 685 -150 715
rect -200 665 -185 685
rect -165 665 -150 685
rect -200 635 -150 665
rect -200 615 -185 635
rect -165 615 -150 635
rect -200 585 -150 615
rect -200 565 -185 585
rect -165 565 -150 585
rect -200 535 -150 565
rect -200 515 -185 535
rect -165 515 -150 535
rect -200 485 -150 515
rect -200 465 -185 485
rect -165 465 -150 485
rect -200 435 -150 465
rect -200 415 -185 435
rect -165 415 -150 435
rect -200 385 -150 415
rect -200 365 -185 385
rect -165 365 -150 385
rect -200 335 -150 365
rect -200 315 -185 335
rect -165 315 -150 335
rect -200 285 -150 315
rect -200 265 -185 285
rect -165 265 -150 285
rect -200 235 -150 265
rect -200 215 -185 235
rect -165 215 -150 235
rect -200 185 -150 215
rect -200 165 -185 185
rect -165 165 -150 185
rect -200 135 -150 165
rect -200 115 -185 135
rect -165 115 -150 135
rect -200 85 -150 115
rect -200 65 -185 85
rect -165 65 -150 85
rect -200 50 -150 65
rect -50 740 0 910
rect 1150 1585 7200 1600
rect 1150 1565 1165 1585
rect 1185 1565 1765 1585
rect 1785 1565 2365 1585
rect 2385 1565 2965 1585
rect 2985 1565 3565 1585
rect 3585 1565 3865 1585
rect 3885 1565 4165 1585
rect 4185 1565 4465 1585
rect 4485 1565 4765 1585
rect 4785 1565 5365 1585
rect 5385 1565 5965 1585
rect 5985 1565 6565 1585
rect 6585 1565 7165 1585
rect 7185 1565 7200 1585
rect 1150 1550 7200 1565
rect 1150 1535 1200 1550
rect 1150 1515 1165 1535
rect 1185 1515 1200 1535
rect 1150 1485 1200 1515
rect 1750 1535 1800 1550
rect 1750 1515 1765 1535
rect 1785 1515 1800 1535
rect 1150 1465 1165 1485
rect 1185 1465 1200 1485
rect 1150 1435 1200 1465
rect 1150 1415 1165 1435
rect 1185 1415 1200 1435
rect 1150 1385 1200 1415
rect 1150 1365 1165 1385
rect 1185 1365 1200 1385
rect 1150 1335 1200 1365
rect 1150 1315 1165 1335
rect 1185 1315 1200 1335
rect 1150 1285 1200 1315
rect 1150 1265 1165 1285
rect 1185 1265 1200 1285
rect 1150 1235 1200 1265
rect 1150 1215 1165 1235
rect 1185 1215 1200 1235
rect 1150 1185 1200 1215
rect 1150 1165 1165 1185
rect 1185 1165 1200 1185
rect 1150 1135 1200 1165
rect 1150 1115 1165 1135
rect 1185 1115 1200 1135
rect 1150 1085 1200 1115
rect 1150 1065 1165 1085
rect 1185 1065 1200 1085
rect 1150 1035 1200 1065
rect 1150 1015 1165 1035
rect 1185 1015 1200 1035
rect 1150 985 1200 1015
rect 1150 965 1165 985
rect 1185 965 1200 985
rect 1150 935 1200 965
rect 1150 915 1165 935
rect 1185 915 1200 935
rect 1150 900 1200 915
rect 1450 1485 1500 1500
rect 1450 1465 1465 1485
rect 1485 1465 1500 1485
rect 1450 1435 1500 1465
rect 1450 1415 1465 1435
rect 1485 1415 1500 1435
rect 1450 1385 1500 1415
rect 1450 1365 1465 1385
rect 1485 1365 1500 1385
rect 1450 1335 1500 1365
rect 1450 1315 1465 1335
rect 1485 1315 1500 1335
rect 1450 1285 1500 1315
rect 1450 1265 1465 1285
rect 1485 1265 1500 1285
rect 1450 1235 1500 1265
rect 1450 1215 1465 1235
rect 1485 1215 1500 1235
rect 1450 1185 1500 1215
rect 1450 1165 1465 1185
rect 1485 1165 1500 1185
rect 1450 1135 1500 1165
rect 1450 1115 1465 1135
rect 1485 1115 1500 1135
rect 1450 1085 1500 1115
rect 1450 1065 1465 1085
rect 1485 1065 1500 1085
rect 1450 1035 1500 1065
rect 1450 1015 1465 1035
rect 1485 1015 1500 1035
rect 1450 985 1500 1015
rect 1750 1485 1800 1515
rect 2350 1535 2400 1550
rect 2350 1515 2365 1535
rect 2385 1515 2400 1535
rect 1750 1465 1765 1485
rect 1785 1465 1800 1485
rect 1750 1435 1800 1465
rect 1750 1415 1765 1435
rect 1785 1415 1800 1435
rect 1750 1385 1800 1415
rect 1750 1365 1765 1385
rect 1785 1365 1800 1385
rect 1750 1335 1800 1365
rect 1750 1315 1765 1335
rect 1785 1315 1800 1335
rect 1750 1285 1800 1315
rect 1750 1265 1765 1285
rect 1785 1265 1800 1285
rect 1750 1235 1800 1265
rect 1750 1215 1765 1235
rect 1785 1215 1800 1235
rect 1750 1185 1800 1215
rect 1750 1165 1765 1185
rect 1785 1165 1800 1185
rect 1750 1135 1800 1165
rect 1750 1115 1765 1135
rect 1785 1115 1800 1135
rect 1750 1085 1800 1115
rect 1750 1065 1765 1085
rect 1785 1065 1800 1085
rect 1750 1035 1800 1065
rect 1750 1015 1765 1035
rect 1785 1015 1800 1035
rect 1750 1000 1800 1015
rect 2050 1485 2100 1500
rect 2050 1465 2065 1485
rect 2085 1465 2100 1485
rect 2050 1435 2100 1465
rect 2050 1415 2065 1435
rect 2085 1415 2100 1435
rect 2050 1385 2100 1415
rect 2050 1365 2065 1385
rect 2085 1365 2100 1385
rect 2050 1335 2100 1365
rect 2050 1315 2065 1335
rect 2085 1315 2100 1335
rect 2050 1285 2100 1315
rect 2050 1265 2065 1285
rect 2085 1265 2100 1285
rect 2050 1235 2100 1265
rect 2050 1215 2065 1235
rect 2085 1215 2100 1235
rect 2050 1185 2100 1215
rect 2050 1165 2065 1185
rect 2085 1165 2100 1185
rect 2050 1135 2100 1165
rect 2050 1115 2065 1135
rect 2085 1115 2100 1135
rect 2050 1085 2100 1115
rect 2050 1065 2065 1085
rect 2085 1065 2100 1085
rect 2050 1035 2100 1065
rect 2050 1015 2065 1035
rect 2085 1015 2100 1035
rect 1450 965 1465 985
rect 1485 965 1500 985
rect 1450 950 1500 965
rect 2050 985 2100 1015
rect 2350 1485 2400 1515
rect 2950 1535 3000 1550
rect 2950 1515 2965 1535
rect 2985 1515 3000 1535
rect 2350 1465 2365 1485
rect 2385 1465 2400 1485
rect 2350 1435 2400 1465
rect 2350 1415 2365 1435
rect 2385 1415 2400 1435
rect 2350 1385 2400 1415
rect 2350 1365 2365 1385
rect 2385 1365 2400 1385
rect 2350 1335 2400 1365
rect 2350 1315 2365 1335
rect 2385 1315 2400 1335
rect 2350 1285 2400 1315
rect 2350 1265 2365 1285
rect 2385 1265 2400 1285
rect 2350 1235 2400 1265
rect 2350 1215 2365 1235
rect 2385 1215 2400 1235
rect 2350 1185 2400 1215
rect 2350 1165 2365 1185
rect 2385 1165 2400 1185
rect 2350 1135 2400 1165
rect 2350 1115 2365 1135
rect 2385 1115 2400 1135
rect 2350 1085 2400 1115
rect 2350 1065 2365 1085
rect 2385 1065 2400 1085
rect 2350 1035 2400 1065
rect 2350 1015 2365 1035
rect 2385 1015 2400 1035
rect 2350 1000 2400 1015
rect 2650 1485 2700 1500
rect 2650 1465 2665 1485
rect 2685 1465 2700 1485
rect 2650 1435 2700 1465
rect 2650 1415 2665 1435
rect 2685 1415 2700 1435
rect 2650 1385 2700 1415
rect 2650 1365 2665 1385
rect 2685 1365 2700 1385
rect 2650 1335 2700 1365
rect 2650 1315 2665 1335
rect 2685 1315 2700 1335
rect 2650 1285 2700 1315
rect 2650 1265 2665 1285
rect 2685 1265 2700 1285
rect 2650 1235 2700 1265
rect 2650 1215 2665 1235
rect 2685 1215 2700 1235
rect 2650 1185 2700 1215
rect 2650 1165 2665 1185
rect 2685 1165 2700 1185
rect 2650 1135 2700 1165
rect 2650 1115 2665 1135
rect 2685 1115 2700 1135
rect 2650 1085 2700 1115
rect 2650 1065 2665 1085
rect 2685 1065 2700 1085
rect 2650 1035 2700 1065
rect 2650 1015 2665 1035
rect 2685 1015 2700 1035
rect 2050 965 2065 985
rect 2085 965 2100 985
rect 2050 950 2100 965
rect 2650 985 2700 1015
rect 2950 1485 3000 1515
rect 3550 1535 3600 1550
rect 3550 1515 3565 1535
rect 3585 1515 3600 1535
rect 2950 1465 2965 1485
rect 2985 1465 3000 1485
rect 2950 1435 3000 1465
rect 2950 1415 2965 1435
rect 2985 1415 3000 1435
rect 2950 1385 3000 1415
rect 2950 1365 2965 1385
rect 2985 1365 3000 1385
rect 2950 1335 3000 1365
rect 2950 1315 2965 1335
rect 2985 1315 3000 1335
rect 2950 1285 3000 1315
rect 2950 1265 2965 1285
rect 2985 1265 3000 1285
rect 2950 1235 3000 1265
rect 2950 1215 2965 1235
rect 2985 1215 3000 1235
rect 2950 1185 3000 1215
rect 2950 1165 2965 1185
rect 2985 1165 3000 1185
rect 2950 1135 3000 1165
rect 2950 1115 2965 1135
rect 2985 1115 3000 1135
rect 2950 1085 3000 1115
rect 2950 1065 2965 1085
rect 2985 1065 3000 1085
rect 2950 1035 3000 1065
rect 2950 1015 2965 1035
rect 2985 1015 3000 1035
rect 2950 1000 3000 1015
rect 3250 1485 3300 1500
rect 3250 1465 3265 1485
rect 3285 1465 3300 1485
rect 3250 1435 3300 1465
rect 3250 1415 3265 1435
rect 3285 1415 3300 1435
rect 3250 1385 3300 1415
rect 3250 1365 3265 1385
rect 3285 1365 3300 1385
rect 3250 1335 3300 1365
rect 3250 1315 3265 1335
rect 3285 1315 3300 1335
rect 3250 1285 3300 1315
rect 3250 1265 3265 1285
rect 3285 1265 3300 1285
rect 3250 1235 3300 1265
rect 3250 1215 3265 1235
rect 3285 1215 3300 1235
rect 3250 1185 3300 1215
rect 3250 1165 3265 1185
rect 3285 1165 3300 1185
rect 3250 1135 3300 1165
rect 3250 1115 3265 1135
rect 3285 1115 3300 1135
rect 3250 1085 3300 1115
rect 3250 1065 3265 1085
rect 3285 1065 3300 1085
rect 3250 1035 3300 1065
rect 3250 1015 3265 1035
rect 3285 1015 3300 1035
rect 2650 965 2665 985
rect 2685 965 2700 985
rect 2650 950 2700 965
rect 3250 985 3300 1015
rect 3250 965 3265 985
rect 3285 965 3300 985
rect 3250 950 3300 965
rect 1450 935 3300 950
rect 1450 915 1465 935
rect 1485 915 2065 935
rect 2085 915 2665 935
rect 2685 915 3265 935
rect 3285 915 3300 935
rect 1450 900 3300 915
rect 3550 1485 3600 1515
rect 3850 1535 3900 1550
rect 3850 1515 3865 1535
rect 3885 1515 3900 1535
rect 3550 1465 3565 1485
rect 3585 1465 3600 1485
rect 3550 1435 3600 1465
rect 3550 1415 3565 1435
rect 3585 1415 3600 1435
rect 3550 1385 3600 1415
rect 3550 1365 3565 1385
rect 3585 1365 3600 1385
rect 3550 1335 3600 1365
rect 3550 1315 3565 1335
rect 3585 1315 3600 1335
rect 3550 1285 3600 1315
rect 3550 1265 3565 1285
rect 3585 1265 3600 1285
rect 3550 1235 3600 1265
rect 3550 1215 3565 1235
rect 3585 1215 3600 1235
rect 3550 1185 3600 1215
rect 3550 1165 3565 1185
rect 3585 1165 3600 1185
rect 3550 1135 3600 1165
rect 3550 1115 3565 1135
rect 3585 1115 3600 1135
rect 3550 1085 3600 1115
rect 3550 1065 3565 1085
rect 3585 1065 3600 1085
rect 3550 1035 3600 1065
rect 3550 1015 3565 1035
rect 3585 1015 3600 1035
rect 3550 985 3600 1015
rect 3550 965 3565 985
rect 3585 965 3600 985
rect 3550 935 3600 965
rect 3550 915 3565 935
rect 3585 915 3600 935
rect 3550 900 3600 915
rect 3700 1485 3750 1500
rect 3700 1465 3715 1485
rect 3735 1465 3750 1485
rect 3700 1435 3750 1465
rect 3700 1415 3715 1435
rect 3735 1415 3750 1435
rect 3700 1385 3750 1415
rect 3700 1365 3715 1385
rect 3735 1365 3750 1385
rect 3700 1335 3750 1365
rect 3700 1315 3715 1335
rect 3735 1315 3750 1335
rect 3700 1285 3750 1315
rect 3700 1265 3715 1285
rect 3735 1265 3750 1285
rect 3700 1235 3750 1265
rect 3700 1215 3715 1235
rect 3735 1215 3750 1235
rect 3700 1185 3750 1215
rect 3700 1165 3715 1185
rect 3735 1165 3750 1185
rect 3700 1135 3750 1165
rect 3700 1115 3715 1135
rect 3735 1115 3750 1135
rect 3700 1085 3750 1115
rect 3700 1065 3715 1085
rect 3735 1065 3750 1085
rect 3700 1035 3750 1065
rect 3700 1015 3715 1035
rect 3735 1015 3750 1035
rect 3700 985 3750 1015
rect 3850 1485 3900 1515
rect 4150 1535 4200 1550
rect 4150 1515 4165 1535
rect 4185 1515 4200 1535
rect 3850 1465 3865 1485
rect 3885 1465 3900 1485
rect 3850 1435 3900 1465
rect 3850 1415 3865 1435
rect 3885 1415 3900 1435
rect 3850 1385 3900 1415
rect 3850 1365 3865 1385
rect 3885 1365 3900 1385
rect 3850 1335 3900 1365
rect 3850 1315 3865 1335
rect 3885 1315 3900 1335
rect 3850 1285 3900 1315
rect 3850 1265 3865 1285
rect 3885 1265 3900 1285
rect 3850 1235 3900 1265
rect 3850 1215 3865 1235
rect 3885 1215 3900 1235
rect 3850 1185 3900 1215
rect 3850 1165 3865 1185
rect 3885 1165 3900 1185
rect 3850 1135 3900 1165
rect 3850 1115 3865 1135
rect 3885 1115 3900 1135
rect 3850 1085 3900 1115
rect 3850 1065 3865 1085
rect 3885 1065 3900 1085
rect 3850 1035 3900 1065
rect 3850 1015 3865 1035
rect 3885 1015 3900 1035
rect 3850 1000 3900 1015
rect 4000 1485 4050 1500
rect 4000 1465 4015 1485
rect 4035 1465 4050 1485
rect 4000 1435 4050 1465
rect 4000 1415 4015 1435
rect 4035 1415 4050 1435
rect 4000 1385 4050 1415
rect 4000 1365 4015 1385
rect 4035 1365 4050 1385
rect 4000 1335 4050 1365
rect 4000 1315 4015 1335
rect 4035 1315 4050 1335
rect 4000 1285 4050 1315
rect 4000 1265 4015 1285
rect 4035 1265 4050 1285
rect 4000 1235 4050 1265
rect 4000 1215 4015 1235
rect 4035 1215 4050 1235
rect 4000 1185 4050 1215
rect 4000 1165 4015 1185
rect 4035 1165 4050 1185
rect 4000 1135 4050 1165
rect 4000 1115 4015 1135
rect 4035 1115 4050 1135
rect 4000 1085 4050 1115
rect 4000 1065 4015 1085
rect 4035 1065 4050 1085
rect 4000 1035 4050 1065
rect 4000 1015 4015 1035
rect 4035 1015 4050 1035
rect 3700 965 3715 985
rect 3735 965 3750 985
rect 3700 950 3750 965
rect 4000 985 4050 1015
rect 4000 965 4015 985
rect 4035 965 4050 985
rect 4000 950 4050 965
rect 3700 935 4050 950
rect 3700 915 3715 935
rect 3735 915 4015 935
rect 4035 915 4050 935
rect 3700 900 4050 915
rect 4150 1485 4200 1515
rect 4450 1535 4500 1550
rect 4450 1515 4465 1535
rect 4485 1515 4500 1535
rect 4150 1465 4165 1485
rect 4185 1465 4200 1485
rect 4150 1435 4200 1465
rect 4150 1415 4165 1435
rect 4185 1415 4200 1435
rect 4150 1385 4200 1415
rect 4150 1365 4165 1385
rect 4185 1365 4200 1385
rect 4150 1335 4200 1365
rect 4150 1315 4165 1335
rect 4185 1315 4200 1335
rect 4150 1285 4200 1315
rect 4150 1265 4165 1285
rect 4185 1265 4200 1285
rect 4150 1235 4200 1265
rect 4150 1215 4165 1235
rect 4185 1215 4200 1235
rect 4150 1185 4200 1215
rect 4150 1165 4165 1185
rect 4185 1165 4200 1185
rect 4150 1135 4200 1165
rect 4150 1115 4165 1135
rect 4185 1115 4200 1135
rect 4150 1085 4200 1115
rect 4150 1065 4165 1085
rect 4185 1065 4200 1085
rect 4150 1035 4200 1065
rect 4150 1015 4165 1035
rect 4185 1015 4200 1035
rect 4150 985 4200 1015
rect 4150 965 4165 985
rect 4185 965 4200 985
rect 4150 935 4200 965
rect 4150 915 4165 935
rect 4185 915 4200 935
rect 4150 900 4200 915
rect 4300 1485 4350 1500
rect 4300 1465 4315 1485
rect 4335 1465 4350 1485
rect 4300 1435 4350 1465
rect 4300 1415 4315 1435
rect 4335 1415 4350 1435
rect 4300 1385 4350 1415
rect 4300 1365 4315 1385
rect 4335 1365 4350 1385
rect 4300 1335 4350 1365
rect 4300 1315 4315 1335
rect 4335 1315 4350 1335
rect 4300 1285 4350 1315
rect 4300 1265 4315 1285
rect 4335 1265 4350 1285
rect 4300 1235 4350 1265
rect 4300 1215 4315 1235
rect 4335 1215 4350 1235
rect 4300 1185 4350 1215
rect 4300 1165 4315 1185
rect 4335 1165 4350 1185
rect 4300 1135 4350 1165
rect 4300 1115 4315 1135
rect 4335 1115 4350 1135
rect 4300 1085 4350 1115
rect 4300 1065 4315 1085
rect 4335 1065 4350 1085
rect 4300 1035 4350 1065
rect 4300 1015 4315 1035
rect 4335 1015 4350 1035
rect 4300 985 4350 1015
rect 4450 1485 4500 1515
rect 4750 1535 4800 1550
rect 4750 1515 4765 1535
rect 4785 1515 4800 1535
rect 4450 1465 4465 1485
rect 4485 1465 4500 1485
rect 4450 1435 4500 1465
rect 4450 1415 4465 1435
rect 4485 1415 4500 1435
rect 4450 1385 4500 1415
rect 4450 1365 4465 1385
rect 4485 1365 4500 1385
rect 4450 1335 4500 1365
rect 4450 1315 4465 1335
rect 4485 1315 4500 1335
rect 4450 1285 4500 1315
rect 4450 1265 4465 1285
rect 4485 1265 4500 1285
rect 4450 1235 4500 1265
rect 4450 1215 4465 1235
rect 4485 1215 4500 1235
rect 4450 1185 4500 1215
rect 4450 1165 4465 1185
rect 4485 1165 4500 1185
rect 4450 1135 4500 1165
rect 4450 1115 4465 1135
rect 4485 1115 4500 1135
rect 4450 1085 4500 1115
rect 4450 1065 4465 1085
rect 4485 1065 4500 1085
rect 4450 1035 4500 1065
rect 4450 1015 4465 1035
rect 4485 1015 4500 1035
rect 4450 1000 4500 1015
rect 4600 1485 4650 1500
rect 4600 1465 4615 1485
rect 4635 1465 4650 1485
rect 4600 1435 4650 1465
rect 4600 1415 4615 1435
rect 4635 1415 4650 1435
rect 4600 1385 4650 1415
rect 4600 1365 4615 1385
rect 4635 1365 4650 1385
rect 4600 1335 4650 1365
rect 4600 1315 4615 1335
rect 4635 1315 4650 1335
rect 4600 1285 4650 1315
rect 4600 1265 4615 1285
rect 4635 1265 4650 1285
rect 4600 1235 4650 1265
rect 4600 1215 4615 1235
rect 4635 1215 4650 1235
rect 4600 1185 4650 1215
rect 4600 1165 4615 1185
rect 4635 1165 4650 1185
rect 4600 1135 4650 1165
rect 4600 1115 4615 1135
rect 4635 1115 4650 1135
rect 4600 1085 4650 1115
rect 4600 1065 4615 1085
rect 4635 1065 4650 1085
rect 4600 1035 4650 1065
rect 4600 1015 4615 1035
rect 4635 1015 4650 1035
rect 4300 965 4315 985
rect 4335 965 4350 985
rect 4300 950 4350 965
rect 4600 985 4650 1015
rect 4600 965 4615 985
rect 4635 965 4650 985
rect 4600 950 4650 965
rect 4300 935 4650 950
rect 4300 915 4315 935
rect 4335 915 4615 935
rect 4635 915 4650 935
rect 4300 900 4650 915
rect 4750 1485 4800 1515
rect 5350 1535 5400 1550
rect 5350 1515 5365 1535
rect 5385 1515 5400 1535
rect 4750 1465 4765 1485
rect 4785 1465 4800 1485
rect 4750 1435 4800 1465
rect 4750 1415 4765 1435
rect 4785 1415 4800 1435
rect 4750 1385 4800 1415
rect 4750 1365 4765 1385
rect 4785 1365 4800 1385
rect 4750 1335 4800 1365
rect 4750 1315 4765 1335
rect 4785 1315 4800 1335
rect 4750 1285 4800 1315
rect 4750 1265 4765 1285
rect 4785 1265 4800 1285
rect 4750 1235 4800 1265
rect 4750 1215 4765 1235
rect 4785 1215 4800 1235
rect 4750 1185 4800 1215
rect 4750 1165 4765 1185
rect 4785 1165 4800 1185
rect 4750 1135 4800 1165
rect 4750 1115 4765 1135
rect 4785 1115 4800 1135
rect 4750 1085 4800 1115
rect 4750 1065 4765 1085
rect 4785 1065 4800 1085
rect 4750 1035 4800 1065
rect 4750 1015 4765 1035
rect 4785 1015 4800 1035
rect 4750 985 4800 1015
rect 4750 965 4765 985
rect 4785 965 4800 985
rect 4750 935 4800 965
rect 4750 915 4765 935
rect 4785 915 4800 935
rect 4750 900 4800 915
rect 5050 1485 5100 1500
rect 5050 1465 5065 1485
rect 5085 1465 5100 1485
rect 5050 1435 5100 1465
rect 5050 1415 5065 1435
rect 5085 1415 5100 1435
rect 5050 1385 5100 1415
rect 5050 1365 5065 1385
rect 5085 1365 5100 1385
rect 5050 1335 5100 1365
rect 5050 1315 5065 1335
rect 5085 1315 5100 1335
rect 5050 1285 5100 1315
rect 5050 1265 5065 1285
rect 5085 1265 5100 1285
rect 5050 1235 5100 1265
rect 5050 1215 5065 1235
rect 5085 1215 5100 1235
rect 5050 1185 5100 1215
rect 5050 1165 5065 1185
rect 5085 1165 5100 1185
rect 5050 1135 5100 1165
rect 5050 1115 5065 1135
rect 5085 1115 5100 1135
rect 5050 1085 5100 1115
rect 5050 1065 5065 1085
rect 5085 1065 5100 1085
rect 5050 1035 5100 1065
rect 5050 1015 5065 1035
rect 5085 1015 5100 1035
rect 5050 985 5100 1015
rect 5350 1485 5400 1515
rect 5950 1535 6000 1550
rect 5950 1515 5965 1535
rect 5985 1515 6000 1535
rect 5350 1465 5365 1485
rect 5385 1465 5400 1485
rect 5350 1435 5400 1465
rect 5350 1415 5365 1435
rect 5385 1415 5400 1435
rect 5350 1385 5400 1415
rect 5350 1365 5365 1385
rect 5385 1365 5400 1385
rect 5350 1335 5400 1365
rect 5350 1315 5365 1335
rect 5385 1315 5400 1335
rect 5350 1285 5400 1315
rect 5350 1265 5365 1285
rect 5385 1265 5400 1285
rect 5350 1235 5400 1265
rect 5350 1215 5365 1235
rect 5385 1215 5400 1235
rect 5350 1185 5400 1215
rect 5350 1165 5365 1185
rect 5385 1165 5400 1185
rect 5350 1135 5400 1165
rect 5350 1115 5365 1135
rect 5385 1115 5400 1135
rect 5350 1085 5400 1115
rect 5350 1065 5365 1085
rect 5385 1065 5400 1085
rect 5350 1035 5400 1065
rect 5350 1015 5365 1035
rect 5385 1015 5400 1035
rect 5350 1000 5400 1015
rect 5650 1485 5700 1500
rect 5650 1465 5665 1485
rect 5685 1465 5700 1485
rect 5650 1435 5700 1465
rect 5650 1415 5665 1435
rect 5685 1415 5700 1435
rect 5650 1385 5700 1415
rect 5650 1365 5665 1385
rect 5685 1365 5700 1385
rect 5650 1335 5700 1365
rect 5650 1315 5665 1335
rect 5685 1315 5700 1335
rect 5650 1285 5700 1315
rect 5650 1265 5665 1285
rect 5685 1265 5700 1285
rect 5650 1235 5700 1265
rect 5650 1215 5665 1235
rect 5685 1215 5700 1235
rect 5650 1185 5700 1215
rect 5650 1165 5665 1185
rect 5685 1165 5700 1185
rect 5650 1135 5700 1165
rect 5650 1115 5665 1135
rect 5685 1115 5700 1135
rect 5650 1085 5700 1115
rect 5650 1065 5665 1085
rect 5685 1065 5700 1085
rect 5650 1035 5700 1065
rect 5650 1015 5665 1035
rect 5685 1015 5700 1035
rect 5050 965 5065 985
rect 5085 965 5100 985
rect 5050 950 5100 965
rect 5650 985 5700 1015
rect 5950 1485 6000 1515
rect 6550 1535 6600 1550
rect 6550 1515 6565 1535
rect 6585 1515 6600 1535
rect 5950 1465 5965 1485
rect 5985 1465 6000 1485
rect 5950 1435 6000 1465
rect 5950 1415 5965 1435
rect 5985 1415 6000 1435
rect 5950 1385 6000 1415
rect 5950 1365 5965 1385
rect 5985 1365 6000 1385
rect 5950 1335 6000 1365
rect 5950 1315 5965 1335
rect 5985 1315 6000 1335
rect 5950 1285 6000 1315
rect 5950 1265 5965 1285
rect 5985 1265 6000 1285
rect 5950 1235 6000 1265
rect 5950 1215 5965 1235
rect 5985 1215 6000 1235
rect 5950 1185 6000 1215
rect 5950 1165 5965 1185
rect 5985 1165 6000 1185
rect 5950 1135 6000 1165
rect 5950 1115 5965 1135
rect 5985 1115 6000 1135
rect 5950 1085 6000 1115
rect 5950 1065 5965 1085
rect 5985 1065 6000 1085
rect 5950 1035 6000 1065
rect 5950 1015 5965 1035
rect 5985 1015 6000 1035
rect 5950 1000 6000 1015
rect 6250 1485 6300 1500
rect 6250 1465 6265 1485
rect 6285 1465 6300 1485
rect 6250 1435 6300 1465
rect 6250 1415 6265 1435
rect 6285 1415 6300 1435
rect 6250 1385 6300 1415
rect 6250 1365 6265 1385
rect 6285 1365 6300 1385
rect 6250 1335 6300 1365
rect 6250 1315 6265 1335
rect 6285 1315 6300 1335
rect 6250 1285 6300 1315
rect 6250 1265 6265 1285
rect 6285 1265 6300 1285
rect 6250 1235 6300 1265
rect 6250 1215 6265 1235
rect 6285 1215 6300 1235
rect 6250 1185 6300 1215
rect 6250 1165 6265 1185
rect 6285 1165 6300 1185
rect 6250 1135 6300 1165
rect 6250 1115 6265 1135
rect 6285 1115 6300 1135
rect 6250 1085 6300 1115
rect 6250 1065 6265 1085
rect 6285 1065 6300 1085
rect 6250 1035 6300 1065
rect 6250 1015 6265 1035
rect 6285 1015 6300 1035
rect 5650 965 5665 985
rect 5685 965 5700 985
rect 5650 950 5700 965
rect 6250 985 6300 1015
rect 6550 1485 6600 1515
rect 7150 1535 7200 1550
rect 7150 1515 7165 1535
rect 7185 1515 7200 1535
rect 6550 1465 6565 1485
rect 6585 1465 6600 1485
rect 6550 1435 6600 1465
rect 6550 1415 6565 1435
rect 6585 1415 6600 1435
rect 6550 1385 6600 1415
rect 6550 1365 6565 1385
rect 6585 1365 6600 1385
rect 6550 1335 6600 1365
rect 6550 1315 6565 1335
rect 6585 1315 6600 1335
rect 6550 1285 6600 1315
rect 6550 1265 6565 1285
rect 6585 1265 6600 1285
rect 6550 1235 6600 1265
rect 6550 1215 6565 1235
rect 6585 1215 6600 1235
rect 6550 1185 6600 1215
rect 6550 1165 6565 1185
rect 6585 1165 6600 1185
rect 6550 1135 6600 1165
rect 6550 1115 6565 1135
rect 6585 1115 6600 1135
rect 6550 1085 6600 1115
rect 6550 1065 6565 1085
rect 6585 1065 6600 1085
rect 6550 1035 6600 1065
rect 6550 1015 6565 1035
rect 6585 1015 6600 1035
rect 6550 1000 6600 1015
rect 6850 1485 6900 1500
rect 6850 1465 6865 1485
rect 6885 1465 6900 1485
rect 6850 1435 6900 1465
rect 6850 1415 6865 1435
rect 6885 1415 6900 1435
rect 6850 1385 6900 1415
rect 6850 1365 6865 1385
rect 6885 1365 6900 1385
rect 6850 1335 6900 1365
rect 6850 1315 6865 1335
rect 6885 1315 6900 1335
rect 6850 1285 6900 1315
rect 6850 1265 6865 1285
rect 6885 1265 6900 1285
rect 6850 1235 6900 1265
rect 6850 1215 6865 1235
rect 6885 1215 6900 1235
rect 6850 1185 6900 1215
rect 6850 1165 6865 1185
rect 6885 1165 6900 1185
rect 6850 1135 6900 1165
rect 6850 1115 6865 1135
rect 6885 1115 6900 1135
rect 6850 1085 6900 1115
rect 6850 1065 6865 1085
rect 6885 1065 6900 1085
rect 6850 1035 6900 1065
rect 6850 1015 6865 1035
rect 6885 1015 6900 1035
rect 6250 965 6265 985
rect 6285 965 6300 985
rect 6250 950 6300 965
rect 6850 985 6900 1015
rect 6850 965 6865 985
rect 6885 965 6900 985
rect 6850 950 6900 965
rect 5050 935 6900 950
rect 5050 915 5065 935
rect 5085 915 5665 935
rect 5685 915 6265 935
rect 6285 915 6865 935
rect 6885 915 6900 935
rect 5050 900 6900 915
rect 7150 1485 7200 1515
rect 7150 1465 7165 1485
rect 7185 1465 7200 1485
rect 7150 1435 7200 1465
rect 7150 1415 7165 1435
rect 7185 1415 7200 1435
rect 7150 1385 7200 1415
rect 7150 1365 7165 1385
rect 7185 1365 7200 1385
rect 7150 1335 7200 1365
rect 7150 1315 7165 1335
rect 7185 1315 7200 1335
rect 7150 1285 7200 1315
rect 7150 1265 7165 1285
rect 7185 1265 7200 1285
rect 7150 1235 7200 1265
rect 7150 1215 7165 1235
rect 7185 1215 7200 1235
rect 7150 1185 7200 1215
rect 7150 1165 7165 1185
rect 7185 1165 7200 1185
rect 7150 1135 7200 1165
rect 7150 1115 7165 1135
rect 7185 1115 7200 1135
rect 7150 1085 7200 1115
rect 7150 1065 7165 1085
rect 7185 1065 7200 1085
rect 7150 1035 7200 1065
rect 7150 1015 7165 1035
rect 7185 1015 7200 1035
rect 7150 985 7200 1015
rect 7150 965 7165 985
rect 7185 965 7200 985
rect 7150 935 7200 965
rect 7150 915 7165 935
rect 7185 915 7200 935
rect 7150 900 7200 915
rect 8350 1585 8400 1660
rect 10750 1690 10800 1700
rect 10750 1660 10760 1690
rect 10790 1660 10800 1690
rect 8350 1565 8365 1585
rect 8385 1565 8400 1585
rect 8350 1540 8400 1565
rect 8350 1510 8360 1540
rect 8390 1510 8400 1540
rect 8350 1485 8400 1510
rect 8350 1465 8365 1485
rect 8385 1465 8400 1485
rect 8350 1440 8400 1465
rect 8350 1410 8360 1440
rect 8390 1410 8400 1440
rect 8350 1385 8400 1410
rect 8350 1365 8365 1385
rect 8385 1365 8400 1385
rect 8350 1340 8400 1365
rect 8350 1310 8360 1340
rect 8390 1310 8400 1340
rect 8350 1285 8400 1310
rect 8350 1265 8365 1285
rect 8385 1265 8400 1285
rect 8350 1240 8400 1265
rect 8350 1210 8360 1240
rect 8390 1210 8400 1240
rect 8350 1185 8400 1210
rect 8350 1165 8365 1185
rect 8385 1165 8400 1185
rect 8350 1140 8400 1165
rect 8350 1110 8360 1140
rect 8390 1110 8400 1140
rect 8350 1085 8400 1110
rect 8350 1065 8365 1085
rect 8385 1065 8400 1085
rect 8350 1040 8400 1065
rect 8350 1010 8360 1040
rect 8390 1010 8400 1040
rect 8350 985 8400 1010
rect 8350 965 8365 985
rect 8385 965 8400 985
rect 8350 940 8400 965
rect 8350 910 8360 940
rect 8390 910 8400 940
rect 100 840 150 850
rect 100 810 110 840
rect 140 810 150 840
rect 100 800 150 810
rect 400 840 450 850
rect 400 810 410 840
rect 440 810 450 840
rect 400 800 450 810
rect 700 840 750 850
rect 700 810 710 840
rect 740 810 750 840
rect 700 800 750 810
rect 1000 840 1050 850
rect 1000 810 1010 840
rect 1040 810 1050 840
rect 1000 800 1050 810
rect 1300 840 1350 850
rect 1300 810 1310 840
rect 1340 810 1350 840
rect 1300 800 1350 810
rect 1600 840 1650 850
rect 1600 810 1610 840
rect 1640 810 1650 840
rect 1600 800 1650 810
rect 1900 840 1950 850
rect 1900 810 1910 840
rect 1940 810 1950 840
rect 1900 800 1950 810
rect 2200 840 2250 850
rect 2200 810 2210 840
rect 2240 810 2250 840
rect 2200 800 2250 810
rect 2350 840 2400 900
rect 2350 810 2360 840
rect 2390 810 2400 840
rect 2350 750 2400 810
rect 2500 840 2550 850
rect 2500 810 2510 840
rect 2540 810 2550 840
rect 2500 800 2550 810
rect 2800 840 2850 850
rect 2800 810 2810 840
rect 2840 810 2850 840
rect 2800 800 2850 810
rect 3100 840 3150 850
rect 3100 810 3110 840
rect 3140 810 3150 840
rect 3100 800 3150 810
rect 3400 840 3450 850
rect 3400 810 3410 840
rect 3440 810 3450 840
rect 3400 800 3450 810
rect 3700 840 3750 850
rect 3700 810 3710 840
rect 3740 810 3750 840
rect 3700 800 3750 810
rect 3850 840 3900 900
rect 3850 810 3860 840
rect 3890 810 3900 840
rect 3850 750 3900 810
rect 4000 840 4050 850
rect 4000 810 4010 840
rect 4040 810 4050 840
rect 4000 800 4050 810
rect 4300 840 4350 850
rect 4300 810 4310 840
rect 4340 810 4350 840
rect 4300 800 4350 810
rect 4450 840 4500 900
rect 4450 810 4460 840
rect 4490 810 4500 840
rect 4450 750 4500 810
rect 4600 840 4650 850
rect 4600 810 4610 840
rect 4640 810 4650 840
rect 4600 800 4650 810
rect 4900 840 4950 850
rect 4900 810 4910 840
rect 4940 810 4950 840
rect 4900 800 4950 810
rect 5200 840 5250 850
rect 5200 810 5210 840
rect 5240 810 5250 840
rect 5200 800 5250 810
rect 5500 840 5550 850
rect 5500 810 5510 840
rect 5540 810 5550 840
rect 5500 800 5550 810
rect 5800 840 5850 850
rect 5800 810 5810 840
rect 5840 810 5850 840
rect 5800 800 5850 810
rect 5950 840 6000 900
rect 5950 810 5960 840
rect 5990 810 6000 840
rect 5950 750 6000 810
rect 6100 840 6150 850
rect 6100 810 6110 840
rect 6140 810 6150 840
rect 6100 800 6150 810
rect 6400 840 6450 850
rect 6400 810 6410 840
rect 6440 810 6450 840
rect 6400 800 6450 810
rect 6700 840 6750 850
rect 6700 810 6710 840
rect 6740 810 6750 840
rect 6700 800 6750 810
rect 7000 840 7050 850
rect 7000 810 7010 840
rect 7040 810 7050 840
rect 7000 800 7050 810
rect 7300 840 7350 850
rect 7300 810 7310 840
rect 7340 810 7350 840
rect 7300 800 7350 810
rect 7600 840 7650 850
rect 7600 810 7610 840
rect 7640 810 7650 840
rect 7600 800 7650 810
rect 7900 840 7950 850
rect 7900 810 7910 840
rect 7940 810 7950 840
rect 7900 800 7950 810
rect 8200 840 8250 850
rect 8200 810 8210 840
rect 8240 810 8250 840
rect 8200 800 8250 810
rect -50 710 -40 740
rect -10 710 0 740
rect -50 685 0 710
rect -50 665 -35 685
rect -15 665 0 685
rect -50 640 0 665
rect -50 610 -40 640
rect -10 610 0 640
rect -50 585 0 610
rect -50 565 -35 585
rect -15 565 0 585
rect -50 540 0 565
rect -50 510 -40 540
rect -10 510 0 540
rect -50 485 0 510
rect -50 465 -35 485
rect -15 465 0 485
rect -50 440 0 465
rect -50 410 -40 440
rect -10 410 0 440
rect -50 385 0 410
rect -50 365 -35 385
rect -15 365 0 385
rect -50 340 0 365
rect -50 310 -40 340
rect -10 310 0 340
rect -50 285 0 310
rect -50 265 -35 285
rect -15 265 0 285
rect -50 240 0 265
rect -50 210 -40 240
rect -10 210 0 240
rect -50 185 0 210
rect -50 165 -35 185
rect -15 165 0 185
rect -50 140 0 165
rect -50 110 -40 140
rect -10 110 0 140
rect -50 85 0 110
rect -50 65 -35 85
rect -15 65 0 85
rect -650 -40 -640 -10
rect -610 -40 -600 -10
rect -650 -115 -600 -40
rect -50 -10 0 65
rect 1150 735 1200 750
rect 1150 715 1165 735
rect 1185 715 1200 735
rect 1150 685 1200 715
rect 1150 665 1165 685
rect 1185 665 1200 685
rect 1150 635 1200 665
rect 1150 615 1165 635
rect 1185 615 1200 635
rect 1150 585 1200 615
rect 1150 565 1165 585
rect 1185 565 1200 585
rect 1150 535 1200 565
rect 1150 515 1165 535
rect 1185 515 1200 535
rect 1150 485 1200 515
rect 1150 465 1165 485
rect 1185 465 1200 485
rect 1150 435 1200 465
rect 1150 415 1165 435
rect 1185 415 1200 435
rect 1150 385 1200 415
rect 1150 365 1165 385
rect 1185 365 1200 385
rect 1150 335 1200 365
rect 1150 315 1165 335
rect 1185 315 1200 335
rect 1150 285 1200 315
rect 1150 265 1165 285
rect 1185 265 1200 285
rect 1150 235 1200 265
rect 1150 215 1165 235
rect 1185 215 1200 235
rect 1150 185 1200 215
rect 1150 165 1165 185
rect 1185 165 1200 185
rect 1150 135 1200 165
rect 1450 735 3300 750
rect 1450 715 1465 735
rect 1485 715 2065 735
rect 2085 715 2665 735
rect 2685 715 3265 735
rect 3285 715 3300 735
rect 1450 700 3300 715
rect 1450 685 1500 700
rect 1450 665 1465 685
rect 1485 665 1500 685
rect 1450 635 1500 665
rect 2050 685 2100 700
rect 2050 665 2065 685
rect 2085 665 2100 685
rect 1450 615 1465 635
rect 1485 615 1500 635
rect 1450 585 1500 615
rect 1450 565 1465 585
rect 1485 565 1500 585
rect 1450 535 1500 565
rect 1450 515 1465 535
rect 1485 515 1500 535
rect 1450 485 1500 515
rect 1450 465 1465 485
rect 1485 465 1500 485
rect 1450 435 1500 465
rect 1450 415 1465 435
rect 1485 415 1500 435
rect 1450 385 1500 415
rect 1450 365 1465 385
rect 1485 365 1500 385
rect 1450 335 1500 365
rect 1450 315 1465 335
rect 1485 315 1500 335
rect 1450 285 1500 315
rect 1450 265 1465 285
rect 1485 265 1500 285
rect 1450 235 1500 265
rect 1450 215 1465 235
rect 1485 215 1500 235
rect 1450 185 1500 215
rect 1450 165 1465 185
rect 1485 165 1500 185
rect 1450 150 1500 165
rect 1750 635 1800 650
rect 1750 615 1765 635
rect 1785 615 1800 635
rect 1750 585 1800 615
rect 1750 565 1765 585
rect 1785 565 1800 585
rect 1750 535 1800 565
rect 1750 515 1765 535
rect 1785 515 1800 535
rect 1750 485 1800 515
rect 1750 465 1765 485
rect 1785 465 1800 485
rect 1750 435 1800 465
rect 1750 415 1765 435
rect 1785 415 1800 435
rect 1750 385 1800 415
rect 1750 365 1765 385
rect 1785 365 1800 385
rect 1750 335 1800 365
rect 1750 315 1765 335
rect 1785 315 1800 335
rect 1750 285 1800 315
rect 1750 265 1765 285
rect 1785 265 1800 285
rect 1750 235 1800 265
rect 1750 215 1765 235
rect 1785 215 1800 235
rect 1750 185 1800 215
rect 1750 165 1765 185
rect 1785 165 1800 185
rect 1150 115 1165 135
rect 1185 115 1200 135
rect 1150 100 1200 115
rect 1750 135 1800 165
rect 2050 635 2100 665
rect 2650 685 2700 700
rect 2650 665 2665 685
rect 2685 665 2700 685
rect 2050 615 2065 635
rect 2085 615 2100 635
rect 2050 585 2100 615
rect 2050 565 2065 585
rect 2085 565 2100 585
rect 2050 535 2100 565
rect 2050 515 2065 535
rect 2085 515 2100 535
rect 2050 485 2100 515
rect 2050 465 2065 485
rect 2085 465 2100 485
rect 2050 435 2100 465
rect 2050 415 2065 435
rect 2085 415 2100 435
rect 2050 385 2100 415
rect 2050 365 2065 385
rect 2085 365 2100 385
rect 2050 335 2100 365
rect 2050 315 2065 335
rect 2085 315 2100 335
rect 2050 285 2100 315
rect 2050 265 2065 285
rect 2085 265 2100 285
rect 2050 235 2100 265
rect 2050 215 2065 235
rect 2085 215 2100 235
rect 2050 185 2100 215
rect 2050 165 2065 185
rect 2085 165 2100 185
rect 2050 150 2100 165
rect 2350 635 2400 650
rect 2350 615 2365 635
rect 2385 615 2400 635
rect 2350 585 2400 615
rect 2350 565 2365 585
rect 2385 565 2400 585
rect 2350 535 2400 565
rect 2350 515 2365 535
rect 2385 515 2400 535
rect 2350 485 2400 515
rect 2350 465 2365 485
rect 2385 465 2400 485
rect 2350 435 2400 465
rect 2350 415 2365 435
rect 2385 415 2400 435
rect 2350 385 2400 415
rect 2350 365 2365 385
rect 2385 365 2400 385
rect 2350 335 2400 365
rect 2350 315 2365 335
rect 2385 315 2400 335
rect 2350 285 2400 315
rect 2350 265 2365 285
rect 2385 265 2400 285
rect 2350 235 2400 265
rect 2350 215 2365 235
rect 2385 215 2400 235
rect 2350 185 2400 215
rect 2350 165 2365 185
rect 2385 165 2400 185
rect 1750 115 1765 135
rect 1785 115 1800 135
rect 1750 100 1800 115
rect 2350 135 2400 165
rect 2650 635 2700 665
rect 3250 685 3300 700
rect 3250 665 3265 685
rect 3285 665 3300 685
rect 2650 615 2665 635
rect 2685 615 2700 635
rect 2650 585 2700 615
rect 2650 565 2665 585
rect 2685 565 2700 585
rect 2650 535 2700 565
rect 2650 515 2665 535
rect 2685 515 2700 535
rect 2650 485 2700 515
rect 2650 465 2665 485
rect 2685 465 2700 485
rect 2650 435 2700 465
rect 2650 415 2665 435
rect 2685 415 2700 435
rect 2650 385 2700 415
rect 2650 365 2665 385
rect 2685 365 2700 385
rect 2650 335 2700 365
rect 2650 315 2665 335
rect 2685 315 2700 335
rect 2650 285 2700 315
rect 2650 265 2665 285
rect 2685 265 2700 285
rect 2650 235 2700 265
rect 2650 215 2665 235
rect 2685 215 2700 235
rect 2650 185 2700 215
rect 2650 165 2665 185
rect 2685 165 2700 185
rect 2650 150 2700 165
rect 2950 635 3000 650
rect 2950 615 2965 635
rect 2985 615 3000 635
rect 2950 585 3000 615
rect 2950 565 2965 585
rect 2985 565 3000 585
rect 2950 535 3000 565
rect 2950 515 2965 535
rect 2985 515 3000 535
rect 2950 485 3000 515
rect 2950 465 2965 485
rect 2985 465 3000 485
rect 2950 435 3000 465
rect 2950 415 2965 435
rect 2985 415 3000 435
rect 2950 385 3000 415
rect 2950 365 2965 385
rect 2985 365 3000 385
rect 2950 335 3000 365
rect 2950 315 2965 335
rect 2985 315 3000 335
rect 2950 285 3000 315
rect 2950 265 2965 285
rect 2985 265 3000 285
rect 2950 235 3000 265
rect 2950 215 2965 235
rect 2985 215 3000 235
rect 2950 185 3000 215
rect 2950 165 2965 185
rect 2985 165 3000 185
rect 2350 115 2365 135
rect 2385 115 2400 135
rect 2350 100 2400 115
rect 2950 135 3000 165
rect 3250 635 3300 665
rect 3250 615 3265 635
rect 3285 615 3300 635
rect 3250 585 3300 615
rect 3250 565 3265 585
rect 3285 565 3300 585
rect 3250 535 3300 565
rect 3250 515 3265 535
rect 3285 515 3300 535
rect 3250 485 3300 515
rect 3250 465 3265 485
rect 3285 465 3300 485
rect 3250 435 3300 465
rect 3250 415 3265 435
rect 3285 415 3300 435
rect 3250 385 3300 415
rect 3250 365 3265 385
rect 3285 365 3300 385
rect 3250 335 3300 365
rect 3250 315 3265 335
rect 3285 315 3300 335
rect 3250 285 3300 315
rect 3250 265 3265 285
rect 3285 265 3300 285
rect 3250 235 3300 265
rect 3250 215 3265 235
rect 3285 215 3300 235
rect 3250 185 3300 215
rect 3250 165 3265 185
rect 3285 165 3300 185
rect 3250 150 3300 165
rect 3550 735 3600 750
rect 3550 715 3565 735
rect 3585 715 3600 735
rect 3550 685 3600 715
rect 3550 665 3565 685
rect 3585 665 3600 685
rect 3550 635 3600 665
rect 3550 615 3565 635
rect 3585 615 3600 635
rect 3550 585 3600 615
rect 3550 565 3565 585
rect 3585 565 3600 585
rect 3550 535 3600 565
rect 3550 515 3565 535
rect 3585 515 3600 535
rect 3550 485 3600 515
rect 3550 465 3565 485
rect 3585 465 3600 485
rect 3550 435 3600 465
rect 3550 415 3565 435
rect 3585 415 3600 435
rect 3550 385 3600 415
rect 3550 365 3565 385
rect 3585 365 3600 385
rect 3550 335 3600 365
rect 3550 315 3565 335
rect 3585 315 3600 335
rect 3550 285 3600 315
rect 3550 265 3565 285
rect 3585 265 3600 285
rect 3550 235 3600 265
rect 3550 215 3565 235
rect 3585 215 3600 235
rect 3550 185 3600 215
rect 3550 165 3565 185
rect 3585 165 3600 185
rect 2950 115 2965 135
rect 2985 115 3000 135
rect 2950 100 3000 115
rect 3550 135 3600 165
rect 3700 735 4050 750
rect 3700 715 3715 735
rect 3735 715 4015 735
rect 4035 715 4050 735
rect 3700 700 4050 715
rect 3700 685 3750 700
rect 3700 665 3715 685
rect 3735 665 3750 685
rect 3700 635 3750 665
rect 4000 685 4050 700
rect 4000 665 4015 685
rect 4035 665 4050 685
rect 3700 615 3715 635
rect 3735 615 3750 635
rect 3700 585 3750 615
rect 3700 565 3715 585
rect 3735 565 3750 585
rect 3700 535 3750 565
rect 3700 515 3715 535
rect 3735 515 3750 535
rect 3700 485 3750 515
rect 3700 465 3715 485
rect 3735 465 3750 485
rect 3700 435 3750 465
rect 3700 415 3715 435
rect 3735 415 3750 435
rect 3700 385 3750 415
rect 3700 365 3715 385
rect 3735 365 3750 385
rect 3700 335 3750 365
rect 3700 315 3715 335
rect 3735 315 3750 335
rect 3700 285 3750 315
rect 3700 265 3715 285
rect 3735 265 3750 285
rect 3700 235 3750 265
rect 3700 215 3715 235
rect 3735 215 3750 235
rect 3700 185 3750 215
rect 3700 165 3715 185
rect 3735 165 3750 185
rect 3700 150 3750 165
rect 3850 635 3900 650
rect 3850 615 3865 635
rect 3885 615 3900 635
rect 3850 585 3900 615
rect 3850 565 3865 585
rect 3885 565 3900 585
rect 3850 535 3900 565
rect 3850 515 3865 535
rect 3885 515 3900 535
rect 3850 485 3900 515
rect 3850 465 3865 485
rect 3885 465 3900 485
rect 3850 435 3900 465
rect 3850 415 3865 435
rect 3885 415 3900 435
rect 3850 385 3900 415
rect 3850 365 3865 385
rect 3885 365 3900 385
rect 3850 335 3900 365
rect 3850 315 3865 335
rect 3885 315 3900 335
rect 3850 285 3900 315
rect 3850 265 3865 285
rect 3885 265 3900 285
rect 3850 235 3900 265
rect 3850 215 3865 235
rect 3885 215 3900 235
rect 3850 185 3900 215
rect 3850 165 3865 185
rect 3885 165 3900 185
rect 3550 115 3565 135
rect 3585 115 3600 135
rect 3550 100 3600 115
rect 3850 135 3900 165
rect 4000 635 4050 665
rect 4000 615 4015 635
rect 4035 615 4050 635
rect 4000 585 4050 615
rect 4000 565 4015 585
rect 4035 565 4050 585
rect 4000 535 4050 565
rect 4000 515 4015 535
rect 4035 515 4050 535
rect 4000 485 4050 515
rect 4000 465 4015 485
rect 4035 465 4050 485
rect 4000 435 4050 465
rect 4000 415 4015 435
rect 4035 415 4050 435
rect 4000 385 4050 415
rect 4000 365 4015 385
rect 4035 365 4050 385
rect 4000 335 4050 365
rect 4000 315 4015 335
rect 4035 315 4050 335
rect 4000 285 4050 315
rect 4000 265 4015 285
rect 4035 265 4050 285
rect 4000 235 4050 265
rect 4000 215 4015 235
rect 4035 215 4050 235
rect 4000 185 4050 215
rect 4000 165 4015 185
rect 4035 165 4050 185
rect 4000 150 4050 165
rect 4150 735 4200 750
rect 4150 715 4165 735
rect 4185 715 4200 735
rect 4150 685 4200 715
rect 4150 665 4165 685
rect 4185 665 4200 685
rect 4150 635 4200 665
rect 4150 615 4165 635
rect 4185 615 4200 635
rect 4150 585 4200 615
rect 4150 565 4165 585
rect 4185 565 4200 585
rect 4150 535 4200 565
rect 4150 515 4165 535
rect 4185 515 4200 535
rect 4150 485 4200 515
rect 4150 465 4165 485
rect 4185 465 4200 485
rect 4150 435 4200 465
rect 4150 415 4165 435
rect 4185 415 4200 435
rect 4150 385 4200 415
rect 4150 365 4165 385
rect 4185 365 4200 385
rect 4150 335 4200 365
rect 4150 315 4165 335
rect 4185 315 4200 335
rect 4150 285 4200 315
rect 4150 265 4165 285
rect 4185 265 4200 285
rect 4150 235 4200 265
rect 4150 215 4165 235
rect 4185 215 4200 235
rect 4150 185 4200 215
rect 4150 165 4165 185
rect 4185 165 4200 185
rect 3850 115 3865 135
rect 3885 115 3900 135
rect 3850 100 3900 115
rect 4150 135 4200 165
rect 4300 735 4650 750
rect 4300 715 4315 735
rect 4335 715 4615 735
rect 4635 715 4650 735
rect 4300 700 4650 715
rect 4300 685 4350 700
rect 4300 665 4315 685
rect 4335 665 4350 685
rect 4300 635 4350 665
rect 4600 685 4650 700
rect 4600 665 4615 685
rect 4635 665 4650 685
rect 4300 615 4315 635
rect 4335 615 4350 635
rect 4300 585 4350 615
rect 4300 565 4315 585
rect 4335 565 4350 585
rect 4300 535 4350 565
rect 4300 515 4315 535
rect 4335 515 4350 535
rect 4300 485 4350 515
rect 4300 465 4315 485
rect 4335 465 4350 485
rect 4300 435 4350 465
rect 4300 415 4315 435
rect 4335 415 4350 435
rect 4300 385 4350 415
rect 4300 365 4315 385
rect 4335 365 4350 385
rect 4300 335 4350 365
rect 4300 315 4315 335
rect 4335 315 4350 335
rect 4300 285 4350 315
rect 4300 265 4315 285
rect 4335 265 4350 285
rect 4300 235 4350 265
rect 4300 215 4315 235
rect 4335 215 4350 235
rect 4300 185 4350 215
rect 4300 165 4315 185
rect 4335 165 4350 185
rect 4300 150 4350 165
rect 4450 635 4500 650
rect 4450 615 4465 635
rect 4485 615 4500 635
rect 4450 585 4500 615
rect 4450 565 4465 585
rect 4485 565 4500 585
rect 4450 535 4500 565
rect 4450 515 4465 535
rect 4485 515 4500 535
rect 4450 485 4500 515
rect 4450 465 4465 485
rect 4485 465 4500 485
rect 4450 435 4500 465
rect 4450 415 4465 435
rect 4485 415 4500 435
rect 4450 385 4500 415
rect 4450 365 4465 385
rect 4485 365 4500 385
rect 4450 335 4500 365
rect 4450 315 4465 335
rect 4485 315 4500 335
rect 4450 285 4500 315
rect 4450 265 4465 285
rect 4485 265 4500 285
rect 4450 235 4500 265
rect 4450 215 4465 235
rect 4485 215 4500 235
rect 4450 185 4500 215
rect 4450 165 4465 185
rect 4485 165 4500 185
rect 4150 115 4165 135
rect 4185 115 4200 135
rect 4150 100 4200 115
rect 4450 135 4500 165
rect 4600 635 4650 665
rect 4600 615 4615 635
rect 4635 615 4650 635
rect 4600 585 4650 615
rect 4600 565 4615 585
rect 4635 565 4650 585
rect 4600 535 4650 565
rect 4600 515 4615 535
rect 4635 515 4650 535
rect 4600 485 4650 515
rect 4600 465 4615 485
rect 4635 465 4650 485
rect 4600 435 4650 465
rect 4600 415 4615 435
rect 4635 415 4650 435
rect 4600 385 4650 415
rect 4600 365 4615 385
rect 4635 365 4650 385
rect 4600 335 4650 365
rect 4600 315 4615 335
rect 4635 315 4650 335
rect 4600 285 4650 315
rect 4600 265 4615 285
rect 4635 265 4650 285
rect 4600 235 4650 265
rect 4600 215 4615 235
rect 4635 215 4650 235
rect 4600 185 4650 215
rect 4600 165 4615 185
rect 4635 165 4650 185
rect 4600 150 4650 165
rect 4750 735 4800 750
rect 4750 715 4765 735
rect 4785 715 4800 735
rect 4750 685 4800 715
rect 4750 665 4765 685
rect 4785 665 4800 685
rect 4750 635 4800 665
rect 4750 615 4765 635
rect 4785 615 4800 635
rect 4750 585 4800 615
rect 4750 565 4765 585
rect 4785 565 4800 585
rect 4750 535 4800 565
rect 4750 515 4765 535
rect 4785 515 4800 535
rect 4750 485 4800 515
rect 4750 465 4765 485
rect 4785 465 4800 485
rect 4750 435 4800 465
rect 4750 415 4765 435
rect 4785 415 4800 435
rect 4750 385 4800 415
rect 4750 365 4765 385
rect 4785 365 4800 385
rect 4750 335 4800 365
rect 4750 315 4765 335
rect 4785 315 4800 335
rect 4750 285 4800 315
rect 4750 265 4765 285
rect 4785 265 4800 285
rect 4750 235 4800 265
rect 4750 215 4765 235
rect 4785 215 4800 235
rect 4750 185 4800 215
rect 4750 165 4765 185
rect 4785 165 4800 185
rect 4450 115 4465 135
rect 4485 115 4500 135
rect 4450 100 4500 115
rect 4750 135 4800 165
rect 5050 735 6900 750
rect 5050 715 5065 735
rect 5085 715 5665 735
rect 5685 715 6265 735
rect 6285 715 6865 735
rect 6885 715 6900 735
rect 5050 700 6900 715
rect 5050 685 5100 700
rect 5050 665 5065 685
rect 5085 665 5100 685
rect 5050 635 5100 665
rect 5650 685 5700 700
rect 5650 665 5665 685
rect 5685 665 5700 685
rect 5050 615 5065 635
rect 5085 615 5100 635
rect 5050 585 5100 615
rect 5050 565 5065 585
rect 5085 565 5100 585
rect 5050 535 5100 565
rect 5050 515 5065 535
rect 5085 515 5100 535
rect 5050 485 5100 515
rect 5050 465 5065 485
rect 5085 465 5100 485
rect 5050 435 5100 465
rect 5050 415 5065 435
rect 5085 415 5100 435
rect 5050 385 5100 415
rect 5050 365 5065 385
rect 5085 365 5100 385
rect 5050 335 5100 365
rect 5050 315 5065 335
rect 5085 315 5100 335
rect 5050 285 5100 315
rect 5050 265 5065 285
rect 5085 265 5100 285
rect 5050 235 5100 265
rect 5050 215 5065 235
rect 5085 215 5100 235
rect 5050 185 5100 215
rect 5050 165 5065 185
rect 5085 165 5100 185
rect 5050 150 5100 165
rect 5350 635 5400 650
rect 5350 615 5365 635
rect 5385 615 5400 635
rect 5350 585 5400 615
rect 5350 565 5365 585
rect 5385 565 5400 585
rect 5350 535 5400 565
rect 5350 515 5365 535
rect 5385 515 5400 535
rect 5350 485 5400 515
rect 5350 465 5365 485
rect 5385 465 5400 485
rect 5350 435 5400 465
rect 5350 415 5365 435
rect 5385 415 5400 435
rect 5350 385 5400 415
rect 5350 365 5365 385
rect 5385 365 5400 385
rect 5350 335 5400 365
rect 5350 315 5365 335
rect 5385 315 5400 335
rect 5350 285 5400 315
rect 5350 265 5365 285
rect 5385 265 5400 285
rect 5350 235 5400 265
rect 5350 215 5365 235
rect 5385 215 5400 235
rect 5350 185 5400 215
rect 5350 165 5365 185
rect 5385 165 5400 185
rect 4750 115 4765 135
rect 4785 115 4800 135
rect 4750 100 4800 115
rect 5350 135 5400 165
rect 5650 635 5700 665
rect 6250 685 6300 700
rect 6250 665 6265 685
rect 6285 665 6300 685
rect 5650 615 5665 635
rect 5685 615 5700 635
rect 5650 585 5700 615
rect 5650 565 5665 585
rect 5685 565 5700 585
rect 5650 535 5700 565
rect 5650 515 5665 535
rect 5685 515 5700 535
rect 5650 485 5700 515
rect 5650 465 5665 485
rect 5685 465 5700 485
rect 5650 435 5700 465
rect 5650 415 5665 435
rect 5685 415 5700 435
rect 5650 385 5700 415
rect 5650 365 5665 385
rect 5685 365 5700 385
rect 5650 335 5700 365
rect 5650 315 5665 335
rect 5685 315 5700 335
rect 5650 285 5700 315
rect 5650 265 5665 285
rect 5685 265 5700 285
rect 5650 235 5700 265
rect 5650 215 5665 235
rect 5685 215 5700 235
rect 5650 185 5700 215
rect 5650 165 5665 185
rect 5685 165 5700 185
rect 5650 150 5700 165
rect 5950 635 6000 650
rect 5950 615 5965 635
rect 5985 615 6000 635
rect 5950 585 6000 615
rect 5950 565 5965 585
rect 5985 565 6000 585
rect 5950 535 6000 565
rect 5950 515 5965 535
rect 5985 515 6000 535
rect 5950 485 6000 515
rect 5950 465 5965 485
rect 5985 465 6000 485
rect 5950 435 6000 465
rect 5950 415 5965 435
rect 5985 415 6000 435
rect 5950 385 6000 415
rect 5950 365 5965 385
rect 5985 365 6000 385
rect 5950 335 6000 365
rect 5950 315 5965 335
rect 5985 315 6000 335
rect 5950 285 6000 315
rect 5950 265 5965 285
rect 5985 265 6000 285
rect 5950 235 6000 265
rect 5950 215 5965 235
rect 5985 215 6000 235
rect 5950 185 6000 215
rect 5950 165 5965 185
rect 5985 165 6000 185
rect 5350 115 5365 135
rect 5385 115 5400 135
rect 5350 100 5400 115
rect 5950 135 6000 165
rect 6250 635 6300 665
rect 6850 685 6900 700
rect 6850 665 6865 685
rect 6885 665 6900 685
rect 6250 615 6265 635
rect 6285 615 6300 635
rect 6250 585 6300 615
rect 6250 565 6265 585
rect 6285 565 6300 585
rect 6250 535 6300 565
rect 6250 515 6265 535
rect 6285 515 6300 535
rect 6250 485 6300 515
rect 6250 465 6265 485
rect 6285 465 6300 485
rect 6250 435 6300 465
rect 6250 415 6265 435
rect 6285 415 6300 435
rect 6250 385 6300 415
rect 6250 365 6265 385
rect 6285 365 6300 385
rect 6250 335 6300 365
rect 6250 315 6265 335
rect 6285 315 6300 335
rect 6250 285 6300 315
rect 6250 265 6265 285
rect 6285 265 6300 285
rect 6250 235 6300 265
rect 6250 215 6265 235
rect 6285 215 6300 235
rect 6250 185 6300 215
rect 6250 165 6265 185
rect 6285 165 6300 185
rect 6250 150 6300 165
rect 6550 635 6600 650
rect 6550 615 6565 635
rect 6585 615 6600 635
rect 6550 585 6600 615
rect 6550 565 6565 585
rect 6585 565 6600 585
rect 6550 535 6600 565
rect 6550 515 6565 535
rect 6585 515 6600 535
rect 6550 485 6600 515
rect 6550 465 6565 485
rect 6585 465 6600 485
rect 6550 435 6600 465
rect 6550 415 6565 435
rect 6585 415 6600 435
rect 6550 385 6600 415
rect 6550 365 6565 385
rect 6585 365 6600 385
rect 6550 335 6600 365
rect 6550 315 6565 335
rect 6585 315 6600 335
rect 6550 285 6600 315
rect 6550 265 6565 285
rect 6585 265 6600 285
rect 6550 235 6600 265
rect 6550 215 6565 235
rect 6585 215 6600 235
rect 6550 185 6600 215
rect 6550 165 6565 185
rect 6585 165 6600 185
rect 5950 115 5965 135
rect 5985 115 6000 135
rect 5950 100 6000 115
rect 6550 135 6600 165
rect 6850 635 6900 665
rect 6850 615 6865 635
rect 6885 615 6900 635
rect 6850 585 6900 615
rect 6850 565 6865 585
rect 6885 565 6900 585
rect 6850 535 6900 565
rect 6850 515 6865 535
rect 6885 515 6900 535
rect 6850 485 6900 515
rect 6850 465 6865 485
rect 6885 465 6900 485
rect 6850 435 6900 465
rect 6850 415 6865 435
rect 6885 415 6900 435
rect 6850 385 6900 415
rect 6850 365 6865 385
rect 6885 365 6900 385
rect 6850 335 6900 365
rect 6850 315 6865 335
rect 6885 315 6900 335
rect 6850 285 6900 315
rect 6850 265 6865 285
rect 6885 265 6900 285
rect 6850 235 6900 265
rect 6850 215 6865 235
rect 6885 215 6900 235
rect 6850 185 6900 215
rect 6850 165 6865 185
rect 6885 165 6900 185
rect 6850 150 6900 165
rect 7150 735 7200 750
rect 7150 715 7165 735
rect 7185 715 7200 735
rect 7150 685 7200 715
rect 7150 665 7165 685
rect 7185 665 7200 685
rect 7150 635 7200 665
rect 7150 615 7165 635
rect 7185 615 7200 635
rect 7150 585 7200 615
rect 7150 565 7165 585
rect 7185 565 7200 585
rect 7150 535 7200 565
rect 7150 515 7165 535
rect 7185 515 7200 535
rect 7150 485 7200 515
rect 7150 465 7165 485
rect 7185 465 7200 485
rect 7150 435 7200 465
rect 7150 415 7165 435
rect 7185 415 7200 435
rect 7150 385 7200 415
rect 7150 365 7165 385
rect 7185 365 7200 385
rect 7150 335 7200 365
rect 7150 315 7165 335
rect 7185 315 7200 335
rect 7150 285 7200 315
rect 7150 265 7165 285
rect 7185 265 7200 285
rect 7150 235 7200 265
rect 7150 215 7165 235
rect 7185 215 7200 235
rect 7150 185 7200 215
rect 7150 165 7165 185
rect 7185 165 7200 185
rect 6550 115 6565 135
rect 6585 115 6600 135
rect 6550 100 6600 115
rect 7150 135 7200 165
rect 7150 115 7165 135
rect 7185 115 7200 135
rect 7150 100 7200 115
rect 1150 85 7200 100
rect 1150 65 1165 85
rect 1185 65 1765 85
rect 1785 65 2365 85
rect 2385 65 2965 85
rect 2985 65 3565 85
rect 3585 65 3865 85
rect 3885 65 4165 85
rect 4185 65 4465 85
rect 4485 65 4765 85
rect 4785 65 5365 85
rect 5385 65 5965 85
rect 5985 65 6565 85
rect 6585 65 7165 85
rect 7185 65 7200 85
rect 1150 50 7200 65
rect 8350 740 8400 910
rect 9550 1585 9600 1600
rect 9550 1565 9565 1585
rect 9585 1565 9600 1585
rect 9550 1535 9600 1565
rect 9550 1515 9565 1535
rect 9585 1515 9600 1535
rect 9550 1485 9600 1515
rect 9550 1465 9565 1485
rect 9585 1465 9600 1485
rect 9550 1435 9600 1465
rect 9550 1415 9565 1435
rect 9585 1415 9600 1435
rect 9550 1385 9600 1415
rect 9550 1365 9565 1385
rect 9585 1365 9600 1385
rect 9550 1335 9600 1365
rect 9550 1315 9565 1335
rect 9585 1315 9600 1335
rect 9550 1285 9600 1315
rect 9550 1265 9565 1285
rect 9585 1265 9600 1285
rect 9550 1235 9600 1265
rect 9550 1215 9565 1235
rect 9585 1215 9600 1235
rect 9550 1185 9600 1215
rect 9550 1165 9565 1185
rect 9585 1165 9600 1185
rect 9550 1135 9600 1165
rect 9550 1115 9565 1135
rect 9585 1115 9600 1135
rect 9550 1085 9600 1115
rect 9550 1065 9565 1085
rect 9585 1065 9600 1085
rect 9550 1035 9600 1065
rect 9550 1015 9565 1035
rect 9585 1015 9600 1035
rect 9550 985 9600 1015
rect 9550 965 9565 985
rect 9585 965 9600 985
rect 9550 935 9600 965
rect 9550 915 9565 935
rect 9585 915 9600 935
rect 8500 840 8550 850
rect 8500 810 8510 840
rect 8540 810 8550 840
rect 8500 800 8550 810
rect 8800 840 8850 850
rect 8800 810 8810 840
rect 8840 810 8850 840
rect 8800 800 8850 810
rect 9100 840 9150 850
rect 9100 810 9110 840
rect 9140 810 9150 840
rect 9100 800 9150 810
rect 9400 840 9450 850
rect 9400 810 9410 840
rect 9440 810 9450 840
rect 9400 800 9450 810
rect 9550 840 9600 915
rect 10750 1585 10800 1660
rect 15550 1690 15600 1700
rect 15550 1660 15560 1690
rect 15590 1660 15600 1690
rect 10750 1565 10765 1585
rect 10785 1565 10800 1585
rect 10750 1540 10800 1565
rect 10750 1510 10760 1540
rect 10790 1510 10800 1540
rect 10750 1485 10800 1510
rect 10750 1465 10765 1485
rect 10785 1465 10800 1485
rect 10750 1440 10800 1465
rect 10750 1410 10760 1440
rect 10790 1410 10800 1440
rect 10750 1385 10800 1410
rect 10750 1365 10765 1385
rect 10785 1365 10800 1385
rect 10750 1340 10800 1365
rect 10750 1310 10760 1340
rect 10790 1310 10800 1340
rect 10750 1285 10800 1310
rect 10750 1265 10765 1285
rect 10785 1265 10800 1285
rect 10750 1240 10800 1265
rect 10750 1210 10760 1240
rect 10790 1210 10800 1240
rect 10750 1185 10800 1210
rect 10750 1165 10765 1185
rect 10785 1165 10800 1185
rect 10750 1140 10800 1165
rect 10750 1110 10760 1140
rect 10790 1110 10800 1140
rect 10750 1085 10800 1110
rect 10750 1065 10765 1085
rect 10785 1065 10800 1085
rect 10750 1040 10800 1065
rect 10750 1010 10760 1040
rect 10790 1010 10800 1040
rect 10750 985 10800 1010
rect 10750 965 10765 985
rect 10785 965 10800 985
rect 10750 940 10800 965
rect 10750 910 10760 940
rect 10790 910 10800 940
rect 9550 810 9560 840
rect 9590 810 9600 840
rect 8350 710 8360 740
rect 8390 710 8400 740
rect 8350 685 8400 710
rect 8350 665 8365 685
rect 8385 665 8400 685
rect 8350 640 8400 665
rect 8350 610 8360 640
rect 8390 610 8400 640
rect 8350 585 8400 610
rect 8350 565 8365 585
rect 8385 565 8400 585
rect 8350 540 8400 565
rect 8350 510 8360 540
rect 8390 510 8400 540
rect 8350 485 8400 510
rect 8350 465 8365 485
rect 8385 465 8400 485
rect 8350 440 8400 465
rect 8350 410 8360 440
rect 8390 410 8400 440
rect 8350 385 8400 410
rect 8350 365 8365 385
rect 8385 365 8400 385
rect 8350 340 8400 365
rect 8350 310 8360 340
rect 8390 310 8400 340
rect 8350 285 8400 310
rect 8350 265 8365 285
rect 8385 265 8400 285
rect 8350 240 8400 265
rect 8350 210 8360 240
rect 8390 210 8400 240
rect 8350 185 8400 210
rect 8350 165 8365 185
rect 8385 165 8400 185
rect 8350 140 8400 165
rect 8350 110 8360 140
rect 8390 110 8400 140
rect 8350 85 8400 110
rect 8350 65 8365 85
rect 8385 65 8400 85
rect -50 -40 -40 -10
rect -10 -40 0 -10
rect -650 -135 -635 -115
rect -615 -135 -600 -115
rect -650 -160 -600 -135
rect -650 -190 -640 -160
rect -610 -190 -600 -160
rect -650 -215 -600 -190
rect -650 -235 -635 -215
rect -615 -235 -600 -215
rect -650 -260 -600 -235
rect -650 -290 -640 -260
rect -610 -290 -600 -260
rect -650 -315 -600 -290
rect -650 -335 -635 -315
rect -615 -335 -600 -315
rect -650 -360 -600 -335
rect -650 -390 -640 -360
rect -610 -390 -600 -360
rect -650 -415 -600 -390
rect -650 -435 -635 -415
rect -615 -435 -600 -415
rect -650 -460 -600 -435
rect -650 -490 -640 -460
rect -610 -490 -600 -460
rect -650 -515 -600 -490
rect -650 -535 -635 -515
rect -615 -535 -600 -515
rect -650 -560 -600 -535
rect -650 -590 -640 -560
rect -610 -590 -600 -560
rect -650 -615 -600 -590
rect -650 -635 -635 -615
rect -615 -635 -600 -615
rect -650 -660 -600 -635
rect -650 -690 -640 -660
rect -610 -690 -600 -660
rect -650 -715 -600 -690
rect -650 -735 -635 -715
rect -615 -735 -600 -715
rect -650 -760 -600 -735
rect -650 -790 -640 -760
rect -610 -790 -600 -760
rect -650 -960 -600 -790
rect -500 -115 -450 -100
rect -500 -135 -485 -115
rect -465 -135 -450 -115
rect -500 -165 -450 -135
rect -500 -185 -485 -165
rect -465 -185 -450 -165
rect -500 -215 -450 -185
rect -500 -235 -485 -215
rect -465 -235 -450 -215
rect -500 -265 -450 -235
rect -500 -285 -485 -265
rect -465 -285 -450 -265
rect -500 -315 -450 -285
rect -500 -335 -485 -315
rect -465 -335 -450 -315
rect -500 -365 -450 -335
rect -500 -385 -485 -365
rect -465 -385 -450 -365
rect -500 -415 -450 -385
rect -500 -435 -485 -415
rect -465 -435 -450 -415
rect -500 -465 -450 -435
rect -500 -485 -485 -465
rect -465 -485 -450 -465
rect -500 -515 -450 -485
rect -500 -535 -485 -515
rect -465 -535 -450 -515
rect -500 -565 -450 -535
rect -500 -585 -485 -565
rect -465 -585 -450 -565
rect -500 -615 -450 -585
rect -500 -635 -485 -615
rect -465 -635 -450 -615
rect -500 -665 -450 -635
rect -500 -685 -485 -665
rect -465 -685 -450 -665
rect -500 -715 -450 -685
rect -500 -735 -485 -715
rect -465 -735 -450 -715
rect -500 -765 -450 -735
rect -500 -785 -485 -765
rect -465 -785 -450 -765
rect -500 -800 -450 -785
rect -350 -115 -300 -100
rect -350 -135 -335 -115
rect -315 -135 -300 -115
rect -350 -165 -300 -135
rect -350 -185 -335 -165
rect -315 -185 -300 -165
rect -350 -215 -300 -185
rect -350 -235 -335 -215
rect -315 -235 -300 -215
rect -350 -265 -300 -235
rect -350 -285 -335 -265
rect -315 -285 -300 -265
rect -350 -315 -300 -285
rect -350 -335 -335 -315
rect -315 -335 -300 -315
rect -350 -365 -300 -335
rect -350 -385 -335 -365
rect -315 -385 -300 -365
rect -350 -415 -300 -385
rect -350 -435 -335 -415
rect -315 -435 -300 -415
rect -350 -465 -300 -435
rect -350 -485 -335 -465
rect -315 -485 -300 -465
rect -350 -515 -300 -485
rect -350 -535 -335 -515
rect -315 -535 -300 -515
rect -350 -565 -300 -535
rect -350 -585 -335 -565
rect -315 -585 -300 -565
rect -350 -615 -300 -585
rect -350 -635 -335 -615
rect -315 -635 -300 -615
rect -350 -665 -300 -635
rect -350 -685 -335 -665
rect -315 -685 -300 -665
rect -350 -715 -300 -685
rect -350 -735 -335 -715
rect -315 -735 -300 -715
rect -350 -765 -300 -735
rect -350 -785 -335 -765
rect -315 -785 -300 -765
rect -500 -860 -450 -850
rect -500 -890 -490 -860
rect -460 -890 -450 -860
rect -500 -900 -450 -890
rect -350 -860 -300 -785
rect -200 -115 -150 -100
rect -200 -135 -185 -115
rect -165 -135 -150 -115
rect -200 -165 -150 -135
rect -200 -185 -185 -165
rect -165 -185 -150 -165
rect -200 -215 -150 -185
rect -200 -235 -185 -215
rect -165 -235 -150 -215
rect -200 -265 -150 -235
rect -200 -285 -185 -265
rect -165 -285 -150 -265
rect -200 -315 -150 -285
rect -200 -335 -185 -315
rect -165 -335 -150 -315
rect -200 -365 -150 -335
rect -200 -385 -185 -365
rect -165 -385 -150 -365
rect -200 -415 -150 -385
rect -200 -435 -185 -415
rect -165 -435 -150 -415
rect -200 -465 -150 -435
rect -200 -485 -185 -465
rect -165 -485 -150 -465
rect -200 -515 -150 -485
rect -200 -535 -185 -515
rect -165 -535 -150 -515
rect -200 -565 -150 -535
rect -200 -585 -185 -565
rect -165 -585 -150 -565
rect -200 -615 -150 -585
rect -200 -635 -185 -615
rect -165 -635 -150 -615
rect -200 -665 -150 -635
rect -200 -685 -185 -665
rect -165 -685 -150 -665
rect -200 -715 -150 -685
rect -200 -735 -185 -715
rect -165 -735 -150 -715
rect -200 -765 -150 -735
rect -200 -785 -185 -765
rect -165 -785 -150 -765
rect -200 -800 -150 -785
rect -50 -115 0 -40
rect 8350 -10 8400 65
rect 9550 735 9600 810
rect 9700 840 9750 850
rect 9700 810 9710 840
rect 9740 810 9750 840
rect 9700 800 9750 810
rect 10000 840 10050 850
rect 10000 810 10010 840
rect 10040 810 10050 840
rect 10000 800 10050 810
rect 10300 840 10350 850
rect 10300 810 10310 840
rect 10340 810 10350 840
rect 10300 800 10350 810
rect 10600 840 10650 850
rect 10600 810 10610 840
rect 10640 810 10650 840
rect 10600 800 10650 810
rect 9550 715 9565 735
rect 9585 715 9600 735
rect 9550 685 9600 715
rect 9550 665 9565 685
rect 9585 665 9600 685
rect 9550 635 9600 665
rect 9550 615 9565 635
rect 9585 615 9600 635
rect 9550 585 9600 615
rect 9550 565 9565 585
rect 9585 565 9600 585
rect 9550 535 9600 565
rect 9550 515 9565 535
rect 9585 515 9600 535
rect 9550 485 9600 515
rect 9550 465 9565 485
rect 9585 465 9600 485
rect 9550 435 9600 465
rect 9550 415 9565 435
rect 9585 415 9600 435
rect 9550 385 9600 415
rect 9550 365 9565 385
rect 9585 365 9600 385
rect 9550 335 9600 365
rect 9550 315 9565 335
rect 9585 315 9600 335
rect 9550 285 9600 315
rect 9550 265 9565 285
rect 9585 265 9600 285
rect 9550 235 9600 265
rect 9550 215 9565 235
rect 9585 215 9600 235
rect 9550 185 9600 215
rect 9550 165 9565 185
rect 9585 165 9600 185
rect 9550 135 9600 165
rect 9550 115 9565 135
rect 9585 115 9600 135
rect 9550 85 9600 115
rect 9550 65 9565 85
rect 9585 65 9600 85
rect 9550 50 9600 65
rect 10750 740 10800 910
rect 11950 1585 14400 1600
rect 11950 1565 11965 1585
rect 11985 1565 12565 1585
rect 12585 1565 13165 1585
rect 13185 1565 13765 1585
rect 13785 1565 14365 1585
rect 14385 1565 14400 1585
rect 11950 1550 14400 1565
rect 11950 1535 12000 1550
rect 11950 1515 11965 1535
rect 11985 1515 12000 1535
rect 11950 1485 12000 1515
rect 12550 1535 12600 1550
rect 12550 1515 12565 1535
rect 12585 1515 12600 1535
rect 11950 1465 11965 1485
rect 11985 1465 12000 1485
rect 11950 1435 12000 1465
rect 11950 1415 11965 1435
rect 11985 1415 12000 1435
rect 11950 1385 12000 1415
rect 11950 1365 11965 1385
rect 11985 1365 12000 1385
rect 11950 1335 12000 1365
rect 11950 1315 11965 1335
rect 11985 1315 12000 1335
rect 11950 1285 12000 1315
rect 11950 1265 11965 1285
rect 11985 1265 12000 1285
rect 11950 1235 12000 1265
rect 11950 1215 11965 1235
rect 11985 1215 12000 1235
rect 11950 1185 12000 1215
rect 11950 1165 11965 1185
rect 11985 1165 12000 1185
rect 11950 1135 12000 1165
rect 11950 1115 11965 1135
rect 11985 1115 12000 1135
rect 11950 1085 12000 1115
rect 11950 1065 11965 1085
rect 11985 1065 12000 1085
rect 11950 1035 12000 1065
rect 11950 1015 11965 1035
rect 11985 1015 12000 1035
rect 11950 985 12000 1015
rect 11950 965 11965 985
rect 11985 965 12000 985
rect 11950 935 12000 965
rect 11950 915 11965 935
rect 11985 915 12000 935
rect 10900 840 10950 850
rect 10900 810 10910 840
rect 10940 810 10950 840
rect 10900 800 10950 810
rect 11200 840 11250 850
rect 11200 810 11210 840
rect 11240 810 11250 840
rect 11200 800 11250 810
rect 11500 840 11550 850
rect 11500 810 11510 840
rect 11540 810 11550 840
rect 11500 800 11550 810
rect 11800 840 11850 850
rect 11800 810 11810 840
rect 11840 810 11850 840
rect 11800 800 11850 810
rect 10750 710 10760 740
rect 10790 710 10800 740
rect 10750 685 10800 710
rect 10750 665 10765 685
rect 10785 665 10800 685
rect 10750 640 10800 665
rect 10750 610 10760 640
rect 10790 610 10800 640
rect 10750 585 10800 610
rect 10750 565 10765 585
rect 10785 565 10800 585
rect 10750 540 10800 565
rect 10750 510 10760 540
rect 10790 510 10800 540
rect 10750 485 10800 510
rect 10750 465 10765 485
rect 10785 465 10800 485
rect 10750 440 10800 465
rect 10750 410 10760 440
rect 10790 410 10800 440
rect 10750 385 10800 410
rect 10750 365 10765 385
rect 10785 365 10800 385
rect 10750 340 10800 365
rect 10750 310 10760 340
rect 10790 310 10800 340
rect 10750 285 10800 310
rect 10750 265 10765 285
rect 10785 265 10800 285
rect 10750 240 10800 265
rect 10750 210 10760 240
rect 10790 210 10800 240
rect 10750 185 10800 210
rect 10750 165 10765 185
rect 10785 165 10800 185
rect 10750 140 10800 165
rect 10750 110 10760 140
rect 10790 110 10800 140
rect 10750 85 10800 110
rect 10750 65 10765 85
rect 10785 65 10800 85
rect 8350 -40 8360 -10
rect 8390 -40 8400 -10
rect -50 -135 -35 -115
rect -15 -135 0 -115
rect -50 -160 0 -135
rect -50 -190 -40 -160
rect -10 -190 0 -160
rect -50 -215 0 -190
rect -50 -235 -35 -215
rect -15 -235 0 -215
rect -50 -260 0 -235
rect -50 -290 -40 -260
rect -10 -290 0 -260
rect -50 -315 0 -290
rect -50 -335 -35 -315
rect -15 -335 0 -315
rect -50 -360 0 -335
rect -50 -390 -40 -360
rect -10 -390 0 -360
rect -50 -415 0 -390
rect -50 -435 -35 -415
rect -15 -435 0 -415
rect -50 -460 0 -435
rect -50 -490 -40 -460
rect -10 -490 0 -460
rect -50 -515 0 -490
rect -50 -535 -35 -515
rect -15 -535 0 -515
rect -50 -560 0 -535
rect -50 -590 -40 -560
rect -10 -590 0 -560
rect -50 -615 0 -590
rect -50 -635 -35 -615
rect -15 -635 0 -615
rect -50 -660 0 -635
rect -50 -690 -40 -660
rect -10 -690 0 -660
rect -50 -715 0 -690
rect -50 -735 -35 -715
rect -15 -735 0 -715
rect -50 -760 0 -735
rect -50 -790 -40 -760
rect -10 -790 0 -760
rect -350 -890 -340 -860
rect -310 -890 -300 -860
rect -650 -990 -640 -960
rect -610 -990 -600 -960
rect -650 -1015 -600 -990
rect -650 -1035 -635 -1015
rect -615 -1035 -600 -1015
rect -650 -1060 -600 -1035
rect -650 -1090 -640 -1060
rect -610 -1090 -600 -1060
rect -650 -1115 -600 -1090
rect -650 -1135 -635 -1115
rect -615 -1135 -600 -1115
rect -650 -1160 -600 -1135
rect -650 -1190 -640 -1160
rect -610 -1190 -600 -1160
rect -650 -1215 -600 -1190
rect -650 -1235 -635 -1215
rect -615 -1235 -600 -1215
rect -650 -1260 -600 -1235
rect -650 -1290 -640 -1260
rect -610 -1290 -600 -1260
rect -650 -1315 -600 -1290
rect -650 -1335 -635 -1315
rect -615 -1335 -600 -1315
rect -650 -1360 -600 -1335
rect -650 -1390 -640 -1360
rect -610 -1390 -600 -1360
rect -650 -1415 -600 -1390
rect -650 -1435 -635 -1415
rect -615 -1435 -600 -1415
rect -650 -1460 -600 -1435
rect -650 -1490 -640 -1460
rect -610 -1490 -600 -1460
rect -650 -1515 -600 -1490
rect -650 -1535 -635 -1515
rect -615 -1535 -600 -1515
rect -650 -1560 -600 -1535
rect -650 -1590 -640 -1560
rect -610 -1590 -600 -1560
rect -650 -1615 -600 -1590
rect -650 -1635 -635 -1615
rect -615 -1635 -600 -1615
rect -650 -1710 -600 -1635
rect -500 -965 -450 -950
rect -500 -985 -485 -965
rect -465 -985 -450 -965
rect -500 -1015 -450 -985
rect -500 -1035 -485 -1015
rect -465 -1035 -450 -1015
rect -500 -1065 -450 -1035
rect -500 -1085 -485 -1065
rect -465 -1085 -450 -1065
rect -500 -1115 -450 -1085
rect -500 -1135 -485 -1115
rect -465 -1135 -450 -1115
rect -500 -1165 -450 -1135
rect -500 -1185 -485 -1165
rect -465 -1185 -450 -1165
rect -500 -1215 -450 -1185
rect -500 -1235 -485 -1215
rect -465 -1235 -450 -1215
rect -500 -1265 -450 -1235
rect -500 -1285 -485 -1265
rect -465 -1285 -450 -1265
rect -500 -1315 -450 -1285
rect -500 -1335 -485 -1315
rect -465 -1335 -450 -1315
rect -500 -1365 -450 -1335
rect -500 -1385 -485 -1365
rect -465 -1385 -450 -1365
rect -500 -1415 -450 -1385
rect -500 -1435 -485 -1415
rect -465 -1435 -450 -1415
rect -500 -1465 -450 -1435
rect -500 -1485 -485 -1465
rect -465 -1485 -450 -1465
rect -500 -1515 -450 -1485
rect -500 -1535 -485 -1515
rect -465 -1535 -450 -1515
rect -500 -1565 -450 -1535
rect -500 -1585 -485 -1565
rect -465 -1585 -450 -1565
rect -500 -1615 -450 -1585
rect -500 -1635 -485 -1615
rect -465 -1635 -450 -1615
rect -500 -1650 -450 -1635
rect -350 -965 -300 -890
rect -200 -860 -150 -850
rect -200 -890 -190 -860
rect -160 -890 -150 -860
rect -200 -900 -150 -890
rect -350 -985 -335 -965
rect -315 -985 -300 -965
rect -350 -1015 -300 -985
rect -350 -1035 -335 -1015
rect -315 -1035 -300 -1015
rect -350 -1065 -300 -1035
rect -350 -1085 -335 -1065
rect -315 -1085 -300 -1065
rect -350 -1115 -300 -1085
rect -350 -1135 -335 -1115
rect -315 -1135 -300 -1115
rect -350 -1165 -300 -1135
rect -350 -1185 -335 -1165
rect -315 -1185 -300 -1165
rect -350 -1215 -300 -1185
rect -350 -1235 -335 -1215
rect -315 -1235 -300 -1215
rect -350 -1265 -300 -1235
rect -350 -1285 -335 -1265
rect -315 -1285 -300 -1265
rect -350 -1315 -300 -1285
rect -350 -1335 -335 -1315
rect -315 -1335 -300 -1315
rect -350 -1365 -300 -1335
rect -350 -1385 -335 -1365
rect -315 -1385 -300 -1365
rect -350 -1415 -300 -1385
rect -350 -1435 -335 -1415
rect -315 -1435 -300 -1415
rect -350 -1465 -300 -1435
rect -350 -1485 -335 -1465
rect -315 -1485 -300 -1465
rect -350 -1515 -300 -1485
rect -350 -1535 -335 -1515
rect -315 -1535 -300 -1515
rect -350 -1565 -300 -1535
rect -350 -1585 -335 -1565
rect -315 -1585 -300 -1565
rect -350 -1615 -300 -1585
rect -350 -1635 -335 -1615
rect -315 -1635 -300 -1615
rect -350 -1650 -300 -1635
rect -200 -965 -150 -950
rect -200 -985 -185 -965
rect -165 -985 -150 -965
rect -200 -1015 -150 -985
rect -200 -1035 -185 -1015
rect -165 -1035 -150 -1015
rect -200 -1065 -150 -1035
rect -200 -1085 -185 -1065
rect -165 -1085 -150 -1065
rect -200 -1115 -150 -1085
rect -200 -1135 -185 -1115
rect -165 -1135 -150 -1115
rect -200 -1165 -150 -1135
rect -200 -1185 -185 -1165
rect -165 -1185 -150 -1165
rect -200 -1215 -150 -1185
rect -200 -1235 -185 -1215
rect -165 -1235 -150 -1215
rect -200 -1265 -150 -1235
rect -200 -1285 -185 -1265
rect -165 -1285 -150 -1265
rect -200 -1315 -150 -1285
rect -200 -1335 -185 -1315
rect -165 -1335 -150 -1315
rect -200 -1365 -150 -1335
rect -200 -1385 -185 -1365
rect -165 -1385 -150 -1365
rect -200 -1415 -150 -1385
rect -200 -1435 -185 -1415
rect -165 -1435 -150 -1415
rect -200 -1465 -150 -1435
rect -200 -1485 -185 -1465
rect -165 -1485 -150 -1465
rect -200 -1515 -150 -1485
rect -200 -1535 -185 -1515
rect -165 -1535 -150 -1515
rect -200 -1565 -150 -1535
rect -200 -1585 -185 -1565
rect -165 -1585 -150 -1565
rect -200 -1615 -150 -1585
rect -200 -1635 -185 -1615
rect -165 -1635 -150 -1615
rect -200 -1650 -150 -1635
rect -50 -960 0 -790
rect 1150 -115 7200 -100
rect 1150 -135 1165 -115
rect 1185 -135 1765 -115
rect 1785 -135 2365 -115
rect 2385 -135 2965 -115
rect 2985 -135 3565 -115
rect 3585 -135 3865 -115
rect 3885 -135 4165 -115
rect 4185 -135 4465 -115
rect 4485 -135 4765 -115
rect 4785 -135 5365 -115
rect 5385 -135 5965 -115
rect 5985 -135 6565 -115
rect 6585 -135 7165 -115
rect 7185 -135 7200 -115
rect 1150 -150 7200 -135
rect 1150 -165 1200 -150
rect 1150 -185 1165 -165
rect 1185 -185 1200 -165
rect 1150 -215 1200 -185
rect 1750 -165 1800 -150
rect 1750 -185 1765 -165
rect 1785 -185 1800 -165
rect 1150 -235 1165 -215
rect 1185 -235 1200 -215
rect 1150 -265 1200 -235
rect 1150 -285 1165 -265
rect 1185 -285 1200 -265
rect 1150 -315 1200 -285
rect 1150 -335 1165 -315
rect 1185 -335 1200 -315
rect 1150 -365 1200 -335
rect 1150 -385 1165 -365
rect 1185 -385 1200 -365
rect 1150 -415 1200 -385
rect 1150 -435 1165 -415
rect 1185 -435 1200 -415
rect 1150 -465 1200 -435
rect 1150 -485 1165 -465
rect 1185 -485 1200 -465
rect 1150 -515 1200 -485
rect 1150 -535 1165 -515
rect 1185 -535 1200 -515
rect 1150 -565 1200 -535
rect 1150 -585 1165 -565
rect 1185 -585 1200 -565
rect 1150 -615 1200 -585
rect 1150 -635 1165 -615
rect 1185 -635 1200 -615
rect 1150 -665 1200 -635
rect 1150 -685 1165 -665
rect 1185 -685 1200 -665
rect 1150 -715 1200 -685
rect 1150 -735 1165 -715
rect 1185 -735 1200 -715
rect 1150 -765 1200 -735
rect 1150 -785 1165 -765
rect 1185 -785 1200 -765
rect 1150 -800 1200 -785
rect 1450 -215 1500 -200
rect 1450 -235 1465 -215
rect 1485 -235 1500 -215
rect 1450 -265 1500 -235
rect 1450 -285 1465 -265
rect 1485 -285 1500 -265
rect 1450 -315 1500 -285
rect 1450 -335 1465 -315
rect 1485 -335 1500 -315
rect 1450 -365 1500 -335
rect 1450 -385 1465 -365
rect 1485 -385 1500 -365
rect 1450 -415 1500 -385
rect 1450 -435 1465 -415
rect 1485 -435 1500 -415
rect 1450 -465 1500 -435
rect 1450 -485 1465 -465
rect 1485 -485 1500 -465
rect 1450 -515 1500 -485
rect 1450 -535 1465 -515
rect 1485 -535 1500 -515
rect 1450 -565 1500 -535
rect 1450 -585 1465 -565
rect 1485 -585 1500 -565
rect 1450 -615 1500 -585
rect 1450 -635 1465 -615
rect 1485 -635 1500 -615
rect 1450 -665 1500 -635
rect 1450 -685 1465 -665
rect 1485 -685 1500 -665
rect 1450 -715 1500 -685
rect 1750 -215 1800 -185
rect 2350 -165 2400 -150
rect 2350 -185 2365 -165
rect 2385 -185 2400 -165
rect 1750 -235 1765 -215
rect 1785 -235 1800 -215
rect 1750 -265 1800 -235
rect 1750 -285 1765 -265
rect 1785 -285 1800 -265
rect 1750 -315 1800 -285
rect 1750 -335 1765 -315
rect 1785 -335 1800 -315
rect 1750 -365 1800 -335
rect 1750 -385 1765 -365
rect 1785 -385 1800 -365
rect 1750 -415 1800 -385
rect 1750 -435 1765 -415
rect 1785 -435 1800 -415
rect 1750 -465 1800 -435
rect 1750 -485 1765 -465
rect 1785 -485 1800 -465
rect 1750 -515 1800 -485
rect 1750 -535 1765 -515
rect 1785 -535 1800 -515
rect 1750 -565 1800 -535
rect 1750 -585 1765 -565
rect 1785 -585 1800 -565
rect 1750 -615 1800 -585
rect 1750 -635 1765 -615
rect 1785 -635 1800 -615
rect 1750 -665 1800 -635
rect 1750 -685 1765 -665
rect 1785 -685 1800 -665
rect 1750 -700 1800 -685
rect 2050 -215 2100 -200
rect 2050 -235 2065 -215
rect 2085 -235 2100 -215
rect 2050 -265 2100 -235
rect 2050 -285 2065 -265
rect 2085 -285 2100 -265
rect 2050 -315 2100 -285
rect 2050 -335 2065 -315
rect 2085 -335 2100 -315
rect 2050 -365 2100 -335
rect 2050 -385 2065 -365
rect 2085 -385 2100 -365
rect 2050 -415 2100 -385
rect 2050 -435 2065 -415
rect 2085 -435 2100 -415
rect 2050 -465 2100 -435
rect 2050 -485 2065 -465
rect 2085 -485 2100 -465
rect 2050 -515 2100 -485
rect 2050 -535 2065 -515
rect 2085 -535 2100 -515
rect 2050 -565 2100 -535
rect 2050 -585 2065 -565
rect 2085 -585 2100 -565
rect 2050 -615 2100 -585
rect 2050 -635 2065 -615
rect 2085 -635 2100 -615
rect 2050 -665 2100 -635
rect 2050 -685 2065 -665
rect 2085 -685 2100 -665
rect 1450 -735 1465 -715
rect 1485 -735 1500 -715
rect 1450 -750 1500 -735
rect 2050 -715 2100 -685
rect 2350 -215 2400 -185
rect 2950 -165 3000 -150
rect 2950 -185 2965 -165
rect 2985 -185 3000 -165
rect 2350 -235 2365 -215
rect 2385 -235 2400 -215
rect 2350 -265 2400 -235
rect 2350 -285 2365 -265
rect 2385 -285 2400 -265
rect 2350 -315 2400 -285
rect 2350 -335 2365 -315
rect 2385 -335 2400 -315
rect 2350 -365 2400 -335
rect 2350 -385 2365 -365
rect 2385 -385 2400 -365
rect 2350 -415 2400 -385
rect 2350 -435 2365 -415
rect 2385 -435 2400 -415
rect 2350 -465 2400 -435
rect 2350 -485 2365 -465
rect 2385 -485 2400 -465
rect 2350 -515 2400 -485
rect 2350 -535 2365 -515
rect 2385 -535 2400 -515
rect 2350 -565 2400 -535
rect 2350 -585 2365 -565
rect 2385 -585 2400 -565
rect 2350 -615 2400 -585
rect 2350 -635 2365 -615
rect 2385 -635 2400 -615
rect 2350 -665 2400 -635
rect 2350 -685 2365 -665
rect 2385 -685 2400 -665
rect 2350 -700 2400 -685
rect 2650 -215 2700 -200
rect 2650 -235 2665 -215
rect 2685 -235 2700 -215
rect 2650 -265 2700 -235
rect 2650 -285 2665 -265
rect 2685 -285 2700 -265
rect 2650 -315 2700 -285
rect 2650 -335 2665 -315
rect 2685 -335 2700 -315
rect 2650 -365 2700 -335
rect 2650 -385 2665 -365
rect 2685 -385 2700 -365
rect 2650 -415 2700 -385
rect 2650 -435 2665 -415
rect 2685 -435 2700 -415
rect 2650 -465 2700 -435
rect 2650 -485 2665 -465
rect 2685 -485 2700 -465
rect 2650 -515 2700 -485
rect 2650 -535 2665 -515
rect 2685 -535 2700 -515
rect 2650 -565 2700 -535
rect 2650 -585 2665 -565
rect 2685 -585 2700 -565
rect 2650 -615 2700 -585
rect 2650 -635 2665 -615
rect 2685 -635 2700 -615
rect 2650 -665 2700 -635
rect 2650 -685 2665 -665
rect 2685 -685 2700 -665
rect 2050 -735 2065 -715
rect 2085 -735 2100 -715
rect 2050 -750 2100 -735
rect 2650 -715 2700 -685
rect 2950 -215 3000 -185
rect 3550 -165 3600 -150
rect 3550 -185 3565 -165
rect 3585 -185 3600 -165
rect 2950 -235 2965 -215
rect 2985 -235 3000 -215
rect 2950 -265 3000 -235
rect 2950 -285 2965 -265
rect 2985 -285 3000 -265
rect 2950 -315 3000 -285
rect 2950 -335 2965 -315
rect 2985 -335 3000 -315
rect 2950 -365 3000 -335
rect 2950 -385 2965 -365
rect 2985 -385 3000 -365
rect 2950 -415 3000 -385
rect 2950 -435 2965 -415
rect 2985 -435 3000 -415
rect 2950 -465 3000 -435
rect 2950 -485 2965 -465
rect 2985 -485 3000 -465
rect 2950 -515 3000 -485
rect 2950 -535 2965 -515
rect 2985 -535 3000 -515
rect 2950 -565 3000 -535
rect 2950 -585 2965 -565
rect 2985 -585 3000 -565
rect 2950 -615 3000 -585
rect 2950 -635 2965 -615
rect 2985 -635 3000 -615
rect 2950 -665 3000 -635
rect 2950 -685 2965 -665
rect 2985 -685 3000 -665
rect 2950 -700 3000 -685
rect 3250 -215 3300 -200
rect 3250 -235 3265 -215
rect 3285 -235 3300 -215
rect 3250 -265 3300 -235
rect 3250 -285 3265 -265
rect 3285 -285 3300 -265
rect 3250 -315 3300 -285
rect 3250 -335 3265 -315
rect 3285 -335 3300 -315
rect 3250 -365 3300 -335
rect 3250 -385 3265 -365
rect 3285 -385 3300 -365
rect 3250 -415 3300 -385
rect 3250 -435 3265 -415
rect 3285 -435 3300 -415
rect 3250 -465 3300 -435
rect 3250 -485 3265 -465
rect 3285 -485 3300 -465
rect 3250 -515 3300 -485
rect 3250 -535 3265 -515
rect 3285 -535 3300 -515
rect 3250 -565 3300 -535
rect 3250 -585 3265 -565
rect 3285 -585 3300 -565
rect 3250 -615 3300 -585
rect 3250 -635 3265 -615
rect 3285 -635 3300 -615
rect 3250 -665 3300 -635
rect 3250 -685 3265 -665
rect 3285 -685 3300 -665
rect 2650 -735 2665 -715
rect 2685 -735 2700 -715
rect 2650 -750 2700 -735
rect 3250 -715 3300 -685
rect 3250 -735 3265 -715
rect 3285 -735 3300 -715
rect 3250 -750 3300 -735
rect 1450 -765 3300 -750
rect 1450 -785 1465 -765
rect 1485 -785 2065 -765
rect 2085 -785 2665 -765
rect 2685 -785 3265 -765
rect 3285 -785 3300 -765
rect 1450 -800 3300 -785
rect 3550 -215 3600 -185
rect 3850 -165 3900 -150
rect 3850 -185 3865 -165
rect 3885 -185 3900 -165
rect 3550 -235 3565 -215
rect 3585 -235 3600 -215
rect 3550 -265 3600 -235
rect 3550 -285 3565 -265
rect 3585 -285 3600 -265
rect 3550 -315 3600 -285
rect 3550 -335 3565 -315
rect 3585 -335 3600 -315
rect 3550 -365 3600 -335
rect 3550 -385 3565 -365
rect 3585 -385 3600 -365
rect 3550 -415 3600 -385
rect 3550 -435 3565 -415
rect 3585 -435 3600 -415
rect 3550 -465 3600 -435
rect 3550 -485 3565 -465
rect 3585 -485 3600 -465
rect 3550 -515 3600 -485
rect 3550 -535 3565 -515
rect 3585 -535 3600 -515
rect 3550 -565 3600 -535
rect 3550 -585 3565 -565
rect 3585 -585 3600 -565
rect 3550 -615 3600 -585
rect 3550 -635 3565 -615
rect 3585 -635 3600 -615
rect 3550 -665 3600 -635
rect 3550 -685 3565 -665
rect 3585 -685 3600 -665
rect 3550 -715 3600 -685
rect 3550 -735 3565 -715
rect 3585 -735 3600 -715
rect 3550 -765 3600 -735
rect 3550 -785 3565 -765
rect 3585 -785 3600 -765
rect 3550 -800 3600 -785
rect 3700 -215 3750 -200
rect 3700 -235 3715 -215
rect 3735 -235 3750 -215
rect 3700 -265 3750 -235
rect 3700 -285 3715 -265
rect 3735 -285 3750 -265
rect 3700 -315 3750 -285
rect 3700 -335 3715 -315
rect 3735 -335 3750 -315
rect 3700 -365 3750 -335
rect 3700 -385 3715 -365
rect 3735 -385 3750 -365
rect 3700 -415 3750 -385
rect 3700 -435 3715 -415
rect 3735 -435 3750 -415
rect 3700 -465 3750 -435
rect 3700 -485 3715 -465
rect 3735 -485 3750 -465
rect 3700 -515 3750 -485
rect 3700 -535 3715 -515
rect 3735 -535 3750 -515
rect 3700 -565 3750 -535
rect 3700 -585 3715 -565
rect 3735 -585 3750 -565
rect 3700 -615 3750 -585
rect 3700 -635 3715 -615
rect 3735 -635 3750 -615
rect 3700 -665 3750 -635
rect 3700 -685 3715 -665
rect 3735 -685 3750 -665
rect 3700 -715 3750 -685
rect 3850 -215 3900 -185
rect 4150 -165 4200 -150
rect 4150 -185 4165 -165
rect 4185 -185 4200 -165
rect 3850 -235 3865 -215
rect 3885 -235 3900 -215
rect 3850 -265 3900 -235
rect 3850 -285 3865 -265
rect 3885 -285 3900 -265
rect 3850 -315 3900 -285
rect 3850 -335 3865 -315
rect 3885 -335 3900 -315
rect 3850 -365 3900 -335
rect 3850 -385 3865 -365
rect 3885 -385 3900 -365
rect 3850 -415 3900 -385
rect 3850 -435 3865 -415
rect 3885 -435 3900 -415
rect 3850 -465 3900 -435
rect 3850 -485 3865 -465
rect 3885 -485 3900 -465
rect 3850 -515 3900 -485
rect 3850 -535 3865 -515
rect 3885 -535 3900 -515
rect 3850 -565 3900 -535
rect 3850 -585 3865 -565
rect 3885 -585 3900 -565
rect 3850 -615 3900 -585
rect 3850 -635 3865 -615
rect 3885 -635 3900 -615
rect 3850 -665 3900 -635
rect 3850 -685 3865 -665
rect 3885 -685 3900 -665
rect 3850 -700 3900 -685
rect 4000 -215 4050 -200
rect 4000 -235 4015 -215
rect 4035 -235 4050 -215
rect 4000 -265 4050 -235
rect 4000 -285 4015 -265
rect 4035 -285 4050 -265
rect 4000 -315 4050 -285
rect 4000 -335 4015 -315
rect 4035 -335 4050 -315
rect 4000 -365 4050 -335
rect 4000 -385 4015 -365
rect 4035 -385 4050 -365
rect 4000 -415 4050 -385
rect 4000 -435 4015 -415
rect 4035 -435 4050 -415
rect 4000 -465 4050 -435
rect 4000 -485 4015 -465
rect 4035 -485 4050 -465
rect 4000 -515 4050 -485
rect 4000 -535 4015 -515
rect 4035 -535 4050 -515
rect 4000 -565 4050 -535
rect 4000 -585 4015 -565
rect 4035 -585 4050 -565
rect 4000 -615 4050 -585
rect 4000 -635 4015 -615
rect 4035 -635 4050 -615
rect 4000 -665 4050 -635
rect 4000 -685 4015 -665
rect 4035 -685 4050 -665
rect 3700 -735 3715 -715
rect 3735 -735 3750 -715
rect 3700 -750 3750 -735
rect 4000 -715 4050 -685
rect 4000 -735 4015 -715
rect 4035 -735 4050 -715
rect 4000 -750 4050 -735
rect 3700 -765 4050 -750
rect 3700 -785 3715 -765
rect 3735 -785 4015 -765
rect 4035 -785 4050 -765
rect 3700 -800 4050 -785
rect 4150 -215 4200 -185
rect 4450 -165 4500 -150
rect 4450 -185 4465 -165
rect 4485 -185 4500 -165
rect 4150 -235 4165 -215
rect 4185 -235 4200 -215
rect 4150 -265 4200 -235
rect 4150 -285 4165 -265
rect 4185 -285 4200 -265
rect 4150 -315 4200 -285
rect 4150 -335 4165 -315
rect 4185 -335 4200 -315
rect 4150 -365 4200 -335
rect 4150 -385 4165 -365
rect 4185 -385 4200 -365
rect 4150 -415 4200 -385
rect 4150 -435 4165 -415
rect 4185 -435 4200 -415
rect 4150 -465 4200 -435
rect 4150 -485 4165 -465
rect 4185 -485 4200 -465
rect 4150 -515 4200 -485
rect 4150 -535 4165 -515
rect 4185 -535 4200 -515
rect 4150 -565 4200 -535
rect 4150 -585 4165 -565
rect 4185 -585 4200 -565
rect 4150 -615 4200 -585
rect 4150 -635 4165 -615
rect 4185 -635 4200 -615
rect 4150 -665 4200 -635
rect 4150 -685 4165 -665
rect 4185 -685 4200 -665
rect 4150 -715 4200 -685
rect 4150 -735 4165 -715
rect 4185 -735 4200 -715
rect 4150 -765 4200 -735
rect 4150 -785 4165 -765
rect 4185 -785 4200 -765
rect 4150 -800 4200 -785
rect 4300 -215 4350 -200
rect 4300 -235 4315 -215
rect 4335 -235 4350 -215
rect 4300 -265 4350 -235
rect 4300 -285 4315 -265
rect 4335 -285 4350 -265
rect 4300 -315 4350 -285
rect 4300 -335 4315 -315
rect 4335 -335 4350 -315
rect 4300 -365 4350 -335
rect 4300 -385 4315 -365
rect 4335 -385 4350 -365
rect 4300 -415 4350 -385
rect 4300 -435 4315 -415
rect 4335 -435 4350 -415
rect 4300 -465 4350 -435
rect 4300 -485 4315 -465
rect 4335 -485 4350 -465
rect 4300 -515 4350 -485
rect 4300 -535 4315 -515
rect 4335 -535 4350 -515
rect 4300 -565 4350 -535
rect 4300 -585 4315 -565
rect 4335 -585 4350 -565
rect 4300 -615 4350 -585
rect 4300 -635 4315 -615
rect 4335 -635 4350 -615
rect 4300 -665 4350 -635
rect 4300 -685 4315 -665
rect 4335 -685 4350 -665
rect 4300 -715 4350 -685
rect 4450 -215 4500 -185
rect 4750 -165 4800 -150
rect 4750 -185 4765 -165
rect 4785 -185 4800 -165
rect 4450 -235 4465 -215
rect 4485 -235 4500 -215
rect 4450 -265 4500 -235
rect 4450 -285 4465 -265
rect 4485 -285 4500 -265
rect 4450 -315 4500 -285
rect 4450 -335 4465 -315
rect 4485 -335 4500 -315
rect 4450 -365 4500 -335
rect 4450 -385 4465 -365
rect 4485 -385 4500 -365
rect 4450 -415 4500 -385
rect 4450 -435 4465 -415
rect 4485 -435 4500 -415
rect 4450 -465 4500 -435
rect 4450 -485 4465 -465
rect 4485 -485 4500 -465
rect 4450 -515 4500 -485
rect 4450 -535 4465 -515
rect 4485 -535 4500 -515
rect 4450 -565 4500 -535
rect 4450 -585 4465 -565
rect 4485 -585 4500 -565
rect 4450 -615 4500 -585
rect 4450 -635 4465 -615
rect 4485 -635 4500 -615
rect 4450 -665 4500 -635
rect 4450 -685 4465 -665
rect 4485 -685 4500 -665
rect 4450 -700 4500 -685
rect 4600 -215 4650 -200
rect 4600 -235 4615 -215
rect 4635 -235 4650 -215
rect 4600 -265 4650 -235
rect 4600 -285 4615 -265
rect 4635 -285 4650 -265
rect 4600 -315 4650 -285
rect 4600 -335 4615 -315
rect 4635 -335 4650 -315
rect 4600 -365 4650 -335
rect 4600 -385 4615 -365
rect 4635 -385 4650 -365
rect 4600 -415 4650 -385
rect 4600 -435 4615 -415
rect 4635 -435 4650 -415
rect 4600 -465 4650 -435
rect 4600 -485 4615 -465
rect 4635 -485 4650 -465
rect 4600 -515 4650 -485
rect 4600 -535 4615 -515
rect 4635 -535 4650 -515
rect 4600 -565 4650 -535
rect 4600 -585 4615 -565
rect 4635 -585 4650 -565
rect 4600 -615 4650 -585
rect 4600 -635 4615 -615
rect 4635 -635 4650 -615
rect 4600 -665 4650 -635
rect 4600 -685 4615 -665
rect 4635 -685 4650 -665
rect 4300 -735 4315 -715
rect 4335 -735 4350 -715
rect 4300 -750 4350 -735
rect 4600 -715 4650 -685
rect 4600 -735 4615 -715
rect 4635 -735 4650 -715
rect 4600 -750 4650 -735
rect 4300 -765 4650 -750
rect 4300 -785 4315 -765
rect 4335 -785 4615 -765
rect 4635 -785 4650 -765
rect 4300 -800 4650 -785
rect 4750 -215 4800 -185
rect 5350 -165 5400 -150
rect 5350 -185 5365 -165
rect 5385 -185 5400 -165
rect 4750 -235 4765 -215
rect 4785 -235 4800 -215
rect 4750 -265 4800 -235
rect 4750 -285 4765 -265
rect 4785 -285 4800 -265
rect 4750 -315 4800 -285
rect 4750 -335 4765 -315
rect 4785 -335 4800 -315
rect 4750 -365 4800 -335
rect 4750 -385 4765 -365
rect 4785 -385 4800 -365
rect 4750 -415 4800 -385
rect 4750 -435 4765 -415
rect 4785 -435 4800 -415
rect 4750 -465 4800 -435
rect 4750 -485 4765 -465
rect 4785 -485 4800 -465
rect 4750 -515 4800 -485
rect 4750 -535 4765 -515
rect 4785 -535 4800 -515
rect 4750 -565 4800 -535
rect 4750 -585 4765 -565
rect 4785 -585 4800 -565
rect 4750 -615 4800 -585
rect 4750 -635 4765 -615
rect 4785 -635 4800 -615
rect 4750 -665 4800 -635
rect 4750 -685 4765 -665
rect 4785 -685 4800 -665
rect 4750 -715 4800 -685
rect 4750 -735 4765 -715
rect 4785 -735 4800 -715
rect 4750 -765 4800 -735
rect 4750 -785 4765 -765
rect 4785 -785 4800 -765
rect 4750 -800 4800 -785
rect 5050 -215 5100 -200
rect 5050 -235 5065 -215
rect 5085 -235 5100 -215
rect 5050 -265 5100 -235
rect 5050 -285 5065 -265
rect 5085 -285 5100 -265
rect 5050 -315 5100 -285
rect 5050 -335 5065 -315
rect 5085 -335 5100 -315
rect 5050 -365 5100 -335
rect 5050 -385 5065 -365
rect 5085 -385 5100 -365
rect 5050 -415 5100 -385
rect 5050 -435 5065 -415
rect 5085 -435 5100 -415
rect 5050 -465 5100 -435
rect 5050 -485 5065 -465
rect 5085 -485 5100 -465
rect 5050 -515 5100 -485
rect 5050 -535 5065 -515
rect 5085 -535 5100 -515
rect 5050 -565 5100 -535
rect 5050 -585 5065 -565
rect 5085 -585 5100 -565
rect 5050 -615 5100 -585
rect 5050 -635 5065 -615
rect 5085 -635 5100 -615
rect 5050 -665 5100 -635
rect 5050 -685 5065 -665
rect 5085 -685 5100 -665
rect 5050 -715 5100 -685
rect 5350 -215 5400 -185
rect 5950 -165 6000 -150
rect 5950 -185 5965 -165
rect 5985 -185 6000 -165
rect 5350 -235 5365 -215
rect 5385 -235 5400 -215
rect 5350 -265 5400 -235
rect 5350 -285 5365 -265
rect 5385 -285 5400 -265
rect 5350 -315 5400 -285
rect 5350 -335 5365 -315
rect 5385 -335 5400 -315
rect 5350 -365 5400 -335
rect 5350 -385 5365 -365
rect 5385 -385 5400 -365
rect 5350 -415 5400 -385
rect 5350 -435 5365 -415
rect 5385 -435 5400 -415
rect 5350 -465 5400 -435
rect 5350 -485 5365 -465
rect 5385 -485 5400 -465
rect 5350 -515 5400 -485
rect 5350 -535 5365 -515
rect 5385 -535 5400 -515
rect 5350 -565 5400 -535
rect 5350 -585 5365 -565
rect 5385 -585 5400 -565
rect 5350 -615 5400 -585
rect 5350 -635 5365 -615
rect 5385 -635 5400 -615
rect 5350 -665 5400 -635
rect 5350 -685 5365 -665
rect 5385 -685 5400 -665
rect 5350 -700 5400 -685
rect 5650 -215 5700 -200
rect 5650 -235 5665 -215
rect 5685 -235 5700 -215
rect 5650 -265 5700 -235
rect 5650 -285 5665 -265
rect 5685 -285 5700 -265
rect 5650 -315 5700 -285
rect 5650 -335 5665 -315
rect 5685 -335 5700 -315
rect 5650 -365 5700 -335
rect 5650 -385 5665 -365
rect 5685 -385 5700 -365
rect 5650 -415 5700 -385
rect 5650 -435 5665 -415
rect 5685 -435 5700 -415
rect 5650 -465 5700 -435
rect 5650 -485 5665 -465
rect 5685 -485 5700 -465
rect 5650 -515 5700 -485
rect 5650 -535 5665 -515
rect 5685 -535 5700 -515
rect 5650 -565 5700 -535
rect 5650 -585 5665 -565
rect 5685 -585 5700 -565
rect 5650 -615 5700 -585
rect 5650 -635 5665 -615
rect 5685 -635 5700 -615
rect 5650 -665 5700 -635
rect 5650 -685 5665 -665
rect 5685 -685 5700 -665
rect 5050 -735 5065 -715
rect 5085 -735 5100 -715
rect 5050 -750 5100 -735
rect 5650 -715 5700 -685
rect 5950 -215 6000 -185
rect 6550 -165 6600 -150
rect 6550 -185 6565 -165
rect 6585 -185 6600 -165
rect 5950 -235 5965 -215
rect 5985 -235 6000 -215
rect 5950 -265 6000 -235
rect 5950 -285 5965 -265
rect 5985 -285 6000 -265
rect 5950 -315 6000 -285
rect 5950 -335 5965 -315
rect 5985 -335 6000 -315
rect 5950 -365 6000 -335
rect 5950 -385 5965 -365
rect 5985 -385 6000 -365
rect 5950 -415 6000 -385
rect 5950 -435 5965 -415
rect 5985 -435 6000 -415
rect 5950 -465 6000 -435
rect 5950 -485 5965 -465
rect 5985 -485 6000 -465
rect 5950 -515 6000 -485
rect 5950 -535 5965 -515
rect 5985 -535 6000 -515
rect 5950 -565 6000 -535
rect 5950 -585 5965 -565
rect 5985 -585 6000 -565
rect 5950 -615 6000 -585
rect 5950 -635 5965 -615
rect 5985 -635 6000 -615
rect 5950 -665 6000 -635
rect 5950 -685 5965 -665
rect 5985 -685 6000 -665
rect 5950 -700 6000 -685
rect 6250 -215 6300 -200
rect 6250 -235 6265 -215
rect 6285 -235 6300 -215
rect 6250 -265 6300 -235
rect 6250 -285 6265 -265
rect 6285 -285 6300 -265
rect 6250 -315 6300 -285
rect 6250 -335 6265 -315
rect 6285 -335 6300 -315
rect 6250 -365 6300 -335
rect 6250 -385 6265 -365
rect 6285 -385 6300 -365
rect 6250 -415 6300 -385
rect 6250 -435 6265 -415
rect 6285 -435 6300 -415
rect 6250 -465 6300 -435
rect 6250 -485 6265 -465
rect 6285 -485 6300 -465
rect 6250 -515 6300 -485
rect 6250 -535 6265 -515
rect 6285 -535 6300 -515
rect 6250 -565 6300 -535
rect 6250 -585 6265 -565
rect 6285 -585 6300 -565
rect 6250 -615 6300 -585
rect 6250 -635 6265 -615
rect 6285 -635 6300 -615
rect 6250 -665 6300 -635
rect 6250 -685 6265 -665
rect 6285 -685 6300 -665
rect 5650 -735 5665 -715
rect 5685 -735 5700 -715
rect 5650 -750 5700 -735
rect 6250 -715 6300 -685
rect 6550 -215 6600 -185
rect 7150 -165 7200 -150
rect 7150 -185 7165 -165
rect 7185 -185 7200 -165
rect 6550 -235 6565 -215
rect 6585 -235 6600 -215
rect 6550 -265 6600 -235
rect 6550 -285 6565 -265
rect 6585 -285 6600 -265
rect 6550 -315 6600 -285
rect 6550 -335 6565 -315
rect 6585 -335 6600 -315
rect 6550 -365 6600 -335
rect 6550 -385 6565 -365
rect 6585 -385 6600 -365
rect 6550 -415 6600 -385
rect 6550 -435 6565 -415
rect 6585 -435 6600 -415
rect 6550 -465 6600 -435
rect 6550 -485 6565 -465
rect 6585 -485 6600 -465
rect 6550 -515 6600 -485
rect 6550 -535 6565 -515
rect 6585 -535 6600 -515
rect 6550 -565 6600 -535
rect 6550 -585 6565 -565
rect 6585 -585 6600 -565
rect 6550 -615 6600 -585
rect 6550 -635 6565 -615
rect 6585 -635 6600 -615
rect 6550 -665 6600 -635
rect 6550 -685 6565 -665
rect 6585 -685 6600 -665
rect 6550 -700 6600 -685
rect 6850 -215 6900 -200
rect 6850 -235 6865 -215
rect 6885 -235 6900 -215
rect 6850 -265 6900 -235
rect 6850 -285 6865 -265
rect 6885 -285 6900 -265
rect 6850 -315 6900 -285
rect 6850 -335 6865 -315
rect 6885 -335 6900 -315
rect 6850 -365 6900 -335
rect 6850 -385 6865 -365
rect 6885 -385 6900 -365
rect 6850 -415 6900 -385
rect 6850 -435 6865 -415
rect 6885 -435 6900 -415
rect 6850 -465 6900 -435
rect 6850 -485 6865 -465
rect 6885 -485 6900 -465
rect 6850 -515 6900 -485
rect 6850 -535 6865 -515
rect 6885 -535 6900 -515
rect 6850 -565 6900 -535
rect 6850 -585 6865 -565
rect 6885 -585 6900 -565
rect 6850 -615 6900 -585
rect 6850 -635 6865 -615
rect 6885 -635 6900 -615
rect 6850 -665 6900 -635
rect 6850 -685 6865 -665
rect 6885 -685 6900 -665
rect 6250 -735 6265 -715
rect 6285 -735 6300 -715
rect 6250 -750 6300 -735
rect 6850 -715 6900 -685
rect 6850 -735 6865 -715
rect 6885 -735 6900 -715
rect 6850 -750 6900 -735
rect 5050 -765 6900 -750
rect 5050 -785 5065 -765
rect 5085 -785 5665 -765
rect 5685 -785 6265 -765
rect 6285 -785 6865 -765
rect 6885 -785 6900 -765
rect 5050 -800 6900 -785
rect 7150 -215 7200 -185
rect 7150 -235 7165 -215
rect 7185 -235 7200 -215
rect 7150 -265 7200 -235
rect 7150 -285 7165 -265
rect 7185 -285 7200 -265
rect 7150 -315 7200 -285
rect 7150 -335 7165 -315
rect 7185 -335 7200 -315
rect 7150 -365 7200 -335
rect 7150 -385 7165 -365
rect 7185 -385 7200 -365
rect 7150 -415 7200 -385
rect 7150 -435 7165 -415
rect 7185 -435 7200 -415
rect 7150 -465 7200 -435
rect 7150 -485 7165 -465
rect 7185 -485 7200 -465
rect 7150 -515 7200 -485
rect 7150 -535 7165 -515
rect 7185 -535 7200 -515
rect 7150 -565 7200 -535
rect 7150 -585 7165 -565
rect 7185 -585 7200 -565
rect 7150 -615 7200 -585
rect 7150 -635 7165 -615
rect 7185 -635 7200 -615
rect 7150 -665 7200 -635
rect 7150 -685 7165 -665
rect 7185 -685 7200 -665
rect 7150 -715 7200 -685
rect 7150 -735 7165 -715
rect 7185 -735 7200 -715
rect 7150 -765 7200 -735
rect 7150 -785 7165 -765
rect 7185 -785 7200 -765
rect 7150 -800 7200 -785
rect 8350 -115 8400 -40
rect 10750 -10 10800 65
rect 10750 -40 10760 -10
rect 10790 -40 10800 -10
rect 8350 -135 8365 -115
rect 8385 -135 8400 -115
rect 8350 -160 8400 -135
rect 8350 -190 8360 -160
rect 8390 -190 8400 -160
rect 8350 -215 8400 -190
rect 8350 -235 8365 -215
rect 8385 -235 8400 -215
rect 8350 -260 8400 -235
rect 8350 -290 8360 -260
rect 8390 -290 8400 -260
rect 8350 -315 8400 -290
rect 8350 -335 8365 -315
rect 8385 -335 8400 -315
rect 8350 -360 8400 -335
rect 8350 -390 8360 -360
rect 8390 -390 8400 -360
rect 8350 -415 8400 -390
rect 8350 -435 8365 -415
rect 8385 -435 8400 -415
rect 8350 -460 8400 -435
rect 8350 -490 8360 -460
rect 8390 -490 8400 -460
rect 8350 -515 8400 -490
rect 8350 -535 8365 -515
rect 8385 -535 8400 -515
rect 8350 -560 8400 -535
rect 8350 -590 8360 -560
rect 8390 -590 8400 -560
rect 8350 -615 8400 -590
rect 8350 -635 8365 -615
rect 8385 -635 8400 -615
rect 8350 -660 8400 -635
rect 8350 -690 8360 -660
rect 8390 -690 8400 -660
rect 8350 -715 8400 -690
rect 8350 -735 8365 -715
rect 8385 -735 8400 -715
rect 8350 -760 8400 -735
rect 8350 -790 8360 -760
rect 8390 -790 8400 -760
rect 100 -860 150 -850
rect 100 -890 110 -860
rect 140 -890 150 -860
rect 100 -900 150 -890
rect 400 -860 450 -850
rect 400 -890 410 -860
rect 440 -890 450 -860
rect 400 -900 450 -890
rect 700 -860 750 -850
rect 700 -890 710 -860
rect 740 -890 750 -860
rect 700 -900 750 -890
rect 1000 -860 1050 -850
rect 1000 -890 1010 -860
rect 1040 -890 1050 -860
rect 1000 -900 1050 -890
rect 1300 -860 1350 -850
rect 1300 -890 1310 -860
rect 1340 -890 1350 -860
rect 1300 -900 1350 -890
rect 1600 -860 1650 -850
rect 1600 -890 1610 -860
rect 1640 -890 1650 -860
rect 1600 -900 1650 -890
rect 1900 -860 1950 -850
rect 1900 -890 1910 -860
rect 1940 -890 1950 -860
rect 1900 -900 1950 -890
rect 2200 -860 2250 -850
rect 2200 -890 2210 -860
rect 2240 -890 2250 -860
rect 2200 -900 2250 -890
rect 2350 -860 2400 -800
rect 2350 -890 2360 -860
rect 2390 -890 2400 -860
rect 2350 -950 2400 -890
rect 2500 -860 2550 -850
rect 2500 -890 2510 -860
rect 2540 -890 2550 -860
rect 2500 -900 2550 -890
rect 2800 -860 2850 -850
rect 2800 -890 2810 -860
rect 2840 -890 2850 -860
rect 2800 -900 2850 -890
rect 3100 -860 3150 -850
rect 3100 -890 3110 -860
rect 3140 -890 3150 -860
rect 3100 -900 3150 -890
rect 3400 -860 3450 -850
rect 3400 -890 3410 -860
rect 3440 -890 3450 -860
rect 3400 -900 3450 -890
rect 3700 -860 3750 -850
rect 3700 -890 3710 -860
rect 3740 -890 3750 -860
rect 3700 -900 3750 -890
rect 3850 -860 3900 -800
rect 3850 -890 3860 -860
rect 3890 -890 3900 -860
rect 3850 -950 3900 -890
rect 4000 -860 4050 -850
rect 4000 -890 4010 -860
rect 4040 -890 4050 -860
rect 4000 -900 4050 -890
rect 4300 -860 4350 -850
rect 4300 -890 4310 -860
rect 4340 -890 4350 -860
rect 4300 -900 4350 -890
rect 4450 -860 4500 -800
rect 4450 -890 4460 -860
rect 4490 -890 4500 -860
rect 4450 -950 4500 -890
rect 4600 -860 4650 -850
rect 4600 -890 4610 -860
rect 4640 -890 4650 -860
rect 4600 -900 4650 -890
rect 4900 -860 4950 -850
rect 4900 -890 4910 -860
rect 4940 -890 4950 -860
rect 4900 -900 4950 -890
rect 5200 -860 5250 -850
rect 5200 -890 5210 -860
rect 5240 -890 5250 -860
rect 5200 -900 5250 -890
rect 5500 -860 5550 -850
rect 5500 -890 5510 -860
rect 5540 -890 5550 -860
rect 5500 -900 5550 -890
rect 5800 -860 5850 -850
rect 5800 -890 5810 -860
rect 5840 -890 5850 -860
rect 5800 -900 5850 -890
rect 5950 -860 6000 -800
rect 5950 -890 5960 -860
rect 5990 -890 6000 -860
rect 5950 -950 6000 -890
rect 6100 -860 6150 -850
rect 6100 -890 6110 -860
rect 6140 -890 6150 -860
rect 6100 -900 6150 -890
rect 6400 -860 6450 -850
rect 6400 -890 6410 -860
rect 6440 -890 6450 -860
rect 6400 -900 6450 -890
rect 6700 -860 6750 -850
rect 6700 -890 6710 -860
rect 6740 -890 6750 -860
rect 6700 -900 6750 -890
rect 7000 -860 7050 -850
rect 7000 -890 7010 -860
rect 7040 -890 7050 -860
rect 7000 -900 7050 -890
rect 7300 -860 7350 -850
rect 7300 -890 7310 -860
rect 7340 -890 7350 -860
rect 7300 -900 7350 -890
rect 7600 -860 7650 -850
rect 7600 -890 7610 -860
rect 7640 -890 7650 -860
rect 7600 -900 7650 -890
rect 7900 -860 7950 -850
rect 7900 -890 7910 -860
rect 7940 -890 7950 -860
rect 7900 -900 7950 -890
rect 8200 -860 8250 -850
rect 8200 -890 8210 -860
rect 8240 -890 8250 -860
rect 8200 -900 8250 -890
rect -50 -990 -40 -960
rect -10 -990 0 -960
rect -50 -1015 0 -990
rect -50 -1035 -35 -1015
rect -15 -1035 0 -1015
rect -50 -1060 0 -1035
rect -50 -1090 -40 -1060
rect -10 -1090 0 -1060
rect -50 -1115 0 -1090
rect -50 -1135 -35 -1115
rect -15 -1135 0 -1115
rect -50 -1160 0 -1135
rect -50 -1190 -40 -1160
rect -10 -1190 0 -1160
rect -50 -1215 0 -1190
rect -50 -1235 -35 -1215
rect -15 -1235 0 -1215
rect -50 -1260 0 -1235
rect -50 -1290 -40 -1260
rect -10 -1290 0 -1260
rect -50 -1315 0 -1290
rect -50 -1335 -35 -1315
rect -15 -1335 0 -1315
rect -50 -1360 0 -1335
rect -50 -1390 -40 -1360
rect -10 -1390 0 -1360
rect -50 -1415 0 -1390
rect -50 -1435 -35 -1415
rect -15 -1435 0 -1415
rect -50 -1460 0 -1435
rect -50 -1490 -40 -1460
rect -10 -1490 0 -1460
rect -50 -1515 0 -1490
rect -50 -1535 -35 -1515
rect -15 -1535 0 -1515
rect -50 -1560 0 -1535
rect -50 -1590 -40 -1560
rect -10 -1590 0 -1560
rect -50 -1615 0 -1590
rect -50 -1635 -35 -1615
rect -15 -1635 0 -1615
rect -650 -1740 -640 -1710
rect -610 -1740 -600 -1710
rect -650 -1750 -600 -1740
rect -50 -1710 0 -1635
rect 1150 -965 1200 -950
rect 1150 -985 1165 -965
rect 1185 -985 1200 -965
rect 1150 -1015 1200 -985
rect 1150 -1035 1165 -1015
rect 1185 -1035 1200 -1015
rect 1150 -1065 1200 -1035
rect 1150 -1085 1165 -1065
rect 1185 -1085 1200 -1065
rect 1150 -1115 1200 -1085
rect 1150 -1135 1165 -1115
rect 1185 -1135 1200 -1115
rect 1150 -1165 1200 -1135
rect 1150 -1185 1165 -1165
rect 1185 -1185 1200 -1165
rect 1150 -1215 1200 -1185
rect 1150 -1235 1165 -1215
rect 1185 -1235 1200 -1215
rect 1150 -1265 1200 -1235
rect 1150 -1285 1165 -1265
rect 1185 -1285 1200 -1265
rect 1150 -1315 1200 -1285
rect 1150 -1335 1165 -1315
rect 1185 -1335 1200 -1315
rect 1150 -1365 1200 -1335
rect 1150 -1385 1165 -1365
rect 1185 -1385 1200 -1365
rect 1150 -1415 1200 -1385
rect 1150 -1435 1165 -1415
rect 1185 -1435 1200 -1415
rect 1150 -1465 1200 -1435
rect 1150 -1485 1165 -1465
rect 1185 -1485 1200 -1465
rect 1150 -1515 1200 -1485
rect 1150 -1535 1165 -1515
rect 1185 -1535 1200 -1515
rect 1150 -1565 1200 -1535
rect 1450 -965 3300 -950
rect 1450 -985 1465 -965
rect 1485 -985 2065 -965
rect 2085 -985 2665 -965
rect 2685 -985 3265 -965
rect 3285 -985 3300 -965
rect 1450 -1000 3300 -985
rect 1450 -1015 1500 -1000
rect 1450 -1035 1465 -1015
rect 1485 -1035 1500 -1015
rect 1450 -1065 1500 -1035
rect 2050 -1015 2100 -1000
rect 2050 -1035 2065 -1015
rect 2085 -1035 2100 -1015
rect 1450 -1085 1465 -1065
rect 1485 -1085 1500 -1065
rect 1450 -1115 1500 -1085
rect 1450 -1135 1465 -1115
rect 1485 -1135 1500 -1115
rect 1450 -1165 1500 -1135
rect 1450 -1185 1465 -1165
rect 1485 -1185 1500 -1165
rect 1450 -1215 1500 -1185
rect 1450 -1235 1465 -1215
rect 1485 -1235 1500 -1215
rect 1450 -1265 1500 -1235
rect 1450 -1285 1465 -1265
rect 1485 -1285 1500 -1265
rect 1450 -1315 1500 -1285
rect 1450 -1335 1465 -1315
rect 1485 -1335 1500 -1315
rect 1450 -1365 1500 -1335
rect 1450 -1385 1465 -1365
rect 1485 -1385 1500 -1365
rect 1450 -1415 1500 -1385
rect 1450 -1435 1465 -1415
rect 1485 -1435 1500 -1415
rect 1450 -1465 1500 -1435
rect 1450 -1485 1465 -1465
rect 1485 -1485 1500 -1465
rect 1450 -1515 1500 -1485
rect 1450 -1535 1465 -1515
rect 1485 -1535 1500 -1515
rect 1450 -1550 1500 -1535
rect 1750 -1065 1800 -1050
rect 1750 -1085 1765 -1065
rect 1785 -1085 1800 -1065
rect 1750 -1115 1800 -1085
rect 1750 -1135 1765 -1115
rect 1785 -1135 1800 -1115
rect 1750 -1165 1800 -1135
rect 1750 -1185 1765 -1165
rect 1785 -1185 1800 -1165
rect 1750 -1215 1800 -1185
rect 1750 -1235 1765 -1215
rect 1785 -1235 1800 -1215
rect 1750 -1265 1800 -1235
rect 1750 -1285 1765 -1265
rect 1785 -1285 1800 -1265
rect 1750 -1315 1800 -1285
rect 1750 -1335 1765 -1315
rect 1785 -1335 1800 -1315
rect 1750 -1365 1800 -1335
rect 1750 -1385 1765 -1365
rect 1785 -1385 1800 -1365
rect 1750 -1415 1800 -1385
rect 1750 -1435 1765 -1415
rect 1785 -1435 1800 -1415
rect 1750 -1465 1800 -1435
rect 1750 -1485 1765 -1465
rect 1785 -1485 1800 -1465
rect 1750 -1515 1800 -1485
rect 1750 -1535 1765 -1515
rect 1785 -1535 1800 -1515
rect 1150 -1585 1165 -1565
rect 1185 -1585 1200 -1565
rect 1150 -1600 1200 -1585
rect 1750 -1565 1800 -1535
rect 2050 -1065 2100 -1035
rect 2650 -1015 2700 -1000
rect 2650 -1035 2665 -1015
rect 2685 -1035 2700 -1015
rect 2050 -1085 2065 -1065
rect 2085 -1085 2100 -1065
rect 2050 -1115 2100 -1085
rect 2050 -1135 2065 -1115
rect 2085 -1135 2100 -1115
rect 2050 -1165 2100 -1135
rect 2050 -1185 2065 -1165
rect 2085 -1185 2100 -1165
rect 2050 -1215 2100 -1185
rect 2050 -1235 2065 -1215
rect 2085 -1235 2100 -1215
rect 2050 -1265 2100 -1235
rect 2050 -1285 2065 -1265
rect 2085 -1285 2100 -1265
rect 2050 -1315 2100 -1285
rect 2050 -1335 2065 -1315
rect 2085 -1335 2100 -1315
rect 2050 -1365 2100 -1335
rect 2050 -1385 2065 -1365
rect 2085 -1385 2100 -1365
rect 2050 -1415 2100 -1385
rect 2050 -1435 2065 -1415
rect 2085 -1435 2100 -1415
rect 2050 -1465 2100 -1435
rect 2050 -1485 2065 -1465
rect 2085 -1485 2100 -1465
rect 2050 -1515 2100 -1485
rect 2050 -1535 2065 -1515
rect 2085 -1535 2100 -1515
rect 2050 -1550 2100 -1535
rect 2350 -1065 2400 -1050
rect 2350 -1085 2365 -1065
rect 2385 -1085 2400 -1065
rect 2350 -1115 2400 -1085
rect 2350 -1135 2365 -1115
rect 2385 -1135 2400 -1115
rect 2350 -1165 2400 -1135
rect 2350 -1185 2365 -1165
rect 2385 -1185 2400 -1165
rect 2350 -1215 2400 -1185
rect 2350 -1235 2365 -1215
rect 2385 -1235 2400 -1215
rect 2350 -1265 2400 -1235
rect 2350 -1285 2365 -1265
rect 2385 -1285 2400 -1265
rect 2350 -1315 2400 -1285
rect 2350 -1335 2365 -1315
rect 2385 -1335 2400 -1315
rect 2350 -1365 2400 -1335
rect 2350 -1385 2365 -1365
rect 2385 -1385 2400 -1365
rect 2350 -1415 2400 -1385
rect 2350 -1435 2365 -1415
rect 2385 -1435 2400 -1415
rect 2350 -1465 2400 -1435
rect 2350 -1485 2365 -1465
rect 2385 -1485 2400 -1465
rect 2350 -1515 2400 -1485
rect 2350 -1535 2365 -1515
rect 2385 -1535 2400 -1515
rect 1750 -1585 1765 -1565
rect 1785 -1585 1800 -1565
rect 1750 -1600 1800 -1585
rect 2350 -1565 2400 -1535
rect 2650 -1065 2700 -1035
rect 3250 -1015 3300 -1000
rect 3250 -1035 3265 -1015
rect 3285 -1035 3300 -1015
rect 2650 -1085 2665 -1065
rect 2685 -1085 2700 -1065
rect 2650 -1115 2700 -1085
rect 2650 -1135 2665 -1115
rect 2685 -1135 2700 -1115
rect 2650 -1165 2700 -1135
rect 2650 -1185 2665 -1165
rect 2685 -1185 2700 -1165
rect 2650 -1215 2700 -1185
rect 2650 -1235 2665 -1215
rect 2685 -1235 2700 -1215
rect 2650 -1265 2700 -1235
rect 2650 -1285 2665 -1265
rect 2685 -1285 2700 -1265
rect 2650 -1315 2700 -1285
rect 2650 -1335 2665 -1315
rect 2685 -1335 2700 -1315
rect 2650 -1365 2700 -1335
rect 2650 -1385 2665 -1365
rect 2685 -1385 2700 -1365
rect 2650 -1415 2700 -1385
rect 2650 -1435 2665 -1415
rect 2685 -1435 2700 -1415
rect 2650 -1465 2700 -1435
rect 2650 -1485 2665 -1465
rect 2685 -1485 2700 -1465
rect 2650 -1515 2700 -1485
rect 2650 -1535 2665 -1515
rect 2685 -1535 2700 -1515
rect 2650 -1550 2700 -1535
rect 2950 -1065 3000 -1050
rect 2950 -1085 2965 -1065
rect 2985 -1085 3000 -1065
rect 2950 -1115 3000 -1085
rect 2950 -1135 2965 -1115
rect 2985 -1135 3000 -1115
rect 2950 -1165 3000 -1135
rect 2950 -1185 2965 -1165
rect 2985 -1185 3000 -1165
rect 2950 -1215 3000 -1185
rect 2950 -1235 2965 -1215
rect 2985 -1235 3000 -1215
rect 2950 -1265 3000 -1235
rect 2950 -1285 2965 -1265
rect 2985 -1285 3000 -1265
rect 2950 -1315 3000 -1285
rect 2950 -1335 2965 -1315
rect 2985 -1335 3000 -1315
rect 2950 -1365 3000 -1335
rect 2950 -1385 2965 -1365
rect 2985 -1385 3000 -1365
rect 2950 -1415 3000 -1385
rect 2950 -1435 2965 -1415
rect 2985 -1435 3000 -1415
rect 2950 -1465 3000 -1435
rect 2950 -1485 2965 -1465
rect 2985 -1485 3000 -1465
rect 2950 -1515 3000 -1485
rect 2950 -1535 2965 -1515
rect 2985 -1535 3000 -1515
rect 2350 -1585 2365 -1565
rect 2385 -1585 2400 -1565
rect 2350 -1600 2400 -1585
rect 2950 -1565 3000 -1535
rect 3250 -1065 3300 -1035
rect 3250 -1085 3265 -1065
rect 3285 -1085 3300 -1065
rect 3250 -1115 3300 -1085
rect 3250 -1135 3265 -1115
rect 3285 -1135 3300 -1115
rect 3250 -1165 3300 -1135
rect 3250 -1185 3265 -1165
rect 3285 -1185 3300 -1165
rect 3250 -1215 3300 -1185
rect 3250 -1235 3265 -1215
rect 3285 -1235 3300 -1215
rect 3250 -1265 3300 -1235
rect 3250 -1285 3265 -1265
rect 3285 -1285 3300 -1265
rect 3250 -1315 3300 -1285
rect 3250 -1335 3265 -1315
rect 3285 -1335 3300 -1315
rect 3250 -1365 3300 -1335
rect 3250 -1385 3265 -1365
rect 3285 -1385 3300 -1365
rect 3250 -1415 3300 -1385
rect 3250 -1435 3265 -1415
rect 3285 -1435 3300 -1415
rect 3250 -1465 3300 -1435
rect 3250 -1485 3265 -1465
rect 3285 -1485 3300 -1465
rect 3250 -1515 3300 -1485
rect 3250 -1535 3265 -1515
rect 3285 -1535 3300 -1515
rect 3250 -1550 3300 -1535
rect 3550 -965 3600 -950
rect 3550 -985 3565 -965
rect 3585 -985 3600 -965
rect 3550 -1015 3600 -985
rect 3550 -1035 3565 -1015
rect 3585 -1035 3600 -1015
rect 3550 -1065 3600 -1035
rect 3550 -1085 3565 -1065
rect 3585 -1085 3600 -1065
rect 3550 -1115 3600 -1085
rect 3550 -1135 3565 -1115
rect 3585 -1135 3600 -1115
rect 3550 -1165 3600 -1135
rect 3550 -1185 3565 -1165
rect 3585 -1185 3600 -1165
rect 3550 -1215 3600 -1185
rect 3550 -1235 3565 -1215
rect 3585 -1235 3600 -1215
rect 3550 -1265 3600 -1235
rect 3550 -1285 3565 -1265
rect 3585 -1285 3600 -1265
rect 3550 -1315 3600 -1285
rect 3550 -1335 3565 -1315
rect 3585 -1335 3600 -1315
rect 3550 -1365 3600 -1335
rect 3550 -1385 3565 -1365
rect 3585 -1385 3600 -1365
rect 3550 -1415 3600 -1385
rect 3550 -1435 3565 -1415
rect 3585 -1435 3600 -1415
rect 3550 -1465 3600 -1435
rect 3550 -1485 3565 -1465
rect 3585 -1485 3600 -1465
rect 3550 -1515 3600 -1485
rect 3550 -1535 3565 -1515
rect 3585 -1535 3600 -1515
rect 2950 -1585 2965 -1565
rect 2985 -1585 3000 -1565
rect 2950 -1600 3000 -1585
rect 3550 -1565 3600 -1535
rect 3700 -965 4050 -950
rect 3700 -985 3715 -965
rect 3735 -985 4015 -965
rect 4035 -985 4050 -965
rect 3700 -1000 4050 -985
rect 3700 -1015 3750 -1000
rect 3700 -1035 3715 -1015
rect 3735 -1035 3750 -1015
rect 3700 -1065 3750 -1035
rect 4000 -1015 4050 -1000
rect 4000 -1035 4015 -1015
rect 4035 -1035 4050 -1015
rect 3700 -1085 3715 -1065
rect 3735 -1085 3750 -1065
rect 3700 -1115 3750 -1085
rect 3700 -1135 3715 -1115
rect 3735 -1135 3750 -1115
rect 3700 -1165 3750 -1135
rect 3700 -1185 3715 -1165
rect 3735 -1185 3750 -1165
rect 3700 -1215 3750 -1185
rect 3700 -1235 3715 -1215
rect 3735 -1235 3750 -1215
rect 3700 -1265 3750 -1235
rect 3700 -1285 3715 -1265
rect 3735 -1285 3750 -1265
rect 3700 -1315 3750 -1285
rect 3700 -1335 3715 -1315
rect 3735 -1335 3750 -1315
rect 3700 -1365 3750 -1335
rect 3700 -1385 3715 -1365
rect 3735 -1385 3750 -1365
rect 3700 -1415 3750 -1385
rect 3700 -1435 3715 -1415
rect 3735 -1435 3750 -1415
rect 3700 -1465 3750 -1435
rect 3700 -1485 3715 -1465
rect 3735 -1485 3750 -1465
rect 3700 -1515 3750 -1485
rect 3700 -1535 3715 -1515
rect 3735 -1535 3750 -1515
rect 3700 -1550 3750 -1535
rect 3850 -1065 3900 -1050
rect 3850 -1085 3865 -1065
rect 3885 -1085 3900 -1065
rect 3850 -1115 3900 -1085
rect 3850 -1135 3865 -1115
rect 3885 -1135 3900 -1115
rect 3850 -1165 3900 -1135
rect 3850 -1185 3865 -1165
rect 3885 -1185 3900 -1165
rect 3850 -1215 3900 -1185
rect 3850 -1235 3865 -1215
rect 3885 -1235 3900 -1215
rect 3850 -1265 3900 -1235
rect 3850 -1285 3865 -1265
rect 3885 -1285 3900 -1265
rect 3850 -1315 3900 -1285
rect 3850 -1335 3865 -1315
rect 3885 -1335 3900 -1315
rect 3850 -1365 3900 -1335
rect 3850 -1385 3865 -1365
rect 3885 -1385 3900 -1365
rect 3850 -1415 3900 -1385
rect 3850 -1435 3865 -1415
rect 3885 -1435 3900 -1415
rect 3850 -1465 3900 -1435
rect 3850 -1485 3865 -1465
rect 3885 -1485 3900 -1465
rect 3850 -1515 3900 -1485
rect 3850 -1535 3865 -1515
rect 3885 -1535 3900 -1515
rect 3550 -1585 3565 -1565
rect 3585 -1585 3600 -1565
rect 3550 -1600 3600 -1585
rect 3850 -1565 3900 -1535
rect 4000 -1065 4050 -1035
rect 4000 -1085 4015 -1065
rect 4035 -1085 4050 -1065
rect 4000 -1115 4050 -1085
rect 4000 -1135 4015 -1115
rect 4035 -1135 4050 -1115
rect 4000 -1165 4050 -1135
rect 4000 -1185 4015 -1165
rect 4035 -1185 4050 -1165
rect 4000 -1215 4050 -1185
rect 4000 -1235 4015 -1215
rect 4035 -1235 4050 -1215
rect 4000 -1265 4050 -1235
rect 4000 -1285 4015 -1265
rect 4035 -1285 4050 -1265
rect 4000 -1315 4050 -1285
rect 4000 -1335 4015 -1315
rect 4035 -1335 4050 -1315
rect 4000 -1365 4050 -1335
rect 4000 -1385 4015 -1365
rect 4035 -1385 4050 -1365
rect 4000 -1415 4050 -1385
rect 4000 -1435 4015 -1415
rect 4035 -1435 4050 -1415
rect 4000 -1465 4050 -1435
rect 4000 -1485 4015 -1465
rect 4035 -1485 4050 -1465
rect 4000 -1515 4050 -1485
rect 4000 -1535 4015 -1515
rect 4035 -1535 4050 -1515
rect 4000 -1550 4050 -1535
rect 4150 -965 4200 -950
rect 4150 -985 4165 -965
rect 4185 -985 4200 -965
rect 4150 -1015 4200 -985
rect 4150 -1035 4165 -1015
rect 4185 -1035 4200 -1015
rect 4150 -1065 4200 -1035
rect 4150 -1085 4165 -1065
rect 4185 -1085 4200 -1065
rect 4150 -1115 4200 -1085
rect 4150 -1135 4165 -1115
rect 4185 -1135 4200 -1115
rect 4150 -1165 4200 -1135
rect 4150 -1185 4165 -1165
rect 4185 -1185 4200 -1165
rect 4150 -1215 4200 -1185
rect 4150 -1235 4165 -1215
rect 4185 -1235 4200 -1215
rect 4150 -1265 4200 -1235
rect 4150 -1285 4165 -1265
rect 4185 -1285 4200 -1265
rect 4150 -1315 4200 -1285
rect 4150 -1335 4165 -1315
rect 4185 -1335 4200 -1315
rect 4150 -1365 4200 -1335
rect 4150 -1385 4165 -1365
rect 4185 -1385 4200 -1365
rect 4150 -1415 4200 -1385
rect 4150 -1435 4165 -1415
rect 4185 -1435 4200 -1415
rect 4150 -1465 4200 -1435
rect 4150 -1485 4165 -1465
rect 4185 -1485 4200 -1465
rect 4150 -1515 4200 -1485
rect 4150 -1535 4165 -1515
rect 4185 -1535 4200 -1515
rect 3850 -1585 3865 -1565
rect 3885 -1585 3900 -1565
rect 3850 -1600 3900 -1585
rect 4150 -1565 4200 -1535
rect 4300 -965 4650 -950
rect 4300 -985 4315 -965
rect 4335 -985 4615 -965
rect 4635 -985 4650 -965
rect 4300 -1000 4650 -985
rect 4300 -1015 4350 -1000
rect 4300 -1035 4315 -1015
rect 4335 -1035 4350 -1015
rect 4300 -1065 4350 -1035
rect 4600 -1015 4650 -1000
rect 4600 -1035 4615 -1015
rect 4635 -1035 4650 -1015
rect 4300 -1085 4315 -1065
rect 4335 -1085 4350 -1065
rect 4300 -1115 4350 -1085
rect 4300 -1135 4315 -1115
rect 4335 -1135 4350 -1115
rect 4300 -1165 4350 -1135
rect 4300 -1185 4315 -1165
rect 4335 -1185 4350 -1165
rect 4300 -1215 4350 -1185
rect 4300 -1235 4315 -1215
rect 4335 -1235 4350 -1215
rect 4300 -1265 4350 -1235
rect 4300 -1285 4315 -1265
rect 4335 -1285 4350 -1265
rect 4300 -1315 4350 -1285
rect 4300 -1335 4315 -1315
rect 4335 -1335 4350 -1315
rect 4300 -1365 4350 -1335
rect 4300 -1385 4315 -1365
rect 4335 -1385 4350 -1365
rect 4300 -1415 4350 -1385
rect 4300 -1435 4315 -1415
rect 4335 -1435 4350 -1415
rect 4300 -1465 4350 -1435
rect 4300 -1485 4315 -1465
rect 4335 -1485 4350 -1465
rect 4300 -1515 4350 -1485
rect 4300 -1535 4315 -1515
rect 4335 -1535 4350 -1515
rect 4300 -1550 4350 -1535
rect 4450 -1065 4500 -1050
rect 4450 -1085 4465 -1065
rect 4485 -1085 4500 -1065
rect 4450 -1115 4500 -1085
rect 4450 -1135 4465 -1115
rect 4485 -1135 4500 -1115
rect 4450 -1165 4500 -1135
rect 4450 -1185 4465 -1165
rect 4485 -1185 4500 -1165
rect 4450 -1215 4500 -1185
rect 4450 -1235 4465 -1215
rect 4485 -1235 4500 -1215
rect 4450 -1265 4500 -1235
rect 4450 -1285 4465 -1265
rect 4485 -1285 4500 -1265
rect 4450 -1315 4500 -1285
rect 4450 -1335 4465 -1315
rect 4485 -1335 4500 -1315
rect 4450 -1365 4500 -1335
rect 4450 -1385 4465 -1365
rect 4485 -1385 4500 -1365
rect 4450 -1415 4500 -1385
rect 4450 -1435 4465 -1415
rect 4485 -1435 4500 -1415
rect 4450 -1465 4500 -1435
rect 4450 -1485 4465 -1465
rect 4485 -1485 4500 -1465
rect 4450 -1515 4500 -1485
rect 4450 -1535 4465 -1515
rect 4485 -1535 4500 -1515
rect 4150 -1585 4165 -1565
rect 4185 -1585 4200 -1565
rect 4150 -1600 4200 -1585
rect 4450 -1565 4500 -1535
rect 4600 -1065 4650 -1035
rect 4600 -1085 4615 -1065
rect 4635 -1085 4650 -1065
rect 4600 -1115 4650 -1085
rect 4600 -1135 4615 -1115
rect 4635 -1135 4650 -1115
rect 4600 -1165 4650 -1135
rect 4600 -1185 4615 -1165
rect 4635 -1185 4650 -1165
rect 4600 -1215 4650 -1185
rect 4600 -1235 4615 -1215
rect 4635 -1235 4650 -1215
rect 4600 -1265 4650 -1235
rect 4600 -1285 4615 -1265
rect 4635 -1285 4650 -1265
rect 4600 -1315 4650 -1285
rect 4600 -1335 4615 -1315
rect 4635 -1335 4650 -1315
rect 4600 -1365 4650 -1335
rect 4600 -1385 4615 -1365
rect 4635 -1385 4650 -1365
rect 4600 -1415 4650 -1385
rect 4600 -1435 4615 -1415
rect 4635 -1435 4650 -1415
rect 4600 -1465 4650 -1435
rect 4600 -1485 4615 -1465
rect 4635 -1485 4650 -1465
rect 4600 -1515 4650 -1485
rect 4600 -1535 4615 -1515
rect 4635 -1535 4650 -1515
rect 4600 -1550 4650 -1535
rect 4750 -965 4800 -950
rect 4750 -985 4765 -965
rect 4785 -985 4800 -965
rect 4750 -1015 4800 -985
rect 4750 -1035 4765 -1015
rect 4785 -1035 4800 -1015
rect 4750 -1065 4800 -1035
rect 4750 -1085 4765 -1065
rect 4785 -1085 4800 -1065
rect 4750 -1115 4800 -1085
rect 4750 -1135 4765 -1115
rect 4785 -1135 4800 -1115
rect 4750 -1165 4800 -1135
rect 4750 -1185 4765 -1165
rect 4785 -1185 4800 -1165
rect 4750 -1215 4800 -1185
rect 4750 -1235 4765 -1215
rect 4785 -1235 4800 -1215
rect 4750 -1265 4800 -1235
rect 4750 -1285 4765 -1265
rect 4785 -1285 4800 -1265
rect 4750 -1315 4800 -1285
rect 4750 -1335 4765 -1315
rect 4785 -1335 4800 -1315
rect 4750 -1365 4800 -1335
rect 4750 -1385 4765 -1365
rect 4785 -1385 4800 -1365
rect 4750 -1415 4800 -1385
rect 4750 -1435 4765 -1415
rect 4785 -1435 4800 -1415
rect 4750 -1465 4800 -1435
rect 4750 -1485 4765 -1465
rect 4785 -1485 4800 -1465
rect 4750 -1515 4800 -1485
rect 4750 -1535 4765 -1515
rect 4785 -1535 4800 -1515
rect 4450 -1585 4465 -1565
rect 4485 -1585 4500 -1565
rect 4450 -1600 4500 -1585
rect 4750 -1565 4800 -1535
rect 5050 -965 6900 -950
rect 5050 -985 5065 -965
rect 5085 -985 5665 -965
rect 5685 -985 6265 -965
rect 6285 -985 6865 -965
rect 6885 -985 6900 -965
rect 5050 -1000 6900 -985
rect 5050 -1015 5100 -1000
rect 5050 -1035 5065 -1015
rect 5085 -1035 5100 -1015
rect 5050 -1065 5100 -1035
rect 5650 -1015 5700 -1000
rect 5650 -1035 5665 -1015
rect 5685 -1035 5700 -1015
rect 5050 -1085 5065 -1065
rect 5085 -1085 5100 -1065
rect 5050 -1115 5100 -1085
rect 5050 -1135 5065 -1115
rect 5085 -1135 5100 -1115
rect 5050 -1165 5100 -1135
rect 5050 -1185 5065 -1165
rect 5085 -1185 5100 -1165
rect 5050 -1215 5100 -1185
rect 5050 -1235 5065 -1215
rect 5085 -1235 5100 -1215
rect 5050 -1265 5100 -1235
rect 5050 -1285 5065 -1265
rect 5085 -1285 5100 -1265
rect 5050 -1315 5100 -1285
rect 5050 -1335 5065 -1315
rect 5085 -1335 5100 -1315
rect 5050 -1365 5100 -1335
rect 5050 -1385 5065 -1365
rect 5085 -1385 5100 -1365
rect 5050 -1415 5100 -1385
rect 5050 -1435 5065 -1415
rect 5085 -1435 5100 -1415
rect 5050 -1465 5100 -1435
rect 5050 -1485 5065 -1465
rect 5085 -1485 5100 -1465
rect 5050 -1515 5100 -1485
rect 5050 -1535 5065 -1515
rect 5085 -1535 5100 -1515
rect 5050 -1550 5100 -1535
rect 5350 -1065 5400 -1050
rect 5350 -1085 5365 -1065
rect 5385 -1085 5400 -1065
rect 5350 -1115 5400 -1085
rect 5350 -1135 5365 -1115
rect 5385 -1135 5400 -1115
rect 5350 -1165 5400 -1135
rect 5350 -1185 5365 -1165
rect 5385 -1185 5400 -1165
rect 5350 -1215 5400 -1185
rect 5350 -1235 5365 -1215
rect 5385 -1235 5400 -1215
rect 5350 -1265 5400 -1235
rect 5350 -1285 5365 -1265
rect 5385 -1285 5400 -1265
rect 5350 -1315 5400 -1285
rect 5350 -1335 5365 -1315
rect 5385 -1335 5400 -1315
rect 5350 -1365 5400 -1335
rect 5350 -1385 5365 -1365
rect 5385 -1385 5400 -1365
rect 5350 -1415 5400 -1385
rect 5350 -1435 5365 -1415
rect 5385 -1435 5400 -1415
rect 5350 -1465 5400 -1435
rect 5350 -1485 5365 -1465
rect 5385 -1485 5400 -1465
rect 5350 -1515 5400 -1485
rect 5350 -1535 5365 -1515
rect 5385 -1535 5400 -1515
rect 4750 -1585 4765 -1565
rect 4785 -1585 4800 -1565
rect 4750 -1600 4800 -1585
rect 5350 -1565 5400 -1535
rect 5650 -1065 5700 -1035
rect 6250 -1015 6300 -1000
rect 6250 -1035 6265 -1015
rect 6285 -1035 6300 -1015
rect 5650 -1085 5665 -1065
rect 5685 -1085 5700 -1065
rect 5650 -1115 5700 -1085
rect 5650 -1135 5665 -1115
rect 5685 -1135 5700 -1115
rect 5650 -1165 5700 -1135
rect 5650 -1185 5665 -1165
rect 5685 -1185 5700 -1165
rect 5650 -1215 5700 -1185
rect 5650 -1235 5665 -1215
rect 5685 -1235 5700 -1215
rect 5650 -1265 5700 -1235
rect 5650 -1285 5665 -1265
rect 5685 -1285 5700 -1265
rect 5650 -1315 5700 -1285
rect 5650 -1335 5665 -1315
rect 5685 -1335 5700 -1315
rect 5650 -1365 5700 -1335
rect 5650 -1385 5665 -1365
rect 5685 -1385 5700 -1365
rect 5650 -1415 5700 -1385
rect 5650 -1435 5665 -1415
rect 5685 -1435 5700 -1415
rect 5650 -1465 5700 -1435
rect 5650 -1485 5665 -1465
rect 5685 -1485 5700 -1465
rect 5650 -1515 5700 -1485
rect 5650 -1535 5665 -1515
rect 5685 -1535 5700 -1515
rect 5650 -1550 5700 -1535
rect 5950 -1065 6000 -1050
rect 5950 -1085 5965 -1065
rect 5985 -1085 6000 -1065
rect 5950 -1115 6000 -1085
rect 5950 -1135 5965 -1115
rect 5985 -1135 6000 -1115
rect 5950 -1165 6000 -1135
rect 5950 -1185 5965 -1165
rect 5985 -1185 6000 -1165
rect 5950 -1215 6000 -1185
rect 5950 -1235 5965 -1215
rect 5985 -1235 6000 -1215
rect 5950 -1265 6000 -1235
rect 5950 -1285 5965 -1265
rect 5985 -1285 6000 -1265
rect 5950 -1315 6000 -1285
rect 5950 -1335 5965 -1315
rect 5985 -1335 6000 -1315
rect 5950 -1365 6000 -1335
rect 5950 -1385 5965 -1365
rect 5985 -1385 6000 -1365
rect 5950 -1415 6000 -1385
rect 5950 -1435 5965 -1415
rect 5985 -1435 6000 -1415
rect 5950 -1465 6000 -1435
rect 5950 -1485 5965 -1465
rect 5985 -1485 6000 -1465
rect 5950 -1515 6000 -1485
rect 5950 -1535 5965 -1515
rect 5985 -1535 6000 -1515
rect 5350 -1585 5365 -1565
rect 5385 -1585 5400 -1565
rect 5350 -1600 5400 -1585
rect 5950 -1565 6000 -1535
rect 6250 -1065 6300 -1035
rect 6850 -1015 6900 -1000
rect 6850 -1035 6865 -1015
rect 6885 -1035 6900 -1015
rect 6250 -1085 6265 -1065
rect 6285 -1085 6300 -1065
rect 6250 -1115 6300 -1085
rect 6250 -1135 6265 -1115
rect 6285 -1135 6300 -1115
rect 6250 -1165 6300 -1135
rect 6250 -1185 6265 -1165
rect 6285 -1185 6300 -1165
rect 6250 -1215 6300 -1185
rect 6250 -1235 6265 -1215
rect 6285 -1235 6300 -1215
rect 6250 -1265 6300 -1235
rect 6250 -1285 6265 -1265
rect 6285 -1285 6300 -1265
rect 6250 -1315 6300 -1285
rect 6250 -1335 6265 -1315
rect 6285 -1335 6300 -1315
rect 6250 -1365 6300 -1335
rect 6250 -1385 6265 -1365
rect 6285 -1385 6300 -1365
rect 6250 -1415 6300 -1385
rect 6250 -1435 6265 -1415
rect 6285 -1435 6300 -1415
rect 6250 -1465 6300 -1435
rect 6250 -1485 6265 -1465
rect 6285 -1485 6300 -1465
rect 6250 -1515 6300 -1485
rect 6250 -1535 6265 -1515
rect 6285 -1535 6300 -1515
rect 6250 -1550 6300 -1535
rect 6550 -1065 6600 -1050
rect 6550 -1085 6565 -1065
rect 6585 -1085 6600 -1065
rect 6550 -1115 6600 -1085
rect 6550 -1135 6565 -1115
rect 6585 -1135 6600 -1115
rect 6550 -1165 6600 -1135
rect 6550 -1185 6565 -1165
rect 6585 -1185 6600 -1165
rect 6550 -1215 6600 -1185
rect 6550 -1235 6565 -1215
rect 6585 -1235 6600 -1215
rect 6550 -1265 6600 -1235
rect 6550 -1285 6565 -1265
rect 6585 -1285 6600 -1265
rect 6550 -1315 6600 -1285
rect 6550 -1335 6565 -1315
rect 6585 -1335 6600 -1315
rect 6550 -1365 6600 -1335
rect 6550 -1385 6565 -1365
rect 6585 -1385 6600 -1365
rect 6550 -1415 6600 -1385
rect 6550 -1435 6565 -1415
rect 6585 -1435 6600 -1415
rect 6550 -1465 6600 -1435
rect 6550 -1485 6565 -1465
rect 6585 -1485 6600 -1465
rect 6550 -1515 6600 -1485
rect 6550 -1535 6565 -1515
rect 6585 -1535 6600 -1515
rect 5950 -1585 5965 -1565
rect 5985 -1585 6000 -1565
rect 5950 -1600 6000 -1585
rect 6550 -1565 6600 -1535
rect 6850 -1065 6900 -1035
rect 6850 -1085 6865 -1065
rect 6885 -1085 6900 -1065
rect 6850 -1115 6900 -1085
rect 6850 -1135 6865 -1115
rect 6885 -1135 6900 -1115
rect 6850 -1165 6900 -1135
rect 6850 -1185 6865 -1165
rect 6885 -1185 6900 -1165
rect 6850 -1215 6900 -1185
rect 6850 -1235 6865 -1215
rect 6885 -1235 6900 -1215
rect 6850 -1265 6900 -1235
rect 6850 -1285 6865 -1265
rect 6885 -1285 6900 -1265
rect 6850 -1315 6900 -1285
rect 6850 -1335 6865 -1315
rect 6885 -1335 6900 -1315
rect 6850 -1365 6900 -1335
rect 6850 -1385 6865 -1365
rect 6885 -1385 6900 -1365
rect 6850 -1415 6900 -1385
rect 6850 -1435 6865 -1415
rect 6885 -1435 6900 -1415
rect 6850 -1465 6900 -1435
rect 6850 -1485 6865 -1465
rect 6885 -1485 6900 -1465
rect 6850 -1515 6900 -1485
rect 6850 -1535 6865 -1515
rect 6885 -1535 6900 -1515
rect 6850 -1550 6900 -1535
rect 7150 -965 7200 -950
rect 7150 -985 7165 -965
rect 7185 -985 7200 -965
rect 7150 -1015 7200 -985
rect 7150 -1035 7165 -1015
rect 7185 -1035 7200 -1015
rect 7150 -1065 7200 -1035
rect 7150 -1085 7165 -1065
rect 7185 -1085 7200 -1065
rect 7150 -1115 7200 -1085
rect 7150 -1135 7165 -1115
rect 7185 -1135 7200 -1115
rect 7150 -1165 7200 -1135
rect 7150 -1185 7165 -1165
rect 7185 -1185 7200 -1165
rect 7150 -1215 7200 -1185
rect 7150 -1235 7165 -1215
rect 7185 -1235 7200 -1215
rect 7150 -1265 7200 -1235
rect 7150 -1285 7165 -1265
rect 7185 -1285 7200 -1265
rect 7150 -1315 7200 -1285
rect 7150 -1335 7165 -1315
rect 7185 -1335 7200 -1315
rect 7150 -1365 7200 -1335
rect 7150 -1385 7165 -1365
rect 7185 -1385 7200 -1365
rect 7150 -1415 7200 -1385
rect 7150 -1435 7165 -1415
rect 7185 -1435 7200 -1415
rect 7150 -1465 7200 -1435
rect 7150 -1485 7165 -1465
rect 7185 -1485 7200 -1465
rect 7150 -1515 7200 -1485
rect 7150 -1535 7165 -1515
rect 7185 -1535 7200 -1515
rect 6550 -1585 6565 -1565
rect 6585 -1585 6600 -1565
rect 6550 -1600 6600 -1585
rect 7150 -1565 7200 -1535
rect 7150 -1585 7165 -1565
rect 7185 -1585 7200 -1565
rect 7150 -1600 7200 -1585
rect 1150 -1615 7200 -1600
rect 1150 -1635 1165 -1615
rect 1185 -1635 1765 -1615
rect 1785 -1635 2365 -1615
rect 2385 -1635 2965 -1615
rect 2985 -1635 3565 -1615
rect 3585 -1635 3865 -1615
rect 3885 -1635 4165 -1615
rect 4185 -1635 4465 -1615
rect 4485 -1635 4765 -1615
rect 4785 -1635 5365 -1615
rect 5385 -1635 5965 -1615
rect 5985 -1635 6565 -1615
rect 6585 -1635 7165 -1615
rect 7185 -1635 7200 -1615
rect 1150 -1650 7200 -1635
rect 8350 -960 8400 -790
rect 9550 -115 9600 -100
rect 9550 -135 9565 -115
rect 9585 -135 9600 -115
rect 9550 -165 9600 -135
rect 9550 -185 9565 -165
rect 9585 -185 9600 -165
rect 9550 -215 9600 -185
rect 9550 -235 9565 -215
rect 9585 -235 9600 -215
rect 9550 -265 9600 -235
rect 9550 -285 9565 -265
rect 9585 -285 9600 -265
rect 9550 -315 9600 -285
rect 9550 -335 9565 -315
rect 9585 -335 9600 -315
rect 9550 -365 9600 -335
rect 9550 -385 9565 -365
rect 9585 -385 9600 -365
rect 9550 -415 9600 -385
rect 9550 -435 9565 -415
rect 9585 -435 9600 -415
rect 9550 -465 9600 -435
rect 9550 -485 9565 -465
rect 9585 -485 9600 -465
rect 9550 -515 9600 -485
rect 9550 -535 9565 -515
rect 9585 -535 9600 -515
rect 9550 -565 9600 -535
rect 9550 -585 9565 -565
rect 9585 -585 9600 -565
rect 9550 -615 9600 -585
rect 9550 -635 9565 -615
rect 9585 -635 9600 -615
rect 9550 -665 9600 -635
rect 9550 -685 9565 -665
rect 9585 -685 9600 -665
rect 9550 -715 9600 -685
rect 9550 -735 9565 -715
rect 9585 -735 9600 -715
rect 9550 -765 9600 -735
rect 9550 -785 9565 -765
rect 9585 -785 9600 -765
rect 8500 -860 8550 -850
rect 8500 -890 8510 -860
rect 8540 -890 8550 -860
rect 8500 -900 8550 -890
rect 8800 -860 8850 -850
rect 8800 -890 8810 -860
rect 8840 -890 8850 -860
rect 8800 -900 8850 -890
rect 9100 -860 9150 -850
rect 9100 -890 9110 -860
rect 9140 -890 9150 -860
rect 9100 -900 9150 -890
rect 9400 -860 9450 -850
rect 9400 -890 9410 -860
rect 9440 -890 9450 -860
rect 9400 -900 9450 -890
rect 9550 -860 9600 -785
rect 10750 -115 10800 -40
rect 10750 -135 10765 -115
rect 10785 -135 10800 -115
rect 10750 -160 10800 -135
rect 10750 -190 10760 -160
rect 10790 -190 10800 -160
rect 10750 -215 10800 -190
rect 10750 -235 10765 -215
rect 10785 -235 10800 -215
rect 10750 -260 10800 -235
rect 10750 -290 10760 -260
rect 10790 -290 10800 -260
rect 10750 -315 10800 -290
rect 10750 -335 10765 -315
rect 10785 -335 10800 -315
rect 10750 -360 10800 -335
rect 10750 -390 10760 -360
rect 10790 -390 10800 -360
rect 10750 -415 10800 -390
rect 10750 -435 10765 -415
rect 10785 -435 10800 -415
rect 10750 -460 10800 -435
rect 10750 -490 10760 -460
rect 10790 -490 10800 -460
rect 10750 -515 10800 -490
rect 10750 -535 10765 -515
rect 10785 -535 10800 -515
rect 10750 -560 10800 -535
rect 10750 -590 10760 -560
rect 10790 -590 10800 -560
rect 10750 -615 10800 -590
rect 10750 -635 10765 -615
rect 10785 -635 10800 -615
rect 10750 -660 10800 -635
rect 10750 -690 10760 -660
rect 10790 -690 10800 -660
rect 10750 -715 10800 -690
rect 10750 -735 10765 -715
rect 10785 -735 10800 -715
rect 10750 -760 10800 -735
rect 10750 -790 10760 -760
rect 10790 -790 10800 -760
rect 9550 -890 9560 -860
rect 9590 -890 9600 -860
rect 8350 -990 8360 -960
rect 8390 -990 8400 -960
rect 8350 -1015 8400 -990
rect 8350 -1035 8365 -1015
rect 8385 -1035 8400 -1015
rect 8350 -1060 8400 -1035
rect 8350 -1090 8360 -1060
rect 8390 -1090 8400 -1060
rect 8350 -1115 8400 -1090
rect 8350 -1135 8365 -1115
rect 8385 -1135 8400 -1115
rect 8350 -1160 8400 -1135
rect 8350 -1190 8360 -1160
rect 8390 -1190 8400 -1160
rect 8350 -1215 8400 -1190
rect 8350 -1235 8365 -1215
rect 8385 -1235 8400 -1215
rect 8350 -1260 8400 -1235
rect 8350 -1290 8360 -1260
rect 8390 -1290 8400 -1260
rect 8350 -1315 8400 -1290
rect 8350 -1335 8365 -1315
rect 8385 -1335 8400 -1315
rect 8350 -1360 8400 -1335
rect 8350 -1390 8360 -1360
rect 8390 -1390 8400 -1360
rect 8350 -1415 8400 -1390
rect 8350 -1435 8365 -1415
rect 8385 -1435 8400 -1415
rect 8350 -1460 8400 -1435
rect 8350 -1490 8360 -1460
rect 8390 -1490 8400 -1460
rect 8350 -1515 8400 -1490
rect 8350 -1535 8365 -1515
rect 8385 -1535 8400 -1515
rect 8350 -1560 8400 -1535
rect 8350 -1590 8360 -1560
rect 8390 -1590 8400 -1560
rect 8350 -1615 8400 -1590
rect 8350 -1635 8365 -1615
rect 8385 -1635 8400 -1615
rect -50 -1740 -40 -1710
rect -10 -1740 0 -1710
rect -50 -1750 0 -1740
rect 8350 -1710 8400 -1635
rect 9550 -965 9600 -890
rect 9700 -860 9750 -850
rect 9700 -890 9710 -860
rect 9740 -890 9750 -860
rect 9700 -900 9750 -890
rect 10000 -860 10050 -850
rect 10000 -890 10010 -860
rect 10040 -890 10050 -860
rect 10000 -900 10050 -890
rect 10300 -860 10350 -850
rect 10300 -890 10310 -860
rect 10340 -890 10350 -860
rect 10300 -900 10350 -890
rect 10600 -860 10650 -850
rect 10600 -890 10610 -860
rect 10640 -890 10650 -860
rect 10600 -900 10650 -890
rect 9550 -985 9565 -965
rect 9585 -985 9600 -965
rect 9550 -1015 9600 -985
rect 9550 -1035 9565 -1015
rect 9585 -1035 9600 -1015
rect 9550 -1065 9600 -1035
rect 9550 -1085 9565 -1065
rect 9585 -1085 9600 -1065
rect 9550 -1115 9600 -1085
rect 9550 -1135 9565 -1115
rect 9585 -1135 9600 -1115
rect 9550 -1165 9600 -1135
rect 9550 -1185 9565 -1165
rect 9585 -1185 9600 -1165
rect 9550 -1215 9600 -1185
rect 9550 -1235 9565 -1215
rect 9585 -1235 9600 -1215
rect 9550 -1265 9600 -1235
rect 9550 -1285 9565 -1265
rect 9585 -1285 9600 -1265
rect 9550 -1315 9600 -1285
rect 9550 -1335 9565 -1315
rect 9585 -1335 9600 -1315
rect 9550 -1365 9600 -1335
rect 9550 -1385 9565 -1365
rect 9585 -1385 9600 -1365
rect 9550 -1415 9600 -1385
rect 9550 -1435 9565 -1415
rect 9585 -1435 9600 -1415
rect 9550 -1465 9600 -1435
rect 9550 -1485 9565 -1465
rect 9585 -1485 9600 -1465
rect 9550 -1515 9600 -1485
rect 9550 -1535 9565 -1515
rect 9585 -1535 9600 -1515
rect 9550 -1565 9600 -1535
rect 9550 -1585 9565 -1565
rect 9585 -1585 9600 -1565
rect 9550 -1615 9600 -1585
rect 9550 -1635 9565 -1615
rect 9585 -1635 9600 -1615
rect 9550 -1650 9600 -1635
rect 10750 -960 10800 -790
rect 11950 735 12000 915
rect 12250 1485 12300 1500
rect 12250 1465 12265 1485
rect 12285 1465 12300 1485
rect 12250 1435 12300 1465
rect 12250 1415 12265 1435
rect 12285 1415 12300 1435
rect 12250 1385 12300 1415
rect 12250 1365 12265 1385
rect 12285 1365 12300 1385
rect 12250 1335 12300 1365
rect 12250 1315 12265 1335
rect 12285 1315 12300 1335
rect 12250 1285 12300 1315
rect 12250 1265 12265 1285
rect 12285 1265 12300 1285
rect 12250 1235 12300 1265
rect 12250 1215 12265 1235
rect 12285 1215 12300 1235
rect 12250 1185 12300 1215
rect 12250 1165 12265 1185
rect 12285 1165 12300 1185
rect 12250 1135 12300 1165
rect 12250 1115 12265 1135
rect 12285 1115 12300 1135
rect 12250 1085 12300 1115
rect 12250 1065 12265 1085
rect 12285 1065 12300 1085
rect 12250 1035 12300 1065
rect 12250 1015 12265 1035
rect 12285 1015 12300 1035
rect 12250 985 12300 1015
rect 12550 1485 12600 1515
rect 13150 1535 13200 1550
rect 13150 1515 13165 1535
rect 13185 1515 13200 1535
rect 12550 1465 12565 1485
rect 12585 1465 12600 1485
rect 12550 1435 12600 1465
rect 12550 1415 12565 1435
rect 12585 1415 12600 1435
rect 12550 1385 12600 1415
rect 12550 1365 12565 1385
rect 12585 1365 12600 1385
rect 12550 1335 12600 1365
rect 12550 1315 12565 1335
rect 12585 1315 12600 1335
rect 12550 1285 12600 1315
rect 12550 1265 12565 1285
rect 12585 1265 12600 1285
rect 12550 1235 12600 1265
rect 12550 1215 12565 1235
rect 12585 1215 12600 1235
rect 12550 1185 12600 1215
rect 12550 1165 12565 1185
rect 12585 1165 12600 1185
rect 12550 1135 12600 1165
rect 12550 1115 12565 1135
rect 12585 1115 12600 1135
rect 12550 1085 12600 1115
rect 12550 1065 12565 1085
rect 12585 1065 12600 1085
rect 12550 1035 12600 1065
rect 12550 1015 12565 1035
rect 12585 1015 12600 1035
rect 12550 1000 12600 1015
rect 12850 1485 12900 1500
rect 12850 1465 12865 1485
rect 12885 1465 12900 1485
rect 12850 1435 12900 1465
rect 12850 1415 12865 1435
rect 12885 1415 12900 1435
rect 12850 1385 12900 1415
rect 12850 1365 12865 1385
rect 12885 1365 12900 1385
rect 12850 1335 12900 1365
rect 12850 1315 12865 1335
rect 12885 1315 12900 1335
rect 12850 1285 12900 1315
rect 12850 1265 12865 1285
rect 12885 1265 12900 1285
rect 12850 1235 12900 1265
rect 12850 1215 12865 1235
rect 12885 1215 12900 1235
rect 12850 1185 12900 1215
rect 12850 1165 12865 1185
rect 12885 1165 12900 1185
rect 12850 1135 12900 1165
rect 12850 1115 12865 1135
rect 12885 1115 12900 1135
rect 12850 1085 12900 1115
rect 12850 1065 12865 1085
rect 12885 1065 12900 1085
rect 12850 1035 12900 1065
rect 12850 1015 12865 1035
rect 12885 1015 12900 1035
rect 12250 965 12265 985
rect 12285 965 12300 985
rect 12250 950 12300 965
rect 12850 985 12900 1015
rect 12850 965 12865 985
rect 12885 965 12900 985
rect 12850 950 12900 965
rect 12250 935 12900 950
rect 12250 915 12265 935
rect 12285 915 12865 935
rect 12885 915 12900 935
rect 12250 900 12900 915
rect 13150 1485 13200 1515
rect 13750 1535 13800 1550
rect 13750 1515 13765 1535
rect 13785 1515 13800 1535
rect 13150 1465 13165 1485
rect 13185 1465 13200 1485
rect 13150 1435 13200 1465
rect 13150 1415 13165 1435
rect 13185 1415 13200 1435
rect 13150 1385 13200 1415
rect 13150 1365 13165 1385
rect 13185 1365 13200 1385
rect 13150 1335 13200 1365
rect 13150 1315 13165 1335
rect 13185 1315 13200 1335
rect 13150 1285 13200 1315
rect 13150 1265 13165 1285
rect 13185 1265 13200 1285
rect 13150 1235 13200 1265
rect 13150 1215 13165 1235
rect 13185 1215 13200 1235
rect 13150 1185 13200 1215
rect 13150 1165 13165 1185
rect 13185 1165 13200 1185
rect 13150 1135 13200 1165
rect 13150 1115 13165 1135
rect 13185 1115 13200 1135
rect 13150 1085 13200 1115
rect 13150 1065 13165 1085
rect 13185 1065 13200 1085
rect 13150 1035 13200 1065
rect 13150 1015 13165 1035
rect 13185 1015 13200 1035
rect 12100 840 12150 850
rect 12100 810 12110 840
rect 12140 810 12150 840
rect 12100 800 12150 810
rect 12400 840 12450 850
rect 12400 810 12410 840
rect 12440 810 12450 840
rect 12400 800 12450 810
rect 12550 840 12600 900
rect 12550 810 12560 840
rect 12590 810 12600 840
rect 12550 750 12600 810
rect 12700 840 12750 850
rect 12700 810 12710 840
rect 12740 810 12750 840
rect 12700 800 12750 810
rect 13000 840 13050 850
rect 13000 810 13010 840
rect 13040 810 13050 840
rect 13000 800 13050 810
rect 13150 840 13200 1015
rect 13450 1485 13500 1500
rect 13450 1465 13465 1485
rect 13485 1465 13500 1485
rect 13450 1435 13500 1465
rect 13450 1415 13465 1435
rect 13485 1415 13500 1435
rect 13450 1385 13500 1415
rect 13450 1365 13465 1385
rect 13485 1365 13500 1385
rect 13450 1335 13500 1365
rect 13450 1315 13465 1335
rect 13485 1315 13500 1335
rect 13450 1285 13500 1315
rect 13450 1265 13465 1285
rect 13485 1265 13500 1285
rect 13450 1235 13500 1265
rect 13450 1215 13465 1235
rect 13485 1215 13500 1235
rect 13450 1185 13500 1215
rect 13450 1165 13465 1185
rect 13485 1165 13500 1185
rect 13450 1135 13500 1165
rect 13450 1115 13465 1135
rect 13485 1115 13500 1135
rect 13450 1085 13500 1115
rect 13450 1065 13465 1085
rect 13485 1065 13500 1085
rect 13450 1035 13500 1065
rect 13450 1015 13465 1035
rect 13485 1015 13500 1035
rect 13450 985 13500 1015
rect 13750 1485 13800 1515
rect 14350 1535 14400 1550
rect 14350 1515 14365 1535
rect 14385 1515 14400 1535
rect 13750 1465 13765 1485
rect 13785 1465 13800 1485
rect 13750 1435 13800 1465
rect 13750 1415 13765 1435
rect 13785 1415 13800 1435
rect 13750 1385 13800 1415
rect 13750 1365 13765 1385
rect 13785 1365 13800 1385
rect 13750 1335 13800 1365
rect 13750 1315 13765 1335
rect 13785 1315 13800 1335
rect 13750 1285 13800 1315
rect 13750 1265 13765 1285
rect 13785 1265 13800 1285
rect 13750 1235 13800 1265
rect 13750 1215 13765 1235
rect 13785 1215 13800 1235
rect 13750 1185 13800 1215
rect 13750 1165 13765 1185
rect 13785 1165 13800 1185
rect 13750 1135 13800 1165
rect 13750 1115 13765 1135
rect 13785 1115 13800 1135
rect 13750 1085 13800 1115
rect 13750 1065 13765 1085
rect 13785 1065 13800 1085
rect 13750 1035 13800 1065
rect 13750 1015 13765 1035
rect 13785 1015 13800 1035
rect 13750 1000 13800 1015
rect 14050 1485 14100 1500
rect 14050 1465 14065 1485
rect 14085 1465 14100 1485
rect 14050 1435 14100 1465
rect 14050 1415 14065 1435
rect 14085 1415 14100 1435
rect 14050 1385 14100 1415
rect 14050 1365 14065 1385
rect 14085 1365 14100 1385
rect 14050 1335 14100 1365
rect 14050 1315 14065 1335
rect 14085 1315 14100 1335
rect 14050 1285 14100 1315
rect 14050 1265 14065 1285
rect 14085 1265 14100 1285
rect 14050 1235 14100 1265
rect 14050 1215 14065 1235
rect 14085 1215 14100 1235
rect 14050 1185 14100 1215
rect 14050 1165 14065 1185
rect 14085 1165 14100 1185
rect 14050 1135 14100 1165
rect 14050 1115 14065 1135
rect 14085 1115 14100 1135
rect 14050 1085 14100 1115
rect 14050 1065 14065 1085
rect 14085 1065 14100 1085
rect 14050 1035 14100 1065
rect 14050 1015 14065 1035
rect 14085 1015 14100 1035
rect 13450 965 13465 985
rect 13485 965 13500 985
rect 13450 950 13500 965
rect 14050 985 14100 1015
rect 14050 965 14065 985
rect 14085 965 14100 985
rect 14050 950 14100 965
rect 13450 935 14100 950
rect 13450 915 13465 935
rect 13485 915 14065 935
rect 14085 915 14100 935
rect 13450 900 14100 915
rect 14350 1485 14400 1515
rect 14350 1465 14365 1485
rect 14385 1465 14400 1485
rect 14350 1435 14400 1465
rect 14350 1415 14365 1435
rect 14385 1415 14400 1435
rect 14350 1385 14400 1415
rect 14350 1365 14365 1385
rect 14385 1365 14400 1385
rect 14350 1335 14400 1365
rect 14350 1315 14365 1335
rect 14385 1315 14400 1335
rect 14350 1285 14400 1315
rect 14350 1265 14365 1285
rect 14385 1265 14400 1285
rect 14350 1235 14400 1265
rect 14350 1215 14365 1235
rect 14385 1215 14400 1235
rect 14350 1185 14400 1215
rect 14350 1165 14365 1185
rect 14385 1165 14400 1185
rect 14350 1135 14400 1165
rect 14350 1115 14365 1135
rect 14385 1115 14400 1135
rect 14350 1085 14400 1115
rect 14350 1065 14365 1085
rect 14385 1065 14400 1085
rect 14350 1035 14400 1065
rect 14350 1015 14365 1035
rect 14385 1015 14400 1035
rect 14350 985 14400 1015
rect 14350 965 14365 985
rect 14385 965 14400 985
rect 14350 935 14400 965
rect 14350 915 14365 935
rect 14385 915 14400 935
rect 13150 810 13160 840
rect 13190 810 13200 840
rect 11950 715 11965 735
rect 11985 715 12000 735
rect 11950 685 12000 715
rect 11950 665 11965 685
rect 11985 665 12000 685
rect 11950 635 12000 665
rect 11950 615 11965 635
rect 11985 615 12000 635
rect 11950 585 12000 615
rect 11950 565 11965 585
rect 11985 565 12000 585
rect 11950 535 12000 565
rect 11950 515 11965 535
rect 11985 515 12000 535
rect 11950 485 12000 515
rect 11950 465 11965 485
rect 11985 465 12000 485
rect 11950 435 12000 465
rect 11950 415 11965 435
rect 11985 415 12000 435
rect 11950 385 12000 415
rect 11950 365 11965 385
rect 11985 365 12000 385
rect 11950 335 12000 365
rect 11950 315 11965 335
rect 11985 315 12000 335
rect 11950 285 12000 315
rect 11950 265 11965 285
rect 11985 265 12000 285
rect 11950 235 12000 265
rect 11950 215 11965 235
rect 11985 215 12000 235
rect 11950 185 12000 215
rect 11950 165 11965 185
rect 11985 165 12000 185
rect 11950 135 12000 165
rect 12250 735 12900 750
rect 12250 715 12265 735
rect 12285 715 12865 735
rect 12885 715 12900 735
rect 12250 700 12900 715
rect 12250 685 12300 700
rect 12250 665 12265 685
rect 12285 665 12300 685
rect 12250 635 12300 665
rect 12850 685 12900 700
rect 12850 665 12865 685
rect 12885 665 12900 685
rect 12250 615 12265 635
rect 12285 615 12300 635
rect 12250 585 12300 615
rect 12250 565 12265 585
rect 12285 565 12300 585
rect 12250 535 12300 565
rect 12250 515 12265 535
rect 12285 515 12300 535
rect 12250 485 12300 515
rect 12250 465 12265 485
rect 12285 465 12300 485
rect 12250 435 12300 465
rect 12250 415 12265 435
rect 12285 415 12300 435
rect 12250 385 12300 415
rect 12250 365 12265 385
rect 12285 365 12300 385
rect 12250 335 12300 365
rect 12250 315 12265 335
rect 12285 315 12300 335
rect 12250 285 12300 315
rect 12250 265 12265 285
rect 12285 265 12300 285
rect 12250 235 12300 265
rect 12250 215 12265 235
rect 12285 215 12300 235
rect 12250 185 12300 215
rect 12250 165 12265 185
rect 12285 165 12300 185
rect 12250 150 12300 165
rect 12550 635 12600 650
rect 12550 615 12565 635
rect 12585 615 12600 635
rect 12550 585 12600 615
rect 12550 565 12565 585
rect 12585 565 12600 585
rect 12550 535 12600 565
rect 12550 515 12565 535
rect 12585 515 12600 535
rect 12550 485 12600 515
rect 12550 465 12565 485
rect 12585 465 12600 485
rect 12550 435 12600 465
rect 12550 415 12565 435
rect 12585 415 12600 435
rect 12550 385 12600 415
rect 12550 365 12565 385
rect 12585 365 12600 385
rect 12550 335 12600 365
rect 12550 315 12565 335
rect 12585 315 12600 335
rect 12550 285 12600 315
rect 12550 265 12565 285
rect 12585 265 12600 285
rect 12550 235 12600 265
rect 12550 215 12565 235
rect 12585 215 12600 235
rect 12550 185 12600 215
rect 12550 165 12565 185
rect 12585 165 12600 185
rect 11950 115 11965 135
rect 11985 115 12000 135
rect 11950 100 12000 115
rect 12550 135 12600 165
rect 12850 635 12900 665
rect 12850 615 12865 635
rect 12885 615 12900 635
rect 12850 585 12900 615
rect 12850 565 12865 585
rect 12885 565 12900 585
rect 12850 535 12900 565
rect 12850 515 12865 535
rect 12885 515 12900 535
rect 12850 485 12900 515
rect 12850 465 12865 485
rect 12885 465 12900 485
rect 12850 435 12900 465
rect 12850 415 12865 435
rect 12885 415 12900 435
rect 12850 385 12900 415
rect 12850 365 12865 385
rect 12885 365 12900 385
rect 12850 335 12900 365
rect 12850 315 12865 335
rect 12885 315 12900 335
rect 12850 285 12900 315
rect 12850 265 12865 285
rect 12885 265 12900 285
rect 12850 235 12900 265
rect 12850 215 12865 235
rect 12885 215 12900 235
rect 12850 185 12900 215
rect 12850 165 12865 185
rect 12885 165 12900 185
rect 12850 150 12900 165
rect 13150 635 13200 810
rect 13300 840 13350 850
rect 13300 810 13310 840
rect 13340 810 13350 840
rect 13300 800 13350 810
rect 13600 840 13650 850
rect 13600 810 13610 840
rect 13640 810 13650 840
rect 13600 800 13650 810
rect 13750 840 13800 900
rect 13750 810 13760 840
rect 13790 810 13800 840
rect 13750 750 13800 810
rect 13900 840 13950 850
rect 13900 810 13910 840
rect 13940 810 13950 840
rect 13900 800 13950 810
rect 14200 840 14250 850
rect 14200 810 14210 840
rect 14240 810 14250 840
rect 14200 800 14250 810
rect 13150 615 13165 635
rect 13185 615 13200 635
rect 13150 585 13200 615
rect 13150 565 13165 585
rect 13185 565 13200 585
rect 13150 535 13200 565
rect 13150 515 13165 535
rect 13185 515 13200 535
rect 13150 485 13200 515
rect 13150 465 13165 485
rect 13185 465 13200 485
rect 13150 435 13200 465
rect 13150 415 13165 435
rect 13185 415 13200 435
rect 13150 385 13200 415
rect 13150 365 13165 385
rect 13185 365 13200 385
rect 13150 335 13200 365
rect 13150 315 13165 335
rect 13185 315 13200 335
rect 13150 285 13200 315
rect 13150 265 13165 285
rect 13185 265 13200 285
rect 13150 235 13200 265
rect 13150 215 13165 235
rect 13185 215 13200 235
rect 13150 185 13200 215
rect 13150 165 13165 185
rect 13185 165 13200 185
rect 12550 115 12565 135
rect 12585 115 12600 135
rect 12550 100 12600 115
rect 13150 135 13200 165
rect 13450 735 14100 750
rect 13450 715 13465 735
rect 13485 715 14065 735
rect 14085 715 14100 735
rect 13450 700 14100 715
rect 13450 685 13500 700
rect 13450 665 13465 685
rect 13485 665 13500 685
rect 13450 635 13500 665
rect 14050 685 14100 700
rect 14050 665 14065 685
rect 14085 665 14100 685
rect 13450 615 13465 635
rect 13485 615 13500 635
rect 13450 585 13500 615
rect 13450 565 13465 585
rect 13485 565 13500 585
rect 13450 535 13500 565
rect 13450 515 13465 535
rect 13485 515 13500 535
rect 13450 485 13500 515
rect 13450 465 13465 485
rect 13485 465 13500 485
rect 13450 435 13500 465
rect 13450 415 13465 435
rect 13485 415 13500 435
rect 13450 385 13500 415
rect 13450 365 13465 385
rect 13485 365 13500 385
rect 13450 335 13500 365
rect 13450 315 13465 335
rect 13485 315 13500 335
rect 13450 285 13500 315
rect 13450 265 13465 285
rect 13485 265 13500 285
rect 13450 235 13500 265
rect 13450 215 13465 235
rect 13485 215 13500 235
rect 13450 185 13500 215
rect 13450 165 13465 185
rect 13485 165 13500 185
rect 13450 150 13500 165
rect 13750 635 13800 650
rect 13750 615 13765 635
rect 13785 615 13800 635
rect 13750 585 13800 615
rect 13750 565 13765 585
rect 13785 565 13800 585
rect 13750 535 13800 565
rect 13750 515 13765 535
rect 13785 515 13800 535
rect 13750 485 13800 515
rect 13750 465 13765 485
rect 13785 465 13800 485
rect 13750 435 13800 465
rect 13750 415 13765 435
rect 13785 415 13800 435
rect 13750 385 13800 415
rect 13750 365 13765 385
rect 13785 365 13800 385
rect 13750 335 13800 365
rect 13750 315 13765 335
rect 13785 315 13800 335
rect 13750 285 13800 315
rect 13750 265 13765 285
rect 13785 265 13800 285
rect 13750 235 13800 265
rect 13750 215 13765 235
rect 13785 215 13800 235
rect 13750 185 13800 215
rect 13750 165 13765 185
rect 13785 165 13800 185
rect 13150 115 13165 135
rect 13185 115 13200 135
rect 13150 100 13200 115
rect 13750 135 13800 165
rect 14050 635 14100 665
rect 14050 615 14065 635
rect 14085 615 14100 635
rect 14050 585 14100 615
rect 14050 565 14065 585
rect 14085 565 14100 585
rect 14050 535 14100 565
rect 14050 515 14065 535
rect 14085 515 14100 535
rect 14050 485 14100 515
rect 14050 465 14065 485
rect 14085 465 14100 485
rect 14050 435 14100 465
rect 14050 415 14065 435
rect 14085 415 14100 435
rect 14050 385 14100 415
rect 14050 365 14065 385
rect 14085 365 14100 385
rect 14050 335 14100 365
rect 14050 315 14065 335
rect 14085 315 14100 335
rect 14050 285 14100 315
rect 14050 265 14065 285
rect 14085 265 14100 285
rect 14050 235 14100 265
rect 14050 215 14065 235
rect 14085 215 14100 235
rect 14050 185 14100 215
rect 14050 165 14065 185
rect 14085 165 14100 185
rect 14050 150 14100 165
rect 14350 735 14400 915
rect 15550 1585 15600 1660
rect 17950 1690 18000 1700
rect 17950 1660 17960 1690
rect 17990 1660 18000 1690
rect 15550 1565 15565 1585
rect 15585 1565 15600 1585
rect 15550 1540 15600 1565
rect 15550 1510 15560 1540
rect 15590 1510 15600 1540
rect 15550 1485 15600 1510
rect 15550 1465 15565 1485
rect 15585 1465 15600 1485
rect 15550 1440 15600 1465
rect 15550 1410 15560 1440
rect 15590 1410 15600 1440
rect 15550 1385 15600 1410
rect 15550 1365 15565 1385
rect 15585 1365 15600 1385
rect 15550 1340 15600 1365
rect 15550 1310 15560 1340
rect 15590 1310 15600 1340
rect 15550 1285 15600 1310
rect 15550 1265 15565 1285
rect 15585 1265 15600 1285
rect 15550 1240 15600 1265
rect 15550 1210 15560 1240
rect 15590 1210 15600 1240
rect 15550 1185 15600 1210
rect 15550 1165 15565 1185
rect 15585 1165 15600 1185
rect 15550 1140 15600 1165
rect 15550 1110 15560 1140
rect 15590 1110 15600 1140
rect 15550 1085 15600 1110
rect 15550 1065 15565 1085
rect 15585 1065 15600 1085
rect 15550 1040 15600 1065
rect 15550 1010 15560 1040
rect 15590 1010 15600 1040
rect 15550 985 15600 1010
rect 15550 965 15565 985
rect 15585 965 15600 985
rect 15550 940 15600 965
rect 15550 910 15560 940
rect 15590 910 15600 940
rect 14500 840 14550 850
rect 14500 810 14510 840
rect 14540 810 14550 840
rect 14500 800 14550 810
rect 14800 840 14850 850
rect 14800 810 14810 840
rect 14840 810 14850 840
rect 14800 800 14850 810
rect 15100 840 15150 850
rect 15100 810 15110 840
rect 15140 810 15150 840
rect 15100 800 15150 810
rect 15400 840 15450 850
rect 15400 810 15410 840
rect 15440 810 15450 840
rect 15400 800 15450 810
rect 14350 715 14365 735
rect 14385 715 14400 735
rect 14350 685 14400 715
rect 14350 665 14365 685
rect 14385 665 14400 685
rect 14350 635 14400 665
rect 14350 615 14365 635
rect 14385 615 14400 635
rect 14350 585 14400 615
rect 14350 565 14365 585
rect 14385 565 14400 585
rect 14350 535 14400 565
rect 14350 515 14365 535
rect 14385 515 14400 535
rect 14350 485 14400 515
rect 14350 465 14365 485
rect 14385 465 14400 485
rect 14350 435 14400 465
rect 14350 415 14365 435
rect 14385 415 14400 435
rect 14350 385 14400 415
rect 14350 365 14365 385
rect 14385 365 14400 385
rect 14350 335 14400 365
rect 14350 315 14365 335
rect 14385 315 14400 335
rect 14350 285 14400 315
rect 14350 265 14365 285
rect 14385 265 14400 285
rect 14350 235 14400 265
rect 14350 215 14365 235
rect 14385 215 14400 235
rect 14350 185 14400 215
rect 14350 165 14365 185
rect 14385 165 14400 185
rect 13750 115 13765 135
rect 13785 115 13800 135
rect 13750 100 13800 115
rect 14350 135 14400 165
rect 14350 115 14365 135
rect 14385 115 14400 135
rect 14350 100 14400 115
rect 11950 85 14400 100
rect 11950 65 11965 85
rect 11985 65 12565 85
rect 12585 65 13165 85
rect 13185 65 13765 85
rect 13785 65 14365 85
rect 14385 65 14400 85
rect 11950 50 14400 65
rect 11950 -100 12000 50
rect 13150 -100 13200 50
rect 14350 -100 14400 50
rect 11950 -115 14400 -100
rect 11950 -135 11965 -115
rect 11985 -135 12565 -115
rect 12585 -135 13165 -115
rect 13185 -135 13765 -115
rect 13785 -135 14365 -115
rect 14385 -135 14400 -115
rect 11950 -150 14400 -135
rect 11950 -165 12000 -150
rect 11950 -185 11965 -165
rect 11985 -185 12000 -165
rect 11950 -215 12000 -185
rect 12550 -165 12600 -150
rect 12550 -185 12565 -165
rect 12585 -185 12600 -165
rect 11950 -235 11965 -215
rect 11985 -235 12000 -215
rect 11950 -265 12000 -235
rect 11950 -285 11965 -265
rect 11985 -285 12000 -265
rect 11950 -315 12000 -285
rect 11950 -335 11965 -315
rect 11985 -335 12000 -315
rect 11950 -365 12000 -335
rect 11950 -385 11965 -365
rect 11985 -385 12000 -365
rect 11950 -415 12000 -385
rect 11950 -435 11965 -415
rect 11985 -435 12000 -415
rect 11950 -465 12000 -435
rect 11950 -485 11965 -465
rect 11985 -485 12000 -465
rect 11950 -515 12000 -485
rect 11950 -535 11965 -515
rect 11985 -535 12000 -515
rect 11950 -565 12000 -535
rect 11950 -585 11965 -565
rect 11985 -585 12000 -565
rect 11950 -615 12000 -585
rect 11950 -635 11965 -615
rect 11985 -635 12000 -615
rect 11950 -665 12000 -635
rect 11950 -685 11965 -665
rect 11985 -685 12000 -665
rect 11950 -715 12000 -685
rect 11950 -735 11965 -715
rect 11985 -735 12000 -715
rect 11950 -765 12000 -735
rect 11950 -785 11965 -765
rect 11985 -785 12000 -765
rect 10900 -860 10950 -850
rect 10900 -890 10910 -860
rect 10940 -890 10950 -860
rect 10900 -900 10950 -890
rect 11200 -860 11250 -850
rect 11200 -890 11210 -860
rect 11240 -890 11250 -860
rect 11200 -900 11250 -890
rect 11500 -860 11550 -850
rect 11500 -890 11510 -860
rect 11540 -890 11550 -860
rect 11500 -900 11550 -890
rect 11800 -860 11850 -850
rect 11800 -890 11810 -860
rect 11840 -890 11850 -860
rect 11800 -900 11850 -890
rect 10750 -990 10760 -960
rect 10790 -990 10800 -960
rect 10750 -1015 10800 -990
rect 10750 -1035 10765 -1015
rect 10785 -1035 10800 -1015
rect 10750 -1060 10800 -1035
rect 10750 -1090 10760 -1060
rect 10790 -1090 10800 -1060
rect 10750 -1115 10800 -1090
rect 10750 -1135 10765 -1115
rect 10785 -1135 10800 -1115
rect 10750 -1160 10800 -1135
rect 10750 -1190 10760 -1160
rect 10790 -1190 10800 -1160
rect 10750 -1215 10800 -1190
rect 10750 -1235 10765 -1215
rect 10785 -1235 10800 -1215
rect 10750 -1260 10800 -1235
rect 10750 -1290 10760 -1260
rect 10790 -1290 10800 -1260
rect 10750 -1315 10800 -1290
rect 10750 -1335 10765 -1315
rect 10785 -1335 10800 -1315
rect 10750 -1360 10800 -1335
rect 10750 -1390 10760 -1360
rect 10790 -1390 10800 -1360
rect 10750 -1415 10800 -1390
rect 10750 -1435 10765 -1415
rect 10785 -1435 10800 -1415
rect 10750 -1460 10800 -1435
rect 10750 -1490 10760 -1460
rect 10790 -1490 10800 -1460
rect 10750 -1515 10800 -1490
rect 10750 -1535 10765 -1515
rect 10785 -1535 10800 -1515
rect 10750 -1560 10800 -1535
rect 10750 -1590 10760 -1560
rect 10790 -1590 10800 -1560
rect 10750 -1615 10800 -1590
rect 10750 -1635 10765 -1615
rect 10785 -1635 10800 -1615
rect 8350 -1740 8360 -1710
rect 8390 -1740 8400 -1710
rect 8350 -1750 8400 -1740
rect 10750 -1710 10800 -1635
rect 11950 -965 12000 -785
rect 12250 -215 12300 -200
rect 12250 -235 12265 -215
rect 12285 -235 12300 -215
rect 12250 -265 12300 -235
rect 12250 -285 12265 -265
rect 12285 -285 12300 -265
rect 12250 -315 12300 -285
rect 12250 -335 12265 -315
rect 12285 -335 12300 -315
rect 12250 -365 12300 -335
rect 12250 -385 12265 -365
rect 12285 -385 12300 -365
rect 12250 -415 12300 -385
rect 12250 -435 12265 -415
rect 12285 -435 12300 -415
rect 12250 -465 12300 -435
rect 12250 -485 12265 -465
rect 12285 -485 12300 -465
rect 12250 -515 12300 -485
rect 12250 -535 12265 -515
rect 12285 -535 12300 -515
rect 12250 -565 12300 -535
rect 12250 -585 12265 -565
rect 12285 -585 12300 -565
rect 12250 -615 12300 -585
rect 12250 -635 12265 -615
rect 12285 -635 12300 -615
rect 12250 -665 12300 -635
rect 12250 -685 12265 -665
rect 12285 -685 12300 -665
rect 12250 -715 12300 -685
rect 12550 -215 12600 -185
rect 13150 -165 13200 -150
rect 13150 -185 13165 -165
rect 13185 -185 13200 -165
rect 12550 -235 12565 -215
rect 12585 -235 12600 -215
rect 12550 -265 12600 -235
rect 12550 -285 12565 -265
rect 12585 -285 12600 -265
rect 12550 -315 12600 -285
rect 12550 -335 12565 -315
rect 12585 -335 12600 -315
rect 12550 -365 12600 -335
rect 12550 -385 12565 -365
rect 12585 -385 12600 -365
rect 12550 -415 12600 -385
rect 12550 -435 12565 -415
rect 12585 -435 12600 -415
rect 12550 -465 12600 -435
rect 12550 -485 12565 -465
rect 12585 -485 12600 -465
rect 12550 -515 12600 -485
rect 12550 -535 12565 -515
rect 12585 -535 12600 -515
rect 12550 -565 12600 -535
rect 12550 -585 12565 -565
rect 12585 -585 12600 -565
rect 12550 -615 12600 -585
rect 12550 -635 12565 -615
rect 12585 -635 12600 -615
rect 12550 -665 12600 -635
rect 12550 -685 12565 -665
rect 12585 -685 12600 -665
rect 12550 -700 12600 -685
rect 12850 -215 12900 -200
rect 12850 -235 12865 -215
rect 12885 -235 12900 -215
rect 12850 -265 12900 -235
rect 12850 -285 12865 -265
rect 12885 -285 12900 -265
rect 12850 -315 12900 -285
rect 12850 -335 12865 -315
rect 12885 -335 12900 -315
rect 12850 -365 12900 -335
rect 12850 -385 12865 -365
rect 12885 -385 12900 -365
rect 12850 -415 12900 -385
rect 12850 -435 12865 -415
rect 12885 -435 12900 -415
rect 12850 -465 12900 -435
rect 12850 -485 12865 -465
rect 12885 -485 12900 -465
rect 12850 -515 12900 -485
rect 12850 -535 12865 -515
rect 12885 -535 12900 -515
rect 12850 -565 12900 -535
rect 12850 -585 12865 -565
rect 12885 -585 12900 -565
rect 12850 -615 12900 -585
rect 12850 -635 12865 -615
rect 12885 -635 12900 -615
rect 12850 -665 12900 -635
rect 12850 -685 12865 -665
rect 12885 -685 12900 -665
rect 12250 -735 12265 -715
rect 12285 -735 12300 -715
rect 12250 -750 12300 -735
rect 12850 -715 12900 -685
rect 12850 -735 12865 -715
rect 12885 -735 12900 -715
rect 12850 -750 12900 -735
rect 12250 -765 12900 -750
rect 12250 -785 12265 -765
rect 12285 -785 12865 -765
rect 12885 -785 12900 -765
rect 12250 -800 12900 -785
rect 13150 -215 13200 -185
rect 13750 -165 13800 -150
rect 13750 -185 13765 -165
rect 13785 -185 13800 -165
rect 13150 -235 13165 -215
rect 13185 -235 13200 -215
rect 13150 -265 13200 -235
rect 13150 -285 13165 -265
rect 13185 -285 13200 -265
rect 13150 -315 13200 -285
rect 13150 -335 13165 -315
rect 13185 -335 13200 -315
rect 13150 -365 13200 -335
rect 13150 -385 13165 -365
rect 13185 -385 13200 -365
rect 13150 -415 13200 -385
rect 13150 -435 13165 -415
rect 13185 -435 13200 -415
rect 13150 -465 13200 -435
rect 13150 -485 13165 -465
rect 13185 -485 13200 -465
rect 13150 -515 13200 -485
rect 13150 -535 13165 -515
rect 13185 -535 13200 -515
rect 13150 -565 13200 -535
rect 13150 -585 13165 -565
rect 13185 -585 13200 -565
rect 13150 -615 13200 -585
rect 13150 -635 13165 -615
rect 13185 -635 13200 -615
rect 13150 -665 13200 -635
rect 13150 -685 13165 -665
rect 13185 -685 13200 -665
rect 12100 -860 12150 -850
rect 12100 -890 12110 -860
rect 12140 -890 12150 -860
rect 12100 -900 12150 -890
rect 12400 -860 12450 -850
rect 12400 -890 12410 -860
rect 12440 -890 12450 -860
rect 12400 -900 12450 -890
rect 12550 -860 12600 -800
rect 12550 -890 12560 -860
rect 12590 -890 12600 -860
rect 12550 -950 12600 -890
rect 12700 -860 12750 -850
rect 12700 -890 12710 -860
rect 12740 -890 12750 -860
rect 12700 -900 12750 -890
rect 13000 -860 13050 -850
rect 13000 -890 13010 -860
rect 13040 -890 13050 -860
rect 13000 -900 13050 -890
rect 13150 -860 13200 -685
rect 13450 -215 13500 -200
rect 13450 -235 13465 -215
rect 13485 -235 13500 -215
rect 13450 -265 13500 -235
rect 13450 -285 13465 -265
rect 13485 -285 13500 -265
rect 13450 -315 13500 -285
rect 13450 -335 13465 -315
rect 13485 -335 13500 -315
rect 13450 -365 13500 -335
rect 13450 -385 13465 -365
rect 13485 -385 13500 -365
rect 13450 -415 13500 -385
rect 13450 -435 13465 -415
rect 13485 -435 13500 -415
rect 13450 -465 13500 -435
rect 13450 -485 13465 -465
rect 13485 -485 13500 -465
rect 13450 -515 13500 -485
rect 13450 -535 13465 -515
rect 13485 -535 13500 -515
rect 13450 -565 13500 -535
rect 13450 -585 13465 -565
rect 13485 -585 13500 -565
rect 13450 -615 13500 -585
rect 13450 -635 13465 -615
rect 13485 -635 13500 -615
rect 13450 -665 13500 -635
rect 13450 -685 13465 -665
rect 13485 -685 13500 -665
rect 13450 -715 13500 -685
rect 13750 -215 13800 -185
rect 14350 -165 14400 -150
rect 14350 -185 14365 -165
rect 14385 -185 14400 -165
rect 13750 -235 13765 -215
rect 13785 -235 13800 -215
rect 13750 -265 13800 -235
rect 13750 -285 13765 -265
rect 13785 -285 13800 -265
rect 13750 -315 13800 -285
rect 13750 -335 13765 -315
rect 13785 -335 13800 -315
rect 13750 -365 13800 -335
rect 13750 -385 13765 -365
rect 13785 -385 13800 -365
rect 13750 -415 13800 -385
rect 13750 -435 13765 -415
rect 13785 -435 13800 -415
rect 13750 -465 13800 -435
rect 13750 -485 13765 -465
rect 13785 -485 13800 -465
rect 13750 -515 13800 -485
rect 13750 -535 13765 -515
rect 13785 -535 13800 -515
rect 13750 -565 13800 -535
rect 13750 -585 13765 -565
rect 13785 -585 13800 -565
rect 13750 -615 13800 -585
rect 13750 -635 13765 -615
rect 13785 -635 13800 -615
rect 13750 -665 13800 -635
rect 13750 -685 13765 -665
rect 13785 -685 13800 -665
rect 13750 -700 13800 -685
rect 14050 -215 14100 -200
rect 14050 -235 14065 -215
rect 14085 -235 14100 -215
rect 14050 -265 14100 -235
rect 14050 -285 14065 -265
rect 14085 -285 14100 -265
rect 14050 -315 14100 -285
rect 14050 -335 14065 -315
rect 14085 -335 14100 -315
rect 14050 -365 14100 -335
rect 14050 -385 14065 -365
rect 14085 -385 14100 -365
rect 14050 -415 14100 -385
rect 14050 -435 14065 -415
rect 14085 -435 14100 -415
rect 14050 -465 14100 -435
rect 14050 -485 14065 -465
rect 14085 -485 14100 -465
rect 14050 -515 14100 -485
rect 14050 -535 14065 -515
rect 14085 -535 14100 -515
rect 14050 -565 14100 -535
rect 14050 -585 14065 -565
rect 14085 -585 14100 -565
rect 14050 -615 14100 -585
rect 14050 -635 14065 -615
rect 14085 -635 14100 -615
rect 14050 -665 14100 -635
rect 14050 -685 14065 -665
rect 14085 -685 14100 -665
rect 13450 -735 13465 -715
rect 13485 -735 13500 -715
rect 13450 -750 13500 -735
rect 14050 -715 14100 -685
rect 14050 -735 14065 -715
rect 14085 -735 14100 -715
rect 14050 -750 14100 -735
rect 13450 -765 14100 -750
rect 13450 -785 13465 -765
rect 13485 -785 14065 -765
rect 14085 -785 14100 -765
rect 13450 -800 14100 -785
rect 14350 -215 14400 -185
rect 14350 -235 14365 -215
rect 14385 -235 14400 -215
rect 14350 -265 14400 -235
rect 14350 -285 14365 -265
rect 14385 -285 14400 -265
rect 14350 -315 14400 -285
rect 14350 -335 14365 -315
rect 14385 -335 14400 -315
rect 14350 -365 14400 -335
rect 14350 -385 14365 -365
rect 14385 -385 14400 -365
rect 14350 -415 14400 -385
rect 14350 -435 14365 -415
rect 14385 -435 14400 -415
rect 14350 -465 14400 -435
rect 14350 -485 14365 -465
rect 14385 -485 14400 -465
rect 14350 -515 14400 -485
rect 14350 -535 14365 -515
rect 14385 -535 14400 -515
rect 14350 -565 14400 -535
rect 14350 -585 14365 -565
rect 14385 -585 14400 -565
rect 14350 -615 14400 -585
rect 14350 -635 14365 -615
rect 14385 -635 14400 -615
rect 14350 -665 14400 -635
rect 14350 -685 14365 -665
rect 14385 -685 14400 -665
rect 14350 -715 14400 -685
rect 14350 -735 14365 -715
rect 14385 -735 14400 -715
rect 14350 -765 14400 -735
rect 14350 -785 14365 -765
rect 14385 -785 14400 -765
rect 13150 -890 13160 -860
rect 13190 -890 13200 -860
rect 11950 -985 11965 -965
rect 11985 -985 12000 -965
rect 11950 -1015 12000 -985
rect 11950 -1035 11965 -1015
rect 11985 -1035 12000 -1015
rect 11950 -1065 12000 -1035
rect 11950 -1085 11965 -1065
rect 11985 -1085 12000 -1065
rect 11950 -1115 12000 -1085
rect 11950 -1135 11965 -1115
rect 11985 -1135 12000 -1115
rect 11950 -1165 12000 -1135
rect 11950 -1185 11965 -1165
rect 11985 -1185 12000 -1165
rect 11950 -1215 12000 -1185
rect 11950 -1235 11965 -1215
rect 11985 -1235 12000 -1215
rect 11950 -1265 12000 -1235
rect 11950 -1285 11965 -1265
rect 11985 -1285 12000 -1265
rect 11950 -1315 12000 -1285
rect 11950 -1335 11965 -1315
rect 11985 -1335 12000 -1315
rect 11950 -1365 12000 -1335
rect 11950 -1385 11965 -1365
rect 11985 -1385 12000 -1365
rect 11950 -1415 12000 -1385
rect 11950 -1435 11965 -1415
rect 11985 -1435 12000 -1415
rect 11950 -1465 12000 -1435
rect 11950 -1485 11965 -1465
rect 11985 -1485 12000 -1465
rect 11950 -1515 12000 -1485
rect 11950 -1535 11965 -1515
rect 11985 -1535 12000 -1515
rect 11950 -1565 12000 -1535
rect 12250 -965 12900 -950
rect 12250 -985 12265 -965
rect 12285 -985 12865 -965
rect 12885 -985 12900 -965
rect 12250 -1000 12900 -985
rect 12250 -1015 12300 -1000
rect 12250 -1035 12265 -1015
rect 12285 -1035 12300 -1015
rect 12250 -1065 12300 -1035
rect 12850 -1015 12900 -1000
rect 12850 -1035 12865 -1015
rect 12885 -1035 12900 -1015
rect 12250 -1085 12265 -1065
rect 12285 -1085 12300 -1065
rect 12250 -1115 12300 -1085
rect 12250 -1135 12265 -1115
rect 12285 -1135 12300 -1115
rect 12250 -1165 12300 -1135
rect 12250 -1185 12265 -1165
rect 12285 -1185 12300 -1165
rect 12250 -1215 12300 -1185
rect 12250 -1235 12265 -1215
rect 12285 -1235 12300 -1215
rect 12250 -1265 12300 -1235
rect 12250 -1285 12265 -1265
rect 12285 -1285 12300 -1265
rect 12250 -1315 12300 -1285
rect 12250 -1335 12265 -1315
rect 12285 -1335 12300 -1315
rect 12250 -1365 12300 -1335
rect 12250 -1385 12265 -1365
rect 12285 -1385 12300 -1365
rect 12250 -1415 12300 -1385
rect 12250 -1435 12265 -1415
rect 12285 -1435 12300 -1415
rect 12250 -1465 12300 -1435
rect 12250 -1485 12265 -1465
rect 12285 -1485 12300 -1465
rect 12250 -1515 12300 -1485
rect 12250 -1535 12265 -1515
rect 12285 -1535 12300 -1515
rect 12250 -1550 12300 -1535
rect 12550 -1065 12600 -1050
rect 12550 -1085 12565 -1065
rect 12585 -1085 12600 -1065
rect 12550 -1115 12600 -1085
rect 12550 -1135 12565 -1115
rect 12585 -1135 12600 -1115
rect 12550 -1165 12600 -1135
rect 12550 -1185 12565 -1165
rect 12585 -1185 12600 -1165
rect 12550 -1215 12600 -1185
rect 12550 -1235 12565 -1215
rect 12585 -1235 12600 -1215
rect 12550 -1265 12600 -1235
rect 12550 -1285 12565 -1265
rect 12585 -1285 12600 -1265
rect 12550 -1315 12600 -1285
rect 12550 -1335 12565 -1315
rect 12585 -1335 12600 -1315
rect 12550 -1365 12600 -1335
rect 12550 -1385 12565 -1365
rect 12585 -1385 12600 -1365
rect 12550 -1415 12600 -1385
rect 12550 -1435 12565 -1415
rect 12585 -1435 12600 -1415
rect 12550 -1465 12600 -1435
rect 12550 -1485 12565 -1465
rect 12585 -1485 12600 -1465
rect 12550 -1515 12600 -1485
rect 12550 -1535 12565 -1515
rect 12585 -1535 12600 -1515
rect 11950 -1585 11965 -1565
rect 11985 -1585 12000 -1565
rect 11950 -1600 12000 -1585
rect 12550 -1565 12600 -1535
rect 12850 -1065 12900 -1035
rect 12850 -1085 12865 -1065
rect 12885 -1085 12900 -1065
rect 12850 -1115 12900 -1085
rect 12850 -1135 12865 -1115
rect 12885 -1135 12900 -1115
rect 12850 -1165 12900 -1135
rect 12850 -1185 12865 -1165
rect 12885 -1185 12900 -1165
rect 12850 -1215 12900 -1185
rect 12850 -1235 12865 -1215
rect 12885 -1235 12900 -1215
rect 12850 -1265 12900 -1235
rect 12850 -1285 12865 -1265
rect 12885 -1285 12900 -1265
rect 12850 -1315 12900 -1285
rect 12850 -1335 12865 -1315
rect 12885 -1335 12900 -1315
rect 12850 -1365 12900 -1335
rect 12850 -1385 12865 -1365
rect 12885 -1385 12900 -1365
rect 12850 -1415 12900 -1385
rect 12850 -1435 12865 -1415
rect 12885 -1435 12900 -1415
rect 12850 -1465 12900 -1435
rect 12850 -1485 12865 -1465
rect 12885 -1485 12900 -1465
rect 12850 -1515 12900 -1485
rect 12850 -1535 12865 -1515
rect 12885 -1535 12900 -1515
rect 12850 -1550 12900 -1535
rect 13150 -1065 13200 -890
rect 13300 -860 13350 -850
rect 13300 -890 13310 -860
rect 13340 -890 13350 -860
rect 13300 -900 13350 -890
rect 13600 -860 13650 -850
rect 13600 -890 13610 -860
rect 13640 -890 13650 -860
rect 13600 -900 13650 -890
rect 13750 -860 13800 -800
rect 13750 -890 13760 -860
rect 13790 -890 13800 -860
rect 13750 -950 13800 -890
rect 13900 -860 13950 -850
rect 13900 -890 13910 -860
rect 13940 -890 13950 -860
rect 13900 -900 13950 -890
rect 14200 -860 14250 -850
rect 14200 -890 14210 -860
rect 14240 -890 14250 -860
rect 14200 -900 14250 -890
rect 13150 -1085 13165 -1065
rect 13185 -1085 13200 -1065
rect 13150 -1115 13200 -1085
rect 13150 -1135 13165 -1115
rect 13185 -1135 13200 -1115
rect 13150 -1165 13200 -1135
rect 13150 -1185 13165 -1165
rect 13185 -1185 13200 -1165
rect 13150 -1215 13200 -1185
rect 13150 -1235 13165 -1215
rect 13185 -1235 13200 -1215
rect 13150 -1265 13200 -1235
rect 13150 -1285 13165 -1265
rect 13185 -1285 13200 -1265
rect 13150 -1315 13200 -1285
rect 13150 -1335 13165 -1315
rect 13185 -1335 13200 -1315
rect 13150 -1365 13200 -1335
rect 13150 -1385 13165 -1365
rect 13185 -1385 13200 -1365
rect 13150 -1415 13200 -1385
rect 13150 -1435 13165 -1415
rect 13185 -1435 13200 -1415
rect 13150 -1465 13200 -1435
rect 13150 -1485 13165 -1465
rect 13185 -1485 13200 -1465
rect 13150 -1515 13200 -1485
rect 13150 -1535 13165 -1515
rect 13185 -1535 13200 -1515
rect 12550 -1585 12565 -1565
rect 12585 -1585 12600 -1565
rect 12550 -1600 12600 -1585
rect 13150 -1565 13200 -1535
rect 13450 -965 14100 -950
rect 13450 -985 13465 -965
rect 13485 -985 14065 -965
rect 14085 -985 14100 -965
rect 13450 -1000 14100 -985
rect 13450 -1015 13500 -1000
rect 13450 -1035 13465 -1015
rect 13485 -1035 13500 -1015
rect 13450 -1065 13500 -1035
rect 14050 -1015 14100 -1000
rect 14050 -1035 14065 -1015
rect 14085 -1035 14100 -1015
rect 13450 -1085 13465 -1065
rect 13485 -1085 13500 -1065
rect 13450 -1115 13500 -1085
rect 13450 -1135 13465 -1115
rect 13485 -1135 13500 -1115
rect 13450 -1165 13500 -1135
rect 13450 -1185 13465 -1165
rect 13485 -1185 13500 -1165
rect 13450 -1215 13500 -1185
rect 13450 -1235 13465 -1215
rect 13485 -1235 13500 -1215
rect 13450 -1265 13500 -1235
rect 13450 -1285 13465 -1265
rect 13485 -1285 13500 -1265
rect 13450 -1315 13500 -1285
rect 13450 -1335 13465 -1315
rect 13485 -1335 13500 -1315
rect 13450 -1365 13500 -1335
rect 13450 -1385 13465 -1365
rect 13485 -1385 13500 -1365
rect 13450 -1415 13500 -1385
rect 13450 -1435 13465 -1415
rect 13485 -1435 13500 -1415
rect 13450 -1465 13500 -1435
rect 13450 -1485 13465 -1465
rect 13485 -1485 13500 -1465
rect 13450 -1515 13500 -1485
rect 13450 -1535 13465 -1515
rect 13485 -1535 13500 -1515
rect 13450 -1550 13500 -1535
rect 13750 -1065 13800 -1050
rect 13750 -1085 13765 -1065
rect 13785 -1085 13800 -1065
rect 13750 -1115 13800 -1085
rect 13750 -1135 13765 -1115
rect 13785 -1135 13800 -1115
rect 13750 -1165 13800 -1135
rect 13750 -1185 13765 -1165
rect 13785 -1185 13800 -1165
rect 13750 -1215 13800 -1185
rect 13750 -1235 13765 -1215
rect 13785 -1235 13800 -1215
rect 13750 -1265 13800 -1235
rect 13750 -1285 13765 -1265
rect 13785 -1285 13800 -1265
rect 13750 -1315 13800 -1285
rect 13750 -1335 13765 -1315
rect 13785 -1335 13800 -1315
rect 13750 -1365 13800 -1335
rect 13750 -1385 13765 -1365
rect 13785 -1385 13800 -1365
rect 13750 -1415 13800 -1385
rect 13750 -1435 13765 -1415
rect 13785 -1435 13800 -1415
rect 13750 -1465 13800 -1435
rect 13750 -1485 13765 -1465
rect 13785 -1485 13800 -1465
rect 13750 -1515 13800 -1485
rect 13750 -1535 13765 -1515
rect 13785 -1535 13800 -1515
rect 13150 -1585 13165 -1565
rect 13185 -1585 13200 -1565
rect 13150 -1600 13200 -1585
rect 13750 -1565 13800 -1535
rect 14050 -1065 14100 -1035
rect 14050 -1085 14065 -1065
rect 14085 -1085 14100 -1065
rect 14050 -1115 14100 -1085
rect 14050 -1135 14065 -1115
rect 14085 -1135 14100 -1115
rect 14050 -1165 14100 -1135
rect 14050 -1185 14065 -1165
rect 14085 -1185 14100 -1165
rect 14050 -1215 14100 -1185
rect 14050 -1235 14065 -1215
rect 14085 -1235 14100 -1215
rect 14050 -1265 14100 -1235
rect 14050 -1285 14065 -1265
rect 14085 -1285 14100 -1265
rect 14050 -1315 14100 -1285
rect 14050 -1335 14065 -1315
rect 14085 -1335 14100 -1315
rect 14050 -1365 14100 -1335
rect 14050 -1385 14065 -1365
rect 14085 -1385 14100 -1365
rect 14050 -1415 14100 -1385
rect 14050 -1435 14065 -1415
rect 14085 -1435 14100 -1415
rect 14050 -1465 14100 -1435
rect 14050 -1485 14065 -1465
rect 14085 -1485 14100 -1465
rect 14050 -1515 14100 -1485
rect 14050 -1535 14065 -1515
rect 14085 -1535 14100 -1515
rect 14050 -1550 14100 -1535
rect 14350 -965 14400 -785
rect 15550 740 15600 910
rect 16750 1585 16800 1600
rect 16750 1565 16765 1585
rect 16785 1565 16800 1585
rect 16750 1535 16800 1565
rect 16750 1515 16765 1535
rect 16785 1515 16800 1535
rect 16750 1485 16800 1515
rect 16750 1465 16765 1485
rect 16785 1465 16800 1485
rect 16750 1435 16800 1465
rect 16750 1415 16765 1435
rect 16785 1415 16800 1435
rect 16750 1385 16800 1415
rect 16750 1365 16765 1385
rect 16785 1365 16800 1385
rect 16750 1335 16800 1365
rect 16750 1315 16765 1335
rect 16785 1315 16800 1335
rect 16750 1285 16800 1315
rect 16750 1265 16765 1285
rect 16785 1265 16800 1285
rect 16750 1235 16800 1265
rect 16750 1215 16765 1235
rect 16785 1215 16800 1235
rect 16750 1185 16800 1215
rect 16750 1165 16765 1185
rect 16785 1165 16800 1185
rect 16750 1135 16800 1165
rect 16750 1115 16765 1135
rect 16785 1115 16800 1135
rect 16750 1085 16800 1115
rect 16750 1065 16765 1085
rect 16785 1065 16800 1085
rect 16750 1035 16800 1065
rect 16750 1015 16765 1035
rect 16785 1015 16800 1035
rect 16750 985 16800 1015
rect 16750 965 16765 985
rect 16785 965 16800 985
rect 16750 935 16800 965
rect 16750 915 16765 935
rect 16785 915 16800 935
rect 15700 840 15750 850
rect 15700 810 15710 840
rect 15740 810 15750 840
rect 15700 800 15750 810
rect 16000 840 16050 850
rect 16000 810 16010 840
rect 16040 810 16050 840
rect 16000 800 16050 810
rect 16300 840 16350 850
rect 16300 810 16310 840
rect 16340 810 16350 840
rect 16300 800 16350 810
rect 16600 840 16650 850
rect 16600 810 16610 840
rect 16640 810 16650 840
rect 16600 800 16650 810
rect 16750 840 16800 915
rect 17950 1585 18000 1660
rect 20350 1690 20400 1700
rect 20350 1660 20360 1690
rect 20390 1660 20400 1690
rect 17950 1565 17965 1585
rect 17985 1565 18000 1585
rect 17950 1540 18000 1565
rect 17950 1510 17960 1540
rect 17990 1510 18000 1540
rect 17950 1485 18000 1510
rect 17950 1465 17965 1485
rect 17985 1465 18000 1485
rect 17950 1440 18000 1465
rect 17950 1410 17960 1440
rect 17990 1410 18000 1440
rect 17950 1385 18000 1410
rect 17950 1365 17965 1385
rect 17985 1365 18000 1385
rect 17950 1340 18000 1365
rect 17950 1310 17960 1340
rect 17990 1310 18000 1340
rect 17950 1285 18000 1310
rect 17950 1265 17965 1285
rect 17985 1265 18000 1285
rect 17950 1240 18000 1265
rect 17950 1210 17960 1240
rect 17990 1210 18000 1240
rect 17950 1185 18000 1210
rect 17950 1165 17965 1185
rect 17985 1165 18000 1185
rect 17950 1140 18000 1165
rect 17950 1110 17960 1140
rect 17990 1110 18000 1140
rect 17950 1085 18000 1110
rect 17950 1065 17965 1085
rect 17985 1065 18000 1085
rect 17950 1040 18000 1065
rect 17950 1010 17960 1040
rect 17990 1010 18000 1040
rect 17950 985 18000 1010
rect 17950 965 17965 985
rect 17985 965 18000 985
rect 17950 940 18000 965
rect 17950 910 17960 940
rect 17990 910 18000 940
rect 16750 810 16760 840
rect 16790 810 16800 840
rect 15550 710 15560 740
rect 15590 710 15600 740
rect 15550 685 15600 710
rect 15550 665 15565 685
rect 15585 665 15600 685
rect 15550 640 15600 665
rect 15550 610 15560 640
rect 15590 610 15600 640
rect 15550 585 15600 610
rect 15550 565 15565 585
rect 15585 565 15600 585
rect 15550 540 15600 565
rect 15550 510 15560 540
rect 15590 510 15600 540
rect 15550 485 15600 510
rect 15550 465 15565 485
rect 15585 465 15600 485
rect 15550 440 15600 465
rect 15550 410 15560 440
rect 15590 410 15600 440
rect 15550 385 15600 410
rect 15550 365 15565 385
rect 15585 365 15600 385
rect 15550 340 15600 365
rect 15550 310 15560 340
rect 15590 310 15600 340
rect 15550 285 15600 310
rect 15550 265 15565 285
rect 15585 265 15600 285
rect 15550 240 15600 265
rect 15550 210 15560 240
rect 15590 210 15600 240
rect 15550 185 15600 210
rect 15550 165 15565 185
rect 15585 165 15600 185
rect 15550 140 15600 165
rect 15550 110 15560 140
rect 15590 110 15600 140
rect 15550 85 15600 110
rect 15550 65 15565 85
rect 15585 65 15600 85
rect 15550 -10 15600 65
rect 16750 735 16800 810
rect 16900 840 16950 850
rect 16900 810 16910 840
rect 16940 810 16950 840
rect 16900 800 16950 810
rect 17200 840 17250 850
rect 17200 810 17210 840
rect 17240 810 17250 840
rect 17200 800 17250 810
rect 17500 840 17550 850
rect 17500 810 17510 840
rect 17540 810 17550 840
rect 17500 800 17550 810
rect 17800 840 17850 850
rect 17800 810 17810 840
rect 17840 810 17850 840
rect 17800 800 17850 810
rect 16750 715 16765 735
rect 16785 715 16800 735
rect 16750 685 16800 715
rect 16750 665 16765 685
rect 16785 665 16800 685
rect 16750 635 16800 665
rect 16750 615 16765 635
rect 16785 615 16800 635
rect 16750 585 16800 615
rect 16750 565 16765 585
rect 16785 565 16800 585
rect 16750 535 16800 565
rect 16750 515 16765 535
rect 16785 515 16800 535
rect 16750 485 16800 515
rect 16750 465 16765 485
rect 16785 465 16800 485
rect 16750 435 16800 465
rect 16750 415 16765 435
rect 16785 415 16800 435
rect 16750 385 16800 415
rect 16750 365 16765 385
rect 16785 365 16800 385
rect 16750 335 16800 365
rect 16750 315 16765 335
rect 16785 315 16800 335
rect 16750 285 16800 315
rect 16750 265 16765 285
rect 16785 265 16800 285
rect 16750 235 16800 265
rect 16750 215 16765 235
rect 16785 215 16800 235
rect 16750 185 16800 215
rect 16750 165 16765 185
rect 16785 165 16800 185
rect 16750 135 16800 165
rect 16750 115 16765 135
rect 16785 115 16800 135
rect 16750 85 16800 115
rect 16750 65 16765 85
rect 16785 65 16800 85
rect 16750 50 16800 65
rect 17950 740 18000 910
rect 19150 1585 19200 1600
rect 19150 1565 19165 1585
rect 19185 1565 19200 1585
rect 19150 1535 19200 1565
rect 19150 1515 19165 1535
rect 19185 1515 19200 1535
rect 19150 1485 19200 1515
rect 19150 1465 19165 1485
rect 19185 1465 19200 1485
rect 19150 1435 19200 1465
rect 19150 1415 19165 1435
rect 19185 1415 19200 1435
rect 19150 1385 19200 1415
rect 19150 1365 19165 1385
rect 19185 1365 19200 1385
rect 19150 1335 19200 1365
rect 19150 1315 19165 1335
rect 19185 1315 19200 1335
rect 19150 1285 19200 1315
rect 19150 1265 19165 1285
rect 19185 1265 19200 1285
rect 19150 1235 19200 1265
rect 19150 1215 19165 1235
rect 19185 1215 19200 1235
rect 19150 1185 19200 1215
rect 19150 1165 19165 1185
rect 19185 1165 19200 1185
rect 19150 1135 19200 1165
rect 19150 1115 19165 1135
rect 19185 1115 19200 1135
rect 19150 1085 19200 1115
rect 19150 1065 19165 1085
rect 19185 1065 19200 1085
rect 19150 1035 19200 1065
rect 19150 1015 19165 1035
rect 19185 1015 19200 1035
rect 19150 985 19200 1015
rect 19150 965 19165 985
rect 19185 965 19200 985
rect 19150 935 19200 965
rect 19150 915 19165 935
rect 19185 915 19200 935
rect 18100 840 18150 850
rect 18100 810 18110 840
rect 18140 810 18150 840
rect 18100 800 18150 810
rect 18400 840 18450 850
rect 18400 810 18410 840
rect 18440 810 18450 840
rect 18400 800 18450 810
rect 18700 840 18750 850
rect 18700 810 18710 840
rect 18740 810 18750 840
rect 18700 800 18750 810
rect 19000 840 19050 850
rect 19000 810 19010 840
rect 19040 810 19050 840
rect 19000 800 19050 810
rect 19150 840 19200 915
rect 20350 1585 20400 1660
rect 20350 1565 20365 1585
rect 20385 1565 20400 1585
rect 20350 1540 20400 1565
rect 20350 1510 20360 1540
rect 20390 1510 20400 1540
rect 20350 1485 20400 1510
rect 20350 1465 20365 1485
rect 20385 1465 20400 1485
rect 20350 1440 20400 1465
rect 20350 1410 20360 1440
rect 20390 1410 20400 1440
rect 20350 1385 20400 1410
rect 20350 1365 20365 1385
rect 20385 1365 20400 1385
rect 20350 1340 20400 1365
rect 20350 1310 20360 1340
rect 20390 1310 20400 1340
rect 20350 1285 20400 1310
rect 20350 1265 20365 1285
rect 20385 1265 20400 1285
rect 20350 1240 20400 1265
rect 20350 1210 20360 1240
rect 20390 1210 20400 1240
rect 20350 1185 20400 1210
rect 20350 1165 20365 1185
rect 20385 1165 20400 1185
rect 20350 1140 20400 1165
rect 20350 1110 20360 1140
rect 20390 1110 20400 1140
rect 20350 1085 20400 1110
rect 20350 1065 20365 1085
rect 20385 1065 20400 1085
rect 20350 1040 20400 1065
rect 20350 1010 20360 1040
rect 20390 1010 20400 1040
rect 20350 985 20400 1010
rect 20350 965 20365 985
rect 20385 965 20400 985
rect 20350 940 20400 965
rect 20350 910 20360 940
rect 20390 910 20400 940
rect 19150 810 19160 840
rect 19190 810 19200 840
rect 17950 710 17960 740
rect 17990 710 18000 740
rect 17950 685 18000 710
rect 17950 665 17965 685
rect 17985 665 18000 685
rect 17950 640 18000 665
rect 17950 610 17960 640
rect 17990 610 18000 640
rect 17950 585 18000 610
rect 17950 565 17965 585
rect 17985 565 18000 585
rect 17950 540 18000 565
rect 17950 510 17960 540
rect 17990 510 18000 540
rect 17950 485 18000 510
rect 17950 465 17965 485
rect 17985 465 18000 485
rect 17950 440 18000 465
rect 17950 410 17960 440
rect 17990 410 18000 440
rect 17950 385 18000 410
rect 17950 365 17965 385
rect 17985 365 18000 385
rect 17950 340 18000 365
rect 17950 310 17960 340
rect 17990 310 18000 340
rect 17950 285 18000 310
rect 17950 265 17965 285
rect 17985 265 18000 285
rect 17950 240 18000 265
rect 17950 210 17960 240
rect 17990 210 18000 240
rect 17950 185 18000 210
rect 17950 165 17965 185
rect 17985 165 18000 185
rect 17950 140 18000 165
rect 17950 110 17960 140
rect 17990 110 18000 140
rect 17950 85 18000 110
rect 17950 65 17965 85
rect 17985 65 18000 85
rect 15550 -40 15560 -10
rect 15590 -40 15600 -10
rect 15550 -115 15600 -40
rect 17950 -10 18000 65
rect 19150 735 19200 810
rect 19300 840 19350 850
rect 19300 810 19310 840
rect 19340 810 19350 840
rect 19300 800 19350 810
rect 19600 840 19650 850
rect 19600 810 19610 840
rect 19640 810 19650 840
rect 19600 800 19650 810
rect 19900 840 19950 850
rect 19900 810 19910 840
rect 19940 810 19950 840
rect 19900 800 19950 810
rect 20200 840 20250 850
rect 20200 810 20210 840
rect 20240 810 20250 840
rect 20200 800 20250 810
rect 19150 715 19165 735
rect 19185 715 19200 735
rect 19150 685 19200 715
rect 19150 665 19165 685
rect 19185 665 19200 685
rect 19150 635 19200 665
rect 19150 615 19165 635
rect 19185 615 19200 635
rect 19150 585 19200 615
rect 19150 565 19165 585
rect 19185 565 19200 585
rect 19150 535 19200 565
rect 19150 515 19165 535
rect 19185 515 19200 535
rect 19150 485 19200 515
rect 19150 465 19165 485
rect 19185 465 19200 485
rect 19150 435 19200 465
rect 19150 415 19165 435
rect 19185 415 19200 435
rect 19150 385 19200 415
rect 19150 365 19165 385
rect 19185 365 19200 385
rect 19150 335 19200 365
rect 19150 315 19165 335
rect 19185 315 19200 335
rect 19150 285 19200 315
rect 19150 265 19165 285
rect 19185 265 19200 285
rect 19150 235 19200 265
rect 19150 215 19165 235
rect 19185 215 19200 235
rect 19150 185 19200 215
rect 19150 165 19165 185
rect 19185 165 19200 185
rect 19150 135 19200 165
rect 19150 115 19165 135
rect 19185 115 19200 135
rect 19150 85 19200 115
rect 19150 65 19165 85
rect 19185 65 19200 85
rect 19150 50 19200 65
rect 20350 740 20400 910
rect 20350 710 20360 740
rect 20390 710 20400 740
rect 20350 685 20400 710
rect 20350 665 20365 685
rect 20385 665 20400 685
rect 20350 640 20400 665
rect 20350 610 20360 640
rect 20390 610 20400 640
rect 20350 585 20400 610
rect 20350 565 20365 585
rect 20385 565 20400 585
rect 20350 540 20400 565
rect 20350 510 20360 540
rect 20390 510 20400 540
rect 20350 485 20400 510
rect 20350 465 20365 485
rect 20385 465 20400 485
rect 20350 440 20400 465
rect 20350 410 20360 440
rect 20390 410 20400 440
rect 20350 385 20400 410
rect 20350 365 20365 385
rect 20385 365 20400 385
rect 20350 340 20400 365
rect 20350 310 20360 340
rect 20390 310 20400 340
rect 20350 285 20400 310
rect 20350 265 20365 285
rect 20385 265 20400 285
rect 20350 240 20400 265
rect 20350 210 20360 240
rect 20390 210 20400 240
rect 20350 185 20400 210
rect 20350 165 20365 185
rect 20385 165 20400 185
rect 20350 140 20400 165
rect 20350 110 20360 140
rect 20390 110 20400 140
rect 20350 85 20400 110
rect 20350 65 20365 85
rect 20385 65 20400 85
rect 17950 -40 17960 -10
rect 17990 -40 18000 -10
rect 15550 -135 15565 -115
rect 15585 -135 15600 -115
rect 15550 -160 15600 -135
rect 15550 -190 15560 -160
rect 15590 -190 15600 -160
rect 15550 -215 15600 -190
rect 15550 -235 15565 -215
rect 15585 -235 15600 -215
rect 15550 -260 15600 -235
rect 15550 -290 15560 -260
rect 15590 -290 15600 -260
rect 15550 -315 15600 -290
rect 15550 -335 15565 -315
rect 15585 -335 15600 -315
rect 15550 -360 15600 -335
rect 15550 -390 15560 -360
rect 15590 -390 15600 -360
rect 15550 -415 15600 -390
rect 15550 -435 15565 -415
rect 15585 -435 15600 -415
rect 15550 -460 15600 -435
rect 15550 -490 15560 -460
rect 15590 -490 15600 -460
rect 15550 -515 15600 -490
rect 15550 -535 15565 -515
rect 15585 -535 15600 -515
rect 15550 -560 15600 -535
rect 15550 -590 15560 -560
rect 15590 -590 15600 -560
rect 15550 -615 15600 -590
rect 15550 -635 15565 -615
rect 15585 -635 15600 -615
rect 15550 -660 15600 -635
rect 15550 -690 15560 -660
rect 15590 -690 15600 -660
rect 15550 -715 15600 -690
rect 15550 -735 15565 -715
rect 15585 -735 15600 -715
rect 15550 -760 15600 -735
rect 15550 -790 15560 -760
rect 15590 -790 15600 -760
rect 14500 -860 14550 -850
rect 14500 -890 14510 -860
rect 14540 -890 14550 -860
rect 14500 -900 14550 -890
rect 14800 -860 14850 -850
rect 14800 -890 14810 -860
rect 14840 -890 14850 -860
rect 14800 -900 14850 -890
rect 15100 -860 15150 -850
rect 15100 -890 15110 -860
rect 15140 -890 15150 -860
rect 15100 -900 15150 -890
rect 15400 -860 15450 -850
rect 15400 -890 15410 -860
rect 15440 -890 15450 -860
rect 15400 -900 15450 -890
rect 14350 -985 14365 -965
rect 14385 -985 14400 -965
rect 14350 -1015 14400 -985
rect 14350 -1035 14365 -1015
rect 14385 -1035 14400 -1015
rect 14350 -1065 14400 -1035
rect 14350 -1085 14365 -1065
rect 14385 -1085 14400 -1065
rect 14350 -1115 14400 -1085
rect 14350 -1135 14365 -1115
rect 14385 -1135 14400 -1115
rect 14350 -1165 14400 -1135
rect 14350 -1185 14365 -1165
rect 14385 -1185 14400 -1165
rect 14350 -1215 14400 -1185
rect 14350 -1235 14365 -1215
rect 14385 -1235 14400 -1215
rect 14350 -1265 14400 -1235
rect 14350 -1285 14365 -1265
rect 14385 -1285 14400 -1265
rect 14350 -1315 14400 -1285
rect 14350 -1335 14365 -1315
rect 14385 -1335 14400 -1315
rect 14350 -1365 14400 -1335
rect 14350 -1385 14365 -1365
rect 14385 -1385 14400 -1365
rect 14350 -1415 14400 -1385
rect 14350 -1435 14365 -1415
rect 14385 -1435 14400 -1415
rect 14350 -1465 14400 -1435
rect 14350 -1485 14365 -1465
rect 14385 -1485 14400 -1465
rect 14350 -1515 14400 -1485
rect 14350 -1535 14365 -1515
rect 14385 -1535 14400 -1515
rect 13750 -1585 13765 -1565
rect 13785 -1585 13800 -1565
rect 13750 -1600 13800 -1585
rect 14350 -1565 14400 -1535
rect 14350 -1585 14365 -1565
rect 14385 -1585 14400 -1565
rect 14350 -1600 14400 -1585
rect 11950 -1615 14400 -1600
rect 11950 -1635 11965 -1615
rect 11985 -1635 12565 -1615
rect 12585 -1635 13165 -1615
rect 13185 -1635 13765 -1615
rect 13785 -1635 14365 -1615
rect 14385 -1635 14400 -1615
rect 11950 -1650 14400 -1635
rect 15550 -960 15600 -790
rect 16750 -115 16800 -100
rect 16750 -135 16765 -115
rect 16785 -135 16800 -115
rect 16750 -165 16800 -135
rect 16750 -185 16765 -165
rect 16785 -185 16800 -165
rect 16750 -215 16800 -185
rect 16750 -235 16765 -215
rect 16785 -235 16800 -215
rect 16750 -265 16800 -235
rect 16750 -285 16765 -265
rect 16785 -285 16800 -265
rect 16750 -315 16800 -285
rect 16750 -335 16765 -315
rect 16785 -335 16800 -315
rect 16750 -365 16800 -335
rect 16750 -385 16765 -365
rect 16785 -385 16800 -365
rect 16750 -415 16800 -385
rect 16750 -435 16765 -415
rect 16785 -435 16800 -415
rect 16750 -465 16800 -435
rect 16750 -485 16765 -465
rect 16785 -485 16800 -465
rect 16750 -515 16800 -485
rect 16750 -535 16765 -515
rect 16785 -535 16800 -515
rect 16750 -565 16800 -535
rect 16750 -585 16765 -565
rect 16785 -585 16800 -565
rect 16750 -615 16800 -585
rect 16750 -635 16765 -615
rect 16785 -635 16800 -615
rect 16750 -665 16800 -635
rect 16750 -685 16765 -665
rect 16785 -685 16800 -665
rect 16750 -715 16800 -685
rect 16750 -735 16765 -715
rect 16785 -735 16800 -715
rect 16750 -765 16800 -735
rect 16750 -785 16765 -765
rect 16785 -785 16800 -765
rect 15700 -860 15750 -850
rect 15700 -890 15710 -860
rect 15740 -890 15750 -860
rect 15700 -900 15750 -890
rect 16000 -860 16050 -850
rect 16000 -890 16010 -860
rect 16040 -890 16050 -860
rect 16000 -900 16050 -890
rect 16300 -860 16350 -850
rect 16300 -890 16310 -860
rect 16340 -890 16350 -860
rect 16300 -900 16350 -890
rect 16600 -860 16650 -850
rect 16600 -890 16610 -860
rect 16640 -890 16650 -860
rect 16600 -900 16650 -890
rect 16750 -860 16800 -785
rect 17950 -115 18000 -40
rect 20350 -10 20400 65
rect 20350 -40 20360 -10
rect 20390 -40 20400 -10
rect 17950 -135 17965 -115
rect 17985 -135 18000 -115
rect 17950 -160 18000 -135
rect 17950 -190 17960 -160
rect 17990 -190 18000 -160
rect 17950 -215 18000 -190
rect 17950 -235 17965 -215
rect 17985 -235 18000 -215
rect 17950 -260 18000 -235
rect 17950 -290 17960 -260
rect 17990 -290 18000 -260
rect 17950 -315 18000 -290
rect 17950 -335 17965 -315
rect 17985 -335 18000 -315
rect 17950 -360 18000 -335
rect 17950 -390 17960 -360
rect 17990 -390 18000 -360
rect 17950 -415 18000 -390
rect 17950 -435 17965 -415
rect 17985 -435 18000 -415
rect 17950 -460 18000 -435
rect 17950 -490 17960 -460
rect 17990 -490 18000 -460
rect 17950 -515 18000 -490
rect 17950 -535 17965 -515
rect 17985 -535 18000 -515
rect 17950 -560 18000 -535
rect 17950 -590 17960 -560
rect 17990 -590 18000 -560
rect 17950 -615 18000 -590
rect 17950 -635 17965 -615
rect 17985 -635 18000 -615
rect 17950 -660 18000 -635
rect 17950 -690 17960 -660
rect 17990 -690 18000 -660
rect 17950 -715 18000 -690
rect 17950 -735 17965 -715
rect 17985 -735 18000 -715
rect 17950 -760 18000 -735
rect 17950 -790 17960 -760
rect 17990 -790 18000 -760
rect 16750 -890 16760 -860
rect 16790 -890 16800 -860
rect 15550 -990 15560 -960
rect 15590 -990 15600 -960
rect 15550 -1015 15600 -990
rect 15550 -1035 15565 -1015
rect 15585 -1035 15600 -1015
rect 15550 -1060 15600 -1035
rect 15550 -1090 15560 -1060
rect 15590 -1090 15600 -1060
rect 15550 -1115 15600 -1090
rect 15550 -1135 15565 -1115
rect 15585 -1135 15600 -1115
rect 15550 -1160 15600 -1135
rect 15550 -1190 15560 -1160
rect 15590 -1190 15600 -1160
rect 15550 -1215 15600 -1190
rect 15550 -1235 15565 -1215
rect 15585 -1235 15600 -1215
rect 15550 -1260 15600 -1235
rect 15550 -1290 15560 -1260
rect 15590 -1290 15600 -1260
rect 15550 -1315 15600 -1290
rect 15550 -1335 15565 -1315
rect 15585 -1335 15600 -1315
rect 15550 -1360 15600 -1335
rect 15550 -1390 15560 -1360
rect 15590 -1390 15600 -1360
rect 15550 -1415 15600 -1390
rect 15550 -1435 15565 -1415
rect 15585 -1435 15600 -1415
rect 15550 -1460 15600 -1435
rect 15550 -1490 15560 -1460
rect 15590 -1490 15600 -1460
rect 15550 -1515 15600 -1490
rect 15550 -1535 15565 -1515
rect 15585 -1535 15600 -1515
rect 15550 -1560 15600 -1535
rect 15550 -1590 15560 -1560
rect 15590 -1590 15600 -1560
rect 15550 -1615 15600 -1590
rect 15550 -1635 15565 -1615
rect 15585 -1635 15600 -1615
rect 10750 -1740 10760 -1710
rect 10790 -1740 10800 -1710
rect 10750 -1750 10800 -1740
rect 15550 -1710 15600 -1635
rect 16750 -965 16800 -890
rect 16900 -860 16950 -850
rect 16900 -890 16910 -860
rect 16940 -890 16950 -860
rect 16900 -900 16950 -890
rect 17200 -860 17250 -850
rect 17200 -890 17210 -860
rect 17240 -890 17250 -860
rect 17200 -900 17250 -890
rect 17500 -860 17550 -850
rect 17500 -890 17510 -860
rect 17540 -890 17550 -860
rect 17500 -900 17550 -890
rect 17800 -860 17850 -850
rect 17800 -890 17810 -860
rect 17840 -890 17850 -860
rect 17800 -900 17850 -890
rect 16750 -985 16765 -965
rect 16785 -985 16800 -965
rect 16750 -1015 16800 -985
rect 16750 -1035 16765 -1015
rect 16785 -1035 16800 -1015
rect 16750 -1065 16800 -1035
rect 16750 -1085 16765 -1065
rect 16785 -1085 16800 -1065
rect 16750 -1115 16800 -1085
rect 16750 -1135 16765 -1115
rect 16785 -1135 16800 -1115
rect 16750 -1165 16800 -1135
rect 16750 -1185 16765 -1165
rect 16785 -1185 16800 -1165
rect 16750 -1215 16800 -1185
rect 16750 -1235 16765 -1215
rect 16785 -1235 16800 -1215
rect 16750 -1265 16800 -1235
rect 16750 -1285 16765 -1265
rect 16785 -1285 16800 -1265
rect 16750 -1315 16800 -1285
rect 16750 -1335 16765 -1315
rect 16785 -1335 16800 -1315
rect 16750 -1365 16800 -1335
rect 16750 -1385 16765 -1365
rect 16785 -1385 16800 -1365
rect 16750 -1415 16800 -1385
rect 16750 -1435 16765 -1415
rect 16785 -1435 16800 -1415
rect 16750 -1465 16800 -1435
rect 16750 -1485 16765 -1465
rect 16785 -1485 16800 -1465
rect 16750 -1515 16800 -1485
rect 16750 -1535 16765 -1515
rect 16785 -1535 16800 -1515
rect 16750 -1565 16800 -1535
rect 16750 -1585 16765 -1565
rect 16785 -1585 16800 -1565
rect 16750 -1615 16800 -1585
rect 16750 -1635 16765 -1615
rect 16785 -1635 16800 -1615
rect 16750 -1650 16800 -1635
rect 17950 -960 18000 -790
rect 19150 -115 19200 -100
rect 19150 -135 19165 -115
rect 19185 -135 19200 -115
rect 19150 -165 19200 -135
rect 19150 -185 19165 -165
rect 19185 -185 19200 -165
rect 19150 -215 19200 -185
rect 19150 -235 19165 -215
rect 19185 -235 19200 -215
rect 19150 -265 19200 -235
rect 19150 -285 19165 -265
rect 19185 -285 19200 -265
rect 19150 -315 19200 -285
rect 19150 -335 19165 -315
rect 19185 -335 19200 -315
rect 19150 -365 19200 -335
rect 19150 -385 19165 -365
rect 19185 -385 19200 -365
rect 19150 -415 19200 -385
rect 19150 -435 19165 -415
rect 19185 -435 19200 -415
rect 19150 -465 19200 -435
rect 19150 -485 19165 -465
rect 19185 -485 19200 -465
rect 19150 -515 19200 -485
rect 19150 -535 19165 -515
rect 19185 -535 19200 -515
rect 19150 -565 19200 -535
rect 19150 -585 19165 -565
rect 19185 -585 19200 -565
rect 19150 -615 19200 -585
rect 19150 -635 19165 -615
rect 19185 -635 19200 -615
rect 19150 -665 19200 -635
rect 19150 -685 19165 -665
rect 19185 -685 19200 -665
rect 19150 -715 19200 -685
rect 19150 -735 19165 -715
rect 19185 -735 19200 -715
rect 19150 -765 19200 -735
rect 19150 -785 19165 -765
rect 19185 -785 19200 -765
rect 18100 -860 18150 -850
rect 18100 -890 18110 -860
rect 18140 -890 18150 -860
rect 18100 -900 18150 -890
rect 18400 -860 18450 -850
rect 18400 -890 18410 -860
rect 18440 -890 18450 -860
rect 18400 -900 18450 -890
rect 18700 -860 18750 -850
rect 18700 -890 18710 -860
rect 18740 -890 18750 -860
rect 18700 -900 18750 -890
rect 19000 -860 19050 -850
rect 19000 -890 19010 -860
rect 19040 -890 19050 -860
rect 19000 -900 19050 -890
rect 19150 -860 19200 -785
rect 20350 -115 20400 -40
rect 20350 -135 20365 -115
rect 20385 -135 20400 -115
rect 20350 -160 20400 -135
rect 20350 -190 20360 -160
rect 20390 -190 20400 -160
rect 20350 -215 20400 -190
rect 20350 -235 20365 -215
rect 20385 -235 20400 -215
rect 20350 -260 20400 -235
rect 20350 -290 20360 -260
rect 20390 -290 20400 -260
rect 20350 -315 20400 -290
rect 20350 -335 20365 -315
rect 20385 -335 20400 -315
rect 20350 -360 20400 -335
rect 20350 -390 20360 -360
rect 20390 -390 20400 -360
rect 20350 -415 20400 -390
rect 20350 -435 20365 -415
rect 20385 -435 20400 -415
rect 20350 -460 20400 -435
rect 20350 -490 20360 -460
rect 20390 -490 20400 -460
rect 20350 -515 20400 -490
rect 20350 -535 20365 -515
rect 20385 -535 20400 -515
rect 20350 -560 20400 -535
rect 20350 -590 20360 -560
rect 20390 -590 20400 -560
rect 20350 -615 20400 -590
rect 20350 -635 20365 -615
rect 20385 -635 20400 -615
rect 20350 -660 20400 -635
rect 20350 -690 20360 -660
rect 20390 -690 20400 -660
rect 20350 -715 20400 -690
rect 20350 -735 20365 -715
rect 20385 -735 20400 -715
rect 20350 -760 20400 -735
rect 20350 -790 20360 -760
rect 20390 -790 20400 -760
rect 19150 -890 19160 -860
rect 19190 -890 19200 -860
rect 17950 -990 17960 -960
rect 17990 -990 18000 -960
rect 17950 -1015 18000 -990
rect 17950 -1035 17965 -1015
rect 17985 -1035 18000 -1015
rect 17950 -1060 18000 -1035
rect 17950 -1090 17960 -1060
rect 17990 -1090 18000 -1060
rect 17950 -1115 18000 -1090
rect 17950 -1135 17965 -1115
rect 17985 -1135 18000 -1115
rect 17950 -1160 18000 -1135
rect 17950 -1190 17960 -1160
rect 17990 -1190 18000 -1160
rect 17950 -1215 18000 -1190
rect 17950 -1235 17965 -1215
rect 17985 -1235 18000 -1215
rect 17950 -1260 18000 -1235
rect 17950 -1290 17960 -1260
rect 17990 -1290 18000 -1260
rect 17950 -1315 18000 -1290
rect 17950 -1335 17965 -1315
rect 17985 -1335 18000 -1315
rect 17950 -1360 18000 -1335
rect 17950 -1390 17960 -1360
rect 17990 -1390 18000 -1360
rect 17950 -1415 18000 -1390
rect 17950 -1435 17965 -1415
rect 17985 -1435 18000 -1415
rect 17950 -1460 18000 -1435
rect 17950 -1490 17960 -1460
rect 17990 -1490 18000 -1460
rect 17950 -1515 18000 -1490
rect 17950 -1535 17965 -1515
rect 17985 -1535 18000 -1515
rect 17950 -1560 18000 -1535
rect 17950 -1590 17960 -1560
rect 17990 -1590 18000 -1560
rect 17950 -1615 18000 -1590
rect 17950 -1635 17965 -1615
rect 17985 -1635 18000 -1615
rect 15550 -1740 15560 -1710
rect 15590 -1740 15600 -1710
rect 15550 -1750 15600 -1740
rect 17950 -1710 18000 -1635
rect 19150 -965 19200 -890
rect 19300 -860 19350 -850
rect 19300 -890 19310 -860
rect 19340 -890 19350 -860
rect 19300 -900 19350 -890
rect 19600 -860 19650 -850
rect 19600 -890 19610 -860
rect 19640 -890 19650 -860
rect 19600 -900 19650 -890
rect 19900 -860 19950 -850
rect 19900 -890 19910 -860
rect 19940 -890 19950 -860
rect 19900 -900 19950 -890
rect 20200 -860 20250 -850
rect 20200 -890 20210 -860
rect 20240 -890 20250 -860
rect 20200 -900 20250 -890
rect 19150 -985 19165 -965
rect 19185 -985 19200 -965
rect 19150 -1015 19200 -985
rect 19150 -1035 19165 -1015
rect 19185 -1035 19200 -1015
rect 19150 -1065 19200 -1035
rect 19150 -1085 19165 -1065
rect 19185 -1085 19200 -1065
rect 19150 -1115 19200 -1085
rect 19150 -1135 19165 -1115
rect 19185 -1135 19200 -1115
rect 19150 -1165 19200 -1135
rect 19150 -1185 19165 -1165
rect 19185 -1185 19200 -1165
rect 19150 -1215 19200 -1185
rect 19150 -1235 19165 -1215
rect 19185 -1235 19200 -1215
rect 19150 -1265 19200 -1235
rect 19150 -1285 19165 -1265
rect 19185 -1285 19200 -1265
rect 19150 -1315 19200 -1285
rect 19150 -1335 19165 -1315
rect 19185 -1335 19200 -1315
rect 19150 -1365 19200 -1335
rect 19150 -1385 19165 -1365
rect 19185 -1385 19200 -1365
rect 19150 -1415 19200 -1385
rect 19150 -1435 19165 -1415
rect 19185 -1435 19200 -1415
rect 19150 -1465 19200 -1435
rect 19150 -1485 19165 -1465
rect 19185 -1485 19200 -1465
rect 19150 -1515 19200 -1485
rect 19150 -1535 19165 -1515
rect 19185 -1535 19200 -1515
rect 19150 -1565 19200 -1535
rect 19150 -1585 19165 -1565
rect 19185 -1585 19200 -1565
rect 19150 -1615 19200 -1585
rect 19150 -1635 19165 -1615
rect 19185 -1635 19200 -1615
rect 19150 -1650 19200 -1635
rect 20350 -960 20400 -790
rect 20350 -990 20360 -960
rect 20390 -990 20400 -960
rect 20350 -1015 20400 -990
rect 20350 -1035 20365 -1015
rect 20385 -1035 20400 -1015
rect 20350 -1060 20400 -1035
rect 20350 -1090 20360 -1060
rect 20390 -1090 20400 -1060
rect 20350 -1115 20400 -1090
rect 20350 -1135 20365 -1115
rect 20385 -1135 20400 -1115
rect 20350 -1160 20400 -1135
rect 20350 -1190 20360 -1160
rect 20390 -1190 20400 -1160
rect 20350 -1215 20400 -1190
rect 20350 -1235 20365 -1215
rect 20385 -1235 20400 -1215
rect 20350 -1260 20400 -1235
rect 20350 -1290 20360 -1260
rect 20390 -1290 20400 -1260
rect 20350 -1315 20400 -1290
rect 20350 -1335 20365 -1315
rect 20385 -1335 20400 -1315
rect 20350 -1360 20400 -1335
rect 20350 -1390 20360 -1360
rect 20390 -1390 20400 -1360
rect 20350 -1415 20400 -1390
rect 20350 -1435 20365 -1415
rect 20385 -1435 20400 -1415
rect 20350 -1460 20400 -1435
rect 20350 -1490 20360 -1460
rect 20390 -1490 20400 -1460
rect 20350 -1515 20400 -1490
rect 20350 -1535 20365 -1515
rect 20385 -1535 20400 -1515
rect 20350 -1560 20400 -1535
rect 20350 -1590 20360 -1560
rect 20390 -1590 20400 -1560
rect 20350 -1615 20400 -1590
rect 20350 -1635 20365 -1615
rect 20385 -1635 20400 -1615
rect 17950 -1740 17960 -1710
rect 17990 -1740 18000 -1710
rect 17950 -1750 18000 -1740
rect 20350 -1710 20400 -1635
rect 20350 -1740 20360 -1710
rect 20390 -1740 20400 -1710
rect 20350 -1750 20400 -1740
<< via1 >>
rect -640 5185 -610 5190
rect -640 5165 -635 5185
rect -635 5165 -615 5185
rect -615 5165 -610 5185
rect -640 5160 -610 5165
rect -40 5160 -10 5190
rect -640 5035 -610 5040
rect -640 5015 -635 5035
rect -635 5015 -615 5035
rect -615 5015 -610 5035
rect -640 5010 -610 5015
rect -640 4935 -610 4940
rect -640 4915 -635 4935
rect -635 4915 -615 4935
rect -615 4915 -610 4935
rect -640 4910 -610 4915
rect -640 4835 -610 4840
rect -640 4815 -635 4835
rect -635 4815 -615 4835
rect -615 4815 -610 4835
rect -640 4810 -610 4815
rect -640 4735 -610 4740
rect -640 4715 -635 4735
rect -635 4715 -615 4735
rect -615 4715 -610 4735
rect -640 4710 -610 4715
rect -640 4635 -610 4640
rect -640 4615 -635 4635
rect -635 4615 -615 4635
rect -615 4615 -610 4635
rect -640 4610 -610 4615
rect 4160 5160 4190 5190
rect -490 4535 -460 4540
rect -490 4515 -485 4535
rect -485 4515 -465 4535
rect -465 4515 -460 4535
rect -490 4510 -460 4515
rect -340 4510 -310 4540
rect -190 4535 -160 4540
rect -190 4515 -185 4535
rect -185 4515 -165 4535
rect -165 4515 -160 4535
rect -190 4510 -160 4515
rect -640 4435 -610 4440
rect -640 4415 -635 4435
rect -635 4415 -615 4435
rect -615 4415 -610 4435
rect -640 4410 -610 4415
rect -640 4335 -610 4340
rect -640 4315 -635 4335
rect -635 4315 -615 4335
rect -615 4315 -610 4335
rect -640 4310 -610 4315
rect -640 4235 -610 4240
rect -640 4215 -635 4235
rect -635 4215 -615 4235
rect -615 4215 -610 4235
rect -640 4210 -610 4215
rect -640 4135 -610 4140
rect -640 4115 -635 4135
rect -635 4115 -615 4135
rect -615 4115 -610 4135
rect -640 4110 -610 4115
rect -640 4035 -610 4040
rect -640 4015 -635 4035
rect -635 4015 -615 4035
rect -615 4015 -610 4035
rect -640 4010 -610 4015
rect 110 4535 140 4540
rect 110 4515 115 4535
rect 115 4515 135 4535
rect 135 4515 140 4535
rect 110 4510 140 4515
rect 410 4535 440 4540
rect 410 4515 415 4535
rect 415 4515 435 4535
rect 435 4515 440 4535
rect 410 4510 440 4515
rect 710 4535 740 4540
rect 710 4515 715 4535
rect 715 4515 735 4535
rect 735 4515 740 4535
rect 710 4510 740 4515
rect 1010 4535 1040 4540
rect 1010 4515 1015 4535
rect 1015 4515 1035 4535
rect 1035 4515 1040 4535
rect 1010 4510 1040 4515
rect 1160 4510 1190 4540
rect 1310 4535 1340 4540
rect 1310 4515 1315 4535
rect 1315 4515 1335 4535
rect 1335 4515 1340 4535
rect 1310 4510 1340 4515
rect 1610 4535 1640 4540
rect 1610 4515 1615 4535
rect 1615 4515 1635 4535
rect 1635 4515 1640 4535
rect 1610 4510 1640 4515
rect -40 4410 -10 4440
rect -40 4335 -10 4340
rect -40 4315 -35 4335
rect -35 4315 -15 4335
rect -15 4315 -10 4335
rect -40 4310 -10 4315
rect -40 4235 -10 4240
rect -40 4215 -35 4235
rect -35 4215 -15 4235
rect -15 4215 -10 4235
rect -40 4210 -10 4215
rect -40 4135 -10 4140
rect -40 4115 -35 4135
rect -35 4115 -15 4135
rect -15 4115 -10 4135
rect -40 4110 -10 4115
rect -40 4035 -10 4040
rect -40 4015 -35 4035
rect -35 4015 -15 4035
rect -15 4015 -10 4035
rect -40 4010 -10 4015
rect -640 3885 -610 3890
rect -640 3865 -635 3885
rect -635 3865 -615 3885
rect -615 3865 -610 3885
rect -640 3860 -610 3865
rect 1910 4535 1940 4540
rect 1910 4515 1915 4535
rect 1915 4515 1935 4535
rect 1935 4515 1940 4535
rect 1910 4510 1940 4515
rect 2060 4510 2090 4540
rect 2210 4535 2240 4540
rect 2210 4515 2215 4535
rect 2215 4515 2235 4535
rect 2235 4515 2240 4535
rect 2210 4510 2240 4515
rect 8360 5185 8390 5190
rect 8360 5165 8365 5185
rect 8365 5165 8385 5185
rect 8385 5165 8390 5185
rect 8360 5160 8390 5165
rect 2510 4535 2540 4540
rect 2510 4515 2515 4535
rect 2515 4515 2535 4535
rect 2535 4515 2540 4535
rect 2510 4510 2540 4515
rect 2810 4535 2840 4540
rect 2810 4515 2815 4535
rect 2815 4515 2835 4535
rect 2835 4515 2840 4535
rect 2810 4510 2840 4515
rect 2960 4510 2990 4540
rect 3110 4535 3140 4540
rect 3110 4515 3115 4535
rect 3115 4515 3135 4535
rect 3135 4515 3140 4535
rect 3110 4510 3140 4515
rect 3410 4535 3440 4540
rect 3410 4515 3415 4535
rect 3415 4515 3435 4535
rect 3435 4515 3440 4535
rect 3410 4510 3440 4515
rect 3710 4535 3740 4540
rect 3710 4515 3715 4535
rect 3715 4515 3735 4535
rect 3735 4515 3740 4535
rect 3710 4510 3740 4515
rect 4010 4535 4040 4540
rect 4010 4515 4015 4535
rect 4015 4515 4035 4535
rect 4035 4515 4040 4535
rect 4010 4510 4040 4515
rect 4310 4535 4340 4540
rect 4310 4515 4315 4535
rect 4315 4515 4335 4535
rect 4335 4515 4340 4535
rect 4310 4510 4340 4515
rect 4610 4535 4640 4540
rect 4610 4515 4615 4535
rect 4615 4515 4635 4535
rect 4635 4515 4640 4535
rect 4610 4510 4640 4515
rect 4910 4535 4940 4540
rect 4910 4515 4915 4535
rect 4915 4515 4935 4535
rect 4935 4515 4940 4535
rect 4910 4510 4940 4515
rect 5210 4535 5240 4540
rect 5210 4515 5215 4535
rect 5215 4515 5235 4535
rect 5235 4515 5240 4535
rect 5210 4510 5240 4515
rect 5360 4510 5390 4540
rect 5510 4535 5540 4540
rect 5510 4515 5515 4535
rect 5515 4515 5535 4535
rect 5535 4515 5540 4535
rect 5510 4510 5540 4515
rect 5810 4535 5840 4540
rect 5810 4515 5815 4535
rect 5815 4515 5835 4535
rect 5835 4515 5840 4535
rect 5810 4510 5840 4515
rect 4160 4410 4190 4440
rect 4160 4335 4190 4340
rect 4160 4315 4165 4335
rect 4165 4315 4185 4335
rect 4185 4315 4190 4335
rect 4160 4310 4190 4315
rect 4160 4235 4190 4240
rect 4160 4215 4165 4235
rect 4165 4215 4185 4235
rect 4185 4215 4190 4235
rect 4160 4210 4190 4215
rect 4160 4135 4190 4140
rect 4160 4115 4165 4135
rect 4165 4115 4185 4135
rect 4185 4115 4190 4135
rect 4160 4110 4190 4115
rect 4160 4035 4190 4040
rect 4160 4015 4165 4035
rect 4165 4015 4185 4035
rect 4185 4015 4190 4035
rect 4160 4010 4190 4015
rect -40 3885 -10 3890
rect -40 3865 -35 3885
rect -35 3865 -15 3885
rect -15 3865 -10 3885
rect -40 3860 -10 3865
rect -640 3735 -610 3740
rect -640 3715 -635 3735
rect -635 3715 -615 3735
rect -615 3715 -610 3735
rect -640 3710 -610 3715
rect -640 3635 -610 3640
rect -640 3615 -635 3635
rect -635 3615 -615 3635
rect -615 3615 -610 3635
rect -640 3610 -610 3615
rect -640 3535 -610 3540
rect -640 3515 -635 3535
rect -635 3515 -615 3535
rect -615 3515 -610 3535
rect -640 3510 -610 3515
rect -640 3435 -610 3440
rect -640 3415 -635 3435
rect -635 3415 -615 3435
rect -615 3415 -610 3435
rect -640 3410 -610 3415
rect -640 3335 -610 3340
rect -640 3315 -635 3335
rect -635 3315 -615 3335
rect -615 3315 -610 3335
rect -640 3310 -610 3315
rect 6110 4535 6140 4540
rect 6110 4515 6115 4535
rect 6115 4515 6135 4535
rect 6135 4515 6140 4535
rect 6110 4510 6140 4515
rect 6260 4510 6290 4540
rect 6410 4535 6440 4540
rect 6410 4515 6415 4535
rect 6415 4515 6435 4535
rect 6435 4515 6440 4535
rect 6410 4510 6440 4515
rect 8660 5185 8690 5190
rect 8660 5165 8665 5185
rect 8665 5165 8685 5185
rect 8685 5165 8690 5185
rect 8660 5160 8690 5165
rect 8360 5035 8390 5040
rect 8360 5015 8365 5035
rect 8365 5015 8385 5035
rect 8385 5015 8390 5035
rect 8360 5010 8390 5015
rect 8360 4935 8390 4940
rect 8360 4915 8365 4935
rect 8365 4915 8385 4935
rect 8385 4915 8390 4935
rect 8360 4910 8390 4915
rect 8360 4835 8390 4840
rect 8360 4815 8365 4835
rect 8365 4815 8385 4835
rect 8385 4815 8390 4835
rect 8360 4810 8390 4815
rect 8360 4735 8390 4740
rect 8360 4715 8365 4735
rect 8365 4715 8385 4735
rect 8385 4715 8390 4735
rect 8360 4710 8390 4715
rect 8360 4635 8390 4640
rect 8360 4615 8365 4635
rect 8365 4615 8385 4635
rect 8385 4615 8390 4635
rect 8360 4610 8390 4615
rect 6710 4535 6740 4540
rect 6710 4515 6715 4535
rect 6715 4515 6735 4535
rect 6735 4515 6740 4535
rect 6710 4510 6740 4515
rect 7010 4535 7040 4540
rect 7010 4515 7015 4535
rect 7015 4515 7035 4535
rect 7035 4515 7040 4535
rect 7010 4510 7040 4515
rect 7160 4510 7190 4540
rect 7310 4535 7340 4540
rect 7310 4515 7315 4535
rect 7315 4515 7335 4535
rect 7335 4515 7340 4535
rect 7310 4510 7340 4515
rect 7610 4535 7640 4540
rect 7610 4515 7615 4535
rect 7615 4515 7635 4535
rect 7635 4515 7640 4535
rect 7610 4510 7640 4515
rect 7910 4535 7940 4540
rect 7910 4515 7915 4535
rect 7915 4515 7935 4535
rect 7935 4515 7940 4535
rect 7910 4510 7940 4515
rect 8210 4535 8240 4540
rect 8210 4515 8215 4535
rect 8215 4515 8235 4535
rect 8235 4515 8240 4535
rect 8210 4510 8240 4515
rect 8960 5185 8990 5190
rect 8960 5165 8965 5185
rect 8965 5165 8985 5185
rect 8985 5165 8990 5185
rect 8960 5160 8990 5165
rect 8660 5035 8690 5040
rect 8660 5015 8665 5035
rect 8665 5015 8685 5035
rect 8685 5015 8690 5035
rect 8660 5010 8690 5015
rect 8660 4935 8690 4940
rect 8660 4915 8665 4935
rect 8665 4915 8685 4935
rect 8685 4915 8690 4935
rect 8660 4910 8690 4915
rect 8660 4835 8690 4840
rect 8660 4815 8665 4835
rect 8665 4815 8685 4835
rect 8685 4815 8690 4835
rect 8660 4810 8690 4815
rect 8660 4735 8690 4740
rect 8660 4715 8665 4735
rect 8665 4715 8685 4735
rect 8685 4715 8690 4735
rect 8660 4710 8690 4715
rect 8660 4635 8690 4640
rect 8660 4615 8665 4635
rect 8665 4615 8685 4635
rect 8685 4615 8690 4635
rect 8660 4610 8690 4615
rect 8510 4535 8540 4540
rect 8510 4515 8515 4535
rect 8515 4515 8535 4535
rect 8535 4515 8540 4535
rect 8510 4510 8540 4515
rect 8360 4435 8390 4440
rect 8360 4415 8365 4435
rect 8365 4415 8385 4435
rect 8385 4415 8390 4435
rect 8360 4410 8390 4415
rect 8360 4335 8390 4340
rect 8360 4315 8365 4335
rect 8365 4315 8385 4335
rect 8385 4315 8390 4335
rect 8360 4310 8390 4315
rect 8360 4235 8390 4240
rect 8360 4215 8365 4235
rect 8365 4215 8385 4235
rect 8385 4215 8390 4235
rect 8360 4210 8390 4215
rect 8360 4135 8390 4140
rect 8360 4115 8365 4135
rect 8365 4115 8385 4135
rect 8385 4115 8390 4135
rect 8360 4110 8390 4115
rect 8360 4035 8390 4040
rect 8360 4015 8365 4035
rect 8365 4015 8385 4035
rect 8385 4015 8390 4035
rect 8360 4010 8390 4015
rect 4160 3885 4190 3890
rect 4160 3865 4165 3885
rect 4165 3865 4185 3885
rect 4185 3865 4190 3885
rect 4160 3860 4190 3865
rect -490 3235 -460 3240
rect -490 3215 -485 3235
rect -485 3215 -465 3235
rect -465 3215 -460 3235
rect -490 3210 -460 3215
rect -340 3210 -310 3240
rect -190 3235 -160 3240
rect -190 3215 -185 3235
rect -185 3215 -165 3235
rect -165 3215 -160 3235
rect -190 3210 -160 3215
rect -640 3135 -610 3140
rect -640 3115 -635 3135
rect -635 3115 -615 3135
rect -615 3115 -610 3135
rect -640 3110 -610 3115
rect -640 3035 -610 3040
rect -640 3015 -635 3035
rect -635 3015 -615 3035
rect -615 3015 -610 3035
rect -640 3010 -610 3015
rect -640 2935 -610 2940
rect -640 2915 -635 2935
rect -635 2915 -615 2935
rect -615 2915 -610 2935
rect -640 2910 -610 2915
rect -640 2835 -610 2840
rect -640 2815 -635 2835
rect -635 2815 -615 2835
rect -615 2815 -610 2835
rect -640 2810 -610 2815
rect -640 2735 -610 2740
rect -640 2715 -635 2735
rect -635 2715 -615 2735
rect -615 2715 -610 2735
rect -640 2710 -610 2715
rect 110 3235 140 3240
rect 110 3215 115 3235
rect 115 3215 135 3235
rect 135 3215 140 3235
rect 110 3210 140 3215
rect 410 3235 440 3240
rect 410 3215 415 3235
rect 415 3215 435 3235
rect 435 3215 440 3235
rect 410 3210 440 3215
rect -40 3110 -10 3140
rect -40 3035 -10 3040
rect -40 3015 -35 3035
rect -35 3015 -15 3035
rect -15 3015 -10 3035
rect -40 3010 -10 3015
rect -40 2935 -10 2940
rect -40 2915 -35 2935
rect -35 2915 -15 2935
rect -15 2915 -10 2935
rect -40 2910 -10 2915
rect -40 2835 -10 2840
rect -40 2815 -35 2835
rect -35 2815 -15 2835
rect -15 2815 -10 2835
rect -40 2810 -10 2815
rect -40 2735 -10 2740
rect -40 2715 -35 2735
rect -35 2715 -15 2735
rect -15 2715 -10 2735
rect -40 2710 -10 2715
rect -640 2585 -610 2590
rect -640 2565 -635 2585
rect -635 2565 -615 2585
rect -615 2565 -610 2585
rect -640 2560 -610 2565
rect 710 3235 740 3240
rect 710 3215 715 3235
rect 715 3215 735 3235
rect 735 3215 740 3235
rect 710 3210 740 3215
rect 1010 3235 1040 3240
rect 1010 3215 1015 3235
rect 1015 3215 1035 3235
rect 1035 3215 1040 3235
rect 1010 3210 1040 3215
rect 1160 3210 1190 3240
rect 1310 3235 1340 3240
rect 1310 3215 1315 3235
rect 1315 3215 1335 3235
rect 1335 3215 1340 3235
rect 1310 3210 1340 3215
rect 1610 3235 1640 3240
rect 1610 3215 1615 3235
rect 1615 3215 1635 3235
rect 1635 3215 1640 3235
rect 1610 3210 1640 3215
rect 1910 3235 1940 3240
rect 1910 3215 1915 3235
rect 1915 3215 1935 3235
rect 1935 3215 1940 3235
rect 1910 3210 1940 3215
rect 2060 3210 2090 3240
rect 2210 3235 2240 3240
rect 2210 3215 2215 3235
rect 2215 3215 2235 3235
rect 2235 3215 2240 3235
rect 2210 3210 2240 3215
rect 2510 3235 2540 3240
rect 2510 3215 2515 3235
rect 2515 3215 2535 3235
rect 2535 3215 2540 3235
rect 2510 3210 2540 3215
rect 2810 3235 2840 3240
rect 2810 3215 2815 3235
rect 2815 3215 2835 3235
rect 2835 3215 2840 3235
rect 2810 3210 2840 3215
rect 2960 3210 2990 3240
rect 3110 3235 3140 3240
rect 3110 3215 3115 3235
rect 3115 3215 3135 3235
rect 3135 3215 3140 3235
rect 3110 3210 3140 3215
rect 3410 3235 3440 3240
rect 3410 3215 3415 3235
rect 3415 3215 3435 3235
rect 3435 3215 3440 3235
rect 3410 3210 3440 3215
rect 9260 5185 9290 5190
rect 9260 5165 9265 5185
rect 9265 5165 9285 5185
rect 9285 5165 9290 5185
rect 9260 5160 9290 5165
rect 8960 5035 8990 5040
rect 8960 5015 8965 5035
rect 8965 5015 8985 5035
rect 8985 5015 8990 5035
rect 8960 5010 8990 5015
rect 8960 4935 8990 4940
rect 8960 4915 8965 4935
rect 8965 4915 8985 4935
rect 8985 4915 8990 4935
rect 8960 4910 8990 4915
rect 8960 4835 8990 4840
rect 8960 4815 8965 4835
rect 8965 4815 8985 4835
rect 8985 4815 8990 4835
rect 8960 4810 8990 4815
rect 8960 4735 8990 4740
rect 8960 4715 8965 4735
rect 8965 4715 8985 4735
rect 8985 4715 8990 4735
rect 8960 4710 8990 4715
rect 8960 4635 8990 4640
rect 8960 4615 8965 4635
rect 8965 4615 8985 4635
rect 8985 4615 8990 4635
rect 8960 4610 8990 4615
rect 8810 4535 8840 4540
rect 8810 4515 8815 4535
rect 8815 4515 8835 4535
rect 8835 4515 8840 4535
rect 8810 4510 8840 4515
rect 8660 4435 8690 4440
rect 8660 4415 8665 4435
rect 8665 4415 8685 4435
rect 8685 4415 8690 4435
rect 8660 4410 8690 4415
rect 8660 4335 8690 4340
rect 8660 4315 8665 4335
rect 8665 4315 8685 4335
rect 8685 4315 8690 4335
rect 8660 4310 8690 4315
rect 8660 4235 8690 4240
rect 8660 4215 8665 4235
rect 8665 4215 8685 4235
rect 8685 4215 8690 4235
rect 8660 4210 8690 4215
rect 8660 4135 8690 4140
rect 8660 4115 8665 4135
rect 8665 4115 8685 4135
rect 8685 4115 8690 4135
rect 8660 4110 8690 4115
rect 8660 4035 8690 4040
rect 8660 4015 8665 4035
rect 8665 4015 8685 4035
rect 8685 4015 8690 4035
rect 8660 4010 8690 4015
rect 8360 3885 8390 3890
rect 8360 3865 8365 3885
rect 8365 3865 8385 3885
rect 8385 3865 8390 3885
rect 8360 3860 8390 3865
rect 3710 3235 3740 3240
rect 3710 3215 3715 3235
rect 3715 3215 3735 3235
rect 3735 3215 3740 3235
rect 3710 3210 3740 3215
rect 4010 3235 4040 3240
rect 4010 3215 4015 3235
rect 4015 3215 4035 3235
rect 4035 3215 4040 3235
rect 4010 3210 4040 3215
rect 4310 3235 4340 3240
rect 4310 3215 4315 3235
rect 4315 3215 4335 3235
rect 4335 3215 4340 3235
rect 4310 3210 4340 3215
rect 4610 3235 4640 3240
rect 4610 3215 4615 3235
rect 4615 3215 4635 3235
rect 4635 3215 4640 3235
rect 4610 3210 4640 3215
rect 4160 3110 4190 3140
rect 4160 3035 4190 3040
rect 4160 3015 4165 3035
rect 4165 3015 4185 3035
rect 4185 3015 4190 3035
rect 4160 3010 4190 3015
rect 4160 2935 4190 2940
rect 4160 2915 4165 2935
rect 4165 2915 4185 2935
rect 4185 2915 4190 2935
rect 4160 2910 4190 2915
rect 4160 2835 4190 2840
rect 4160 2815 4165 2835
rect 4165 2815 4185 2835
rect 4185 2815 4190 2835
rect 4160 2810 4190 2815
rect 4160 2735 4190 2740
rect 4160 2715 4165 2735
rect 4165 2715 4185 2735
rect 4185 2715 4190 2735
rect 4160 2710 4190 2715
rect -40 2585 -10 2590
rect -40 2565 -35 2585
rect -35 2565 -15 2585
rect -15 2565 -10 2585
rect -40 2560 -10 2565
rect 4910 3235 4940 3240
rect 4910 3215 4915 3235
rect 4915 3215 4935 3235
rect 4935 3215 4940 3235
rect 4910 3210 4940 3215
rect 5210 3235 5240 3240
rect 5210 3215 5215 3235
rect 5215 3215 5235 3235
rect 5235 3215 5240 3235
rect 5210 3210 5240 3215
rect 5360 3210 5390 3240
rect 5510 3235 5540 3240
rect 5510 3215 5515 3235
rect 5515 3215 5535 3235
rect 5535 3215 5540 3235
rect 5510 3210 5540 3215
rect 5810 3235 5840 3240
rect 5810 3215 5815 3235
rect 5815 3215 5835 3235
rect 5835 3215 5840 3235
rect 5810 3210 5840 3215
rect 6110 3235 6140 3240
rect 6110 3215 6115 3235
rect 6115 3215 6135 3235
rect 6135 3215 6140 3235
rect 6110 3210 6140 3215
rect 6260 3210 6290 3240
rect 6410 3235 6440 3240
rect 6410 3215 6415 3235
rect 6415 3215 6435 3235
rect 6435 3215 6440 3235
rect 6410 3210 6440 3215
rect 6710 3235 6740 3240
rect 6710 3215 6715 3235
rect 6715 3215 6735 3235
rect 6735 3215 6740 3235
rect 6710 3210 6740 3215
rect 7010 3235 7040 3240
rect 7010 3215 7015 3235
rect 7015 3215 7035 3235
rect 7035 3215 7040 3235
rect 7010 3210 7040 3215
rect 7160 3210 7190 3240
rect 7310 3235 7340 3240
rect 7310 3215 7315 3235
rect 7315 3215 7335 3235
rect 7335 3215 7340 3235
rect 7310 3210 7340 3215
rect 7610 3235 7640 3240
rect 7610 3215 7615 3235
rect 7615 3215 7635 3235
rect 7635 3215 7640 3235
rect 7610 3210 7640 3215
rect 9560 5185 9590 5190
rect 9560 5165 9565 5185
rect 9565 5165 9585 5185
rect 9585 5165 9590 5185
rect 9560 5160 9590 5165
rect 9260 5035 9290 5040
rect 9260 5015 9265 5035
rect 9265 5015 9285 5035
rect 9285 5015 9290 5035
rect 9260 5010 9290 5015
rect 9260 4935 9290 4940
rect 9260 4915 9265 4935
rect 9265 4915 9285 4935
rect 9285 4915 9290 4935
rect 9260 4910 9290 4915
rect 9260 4835 9290 4840
rect 9260 4815 9265 4835
rect 9265 4815 9285 4835
rect 9285 4815 9290 4835
rect 9260 4810 9290 4815
rect 9260 4735 9290 4740
rect 9260 4715 9265 4735
rect 9265 4715 9285 4735
rect 9285 4715 9290 4735
rect 9260 4710 9290 4715
rect 9260 4635 9290 4640
rect 9260 4615 9265 4635
rect 9265 4615 9285 4635
rect 9285 4615 9290 4635
rect 9260 4610 9290 4615
rect 9110 4535 9140 4540
rect 9110 4515 9115 4535
rect 9115 4515 9135 4535
rect 9135 4515 9140 4535
rect 9110 4510 9140 4515
rect 8960 4435 8990 4440
rect 8960 4415 8965 4435
rect 8965 4415 8985 4435
rect 8985 4415 8990 4435
rect 8960 4410 8990 4415
rect 8960 4335 8990 4340
rect 8960 4315 8965 4335
rect 8965 4315 8985 4335
rect 8985 4315 8990 4335
rect 8960 4310 8990 4315
rect 8960 4235 8990 4240
rect 8960 4215 8965 4235
rect 8965 4215 8985 4235
rect 8985 4215 8990 4235
rect 8960 4210 8990 4215
rect 8960 4135 8990 4140
rect 8960 4115 8965 4135
rect 8965 4115 8985 4135
rect 8985 4115 8990 4135
rect 8960 4110 8990 4115
rect 8960 4035 8990 4040
rect 8960 4015 8965 4035
rect 8965 4015 8985 4035
rect 8985 4015 8990 4035
rect 8960 4010 8990 4015
rect 8660 3885 8690 3890
rect 8660 3865 8665 3885
rect 8665 3865 8685 3885
rect 8685 3865 8690 3885
rect 8660 3860 8690 3865
rect 8360 3735 8390 3740
rect 8360 3715 8365 3735
rect 8365 3715 8385 3735
rect 8385 3715 8390 3735
rect 8360 3710 8390 3715
rect 8360 3635 8390 3640
rect 8360 3615 8365 3635
rect 8365 3615 8385 3635
rect 8385 3615 8390 3635
rect 8360 3610 8390 3615
rect 8360 3535 8390 3540
rect 8360 3515 8365 3535
rect 8365 3515 8385 3535
rect 8385 3515 8390 3535
rect 8360 3510 8390 3515
rect 8360 3435 8390 3440
rect 8360 3415 8365 3435
rect 8365 3415 8385 3435
rect 8385 3415 8390 3435
rect 8360 3410 8390 3415
rect 8360 3335 8390 3340
rect 8360 3315 8365 3335
rect 8365 3315 8385 3335
rect 8385 3315 8390 3335
rect 8360 3310 8390 3315
rect 7910 3235 7940 3240
rect 7910 3215 7915 3235
rect 7915 3215 7935 3235
rect 7935 3215 7940 3235
rect 7910 3210 7940 3215
rect 8210 3235 8240 3240
rect 8210 3215 8215 3235
rect 8215 3215 8235 3235
rect 8235 3215 8240 3235
rect 8210 3210 8240 3215
rect 9860 5185 9890 5190
rect 9860 5165 9865 5185
rect 9865 5165 9885 5185
rect 9885 5165 9890 5185
rect 9860 5160 9890 5165
rect 9560 5035 9590 5040
rect 9560 5015 9565 5035
rect 9565 5015 9585 5035
rect 9585 5015 9590 5035
rect 9560 5010 9590 5015
rect 9560 4935 9590 4940
rect 9560 4915 9565 4935
rect 9565 4915 9585 4935
rect 9585 4915 9590 4935
rect 9560 4910 9590 4915
rect 9560 4835 9590 4840
rect 9560 4815 9565 4835
rect 9565 4815 9585 4835
rect 9585 4815 9590 4835
rect 9560 4810 9590 4815
rect 9560 4735 9590 4740
rect 9560 4715 9565 4735
rect 9565 4715 9585 4735
rect 9585 4715 9590 4735
rect 9560 4710 9590 4715
rect 9560 4635 9590 4640
rect 9560 4615 9565 4635
rect 9565 4615 9585 4635
rect 9585 4615 9590 4635
rect 9560 4610 9590 4615
rect 9410 4535 9440 4540
rect 9410 4515 9415 4535
rect 9415 4515 9435 4535
rect 9435 4515 9440 4535
rect 9410 4510 9440 4515
rect 9260 4435 9290 4440
rect 9260 4415 9265 4435
rect 9265 4415 9285 4435
rect 9285 4415 9290 4435
rect 9260 4410 9290 4415
rect 9260 4335 9290 4340
rect 9260 4315 9265 4335
rect 9265 4315 9285 4335
rect 9285 4315 9290 4335
rect 9260 4310 9290 4315
rect 9260 4235 9290 4240
rect 9260 4215 9265 4235
rect 9265 4215 9285 4235
rect 9285 4215 9290 4235
rect 9260 4210 9290 4215
rect 9260 4135 9290 4140
rect 9260 4115 9265 4135
rect 9265 4115 9285 4135
rect 9285 4115 9290 4135
rect 9260 4110 9290 4115
rect 9260 4035 9290 4040
rect 9260 4015 9265 4035
rect 9265 4015 9285 4035
rect 9285 4015 9290 4035
rect 9260 4010 9290 4015
rect 8960 3885 8990 3890
rect 8960 3865 8965 3885
rect 8965 3865 8985 3885
rect 8985 3865 8990 3885
rect 8960 3860 8990 3865
rect 8660 3735 8690 3740
rect 8660 3715 8665 3735
rect 8665 3715 8685 3735
rect 8685 3715 8690 3735
rect 8660 3710 8690 3715
rect 8660 3635 8690 3640
rect 8660 3615 8665 3635
rect 8665 3615 8685 3635
rect 8685 3615 8690 3635
rect 8660 3610 8690 3615
rect 8660 3535 8690 3540
rect 8660 3515 8665 3535
rect 8665 3515 8685 3535
rect 8685 3515 8690 3535
rect 8660 3510 8690 3515
rect 8660 3435 8690 3440
rect 8660 3415 8665 3435
rect 8665 3415 8685 3435
rect 8685 3415 8690 3435
rect 8660 3410 8690 3415
rect 8660 3335 8690 3340
rect 8660 3315 8665 3335
rect 8665 3315 8685 3335
rect 8685 3315 8690 3335
rect 8660 3310 8690 3315
rect 8510 3235 8540 3240
rect 8510 3215 8515 3235
rect 8515 3215 8535 3235
rect 8535 3215 8540 3235
rect 8510 3210 8540 3215
rect 8360 3135 8390 3140
rect 8360 3115 8365 3135
rect 8365 3115 8385 3135
rect 8385 3115 8390 3135
rect 8360 3110 8390 3115
rect 8360 3035 8390 3040
rect 8360 3015 8365 3035
rect 8365 3015 8385 3035
rect 8385 3015 8390 3035
rect 8360 3010 8390 3015
rect 8360 2935 8390 2940
rect 8360 2915 8365 2935
rect 8365 2915 8385 2935
rect 8385 2915 8390 2935
rect 8360 2910 8390 2915
rect 8360 2835 8390 2840
rect 8360 2815 8365 2835
rect 8365 2815 8385 2835
rect 8385 2815 8390 2835
rect 8360 2810 8390 2815
rect 8360 2735 8390 2740
rect 8360 2715 8365 2735
rect 8365 2715 8385 2735
rect 8385 2715 8390 2735
rect 8360 2710 8390 2715
rect 4160 2585 4190 2590
rect 4160 2565 4165 2585
rect 4165 2565 4185 2585
rect 4185 2565 4190 2585
rect 4160 2560 4190 2565
rect 10160 5185 10190 5190
rect 10160 5165 10165 5185
rect 10165 5165 10185 5185
rect 10185 5165 10190 5185
rect 10160 5160 10190 5165
rect 9860 5035 9890 5040
rect 9860 5015 9865 5035
rect 9865 5015 9885 5035
rect 9885 5015 9890 5035
rect 9860 5010 9890 5015
rect 9860 4935 9890 4940
rect 9860 4915 9865 4935
rect 9865 4915 9885 4935
rect 9885 4915 9890 4935
rect 9860 4910 9890 4915
rect 9860 4835 9890 4840
rect 9860 4815 9865 4835
rect 9865 4815 9885 4835
rect 9885 4815 9890 4835
rect 9860 4810 9890 4815
rect 9860 4735 9890 4740
rect 9860 4715 9865 4735
rect 9865 4715 9885 4735
rect 9885 4715 9890 4735
rect 9860 4710 9890 4715
rect 9860 4635 9890 4640
rect 9860 4615 9865 4635
rect 9865 4615 9885 4635
rect 9885 4615 9890 4635
rect 9860 4610 9890 4615
rect 9710 4535 9740 4540
rect 9710 4515 9715 4535
rect 9715 4515 9735 4535
rect 9735 4515 9740 4535
rect 9710 4510 9740 4515
rect 9560 4435 9590 4440
rect 9560 4415 9565 4435
rect 9565 4415 9585 4435
rect 9585 4415 9590 4435
rect 9560 4410 9590 4415
rect 9560 4335 9590 4340
rect 9560 4315 9565 4335
rect 9565 4315 9585 4335
rect 9585 4315 9590 4335
rect 9560 4310 9590 4315
rect 9560 4235 9590 4240
rect 9560 4215 9565 4235
rect 9565 4215 9585 4235
rect 9585 4215 9590 4235
rect 9560 4210 9590 4215
rect 9560 4135 9590 4140
rect 9560 4115 9565 4135
rect 9565 4115 9585 4135
rect 9585 4115 9590 4135
rect 9560 4110 9590 4115
rect 9560 4035 9590 4040
rect 9560 4015 9565 4035
rect 9565 4015 9585 4035
rect 9585 4015 9590 4035
rect 9560 4010 9590 4015
rect 9260 3885 9290 3890
rect 9260 3865 9265 3885
rect 9265 3865 9285 3885
rect 9285 3865 9290 3885
rect 9260 3860 9290 3865
rect 8960 3735 8990 3740
rect 8960 3715 8965 3735
rect 8965 3715 8985 3735
rect 8985 3715 8990 3735
rect 8960 3710 8990 3715
rect 8960 3635 8990 3640
rect 8960 3615 8965 3635
rect 8965 3615 8985 3635
rect 8985 3615 8990 3635
rect 8960 3610 8990 3615
rect 8960 3535 8990 3540
rect 8960 3515 8965 3535
rect 8965 3515 8985 3535
rect 8985 3515 8990 3535
rect 8960 3510 8990 3515
rect 8960 3435 8990 3440
rect 8960 3415 8965 3435
rect 8965 3415 8985 3435
rect 8985 3415 8990 3435
rect 8960 3410 8990 3415
rect 8960 3335 8990 3340
rect 8960 3315 8965 3335
rect 8965 3315 8985 3335
rect 8985 3315 8990 3335
rect 8960 3310 8990 3315
rect 8810 3235 8840 3240
rect 8810 3215 8815 3235
rect 8815 3215 8835 3235
rect 8835 3215 8840 3235
rect 8810 3210 8840 3215
rect 8660 3135 8690 3140
rect 8660 3115 8665 3135
rect 8665 3115 8685 3135
rect 8685 3115 8690 3135
rect 8660 3110 8690 3115
rect 8660 3035 8690 3040
rect 8660 3015 8665 3035
rect 8665 3015 8685 3035
rect 8685 3015 8690 3035
rect 8660 3010 8690 3015
rect 8660 2935 8690 2940
rect 8660 2915 8665 2935
rect 8665 2915 8685 2935
rect 8685 2915 8690 2935
rect 8660 2910 8690 2915
rect 8660 2835 8690 2840
rect 8660 2815 8665 2835
rect 8665 2815 8685 2835
rect 8685 2815 8690 2835
rect 8660 2810 8690 2815
rect 8660 2735 8690 2740
rect 8660 2715 8665 2735
rect 8665 2715 8685 2735
rect 8685 2715 8690 2735
rect 8660 2710 8690 2715
rect 8360 2585 8390 2590
rect 8360 2565 8365 2585
rect 8365 2565 8385 2585
rect 8385 2565 8390 2585
rect 8360 2560 8390 2565
rect 10460 5185 10490 5190
rect 10460 5165 10465 5185
rect 10465 5165 10485 5185
rect 10485 5165 10490 5185
rect 10460 5160 10490 5165
rect 10160 5035 10190 5040
rect 10160 5015 10165 5035
rect 10165 5015 10185 5035
rect 10185 5015 10190 5035
rect 10160 5010 10190 5015
rect 10160 4935 10190 4940
rect 10160 4915 10165 4935
rect 10165 4915 10185 4935
rect 10185 4915 10190 4935
rect 10160 4910 10190 4915
rect 10160 4835 10190 4840
rect 10160 4815 10165 4835
rect 10165 4815 10185 4835
rect 10185 4815 10190 4835
rect 10160 4810 10190 4815
rect 10160 4735 10190 4740
rect 10160 4715 10165 4735
rect 10165 4715 10185 4735
rect 10185 4715 10190 4735
rect 10160 4710 10190 4715
rect 10160 4635 10190 4640
rect 10160 4615 10165 4635
rect 10165 4615 10185 4635
rect 10185 4615 10190 4635
rect 10160 4610 10190 4615
rect 10010 4535 10040 4540
rect 10010 4515 10015 4535
rect 10015 4515 10035 4535
rect 10035 4515 10040 4535
rect 10010 4510 10040 4515
rect 9860 4435 9890 4440
rect 9860 4415 9865 4435
rect 9865 4415 9885 4435
rect 9885 4415 9890 4435
rect 9860 4410 9890 4415
rect 9860 4335 9890 4340
rect 9860 4315 9865 4335
rect 9865 4315 9885 4335
rect 9885 4315 9890 4335
rect 9860 4310 9890 4315
rect 9860 4235 9890 4240
rect 9860 4215 9865 4235
rect 9865 4215 9885 4235
rect 9885 4215 9890 4235
rect 9860 4210 9890 4215
rect 9860 4135 9890 4140
rect 9860 4115 9865 4135
rect 9865 4115 9885 4135
rect 9885 4115 9890 4135
rect 9860 4110 9890 4115
rect 9860 4035 9890 4040
rect 9860 4015 9865 4035
rect 9865 4015 9885 4035
rect 9885 4015 9890 4035
rect 9860 4010 9890 4015
rect 9560 3885 9590 3890
rect 9560 3865 9565 3885
rect 9565 3865 9585 3885
rect 9585 3865 9590 3885
rect 9560 3860 9590 3865
rect 9260 3735 9290 3740
rect 9260 3715 9265 3735
rect 9265 3715 9285 3735
rect 9285 3715 9290 3735
rect 9260 3710 9290 3715
rect 9260 3635 9290 3640
rect 9260 3615 9265 3635
rect 9265 3615 9285 3635
rect 9285 3615 9290 3635
rect 9260 3610 9290 3615
rect 9260 3535 9290 3540
rect 9260 3515 9265 3535
rect 9265 3515 9285 3535
rect 9285 3515 9290 3535
rect 9260 3510 9290 3515
rect 9260 3435 9290 3440
rect 9260 3415 9265 3435
rect 9265 3415 9285 3435
rect 9285 3415 9290 3435
rect 9260 3410 9290 3415
rect 9260 3335 9290 3340
rect 9260 3315 9265 3335
rect 9265 3315 9285 3335
rect 9285 3315 9290 3335
rect 9260 3310 9290 3315
rect 9110 3235 9140 3240
rect 9110 3215 9115 3235
rect 9115 3215 9135 3235
rect 9135 3215 9140 3235
rect 9110 3210 9140 3215
rect 8960 3135 8990 3140
rect 8960 3115 8965 3135
rect 8965 3115 8985 3135
rect 8985 3115 8990 3135
rect 8960 3110 8990 3115
rect 8960 3035 8990 3040
rect 8960 3015 8965 3035
rect 8965 3015 8985 3035
rect 8985 3015 8990 3035
rect 8960 3010 8990 3015
rect 8960 2935 8990 2940
rect 8960 2915 8965 2935
rect 8965 2915 8985 2935
rect 8985 2915 8990 2935
rect 8960 2910 8990 2915
rect 8960 2835 8990 2840
rect 8960 2815 8965 2835
rect 8965 2815 8985 2835
rect 8985 2815 8990 2835
rect 8960 2810 8990 2815
rect 8960 2735 8990 2740
rect 8960 2715 8965 2735
rect 8965 2715 8985 2735
rect 8985 2715 8990 2735
rect 8960 2710 8990 2715
rect 8660 2585 8690 2590
rect 8660 2565 8665 2585
rect 8665 2565 8685 2585
rect 8685 2565 8690 2585
rect 8660 2560 8690 2565
rect 10760 5185 10790 5190
rect 10760 5165 10765 5185
rect 10765 5165 10785 5185
rect 10785 5165 10790 5185
rect 10760 5160 10790 5165
rect 10460 5035 10490 5040
rect 10460 5015 10465 5035
rect 10465 5015 10485 5035
rect 10485 5015 10490 5035
rect 10460 5010 10490 5015
rect 10460 4935 10490 4940
rect 10460 4915 10465 4935
rect 10465 4915 10485 4935
rect 10485 4915 10490 4935
rect 10460 4910 10490 4915
rect 10460 4835 10490 4840
rect 10460 4815 10465 4835
rect 10465 4815 10485 4835
rect 10485 4815 10490 4835
rect 10460 4810 10490 4815
rect 10460 4735 10490 4740
rect 10460 4715 10465 4735
rect 10465 4715 10485 4735
rect 10485 4715 10490 4735
rect 10460 4710 10490 4715
rect 10460 4635 10490 4640
rect 10460 4615 10465 4635
rect 10465 4615 10485 4635
rect 10485 4615 10490 4635
rect 10460 4610 10490 4615
rect 10310 4535 10340 4540
rect 10310 4515 10315 4535
rect 10315 4515 10335 4535
rect 10335 4515 10340 4535
rect 10310 4510 10340 4515
rect 10160 4435 10190 4440
rect 10160 4415 10165 4435
rect 10165 4415 10185 4435
rect 10185 4415 10190 4435
rect 10160 4410 10190 4415
rect 10160 4335 10190 4340
rect 10160 4315 10165 4335
rect 10165 4315 10185 4335
rect 10185 4315 10190 4335
rect 10160 4310 10190 4315
rect 10160 4235 10190 4240
rect 10160 4215 10165 4235
rect 10165 4215 10185 4235
rect 10185 4215 10190 4235
rect 10160 4210 10190 4215
rect 10160 4135 10190 4140
rect 10160 4115 10165 4135
rect 10165 4115 10185 4135
rect 10185 4115 10190 4135
rect 10160 4110 10190 4115
rect 10160 4035 10190 4040
rect 10160 4015 10165 4035
rect 10165 4015 10185 4035
rect 10185 4015 10190 4035
rect 10160 4010 10190 4015
rect 9860 3885 9890 3890
rect 9860 3865 9865 3885
rect 9865 3865 9885 3885
rect 9885 3865 9890 3885
rect 9860 3860 9890 3865
rect 9560 3735 9590 3740
rect 9560 3715 9565 3735
rect 9565 3715 9585 3735
rect 9585 3715 9590 3735
rect 9560 3710 9590 3715
rect 9560 3635 9590 3640
rect 9560 3615 9565 3635
rect 9565 3615 9585 3635
rect 9585 3615 9590 3635
rect 9560 3610 9590 3615
rect 9560 3535 9590 3540
rect 9560 3515 9565 3535
rect 9565 3515 9585 3535
rect 9585 3515 9590 3535
rect 9560 3510 9590 3515
rect 9560 3435 9590 3440
rect 9560 3415 9565 3435
rect 9565 3415 9585 3435
rect 9585 3415 9590 3435
rect 9560 3410 9590 3415
rect 9560 3335 9590 3340
rect 9560 3315 9565 3335
rect 9565 3315 9585 3335
rect 9585 3315 9590 3335
rect 9560 3310 9590 3315
rect 9410 3235 9440 3240
rect 9410 3215 9415 3235
rect 9415 3215 9435 3235
rect 9435 3215 9440 3235
rect 9410 3210 9440 3215
rect 9260 3135 9290 3140
rect 9260 3115 9265 3135
rect 9265 3115 9285 3135
rect 9285 3115 9290 3135
rect 9260 3110 9290 3115
rect 9260 3035 9290 3040
rect 9260 3015 9265 3035
rect 9265 3015 9285 3035
rect 9285 3015 9290 3035
rect 9260 3010 9290 3015
rect 9260 2935 9290 2940
rect 9260 2915 9265 2935
rect 9265 2915 9285 2935
rect 9285 2915 9290 2935
rect 9260 2910 9290 2915
rect 9260 2835 9290 2840
rect 9260 2815 9265 2835
rect 9265 2815 9285 2835
rect 9285 2815 9290 2835
rect 9260 2810 9290 2815
rect 9260 2735 9290 2740
rect 9260 2715 9265 2735
rect 9265 2715 9285 2735
rect 9285 2715 9290 2735
rect 9260 2710 9290 2715
rect 8960 2585 8990 2590
rect 8960 2565 8965 2585
rect 8965 2565 8985 2585
rect 8985 2565 8990 2585
rect 8960 2560 8990 2565
rect 11960 5185 11990 5190
rect 11960 5165 11965 5185
rect 11965 5165 11985 5185
rect 11985 5165 11990 5185
rect 11960 5160 11990 5165
rect 10760 5035 10790 5040
rect 10760 5015 10765 5035
rect 10765 5015 10785 5035
rect 10785 5015 10790 5035
rect 10760 5010 10790 5015
rect 10760 4935 10790 4940
rect 10760 4915 10765 4935
rect 10765 4915 10785 4935
rect 10785 4915 10790 4935
rect 10760 4910 10790 4915
rect 10760 4835 10790 4840
rect 10760 4815 10765 4835
rect 10765 4815 10785 4835
rect 10785 4815 10790 4835
rect 10760 4810 10790 4815
rect 10760 4735 10790 4740
rect 10760 4715 10765 4735
rect 10765 4715 10785 4735
rect 10785 4715 10790 4735
rect 10760 4710 10790 4715
rect 10760 4635 10790 4640
rect 10760 4615 10765 4635
rect 10765 4615 10785 4635
rect 10785 4615 10790 4635
rect 10760 4610 10790 4615
rect 10610 4535 10640 4540
rect 10610 4515 10615 4535
rect 10615 4515 10635 4535
rect 10635 4515 10640 4535
rect 10610 4510 10640 4515
rect 10460 4435 10490 4440
rect 10460 4415 10465 4435
rect 10465 4415 10485 4435
rect 10485 4415 10490 4435
rect 10460 4410 10490 4415
rect 10460 4335 10490 4340
rect 10460 4315 10465 4335
rect 10465 4315 10485 4335
rect 10485 4315 10490 4335
rect 10460 4310 10490 4315
rect 10460 4235 10490 4240
rect 10460 4215 10465 4235
rect 10465 4215 10485 4235
rect 10485 4215 10490 4235
rect 10460 4210 10490 4215
rect 10460 4135 10490 4140
rect 10460 4115 10465 4135
rect 10465 4115 10485 4135
rect 10485 4115 10490 4135
rect 10460 4110 10490 4115
rect 10460 4035 10490 4040
rect 10460 4015 10465 4035
rect 10465 4015 10485 4035
rect 10485 4015 10490 4035
rect 10460 4010 10490 4015
rect 10160 3885 10190 3890
rect 10160 3865 10165 3885
rect 10165 3865 10185 3885
rect 10185 3865 10190 3885
rect 10160 3860 10190 3865
rect 9860 3735 9890 3740
rect 9860 3715 9865 3735
rect 9865 3715 9885 3735
rect 9885 3715 9890 3735
rect 9860 3710 9890 3715
rect 9860 3635 9890 3640
rect 9860 3615 9865 3635
rect 9865 3615 9885 3635
rect 9885 3615 9890 3635
rect 9860 3610 9890 3615
rect 9860 3535 9890 3540
rect 9860 3515 9865 3535
rect 9865 3515 9885 3535
rect 9885 3515 9890 3535
rect 9860 3510 9890 3515
rect 9860 3435 9890 3440
rect 9860 3415 9865 3435
rect 9865 3415 9885 3435
rect 9885 3415 9890 3435
rect 9860 3410 9890 3415
rect 9860 3335 9890 3340
rect 9860 3315 9865 3335
rect 9865 3315 9885 3335
rect 9885 3315 9890 3335
rect 9860 3310 9890 3315
rect 9710 3235 9740 3240
rect 9710 3215 9715 3235
rect 9715 3215 9735 3235
rect 9735 3215 9740 3235
rect 9710 3210 9740 3215
rect 9560 3135 9590 3140
rect 9560 3115 9565 3135
rect 9565 3115 9585 3135
rect 9585 3115 9590 3135
rect 9560 3110 9590 3115
rect 9560 3035 9590 3040
rect 9560 3015 9565 3035
rect 9565 3015 9585 3035
rect 9585 3015 9590 3035
rect 9560 3010 9590 3015
rect 9560 2935 9590 2940
rect 9560 2915 9565 2935
rect 9565 2915 9585 2935
rect 9585 2915 9590 2935
rect 9560 2910 9590 2915
rect 9560 2835 9590 2840
rect 9560 2815 9565 2835
rect 9565 2815 9585 2835
rect 9585 2815 9590 2835
rect 9560 2810 9590 2815
rect 9560 2735 9590 2740
rect 9560 2715 9565 2735
rect 9565 2715 9585 2735
rect 9585 2715 9590 2735
rect 9560 2710 9590 2715
rect 9260 2585 9290 2590
rect 9260 2565 9265 2585
rect 9265 2565 9285 2585
rect 9285 2565 9290 2585
rect 9260 2560 9290 2565
rect 10910 4535 10940 4540
rect 10910 4515 10915 4535
rect 10915 4515 10935 4535
rect 10935 4515 10940 4535
rect 10910 4510 10940 4515
rect 11210 4535 11240 4540
rect 11210 4515 11215 4535
rect 11215 4515 11235 4535
rect 11235 4515 11240 4535
rect 11210 4510 11240 4515
rect 13160 5185 13190 5190
rect 13160 5165 13165 5185
rect 13165 5165 13185 5185
rect 13185 5165 13190 5185
rect 13160 5160 13190 5165
rect 11960 5035 11990 5040
rect 11960 5015 11965 5035
rect 11965 5015 11985 5035
rect 11985 5015 11990 5035
rect 11960 5010 11990 5015
rect 11960 4935 11990 4940
rect 11960 4915 11965 4935
rect 11965 4915 11985 4935
rect 11985 4915 11990 4935
rect 11960 4910 11990 4915
rect 11960 4835 11990 4840
rect 11960 4815 11965 4835
rect 11965 4815 11985 4835
rect 11985 4815 11990 4835
rect 11960 4810 11990 4815
rect 11960 4735 11990 4740
rect 11960 4715 11965 4735
rect 11965 4715 11985 4735
rect 11985 4715 11990 4735
rect 11960 4710 11990 4715
rect 11960 4635 11990 4640
rect 11960 4615 11965 4635
rect 11965 4615 11985 4635
rect 11985 4615 11990 4635
rect 11960 4610 11990 4615
rect 11360 4510 11390 4540
rect 10760 4435 10790 4440
rect 10760 4415 10765 4435
rect 10765 4415 10785 4435
rect 10785 4415 10790 4435
rect 10760 4410 10790 4415
rect 10760 4335 10790 4340
rect 10760 4315 10765 4335
rect 10765 4315 10785 4335
rect 10785 4315 10790 4335
rect 10760 4310 10790 4315
rect 10760 4235 10790 4240
rect 10760 4215 10765 4235
rect 10765 4215 10785 4235
rect 10785 4215 10790 4235
rect 10760 4210 10790 4215
rect 10760 4135 10790 4140
rect 10760 4115 10765 4135
rect 10765 4115 10785 4135
rect 10785 4115 10790 4135
rect 10760 4110 10790 4115
rect 10760 4035 10790 4040
rect 10760 4015 10765 4035
rect 10765 4015 10785 4035
rect 10785 4015 10790 4035
rect 10760 4010 10790 4015
rect 10460 3885 10490 3890
rect 10460 3865 10465 3885
rect 10465 3865 10485 3885
rect 10485 3865 10490 3885
rect 10460 3860 10490 3865
rect 10160 3735 10190 3740
rect 10160 3715 10165 3735
rect 10165 3715 10185 3735
rect 10185 3715 10190 3735
rect 10160 3710 10190 3715
rect 10160 3635 10190 3640
rect 10160 3615 10165 3635
rect 10165 3615 10185 3635
rect 10185 3615 10190 3635
rect 10160 3610 10190 3615
rect 10160 3535 10190 3540
rect 10160 3515 10165 3535
rect 10165 3515 10185 3535
rect 10185 3515 10190 3535
rect 10160 3510 10190 3515
rect 10160 3435 10190 3440
rect 10160 3415 10165 3435
rect 10165 3415 10185 3435
rect 10185 3415 10190 3435
rect 10160 3410 10190 3415
rect 10160 3335 10190 3340
rect 10160 3315 10165 3335
rect 10165 3315 10185 3335
rect 10185 3315 10190 3335
rect 10160 3310 10190 3315
rect 10010 3235 10040 3240
rect 10010 3215 10015 3235
rect 10015 3215 10035 3235
rect 10035 3215 10040 3235
rect 10010 3210 10040 3215
rect 9860 3135 9890 3140
rect 9860 3115 9865 3135
rect 9865 3115 9885 3135
rect 9885 3115 9890 3135
rect 9860 3110 9890 3115
rect 9860 3035 9890 3040
rect 9860 3015 9865 3035
rect 9865 3015 9885 3035
rect 9885 3015 9890 3035
rect 9860 3010 9890 3015
rect 9860 2935 9890 2940
rect 9860 2915 9865 2935
rect 9865 2915 9885 2935
rect 9885 2915 9890 2935
rect 9860 2910 9890 2915
rect 9860 2835 9890 2840
rect 9860 2815 9865 2835
rect 9865 2815 9885 2835
rect 9885 2815 9890 2835
rect 9860 2810 9890 2815
rect 9860 2735 9890 2740
rect 9860 2715 9865 2735
rect 9865 2715 9885 2735
rect 9885 2715 9890 2735
rect 9860 2710 9890 2715
rect 9560 2585 9590 2590
rect 9560 2565 9565 2585
rect 9565 2565 9585 2585
rect 9585 2565 9590 2585
rect 9560 2560 9590 2565
rect 10760 3885 10790 3890
rect 10760 3865 10765 3885
rect 10765 3865 10785 3885
rect 10785 3865 10790 3885
rect 10760 3860 10790 3865
rect 10460 3735 10490 3740
rect 10460 3715 10465 3735
rect 10465 3715 10485 3735
rect 10485 3715 10490 3735
rect 10460 3710 10490 3715
rect 10460 3635 10490 3640
rect 10460 3615 10465 3635
rect 10465 3615 10485 3635
rect 10485 3615 10490 3635
rect 10460 3610 10490 3615
rect 10460 3535 10490 3540
rect 10460 3515 10465 3535
rect 10465 3515 10485 3535
rect 10485 3515 10490 3535
rect 10460 3510 10490 3515
rect 10460 3435 10490 3440
rect 10460 3415 10465 3435
rect 10465 3415 10485 3435
rect 10485 3415 10490 3435
rect 10460 3410 10490 3415
rect 10460 3335 10490 3340
rect 10460 3315 10465 3335
rect 10465 3315 10485 3335
rect 10485 3315 10490 3335
rect 10460 3310 10490 3315
rect 10310 3235 10340 3240
rect 10310 3215 10315 3235
rect 10315 3215 10335 3235
rect 10335 3215 10340 3235
rect 10310 3210 10340 3215
rect 10160 3135 10190 3140
rect 10160 3115 10165 3135
rect 10165 3115 10185 3135
rect 10185 3115 10190 3135
rect 10160 3110 10190 3115
rect 10160 3035 10190 3040
rect 10160 3015 10165 3035
rect 10165 3015 10185 3035
rect 10185 3015 10190 3035
rect 10160 3010 10190 3015
rect 10160 2935 10190 2940
rect 10160 2915 10165 2935
rect 10165 2915 10185 2935
rect 10185 2915 10190 2935
rect 10160 2910 10190 2915
rect 10160 2835 10190 2840
rect 10160 2815 10165 2835
rect 10165 2815 10185 2835
rect 10185 2815 10190 2835
rect 10160 2810 10190 2815
rect 10160 2735 10190 2740
rect 10160 2715 10165 2735
rect 10165 2715 10185 2735
rect 10185 2715 10190 2735
rect 10160 2710 10190 2715
rect 9860 2585 9890 2590
rect 9860 2565 9865 2585
rect 9865 2565 9885 2585
rect 9885 2565 9890 2585
rect 9860 2560 9890 2565
rect 10760 3735 10790 3740
rect 10760 3715 10765 3735
rect 10765 3715 10785 3735
rect 10785 3715 10790 3735
rect 10760 3710 10790 3715
rect 10760 3635 10790 3640
rect 10760 3615 10765 3635
rect 10765 3615 10785 3635
rect 10785 3615 10790 3635
rect 10760 3610 10790 3615
rect 10760 3535 10790 3540
rect 10760 3515 10765 3535
rect 10765 3515 10785 3535
rect 10785 3515 10790 3535
rect 10760 3510 10790 3515
rect 10760 3435 10790 3440
rect 10760 3415 10765 3435
rect 10765 3415 10785 3435
rect 10785 3415 10790 3435
rect 10760 3410 10790 3415
rect 10760 3335 10790 3340
rect 10760 3315 10765 3335
rect 10765 3315 10785 3335
rect 10785 3315 10790 3335
rect 10760 3310 10790 3315
rect 10610 3235 10640 3240
rect 10610 3215 10615 3235
rect 10615 3215 10635 3235
rect 10635 3215 10640 3235
rect 10610 3210 10640 3215
rect 10460 3135 10490 3140
rect 10460 3115 10465 3135
rect 10465 3115 10485 3135
rect 10485 3115 10490 3135
rect 10460 3110 10490 3115
rect 10460 3035 10490 3040
rect 10460 3015 10465 3035
rect 10465 3015 10485 3035
rect 10485 3015 10490 3035
rect 10460 3010 10490 3015
rect 10460 2935 10490 2940
rect 10460 2915 10465 2935
rect 10465 2915 10485 2935
rect 10485 2915 10490 2935
rect 10460 2910 10490 2915
rect 10460 2835 10490 2840
rect 10460 2815 10465 2835
rect 10465 2815 10485 2835
rect 10485 2815 10490 2835
rect 10460 2810 10490 2815
rect 10460 2735 10490 2740
rect 10460 2715 10465 2735
rect 10465 2715 10485 2735
rect 10485 2715 10490 2735
rect 10460 2710 10490 2715
rect 10160 2585 10190 2590
rect 10160 2565 10165 2585
rect 10165 2565 10185 2585
rect 10185 2565 10190 2585
rect 10160 2560 10190 2565
rect 11510 4535 11540 4540
rect 11510 4515 11515 4535
rect 11515 4515 11535 4535
rect 11535 4515 11540 4535
rect 11510 4510 11540 4515
rect 11810 4535 11840 4540
rect 11810 4515 11815 4535
rect 11815 4515 11835 4535
rect 11835 4515 11840 4535
rect 11810 4510 11840 4515
rect 10910 3235 10940 3240
rect 10910 3215 10915 3235
rect 10915 3215 10935 3235
rect 10935 3215 10940 3235
rect 10910 3210 10940 3215
rect 11210 3235 11240 3240
rect 11210 3215 11215 3235
rect 11215 3215 11235 3235
rect 11235 3215 11240 3235
rect 11210 3210 11240 3215
rect 12110 4535 12140 4540
rect 12110 4515 12115 4535
rect 12115 4515 12135 4535
rect 12135 4515 12140 4535
rect 12110 4510 12140 4515
rect 12410 4535 12440 4540
rect 12410 4515 12415 4535
rect 12415 4515 12435 4535
rect 12435 4515 12440 4535
rect 12410 4510 12440 4515
rect 14360 5185 14390 5190
rect 14360 5165 14365 5185
rect 14365 5165 14385 5185
rect 14385 5165 14390 5185
rect 14360 5160 14390 5165
rect 13160 5035 13190 5040
rect 13160 5015 13165 5035
rect 13165 5015 13185 5035
rect 13185 5015 13190 5035
rect 13160 5010 13190 5015
rect 13160 4935 13190 4940
rect 13160 4915 13165 4935
rect 13165 4915 13185 4935
rect 13185 4915 13190 4935
rect 13160 4910 13190 4915
rect 13160 4835 13190 4840
rect 13160 4815 13165 4835
rect 13165 4815 13185 4835
rect 13185 4815 13190 4835
rect 13160 4810 13190 4815
rect 13160 4735 13190 4740
rect 13160 4715 13165 4735
rect 13165 4715 13185 4735
rect 13185 4715 13190 4735
rect 13160 4710 13190 4715
rect 13160 4635 13190 4640
rect 13160 4615 13165 4635
rect 13165 4615 13185 4635
rect 13185 4615 13190 4635
rect 13160 4610 13190 4615
rect 12560 4510 12590 4540
rect 11960 4435 11990 4440
rect 11960 4415 11965 4435
rect 11965 4415 11985 4435
rect 11985 4415 11990 4435
rect 11960 4410 11990 4415
rect 11960 4335 11990 4340
rect 11960 4315 11965 4335
rect 11965 4315 11985 4335
rect 11985 4315 11990 4335
rect 11960 4310 11990 4315
rect 11960 4235 11990 4240
rect 11960 4215 11965 4235
rect 11965 4215 11985 4235
rect 11985 4215 11990 4235
rect 11960 4210 11990 4215
rect 11960 4135 11990 4140
rect 11960 4115 11965 4135
rect 11965 4115 11985 4135
rect 11985 4115 11990 4135
rect 11960 4110 11990 4115
rect 11960 4035 11990 4040
rect 11960 4015 11965 4035
rect 11965 4015 11985 4035
rect 11985 4015 11990 4035
rect 11960 4010 11990 4015
rect 11960 3885 11990 3890
rect 11960 3865 11965 3885
rect 11965 3865 11985 3885
rect 11985 3865 11990 3885
rect 11960 3860 11990 3865
rect 11960 3735 11990 3740
rect 11960 3715 11965 3735
rect 11965 3715 11985 3735
rect 11985 3715 11990 3735
rect 11960 3710 11990 3715
rect 11960 3635 11990 3640
rect 11960 3615 11965 3635
rect 11965 3615 11985 3635
rect 11985 3615 11990 3635
rect 11960 3610 11990 3615
rect 11960 3535 11990 3540
rect 11960 3515 11965 3535
rect 11965 3515 11985 3535
rect 11985 3515 11990 3535
rect 11960 3510 11990 3515
rect 11960 3435 11990 3440
rect 11960 3415 11965 3435
rect 11965 3415 11985 3435
rect 11985 3415 11990 3435
rect 11960 3410 11990 3415
rect 11960 3335 11990 3340
rect 11960 3315 11965 3335
rect 11965 3315 11985 3335
rect 11985 3315 11990 3335
rect 11960 3310 11990 3315
rect 11360 3210 11390 3240
rect 10760 3135 10790 3140
rect 10760 3115 10765 3135
rect 10765 3115 10785 3135
rect 10785 3115 10790 3135
rect 10760 3110 10790 3115
rect 10760 3035 10790 3040
rect 10760 3015 10765 3035
rect 10765 3015 10785 3035
rect 10785 3015 10790 3035
rect 10760 3010 10790 3015
rect 10760 2935 10790 2940
rect 10760 2915 10765 2935
rect 10765 2915 10785 2935
rect 10785 2915 10790 2935
rect 10760 2910 10790 2915
rect 10760 2835 10790 2840
rect 10760 2815 10765 2835
rect 10765 2815 10785 2835
rect 10785 2815 10790 2835
rect 10760 2810 10790 2815
rect 10760 2735 10790 2740
rect 10760 2715 10765 2735
rect 10765 2715 10785 2735
rect 10785 2715 10790 2735
rect 10760 2710 10790 2715
rect 10460 2585 10490 2590
rect 10460 2565 10465 2585
rect 10465 2565 10485 2585
rect 10485 2565 10490 2585
rect 10460 2560 10490 2565
rect 11510 3235 11540 3240
rect 11510 3215 11515 3235
rect 11515 3215 11535 3235
rect 11535 3215 11540 3235
rect 11510 3210 11540 3215
rect 11810 3235 11840 3240
rect 11810 3215 11815 3235
rect 11815 3215 11835 3235
rect 11835 3215 11840 3235
rect 11810 3210 11840 3215
rect 12710 4535 12740 4540
rect 12710 4515 12715 4535
rect 12715 4515 12735 4535
rect 12735 4515 12740 4535
rect 12710 4510 12740 4515
rect 13010 4535 13040 4540
rect 13010 4515 13015 4535
rect 13015 4515 13035 4535
rect 13035 4515 13040 4535
rect 13010 4510 13040 4515
rect 12110 3235 12140 3240
rect 12110 3215 12115 3235
rect 12115 3215 12135 3235
rect 12135 3215 12140 3235
rect 12110 3210 12140 3215
rect 12410 3235 12440 3240
rect 12410 3215 12415 3235
rect 12415 3215 12435 3235
rect 12435 3215 12440 3235
rect 12410 3210 12440 3215
rect 13310 4535 13340 4540
rect 13310 4515 13315 4535
rect 13315 4515 13335 4535
rect 13335 4515 13340 4535
rect 13310 4510 13340 4515
rect 13610 4535 13640 4540
rect 13610 4515 13615 4535
rect 13615 4515 13635 4535
rect 13635 4515 13640 4535
rect 13610 4510 13640 4515
rect 15560 5185 15590 5190
rect 15560 5165 15565 5185
rect 15565 5165 15585 5185
rect 15585 5165 15590 5185
rect 15560 5160 15590 5165
rect 14360 5035 14390 5040
rect 14360 5015 14365 5035
rect 14365 5015 14385 5035
rect 14385 5015 14390 5035
rect 14360 5010 14390 5015
rect 14360 4935 14390 4940
rect 14360 4915 14365 4935
rect 14365 4915 14385 4935
rect 14385 4915 14390 4935
rect 14360 4910 14390 4915
rect 14360 4835 14390 4840
rect 14360 4815 14365 4835
rect 14365 4815 14385 4835
rect 14385 4815 14390 4835
rect 14360 4810 14390 4815
rect 14360 4735 14390 4740
rect 14360 4715 14365 4735
rect 14365 4715 14385 4735
rect 14385 4715 14390 4735
rect 14360 4710 14390 4715
rect 14360 4635 14390 4640
rect 14360 4615 14365 4635
rect 14365 4615 14385 4635
rect 14385 4615 14390 4635
rect 14360 4610 14390 4615
rect 13760 4510 13790 4540
rect 13160 4435 13190 4440
rect 13160 4415 13165 4435
rect 13165 4415 13185 4435
rect 13185 4415 13190 4435
rect 13160 4410 13190 4415
rect 13160 4335 13190 4340
rect 13160 4315 13165 4335
rect 13165 4315 13185 4335
rect 13185 4315 13190 4335
rect 13160 4310 13190 4315
rect 13160 4235 13190 4240
rect 13160 4215 13165 4235
rect 13165 4215 13185 4235
rect 13185 4215 13190 4235
rect 13160 4210 13190 4215
rect 13160 4135 13190 4140
rect 13160 4115 13165 4135
rect 13165 4115 13185 4135
rect 13185 4115 13190 4135
rect 13160 4110 13190 4115
rect 13160 4035 13190 4040
rect 13160 4015 13165 4035
rect 13165 4015 13185 4035
rect 13185 4015 13190 4035
rect 13160 4010 13190 4015
rect 13160 3885 13190 3890
rect 13160 3865 13165 3885
rect 13165 3865 13185 3885
rect 13185 3865 13190 3885
rect 13160 3860 13190 3865
rect 13160 3735 13190 3740
rect 13160 3715 13165 3735
rect 13165 3715 13185 3735
rect 13185 3715 13190 3735
rect 13160 3710 13190 3715
rect 13160 3635 13190 3640
rect 13160 3615 13165 3635
rect 13165 3615 13185 3635
rect 13185 3615 13190 3635
rect 13160 3610 13190 3615
rect 13160 3535 13190 3540
rect 13160 3515 13165 3535
rect 13165 3515 13185 3535
rect 13185 3515 13190 3535
rect 13160 3510 13190 3515
rect 13160 3435 13190 3440
rect 13160 3415 13165 3435
rect 13165 3415 13185 3435
rect 13185 3415 13190 3435
rect 13160 3410 13190 3415
rect 13160 3335 13190 3340
rect 13160 3315 13165 3335
rect 13165 3315 13185 3335
rect 13185 3315 13190 3335
rect 13160 3310 13190 3315
rect 12560 3210 12590 3240
rect 11960 3135 11990 3140
rect 11960 3115 11965 3135
rect 11965 3115 11985 3135
rect 11985 3115 11990 3135
rect 11960 3110 11990 3115
rect 11960 3035 11990 3040
rect 11960 3015 11965 3035
rect 11965 3015 11985 3035
rect 11985 3015 11990 3035
rect 11960 3010 11990 3015
rect 11960 2935 11990 2940
rect 11960 2915 11965 2935
rect 11965 2915 11985 2935
rect 11985 2915 11990 2935
rect 11960 2910 11990 2915
rect 11960 2835 11990 2840
rect 11960 2815 11965 2835
rect 11965 2815 11985 2835
rect 11985 2815 11990 2835
rect 11960 2810 11990 2815
rect 11960 2735 11990 2740
rect 11960 2715 11965 2735
rect 11965 2715 11985 2735
rect 11985 2715 11990 2735
rect 11960 2710 11990 2715
rect 10760 2585 10790 2590
rect 10760 2565 10765 2585
rect 10765 2565 10785 2585
rect 10785 2565 10790 2585
rect 10760 2560 10790 2565
rect 12710 3235 12740 3240
rect 12710 3215 12715 3235
rect 12715 3215 12735 3235
rect 12735 3215 12740 3235
rect 12710 3210 12740 3215
rect 13010 3235 13040 3240
rect 13010 3215 13015 3235
rect 13015 3215 13035 3235
rect 13035 3215 13040 3235
rect 13010 3210 13040 3215
rect 13910 4535 13940 4540
rect 13910 4515 13915 4535
rect 13915 4515 13935 4535
rect 13935 4515 13940 4535
rect 13910 4510 13940 4515
rect 14210 4535 14240 4540
rect 14210 4515 14215 4535
rect 14215 4515 14235 4535
rect 14235 4515 14240 4535
rect 14210 4510 14240 4515
rect 13310 3235 13340 3240
rect 13310 3215 13315 3235
rect 13315 3215 13335 3235
rect 13335 3215 13340 3235
rect 13310 3210 13340 3215
rect 13610 3235 13640 3240
rect 13610 3215 13615 3235
rect 13615 3215 13635 3235
rect 13635 3215 13640 3235
rect 13610 3210 13640 3215
rect 14510 4535 14540 4540
rect 14510 4515 14515 4535
rect 14515 4515 14535 4535
rect 14535 4515 14540 4535
rect 14510 4510 14540 4515
rect 14810 4535 14840 4540
rect 14810 4515 14815 4535
rect 14815 4515 14835 4535
rect 14835 4515 14840 4535
rect 14810 4510 14840 4515
rect 17960 5185 17990 5190
rect 17960 5165 17965 5185
rect 17965 5165 17985 5185
rect 17985 5165 17990 5185
rect 17960 5160 17990 5165
rect 20360 5185 20390 5190
rect 20360 5165 20365 5185
rect 20365 5165 20385 5185
rect 20385 5165 20390 5185
rect 20360 5160 20390 5165
rect 15560 5035 15590 5040
rect 15560 5015 15565 5035
rect 15565 5015 15585 5035
rect 15585 5015 15590 5035
rect 15560 5010 15590 5015
rect 15560 4935 15590 4940
rect 15560 4915 15565 4935
rect 15565 4915 15585 4935
rect 15585 4915 15590 4935
rect 15560 4910 15590 4915
rect 15560 4835 15590 4840
rect 15560 4815 15565 4835
rect 15565 4815 15585 4835
rect 15585 4815 15590 4835
rect 15560 4810 15590 4815
rect 15560 4735 15590 4740
rect 15560 4715 15565 4735
rect 15565 4715 15585 4735
rect 15585 4715 15590 4735
rect 15560 4710 15590 4715
rect 15560 4635 15590 4640
rect 15560 4615 15565 4635
rect 15565 4615 15585 4635
rect 15585 4615 15590 4635
rect 15560 4610 15590 4615
rect 14960 4510 14990 4540
rect 14360 4435 14390 4440
rect 14360 4415 14365 4435
rect 14365 4415 14385 4435
rect 14385 4415 14390 4435
rect 14360 4410 14390 4415
rect 14360 4335 14390 4340
rect 14360 4315 14365 4335
rect 14365 4315 14385 4335
rect 14385 4315 14390 4335
rect 14360 4310 14390 4315
rect 14360 4235 14390 4240
rect 14360 4215 14365 4235
rect 14365 4215 14385 4235
rect 14385 4215 14390 4235
rect 14360 4210 14390 4215
rect 14360 4135 14390 4140
rect 14360 4115 14365 4135
rect 14365 4115 14385 4135
rect 14385 4115 14390 4135
rect 14360 4110 14390 4115
rect 14360 4035 14390 4040
rect 14360 4015 14365 4035
rect 14365 4015 14385 4035
rect 14385 4015 14390 4035
rect 14360 4010 14390 4015
rect 14360 3885 14390 3890
rect 14360 3865 14365 3885
rect 14365 3865 14385 3885
rect 14385 3865 14390 3885
rect 14360 3860 14390 3865
rect 14360 3735 14390 3740
rect 14360 3715 14365 3735
rect 14365 3715 14385 3735
rect 14385 3715 14390 3735
rect 14360 3710 14390 3715
rect 14360 3635 14390 3640
rect 14360 3615 14365 3635
rect 14365 3615 14385 3635
rect 14385 3615 14390 3635
rect 14360 3610 14390 3615
rect 14360 3535 14390 3540
rect 14360 3515 14365 3535
rect 14365 3515 14385 3535
rect 14385 3515 14390 3535
rect 14360 3510 14390 3515
rect 14360 3435 14390 3440
rect 14360 3415 14365 3435
rect 14365 3415 14385 3435
rect 14385 3415 14390 3435
rect 14360 3410 14390 3415
rect 14360 3335 14390 3340
rect 14360 3315 14365 3335
rect 14365 3315 14385 3335
rect 14385 3315 14390 3335
rect 14360 3310 14390 3315
rect 13760 3210 13790 3240
rect 13160 3135 13190 3140
rect 13160 3115 13165 3135
rect 13165 3115 13185 3135
rect 13185 3115 13190 3135
rect 13160 3110 13190 3115
rect 13160 3035 13190 3040
rect 13160 3015 13165 3035
rect 13165 3015 13185 3035
rect 13185 3015 13190 3035
rect 13160 3010 13190 3015
rect 13160 2935 13190 2940
rect 13160 2915 13165 2935
rect 13165 2915 13185 2935
rect 13185 2915 13190 2935
rect 13160 2910 13190 2915
rect 13160 2835 13190 2840
rect 13160 2815 13165 2835
rect 13165 2815 13185 2835
rect 13185 2815 13190 2835
rect 13160 2810 13190 2815
rect 13160 2735 13190 2740
rect 13160 2715 13165 2735
rect 13165 2715 13185 2735
rect 13185 2715 13190 2735
rect 13160 2710 13190 2715
rect 11960 2585 11990 2590
rect 11960 2565 11965 2585
rect 11965 2565 11985 2585
rect 11985 2565 11990 2585
rect 11960 2560 11990 2565
rect 13910 3235 13940 3240
rect 13910 3215 13915 3235
rect 13915 3215 13935 3235
rect 13935 3215 13940 3235
rect 13910 3210 13940 3215
rect 14210 3235 14240 3240
rect 14210 3215 14215 3235
rect 14215 3215 14235 3235
rect 14235 3215 14240 3235
rect 14210 3210 14240 3215
rect 15110 4535 15140 4540
rect 15110 4515 15115 4535
rect 15115 4515 15135 4535
rect 15135 4515 15140 4535
rect 15110 4510 15140 4515
rect 15410 4535 15440 4540
rect 15410 4515 15415 4535
rect 15415 4515 15435 4535
rect 15435 4515 15440 4535
rect 15410 4510 15440 4515
rect 14510 3235 14540 3240
rect 14510 3215 14515 3235
rect 14515 3215 14535 3235
rect 14535 3215 14540 3235
rect 14510 3210 14540 3215
rect 14810 3235 14840 3240
rect 14810 3215 14815 3235
rect 14815 3215 14835 3235
rect 14835 3215 14840 3235
rect 14810 3210 14840 3215
rect 15710 4535 15740 4540
rect 15710 4515 15715 4535
rect 15715 4515 15735 4535
rect 15735 4515 15740 4535
rect 15710 4510 15740 4515
rect 16010 4535 16040 4540
rect 16010 4515 16015 4535
rect 16015 4515 16035 4535
rect 16035 4515 16040 4535
rect 16010 4510 16040 4515
rect 15560 4435 15590 4440
rect 15560 4415 15565 4435
rect 15565 4415 15585 4435
rect 15585 4415 15590 4435
rect 15560 4410 15590 4415
rect 15560 4335 15590 4340
rect 15560 4315 15565 4335
rect 15565 4315 15585 4335
rect 15585 4315 15590 4335
rect 15560 4310 15590 4315
rect 15560 4235 15590 4240
rect 15560 4215 15565 4235
rect 15565 4215 15585 4235
rect 15585 4215 15590 4235
rect 15560 4210 15590 4215
rect 15560 4135 15590 4140
rect 15560 4115 15565 4135
rect 15565 4115 15585 4135
rect 15585 4115 15590 4135
rect 15560 4110 15590 4115
rect 15560 4035 15590 4040
rect 15560 4015 15565 4035
rect 15565 4015 15585 4035
rect 15585 4015 15590 4035
rect 15560 4010 15590 4015
rect 16310 4535 16340 4540
rect 16310 4515 16315 4535
rect 16315 4515 16335 4535
rect 16335 4515 16340 4535
rect 16310 4510 16340 4515
rect 16610 4535 16640 4540
rect 16610 4515 16615 4535
rect 16615 4515 16635 4535
rect 16635 4515 16640 4535
rect 16610 4510 16640 4515
rect 16760 4510 16790 4540
rect 16910 4535 16940 4540
rect 16910 4515 16915 4535
rect 16915 4515 16935 4535
rect 16935 4515 16940 4535
rect 16910 4510 16940 4515
rect 17210 4535 17240 4540
rect 17210 4515 17215 4535
rect 17215 4515 17235 4535
rect 17235 4515 17240 4535
rect 17210 4510 17240 4515
rect 17960 4935 17990 4940
rect 17960 4915 17965 4935
rect 17965 4915 17985 4935
rect 17985 4915 17990 4935
rect 17960 4910 17990 4915
rect 17960 4835 17990 4840
rect 17960 4815 17965 4835
rect 17965 4815 17985 4835
rect 17985 4815 17990 4835
rect 17960 4810 17990 4815
rect 17960 4735 17990 4740
rect 17960 4715 17965 4735
rect 17965 4715 17985 4735
rect 17985 4715 17990 4735
rect 17960 4710 17990 4715
rect 17960 4635 17990 4640
rect 17960 4615 17965 4635
rect 17965 4615 17985 4635
rect 17985 4615 17990 4635
rect 17960 4610 17990 4615
rect 17510 4535 17540 4540
rect 17510 4515 17515 4535
rect 17515 4515 17535 4535
rect 17535 4515 17540 4535
rect 17510 4510 17540 4515
rect 17810 4535 17840 4540
rect 17810 4515 17815 4535
rect 17815 4515 17835 4535
rect 17835 4515 17840 4535
rect 17810 4510 17840 4515
rect 18110 4535 18140 4540
rect 18110 4515 18115 4535
rect 18115 4515 18135 4535
rect 18135 4515 18140 4535
rect 18110 4510 18140 4515
rect 18410 4535 18440 4540
rect 18410 4515 18415 4535
rect 18415 4515 18435 4535
rect 18435 4515 18440 4535
rect 18410 4510 18440 4515
rect 17960 4435 17990 4440
rect 17960 4415 17965 4435
rect 17965 4415 17985 4435
rect 17985 4415 17990 4435
rect 17960 4410 17990 4415
rect 17960 4335 17990 4340
rect 17960 4315 17965 4335
rect 17965 4315 17985 4335
rect 17985 4315 17990 4335
rect 17960 4310 17990 4315
rect 17960 4235 17990 4240
rect 17960 4215 17965 4235
rect 17965 4215 17985 4235
rect 17985 4215 17990 4235
rect 17960 4210 17990 4215
rect 17960 4135 17990 4140
rect 17960 4115 17965 4135
rect 17965 4115 17985 4135
rect 17985 4115 17990 4135
rect 17960 4110 17990 4115
rect 18710 4535 18740 4540
rect 18710 4515 18715 4535
rect 18715 4515 18735 4535
rect 18735 4515 18740 4535
rect 18710 4510 18740 4515
rect 19010 4535 19040 4540
rect 19010 4515 19015 4535
rect 19015 4515 19035 4535
rect 19035 4515 19040 4535
rect 19010 4510 19040 4515
rect 19160 4510 19190 4540
rect 19310 4535 19340 4540
rect 19310 4515 19315 4535
rect 19315 4515 19335 4535
rect 19335 4515 19340 4535
rect 19310 4510 19340 4515
rect 19610 4535 19640 4540
rect 19610 4515 19615 4535
rect 19615 4515 19635 4535
rect 19635 4515 19640 4535
rect 19610 4510 19640 4515
rect 20360 5035 20390 5040
rect 20360 5015 20365 5035
rect 20365 5015 20385 5035
rect 20385 5015 20390 5035
rect 20360 5010 20390 5015
rect 20360 4935 20390 4940
rect 20360 4915 20365 4935
rect 20365 4915 20385 4935
rect 20385 4915 20390 4935
rect 20360 4910 20390 4915
rect 20360 4835 20390 4840
rect 20360 4815 20365 4835
rect 20365 4815 20385 4835
rect 20385 4815 20390 4835
rect 20360 4810 20390 4815
rect 20360 4735 20390 4740
rect 20360 4715 20365 4735
rect 20365 4715 20385 4735
rect 20385 4715 20390 4735
rect 20360 4710 20390 4715
rect 20360 4635 20390 4640
rect 20360 4615 20365 4635
rect 20365 4615 20385 4635
rect 20385 4615 20390 4635
rect 20360 4610 20390 4615
rect 19910 4535 19940 4540
rect 19910 4515 19915 4535
rect 19915 4515 19935 4535
rect 19935 4515 19940 4535
rect 19910 4510 19940 4515
rect 20210 4535 20240 4540
rect 20210 4515 20215 4535
rect 20215 4515 20235 4535
rect 20235 4515 20240 4535
rect 20210 4510 20240 4515
rect 20360 4435 20390 4440
rect 20360 4415 20365 4435
rect 20365 4415 20385 4435
rect 20385 4415 20390 4435
rect 20360 4410 20390 4415
rect 20360 4335 20390 4340
rect 20360 4315 20365 4335
rect 20365 4315 20385 4335
rect 20385 4315 20390 4335
rect 20360 4310 20390 4315
rect 20360 4235 20390 4240
rect 20360 4215 20365 4235
rect 20365 4215 20385 4235
rect 20385 4215 20390 4235
rect 20360 4210 20390 4215
rect 20360 4135 20390 4140
rect 20360 4115 20365 4135
rect 20365 4115 20385 4135
rect 20385 4115 20390 4135
rect 20360 4110 20390 4115
rect 20360 4035 20390 4040
rect 20360 4015 20365 4035
rect 20365 4015 20385 4035
rect 20385 4015 20390 4035
rect 20360 4010 20390 4015
rect 15560 3885 15590 3890
rect 15560 3865 15565 3885
rect 15565 3865 15585 3885
rect 15585 3865 15590 3885
rect 15560 3860 15590 3865
rect 20360 3885 20390 3890
rect 20360 3865 20365 3885
rect 20365 3865 20385 3885
rect 20385 3865 20390 3885
rect 20360 3860 20390 3865
rect 15560 3735 15590 3740
rect 15560 3715 15565 3735
rect 15565 3715 15585 3735
rect 15585 3715 15590 3735
rect 15560 3710 15590 3715
rect 15560 3635 15590 3640
rect 15560 3615 15565 3635
rect 15565 3615 15585 3635
rect 15585 3615 15590 3635
rect 15560 3610 15590 3615
rect 15560 3535 15590 3540
rect 15560 3515 15565 3535
rect 15565 3515 15585 3535
rect 15585 3515 15590 3535
rect 15560 3510 15590 3515
rect 15560 3435 15590 3440
rect 15560 3415 15565 3435
rect 15565 3415 15585 3435
rect 15585 3415 15590 3435
rect 15560 3410 15590 3415
rect 15560 3335 15590 3340
rect 15560 3315 15565 3335
rect 15565 3315 15585 3335
rect 15585 3315 15590 3335
rect 15560 3310 15590 3315
rect 14960 3210 14990 3240
rect 14360 3135 14390 3140
rect 14360 3115 14365 3135
rect 14365 3115 14385 3135
rect 14385 3115 14390 3135
rect 14360 3110 14390 3115
rect 14360 3035 14390 3040
rect 14360 3015 14365 3035
rect 14365 3015 14385 3035
rect 14385 3015 14390 3035
rect 14360 3010 14390 3015
rect 14360 2935 14390 2940
rect 14360 2915 14365 2935
rect 14365 2915 14385 2935
rect 14385 2915 14390 2935
rect 14360 2910 14390 2915
rect 14360 2835 14390 2840
rect 14360 2815 14365 2835
rect 14365 2815 14385 2835
rect 14385 2815 14390 2835
rect 14360 2810 14390 2815
rect 14360 2735 14390 2740
rect 14360 2715 14365 2735
rect 14365 2715 14385 2735
rect 14385 2715 14390 2735
rect 14360 2710 14390 2715
rect 13160 2585 13190 2590
rect 13160 2565 13165 2585
rect 13165 2565 13185 2585
rect 13185 2565 13190 2585
rect 13160 2560 13190 2565
rect 15110 3235 15140 3240
rect 15110 3215 15115 3235
rect 15115 3215 15135 3235
rect 15135 3215 15140 3235
rect 15110 3210 15140 3215
rect 15410 3235 15440 3240
rect 15410 3215 15415 3235
rect 15415 3215 15435 3235
rect 15435 3215 15440 3235
rect 15410 3210 15440 3215
rect 15710 3235 15740 3240
rect 15710 3215 15715 3235
rect 15715 3215 15735 3235
rect 15735 3215 15740 3235
rect 15710 3210 15740 3215
rect 16010 3235 16040 3240
rect 16010 3215 16015 3235
rect 16015 3215 16035 3235
rect 16035 3215 16040 3235
rect 16010 3210 16040 3215
rect 15560 3135 15590 3140
rect 15560 3115 15565 3135
rect 15565 3115 15585 3135
rect 15585 3115 15590 3135
rect 15560 3110 15590 3115
rect 15560 3035 15590 3040
rect 15560 3015 15565 3035
rect 15565 3015 15585 3035
rect 15585 3015 15590 3035
rect 15560 3010 15590 3015
rect 15560 2935 15590 2940
rect 15560 2915 15565 2935
rect 15565 2915 15585 2935
rect 15585 2915 15590 2935
rect 15560 2910 15590 2915
rect 15560 2835 15590 2840
rect 15560 2815 15565 2835
rect 15565 2815 15585 2835
rect 15585 2815 15590 2835
rect 15560 2810 15590 2815
rect 15560 2735 15590 2740
rect 15560 2715 15565 2735
rect 15565 2715 15585 2735
rect 15585 2715 15590 2735
rect 15560 2710 15590 2715
rect 14360 2585 14390 2590
rect 14360 2565 14365 2585
rect 14365 2565 14385 2585
rect 14385 2565 14390 2585
rect 14360 2560 14390 2565
rect 16310 3235 16340 3240
rect 16310 3215 16315 3235
rect 16315 3215 16335 3235
rect 16335 3215 16340 3235
rect 16310 3210 16340 3215
rect 16610 3235 16640 3240
rect 16610 3215 16615 3235
rect 16615 3215 16635 3235
rect 16635 3215 16640 3235
rect 16610 3210 16640 3215
rect 16760 3210 16790 3240
rect 16910 3235 16940 3240
rect 16910 3215 16915 3235
rect 16915 3215 16935 3235
rect 16935 3215 16940 3235
rect 16910 3210 16940 3215
rect 17210 3235 17240 3240
rect 17210 3215 17215 3235
rect 17215 3215 17235 3235
rect 17235 3215 17240 3235
rect 17210 3210 17240 3215
rect 17960 3635 17990 3640
rect 17960 3615 17965 3635
rect 17965 3615 17985 3635
rect 17985 3615 17990 3635
rect 17960 3610 17990 3615
rect 17960 3535 17990 3540
rect 17960 3515 17965 3535
rect 17965 3515 17985 3535
rect 17985 3515 17990 3535
rect 17960 3510 17990 3515
rect 17960 3435 17990 3440
rect 17960 3415 17965 3435
rect 17965 3415 17985 3435
rect 17985 3415 17990 3435
rect 17960 3410 17990 3415
rect 17960 3335 17990 3340
rect 17960 3315 17965 3335
rect 17965 3315 17985 3335
rect 17985 3315 17990 3335
rect 17960 3310 17990 3315
rect 17510 3235 17540 3240
rect 17510 3215 17515 3235
rect 17515 3215 17535 3235
rect 17535 3215 17540 3235
rect 17510 3210 17540 3215
rect 17810 3235 17840 3240
rect 17810 3215 17815 3235
rect 17815 3215 17835 3235
rect 17835 3215 17840 3235
rect 17810 3210 17840 3215
rect 18110 3235 18140 3240
rect 18110 3215 18115 3235
rect 18115 3215 18135 3235
rect 18135 3215 18140 3235
rect 18110 3210 18140 3215
rect 18410 3235 18440 3240
rect 18410 3215 18415 3235
rect 18415 3215 18435 3235
rect 18435 3215 18440 3235
rect 18410 3210 18440 3215
rect 17960 3135 17990 3140
rect 17960 3115 17965 3135
rect 17965 3115 17985 3135
rect 17985 3115 17990 3135
rect 17960 3110 17990 3115
rect 17960 3035 17990 3040
rect 17960 3015 17965 3035
rect 17965 3015 17985 3035
rect 17985 3015 17990 3035
rect 17960 3010 17990 3015
rect 17960 2935 17990 2940
rect 17960 2915 17965 2935
rect 17965 2915 17985 2935
rect 17985 2915 17990 2935
rect 17960 2910 17990 2915
rect 17960 2835 17990 2840
rect 17960 2815 17965 2835
rect 17965 2815 17985 2835
rect 17985 2815 17990 2835
rect 17960 2810 17990 2815
rect 18710 3235 18740 3240
rect 18710 3215 18715 3235
rect 18715 3215 18735 3235
rect 18735 3215 18740 3235
rect 18710 3210 18740 3215
rect 19010 3235 19040 3240
rect 19010 3215 19015 3235
rect 19015 3215 19035 3235
rect 19035 3215 19040 3235
rect 19010 3210 19040 3215
rect 19160 3210 19190 3240
rect 19310 3235 19340 3240
rect 19310 3215 19315 3235
rect 19315 3215 19335 3235
rect 19335 3215 19340 3235
rect 19310 3210 19340 3215
rect 19610 3235 19640 3240
rect 19610 3215 19615 3235
rect 19615 3215 19635 3235
rect 19635 3215 19640 3235
rect 19610 3210 19640 3215
rect 20360 3735 20390 3740
rect 20360 3715 20365 3735
rect 20365 3715 20385 3735
rect 20385 3715 20390 3735
rect 20360 3710 20390 3715
rect 20360 3635 20390 3640
rect 20360 3615 20365 3635
rect 20365 3615 20385 3635
rect 20385 3615 20390 3635
rect 20360 3610 20390 3615
rect 20360 3535 20390 3540
rect 20360 3515 20365 3535
rect 20365 3515 20385 3535
rect 20385 3515 20390 3535
rect 20360 3510 20390 3515
rect 20360 3435 20390 3440
rect 20360 3415 20365 3435
rect 20365 3415 20385 3435
rect 20385 3415 20390 3435
rect 20360 3410 20390 3415
rect 20360 3335 20390 3340
rect 20360 3315 20365 3335
rect 20365 3315 20385 3335
rect 20385 3315 20390 3335
rect 20360 3310 20390 3315
rect 19910 3235 19940 3240
rect 19910 3215 19915 3235
rect 19915 3215 19935 3235
rect 19935 3215 19940 3235
rect 19910 3210 19940 3215
rect 20210 3235 20240 3240
rect 20210 3215 20215 3235
rect 20215 3215 20235 3235
rect 20235 3215 20240 3235
rect 20210 3210 20240 3215
rect 20360 3135 20390 3140
rect 20360 3115 20365 3135
rect 20365 3115 20385 3135
rect 20385 3115 20390 3135
rect 20360 3110 20390 3115
rect 20360 3035 20390 3040
rect 20360 3015 20365 3035
rect 20365 3015 20385 3035
rect 20385 3015 20390 3035
rect 20360 3010 20390 3015
rect 20360 2935 20390 2940
rect 20360 2915 20365 2935
rect 20365 2915 20385 2935
rect 20385 2915 20390 2935
rect 20360 2910 20390 2915
rect 20360 2835 20390 2840
rect 20360 2815 20365 2835
rect 20365 2815 20385 2835
rect 20385 2815 20390 2835
rect 20360 2810 20390 2815
rect 20360 2735 20390 2740
rect 20360 2715 20365 2735
rect 20365 2715 20385 2735
rect 20385 2715 20390 2735
rect 20360 2710 20390 2715
rect 15560 2585 15590 2590
rect 15560 2565 15565 2585
rect 15565 2565 15585 2585
rect 15585 2565 15590 2585
rect 15560 2560 15590 2565
rect 17960 2585 17990 2590
rect 17960 2565 17965 2585
rect 17965 2565 17985 2585
rect 17985 2565 17990 2585
rect 17960 2560 17990 2565
rect 20360 2585 20390 2590
rect 20360 2565 20365 2585
rect 20365 2565 20385 2585
rect 20385 2565 20390 2585
rect 20360 2560 20390 2565
rect -640 1685 -610 1690
rect -640 1665 -635 1685
rect -635 1665 -615 1685
rect -615 1665 -610 1685
rect -640 1660 -610 1665
rect -40 1685 -10 1690
rect -40 1665 -35 1685
rect -35 1665 -15 1685
rect -15 1665 -10 1685
rect -40 1660 -10 1665
rect -640 1535 -610 1540
rect -640 1515 -635 1535
rect -635 1515 -615 1535
rect -615 1515 -610 1535
rect -640 1510 -610 1515
rect -640 1435 -610 1440
rect -640 1415 -635 1435
rect -635 1415 -615 1435
rect -615 1415 -610 1435
rect -640 1410 -610 1415
rect -640 1335 -610 1340
rect -640 1315 -635 1335
rect -635 1315 -615 1335
rect -615 1315 -610 1335
rect -640 1310 -610 1315
rect -640 1235 -610 1240
rect -640 1215 -635 1235
rect -635 1215 -615 1235
rect -615 1215 -610 1235
rect -640 1210 -610 1215
rect -640 1135 -610 1140
rect -640 1115 -635 1135
rect -635 1115 -615 1135
rect -615 1115 -610 1135
rect -640 1110 -610 1115
rect -640 1035 -610 1040
rect -640 1015 -635 1035
rect -635 1015 -615 1035
rect -615 1015 -610 1035
rect -640 1010 -610 1015
rect -640 935 -610 940
rect -640 915 -635 935
rect -635 915 -615 935
rect -615 915 -610 935
rect -640 910 -610 915
rect -490 835 -460 840
rect -490 815 -485 835
rect -485 815 -465 835
rect -465 815 -460 835
rect -490 810 -460 815
rect 8360 1685 8390 1690
rect 8360 1665 8365 1685
rect 8365 1665 8385 1685
rect 8385 1665 8390 1685
rect 8360 1660 8390 1665
rect -40 1535 -10 1540
rect -40 1515 -35 1535
rect -35 1515 -15 1535
rect -15 1515 -10 1535
rect -40 1510 -10 1515
rect -40 1435 -10 1440
rect -40 1415 -35 1435
rect -35 1415 -15 1435
rect -15 1415 -10 1435
rect -40 1410 -10 1415
rect -40 1335 -10 1340
rect -40 1315 -35 1335
rect -35 1315 -15 1335
rect -15 1315 -10 1335
rect -40 1310 -10 1315
rect -40 1235 -10 1240
rect -40 1215 -35 1235
rect -35 1215 -15 1235
rect -15 1215 -10 1235
rect -40 1210 -10 1215
rect -40 1135 -10 1140
rect -40 1115 -35 1135
rect -35 1115 -15 1135
rect -15 1115 -10 1135
rect -40 1110 -10 1115
rect -40 1035 -10 1040
rect -40 1015 -35 1035
rect -35 1015 -15 1035
rect -15 1015 -10 1035
rect -40 1010 -10 1015
rect -40 935 -10 940
rect -40 915 -35 935
rect -35 915 -15 935
rect -15 915 -10 935
rect -40 910 -10 915
rect -340 810 -310 840
rect -640 735 -610 740
rect -640 715 -635 735
rect -635 715 -615 735
rect -615 715 -610 735
rect -640 710 -610 715
rect -640 635 -610 640
rect -640 615 -635 635
rect -635 615 -615 635
rect -615 615 -610 635
rect -640 610 -610 615
rect -640 535 -610 540
rect -640 515 -635 535
rect -635 515 -615 535
rect -615 515 -610 535
rect -640 510 -610 515
rect -640 435 -610 440
rect -640 415 -635 435
rect -635 415 -615 435
rect -615 415 -610 435
rect -640 410 -610 415
rect -640 335 -610 340
rect -640 315 -635 335
rect -635 315 -615 335
rect -615 315 -610 335
rect -640 310 -610 315
rect -640 235 -610 240
rect -640 215 -635 235
rect -635 215 -615 235
rect -615 215 -610 235
rect -640 210 -610 215
rect -640 135 -610 140
rect -640 115 -635 135
rect -635 115 -615 135
rect -615 115 -610 135
rect -640 110 -610 115
rect -190 835 -160 840
rect -190 815 -185 835
rect -185 815 -165 835
rect -165 815 -160 835
rect -190 810 -160 815
rect 10760 1685 10790 1690
rect 10760 1665 10765 1685
rect 10765 1665 10785 1685
rect 10785 1665 10790 1685
rect 10760 1660 10790 1665
rect 8360 1535 8390 1540
rect 8360 1515 8365 1535
rect 8365 1515 8385 1535
rect 8385 1515 8390 1535
rect 8360 1510 8390 1515
rect 8360 1435 8390 1440
rect 8360 1415 8365 1435
rect 8365 1415 8385 1435
rect 8385 1415 8390 1435
rect 8360 1410 8390 1415
rect 8360 1335 8390 1340
rect 8360 1315 8365 1335
rect 8365 1315 8385 1335
rect 8385 1315 8390 1335
rect 8360 1310 8390 1315
rect 8360 1235 8390 1240
rect 8360 1215 8365 1235
rect 8365 1215 8385 1235
rect 8385 1215 8390 1235
rect 8360 1210 8390 1215
rect 8360 1135 8390 1140
rect 8360 1115 8365 1135
rect 8365 1115 8385 1135
rect 8385 1115 8390 1135
rect 8360 1110 8390 1115
rect 8360 1035 8390 1040
rect 8360 1015 8365 1035
rect 8365 1015 8385 1035
rect 8385 1015 8390 1035
rect 8360 1010 8390 1015
rect 8360 935 8390 940
rect 8360 915 8365 935
rect 8365 915 8385 935
rect 8385 915 8390 935
rect 8360 910 8390 915
rect 110 835 140 840
rect 110 815 115 835
rect 115 815 135 835
rect 135 815 140 835
rect 110 810 140 815
rect 410 835 440 840
rect 410 815 415 835
rect 415 815 435 835
rect 435 815 440 835
rect 410 810 440 815
rect 710 835 740 840
rect 710 815 715 835
rect 715 815 735 835
rect 735 815 740 835
rect 710 810 740 815
rect 1010 835 1040 840
rect 1010 815 1015 835
rect 1015 815 1035 835
rect 1035 815 1040 835
rect 1010 810 1040 815
rect 1310 835 1340 840
rect 1310 815 1315 835
rect 1315 815 1335 835
rect 1335 815 1340 835
rect 1310 810 1340 815
rect 1610 835 1640 840
rect 1610 815 1615 835
rect 1615 815 1635 835
rect 1635 815 1640 835
rect 1610 810 1640 815
rect 1910 835 1940 840
rect 1910 815 1915 835
rect 1915 815 1935 835
rect 1935 815 1940 835
rect 1910 810 1940 815
rect 2210 835 2240 840
rect 2210 815 2215 835
rect 2215 815 2235 835
rect 2235 815 2240 835
rect 2210 810 2240 815
rect 2360 810 2390 840
rect 2510 835 2540 840
rect 2510 815 2515 835
rect 2515 815 2535 835
rect 2535 815 2540 835
rect 2510 810 2540 815
rect 2810 835 2840 840
rect 2810 815 2815 835
rect 2815 815 2835 835
rect 2835 815 2840 835
rect 2810 810 2840 815
rect 3110 835 3140 840
rect 3110 815 3115 835
rect 3115 815 3135 835
rect 3135 815 3140 835
rect 3110 810 3140 815
rect 3410 835 3440 840
rect 3410 815 3415 835
rect 3415 815 3435 835
rect 3435 815 3440 835
rect 3410 810 3440 815
rect 3710 835 3740 840
rect 3710 815 3715 835
rect 3715 815 3735 835
rect 3735 815 3740 835
rect 3710 810 3740 815
rect 3860 810 3890 840
rect 4010 835 4040 840
rect 4010 815 4015 835
rect 4015 815 4035 835
rect 4035 815 4040 835
rect 4010 810 4040 815
rect 4310 835 4340 840
rect 4310 815 4315 835
rect 4315 815 4335 835
rect 4335 815 4340 835
rect 4310 810 4340 815
rect 4460 810 4490 840
rect 4610 835 4640 840
rect 4610 815 4615 835
rect 4615 815 4635 835
rect 4635 815 4640 835
rect 4610 810 4640 815
rect 4910 835 4940 840
rect 4910 815 4915 835
rect 4915 815 4935 835
rect 4935 815 4940 835
rect 4910 810 4940 815
rect 5210 835 5240 840
rect 5210 815 5215 835
rect 5215 815 5235 835
rect 5235 815 5240 835
rect 5210 810 5240 815
rect 5510 835 5540 840
rect 5510 815 5515 835
rect 5515 815 5535 835
rect 5535 815 5540 835
rect 5510 810 5540 815
rect 5810 835 5840 840
rect 5810 815 5815 835
rect 5815 815 5835 835
rect 5835 815 5840 835
rect 5810 810 5840 815
rect 5960 810 5990 840
rect 6110 835 6140 840
rect 6110 815 6115 835
rect 6115 815 6135 835
rect 6135 815 6140 835
rect 6110 810 6140 815
rect 6410 835 6440 840
rect 6410 815 6415 835
rect 6415 815 6435 835
rect 6435 815 6440 835
rect 6410 810 6440 815
rect 6710 835 6740 840
rect 6710 815 6715 835
rect 6715 815 6735 835
rect 6735 815 6740 835
rect 6710 810 6740 815
rect 7010 835 7040 840
rect 7010 815 7015 835
rect 7015 815 7035 835
rect 7035 815 7040 835
rect 7010 810 7040 815
rect 7310 835 7340 840
rect 7310 815 7315 835
rect 7315 815 7335 835
rect 7335 815 7340 835
rect 7310 810 7340 815
rect 7610 835 7640 840
rect 7610 815 7615 835
rect 7615 815 7635 835
rect 7635 815 7640 835
rect 7610 810 7640 815
rect 7910 835 7940 840
rect 7910 815 7915 835
rect 7915 815 7935 835
rect 7935 815 7940 835
rect 7910 810 7940 815
rect 8210 835 8240 840
rect 8210 815 8215 835
rect 8215 815 8235 835
rect 8235 815 8240 835
rect 8210 810 8240 815
rect -40 735 -10 740
rect -40 715 -35 735
rect -35 715 -15 735
rect -15 715 -10 735
rect -40 710 -10 715
rect -40 635 -10 640
rect -40 615 -35 635
rect -35 615 -15 635
rect -15 615 -10 635
rect -40 610 -10 615
rect -40 535 -10 540
rect -40 515 -35 535
rect -35 515 -15 535
rect -15 515 -10 535
rect -40 510 -10 515
rect -40 435 -10 440
rect -40 415 -35 435
rect -35 415 -15 435
rect -15 415 -10 435
rect -40 410 -10 415
rect -40 335 -10 340
rect -40 315 -35 335
rect -35 315 -15 335
rect -15 315 -10 335
rect -40 310 -10 315
rect -40 235 -10 240
rect -40 215 -35 235
rect -35 215 -15 235
rect -15 215 -10 235
rect -40 210 -10 215
rect -40 135 -10 140
rect -40 115 -35 135
rect -35 115 -15 135
rect -15 115 -10 135
rect -40 110 -10 115
rect -640 -15 -610 -10
rect -640 -35 -635 -15
rect -635 -35 -615 -15
rect -615 -35 -610 -15
rect -640 -40 -610 -35
rect 8510 835 8540 840
rect 8510 815 8515 835
rect 8515 815 8535 835
rect 8535 815 8540 835
rect 8510 810 8540 815
rect 8810 835 8840 840
rect 8810 815 8815 835
rect 8815 815 8835 835
rect 8835 815 8840 835
rect 8810 810 8840 815
rect 9110 835 9140 840
rect 9110 815 9115 835
rect 9115 815 9135 835
rect 9135 815 9140 835
rect 9110 810 9140 815
rect 9410 835 9440 840
rect 9410 815 9415 835
rect 9415 815 9435 835
rect 9435 815 9440 835
rect 9410 810 9440 815
rect 15560 1685 15590 1690
rect 15560 1665 15565 1685
rect 15565 1665 15585 1685
rect 15585 1665 15590 1685
rect 15560 1660 15590 1665
rect 10760 1535 10790 1540
rect 10760 1515 10765 1535
rect 10765 1515 10785 1535
rect 10785 1515 10790 1535
rect 10760 1510 10790 1515
rect 10760 1435 10790 1440
rect 10760 1415 10765 1435
rect 10765 1415 10785 1435
rect 10785 1415 10790 1435
rect 10760 1410 10790 1415
rect 10760 1335 10790 1340
rect 10760 1315 10765 1335
rect 10765 1315 10785 1335
rect 10785 1315 10790 1335
rect 10760 1310 10790 1315
rect 10760 1235 10790 1240
rect 10760 1215 10765 1235
rect 10765 1215 10785 1235
rect 10785 1215 10790 1235
rect 10760 1210 10790 1215
rect 10760 1135 10790 1140
rect 10760 1115 10765 1135
rect 10765 1115 10785 1135
rect 10785 1115 10790 1135
rect 10760 1110 10790 1115
rect 10760 1035 10790 1040
rect 10760 1015 10765 1035
rect 10765 1015 10785 1035
rect 10785 1015 10790 1035
rect 10760 1010 10790 1015
rect 10760 935 10790 940
rect 10760 915 10765 935
rect 10765 915 10785 935
rect 10785 915 10790 935
rect 10760 910 10790 915
rect 9560 810 9590 840
rect 8360 735 8390 740
rect 8360 715 8365 735
rect 8365 715 8385 735
rect 8385 715 8390 735
rect 8360 710 8390 715
rect 8360 635 8390 640
rect 8360 615 8365 635
rect 8365 615 8385 635
rect 8385 615 8390 635
rect 8360 610 8390 615
rect 8360 535 8390 540
rect 8360 515 8365 535
rect 8365 515 8385 535
rect 8385 515 8390 535
rect 8360 510 8390 515
rect 8360 435 8390 440
rect 8360 415 8365 435
rect 8365 415 8385 435
rect 8385 415 8390 435
rect 8360 410 8390 415
rect 8360 335 8390 340
rect 8360 315 8365 335
rect 8365 315 8385 335
rect 8385 315 8390 335
rect 8360 310 8390 315
rect 8360 235 8390 240
rect 8360 215 8365 235
rect 8365 215 8385 235
rect 8385 215 8390 235
rect 8360 210 8390 215
rect 8360 135 8390 140
rect 8360 115 8365 135
rect 8365 115 8385 135
rect 8385 115 8390 135
rect 8360 110 8390 115
rect -40 -15 -10 -10
rect -40 -35 -35 -15
rect -35 -35 -15 -15
rect -15 -35 -10 -15
rect -40 -40 -10 -35
rect -640 -165 -610 -160
rect -640 -185 -635 -165
rect -635 -185 -615 -165
rect -615 -185 -610 -165
rect -640 -190 -610 -185
rect -640 -265 -610 -260
rect -640 -285 -635 -265
rect -635 -285 -615 -265
rect -615 -285 -610 -265
rect -640 -290 -610 -285
rect -640 -365 -610 -360
rect -640 -385 -635 -365
rect -635 -385 -615 -365
rect -615 -385 -610 -365
rect -640 -390 -610 -385
rect -640 -465 -610 -460
rect -640 -485 -635 -465
rect -635 -485 -615 -465
rect -615 -485 -610 -465
rect -640 -490 -610 -485
rect -640 -565 -610 -560
rect -640 -585 -635 -565
rect -635 -585 -615 -565
rect -615 -585 -610 -565
rect -640 -590 -610 -585
rect -640 -665 -610 -660
rect -640 -685 -635 -665
rect -635 -685 -615 -665
rect -615 -685 -610 -665
rect -640 -690 -610 -685
rect -640 -765 -610 -760
rect -640 -785 -635 -765
rect -635 -785 -615 -765
rect -615 -785 -610 -765
rect -640 -790 -610 -785
rect -490 -865 -460 -860
rect -490 -885 -485 -865
rect -485 -885 -465 -865
rect -465 -885 -460 -865
rect -490 -890 -460 -885
rect 9710 835 9740 840
rect 9710 815 9715 835
rect 9715 815 9735 835
rect 9735 815 9740 835
rect 9710 810 9740 815
rect 10010 835 10040 840
rect 10010 815 10015 835
rect 10015 815 10035 835
rect 10035 815 10040 835
rect 10010 810 10040 815
rect 10310 835 10340 840
rect 10310 815 10315 835
rect 10315 815 10335 835
rect 10335 815 10340 835
rect 10310 810 10340 815
rect 10610 835 10640 840
rect 10610 815 10615 835
rect 10615 815 10635 835
rect 10635 815 10640 835
rect 10610 810 10640 815
rect 10910 835 10940 840
rect 10910 815 10915 835
rect 10915 815 10935 835
rect 10935 815 10940 835
rect 10910 810 10940 815
rect 11210 835 11240 840
rect 11210 815 11215 835
rect 11215 815 11235 835
rect 11235 815 11240 835
rect 11210 810 11240 815
rect 11510 835 11540 840
rect 11510 815 11515 835
rect 11515 815 11535 835
rect 11535 815 11540 835
rect 11510 810 11540 815
rect 11810 835 11840 840
rect 11810 815 11815 835
rect 11815 815 11835 835
rect 11835 815 11840 835
rect 11810 810 11840 815
rect 10760 735 10790 740
rect 10760 715 10765 735
rect 10765 715 10785 735
rect 10785 715 10790 735
rect 10760 710 10790 715
rect 10760 635 10790 640
rect 10760 615 10765 635
rect 10765 615 10785 635
rect 10785 615 10790 635
rect 10760 610 10790 615
rect 10760 535 10790 540
rect 10760 515 10765 535
rect 10765 515 10785 535
rect 10785 515 10790 535
rect 10760 510 10790 515
rect 10760 435 10790 440
rect 10760 415 10765 435
rect 10765 415 10785 435
rect 10785 415 10790 435
rect 10760 410 10790 415
rect 10760 335 10790 340
rect 10760 315 10765 335
rect 10765 315 10785 335
rect 10785 315 10790 335
rect 10760 310 10790 315
rect 10760 235 10790 240
rect 10760 215 10765 235
rect 10765 215 10785 235
rect 10785 215 10790 235
rect 10760 210 10790 215
rect 10760 135 10790 140
rect 10760 115 10765 135
rect 10765 115 10785 135
rect 10785 115 10790 135
rect 10760 110 10790 115
rect 8360 -15 8390 -10
rect 8360 -35 8365 -15
rect 8365 -35 8385 -15
rect 8385 -35 8390 -15
rect 8360 -40 8390 -35
rect -40 -165 -10 -160
rect -40 -185 -35 -165
rect -35 -185 -15 -165
rect -15 -185 -10 -165
rect -40 -190 -10 -185
rect -40 -265 -10 -260
rect -40 -285 -35 -265
rect -35 -285 -15 -265
rect -15 -285 -10 -265
rect -40 -290 -10 -285
rect -40 -365 -10 -360
rect -40 -385 -35 -365
rect -35 -385 -15 -365
rect -15 -385 -10 -365
rect -40 -390 -10 -385
rect -40 -465 -10 -460
rect -40 -485 -35 -465
rect -35 -485 -15 -465
rect -15 -485 -10 -465
rect -40 -490 -10 -485
rect -40 -565 -10 -560
rect -40 -585 -35 -565
rect -35 -585 -15 -565
rect -15 -585 -10 -565
rect -40 -590 -10 -585
rect -40 -665 -10 -660
rect -40 -685 -35 -665
rect -35 -685 -15 -665
rect -15 -685 -10 -665
rect -40 -690 -10 -685
rect -40 -765 -10 -760
rect -40 -785 -35 -765
rect -35 -785 -15 -765
rect -15 -785 -10 -765
rect -40 -790 -10 -785
rect -340 -890 -310 -860
rect -640 -965 -610 -960
rect -640 -985 -635 -965
rect -635 -985 -615 -965
rect -615 -985 -610 -965
rect -640 -990 -610 -985
rect -640 -1065 -610 -1060
rect -640 -1085 -635 -1065
rect -635 -1085 -615 -1065
rect -615 -1085 -610 -1065
rect -640 -1090 -610 -1085
rect -640 -1165 -610 -1160
rect -640 -1185 -635 -1165
rect -635 -1185 -615 -1165
rect -615 -1185 -610 -1165
rect -640 -1190 -610 -1185
rect -640 -1265 -610 -1260
rect -640 -1285 -635 -1265
rect -635 -1285 -615 -1265
rect -615 -1285 -610 -1265
rect -640 -1290 -610 -1285
rect -640 -1365 -610 -1360
rect -640 -1385 -635 -1365
rect -635 -1385 -615 -1365
rect -615 -1385 -610 -1365
rect -640 -1390 -610 -1385
rect -640 -1465 -610 -1460
rect -640 -1485 -635 -1465
rect -635 -1485 -615 -1465
rect -615 -1485 -610 -1465
rect -640 -1490 -610 -1485
rect -640 -1565 -610 -1560
rect -640 -1585 -635 -1565
rect -635 -1585 -615 -1565
rect -615 -1585 -610 -1565
rect -640 -1590 -610 -1585
rect -190 -865 -160 -860
rect -190 -885 -185 -865
rect -185 -885 -165 -865
rect -165 -885 -160 -865
rect -190 -890 -160 -885
rect 10760 -15 10790 -10
rect 10760 -35 10765 -15
rect 10765 -35 10785 -15
rect 10785 -35 10790 -15
rect 10760 -40 10790 -35
rect 8360 -165 8390 -160
rect 8360 -185 8365 -165
rect 8365 -185 8385 -165
rect 8385 -185 8390 -165
rect 8360 -190 8390 -185
rect 8360 -265 8390 -260
rect 8360 -285 8365 -265
rect 8365 -285 8385 -265
rect 8385 -285 8390 -265
rect 8360 -290 8390 -285
rect 8360 -365 8390 -360
rect 8360 -385 8365 -365
rect 8365 -385 8385 -365
rect 8385 -385 8390 -365
rect 8360 -390 8390 -385
rect 8360 -465 8390 -460
rect 8360 -485 8365 -465
rect 8365 -485 8385 -465
rect 8385 -485 8390 -465
rect 8360 -490 8390 -485
rect 8360 -565 8390 -560
rect 8360 -585 8365 -565
rect 8365 -585 8385 -565
rect 8385 -585 8390 -565
rect 8360 -590 8390 -585
rect 8360 -665 8390 -660
rect 8360 -685 8365 -665
rect 8365 -685 8385 -665
rect 8385 -685 8390 -665
rect 8360 -690 8390 -685
rect 8360 -765 8390 -760
rect 8360 -785 8365 -765
rect 8365 -785 8385 -765
rect 8385 -785 8390 -765
rect 8360 -790 8390 -785
rect 110 -865 140 -860
rect 110 -885 115 -865
rect 115 -885 135 -865
rect 135 -885 140 -865
rect 110 -890 140 -885
rect 410 -865 440 -860
rect 410 -885 415 -865
rect 415 -885 435 -865
rect 435 -885 440 -865
rect 410 -890 440 -885
rect 710 -865 740 -860
rect 710 -885 715 -865
rect 715 -885 735 -865
rect 735 -885 740 -865
rect 710 -890 740 -885
rect 1010 -865 1040 -860
rect 1010 -885 1015 -865
rect 1015 -885 1035 -865
rect 1035 -885 1040 -865
rect 1010 -890 1040 -885
rect 1310 -865 1340 -860
rect 1310 -885 1315 -865
rect 1315 -885 1335 -865
rect 1335 -885 1340 -865
rect 1310 -890 1340 -885
rect 1610 -865 1640 -860
rect 1610 -885 1615 -865
rect 1615 -885 1635 -865
rect 1635 -885 1640 -865
rect 1610 -890 1640 -885
rect 1910 -865 1940 -860
rect 1910 -885 1915 -865
rect 1915 -885 1935 -865
rect 1935 -885 1940 -865
rect 1910 -890 1940 -885
rect 2210 -865 2240 -860
rect 2210 -885 2215 -865
rect 2215 -885 2235 -865
rect 2235 -885 2240 -865
rect 2210 -890 2240 -885
rect 2360 -890 2390 -860
rect 2510 -865 2540 -860
rect 2510 -885 2515 -865
rect 2515 -885 2535 -865
rect 2535 -885 2540 -865
rect 2510 -890 2540 -885
rect 2810 -865 2840 -860
rect 2810 -885 2815 -865
rect 2815 -885 2835 -865
rect 2835 -885 2840 -865
rect 2810 -890 2840 -885
rect 3110 -865 3140 -860
rect 3110 -885 3115 -865
rect 3115 -885 3135 -865
rect 3135 -885 3140 -865
rect 3110 -890 3140 -885
rect 3410 -865 3440 -860
rect 3410 -885 3415 -865
rect 3415 -885 3435 -865
rect 3435 -885 3440 -865
rect 3410 -890 3440 -885
rect 3710 -865 3740 -860
rect 3710 -885 3715 -865
rect 3715 -885 3735 -865
rect 3735 -885 3740 -865
rect 3710 -890 3740 -885
rect 3860 -890 3890 -860
rect 4010 -865 4040 -860
rect 4010 -885 4015 -865
rect 4015 -885 4035 -865
rect 4035 -885 4040 -865
rect 4010 -890 4040 -885
rect 4310 -865 4340 -860
rect 4310 -885 4315 -865
rect 4315 -885 4335 -865
rect 4335 -885 4340 -865
rect 4310 -890 4340 -885
rect 4460 -890 4490 -860
rect 4610 -865 4640 -860
rect 4610 -885 4615 -865
rect 4615 -885 4635 -865
rect 4635 -885 4640 -865
rect 4610 -890 4640 -885
rect 4910 -865 4940 -860
rect 4910 -885 4915 -865
rect 4915 -885 4935 -865
rect 4935 -885 4940 -865
rect 4910 -890 4940 -885
rect 5210 -865 5240 -860
rect 5210 -885 5215 -865
rect 5215 -885 5235 -865
rect 5235 -885 5240 -865
rect 5210 -890 5240 -885
rect 5510 -865 5540 -860
rect 5510 -885 5515 -865
rect 5515 -885 5535 -865
rect 5535 -885 5540 -865
rect 5510 -890 5540 -885
rect 5810 -865 5840 -860
rect 5810 -885 5815 -865
rect 5815 -885 5835 -865
rect 5835 -885 5840 -865
rect 5810 -890 5840 -885
rect 5960 -890 5990 -860
rect 6110 -865 6140 -860
rect 6110 -885 6115 -865
rect 6115 -885 6135 -865
rect 6135 -885 6140 -865
rect 6110 -890 6140 -885
rect 6410 -865 6440 -860
rect 6410 -885 6415 -865
rect 6415 -885 6435 -865
rect 6435 -885 6440 -865
rect 6410 -890 6440 -885
rect 6710 -865 6740 -860
rect 6710 -885 6715 -865
rect 6715 -885 6735 -865
rect 6735 -885 6740 -865
rect 6710 -890 6740 -885
rect 7010 -865 7040 -860
rect 7010 -885 7015 -865
rect 7015 -885 7035 -865
rect 7035 -885 7040 -865
rect 7010 -890 7040 -885
rect 7310 -865 7340 -860
rect 7310 -885 7315 -865
rect 7315 -885 7335 -865
rect 7335 -885 7340 -865
rect 7310 -890 7340 -885
rect 7610 -865 7640 -860
rect 7610 -885 7615 -865
rect 7615 -885 7635 -865
rect 7635 -885 7640 -865
rect 7610 -890 7640 -885
rect 7910 -865 7940 -860
rect 7910 -885 7915 -865
rect 7915 -885 7935 -865
rect 7935 -885 7940 -865
rect 7910 -890 7940 -885
rect 8210 -865 8240 -860
rect 8210 -885 8215 -865
rect 8215 -885 8235 -865
rect 8235 -885 8240 -865
rect 8210 -890 8240 -885
rect -40 -965 -10 -960
rect -40 -985 -35 -965
rect -35 -985 -15 -965
rect -15 -985 -10 -965
rect -40 -990 -10 -985
rect -40 -1065 -10 -1060
rect -40 -1085 -35 -1065
rect -35 -1085 -15 -1065
rect -15 -1085 -10 -1065
rect -40 -1090 -10 -1085
rect -40 -1165 -10 -1160
rect -40 -1185 -35 -1165
rect -35 -1185 -15 -1165
rect -15 -1185 -10 -1165
rect -40 -1190 -10 -1185
rect -40 -1265 -10 -1260
rect -40 -1285 -35 -1265
rect -35 -1285 -15 -1265
rect -15 -1285 -10 -1265
rect -40 -1290 -10 -1285
rect -40 -1365 -10 -1360
rect -40 -1385 -35 -1365
rect -35 -1385 -15 -1365
rect -15 -1385 -10 -1365
rect -40 -1390 -10 -1385
rect -40 -1465 -10 -1460
rect -40 -1485 -35 -1465
rect -35 -1485 -15 -1465
rect -15 -1485 -10 -1465
rect -40 -1490 -10 -1485
rect -40 -1565 -10 -1560
rect -40 -1585 -35 -1565
rect -35 -1585 -15 -1565
rect -15 -1585 -10 -1565
rect -40 -1590 -10 -1585
rect -640 -1715 -610 -1710
rect -640 -1735 -635 -1715
rect -635 -1735 -615 -1715
rect -615 -1735 -610 -1715
rect -640 -1740 -610 -1735
rect 8510 -865 8540 -860
rect 8510 -885 8515 -865
rect 8515 -885 8535 -865
rect 8535 -885 8540 -865
rect 8510 -890 8540 -885
rect 8810 -865 8840 -860
rect 8810 -885 8815 -865
rect 8815 -885 8835 -865
rect 8835 -885 8840 -865
rect 8810 -890 8840 -885
rect 9110 -865 9140 -860
rect 9110 -885 9115 -865
rect 9115 -885 9135 -865
rect 9135 -885 9140 -865
rect 9110 -890 9140 -885
rect 9410 -865 9440 -860
rect 9410 -885 9415 -865
rect 9415 -885 9435 -865
rect 9435 -885 9440 -865
rect 9410 -890 9440 -885
rect 10760 -165 10790 -160
rect 10760 -185 10765 -165
rect 10765 -185 10785 -165
rect 10785 -185 10790 -165
rect 10760 -190 10790 -185
rect 10760 -265 10790 -260
rect 10760 -285 10765 -265
rect 10765 -285 10785 -265
rect 10785 -285 10790 -265
rect 10760 -290 10790 -285
rect 10760 -365 10790 -360
rect 10760 -385 10765 -365
rect 10765 -385 10785 -365
rect 10785 -385 10790 -365
rect 10760 -390 10790 -385
rect 10760 -465 10790 -460
rect 10760 -485 10765 -465
rect 10765 -485 10785 -465
rect 10785 -485 10790 -465
rect 10760 -490 10790 -485
rect 10760 -565 10790 -560
rect 10760 -585 10765 -565
rect 10765 -585 10785 -565
rect 10785 -585 10790 -565
rect 10760 -590 10790 -585
rect 10760 -665 10790 -660
rect 10760 -685 10765 -665
rect 10765 -685 10785 -665
rect 10785 -685 10790 -665
rect 10760 -690 10790 -685
rect 10760 -765 10790 -760
rect 10760 -785 10765 -765
rect 10765 -785 10785 -765
rect 10785 -785 10790 -765
rect 10760 -790 10790 -785
rect 9560 -890 9590 -860
rect 8360 -965 8390 -960
rect 8360 -985 8365 -965
rect 8365 -985 8385 -965
rect 8385 -985 8390 -965
rect 8360 -990 8390 -985
rect 8360 -1065 8390 -1060
rect 8360 -1085 8365 -1065
rect 8365 -1085 8385 -1065
rect 8385 -1085 8390 -1065
rect 8360 -1090 8390 -1085
rect 8360 -1165 8390 -1160
rect 8360 -1185 8365 -1165
rect 8365 -1185 8385 -1165
rect 8385 -1185 8390 -1165
rect 8360 -1190 8390 -1185
rect 8360 -1265 8390 -1260
rect 8360 -1285 8365 -1265
rect 8365 -1285 8385 -1265
rect 8385 -1285 8390 -1265
rect 8360 -1290 8390 -1285
rect 8360 -1365 8390 -1360
rect 8360 -1385 8365 -1365
rect 8365 -1385 8385 -1365
rect 8385 -1385 8390 -1365
rect 8360 -1390 8390 -1385
rect 8360 -1465 8390 -1460
rect 8360 -1485 8365 -1465
rect 8365 -1485 8385 -1465
rect 8385 -1485 8390 -1465
rect 8360 -1490 8390 -1485
rect 8360 -1565 8390 -1560
rect 8360 -1585 8365 -1565
rect 8365 -1585 8385 -1565
rect 8385 -1585 8390 -1565
rect 8360 -1590 8390 -1585
rect -40 -1715 -10 -1710
rect -40 -1735 -35 -1715
rect -35 -1735 -15 -1715
rect -15 -1735 -10 -1715
rect -40 -1740 -10 -1735
rect 9710 -865 9740 -860
rect 9710 -885 9715 -865
rect 9715 -885 9735 -865
rect 9735 -885 9740 -865
rect 9710 -890 9740 -885
rect 10010 -865 10040 -860
rect 10010 -885 10015 -865
rect 10015 -885 10035 -865
rect 10035 -885 10040 -865
rect 10010 -890 10040 -885
rect 10310 -865 10340 -860
rect 10310 -885 10315 -865
rect 10315 -885 10335 -865
rect 10335 -885 10340 -865
rect 10310 -890 10340 -885
rect 10610 -865 10640 -860
rect 10610 -885 10615 -865
rect 10615 -885 10635 -865
rect 10635 -885 10640 -865
rect 10610 -890 10640 -885
rect 12110 835 12140 840
rect 12110 815 12115 835
rect 12115 815 12135 835
rect 12135 815 12140 835
rect 12110 810 12140 815
rect 12410 835 12440 840
rect 12410 815 12415 835
rect 12415 815 12435 835
rect 12435 815 12440 835
rect 12410 810 12440 815
rect 12560 810 12590 840
rect 12710 835 12740 840
rect 12710 815 12715 835
rect 12715 815 12735 835
rect 12735 815 12740 835
rect 12710 810 12740 815
rect 13010 835 13040 840
rect 13010 815 13015 835
rect 13015 815 13035 835
rect 13035 815 13040 835
rect 13010 810 13040 815
rect 13160 810 13190 840
rect 13310 835 13340 840
rect 13310 815 13315 835
rect 13315 815 13335 835
rect 13335 815 13340 835
rect 13310 810 13340 815
rect 13610 835 13640 840
rect 13610 815 13615 835
rect 13615 815 13635 835
rect 13635 815 13640 835
rect 13610 810 13640 815
rect 13760 810 13790 840
rect 13910 835 13940 840
rect 13910 815 13915 835
rect 13915 815 13935 835
rect 13935 815 13940 835
rect 13910 810 13940 815
rect 14210 835 14240 840
rect 14210 815 14215 835
rect 14215 815 14235 835
rect 14235 815 14240 835
rect 14210 810 14240 815
rect 17960 1685 17990 1690
rect 17960 1665 17965 1685
rect 17965 1665 17985 1685
rect 17985 1665 17990 1685
rect 17960 1660 17990 1665
rect 15560 1535 15590 1540
rect 15560 1515 15565 1535
rect 15565 1515 15585 1535
rect 15585 1515 15590 1535
rect 15560 1510 15590 1515
rect 15560 1435 15590 1440
rect 15560 1415 15565 1435
rect 15565 1415 15585 1435
rect 15585 1415 15590 1435
rect 15560 1410 15590 1415
rect 15560 1335 15590 1340
rect 15560 1315 15565 1335
rect 15565 1315 15585 1335
rect 15585 1315 15590 1335
rect 15560 1310 15590 1315
rect 15560 1235 15590 1240
rect 15560 1215 15565 1235
rect 15565 1215 15585 1235
rect 15585 1215 15590 1235
rect 15560 1210 15590 1215
rect 15560 1135 15590 1140
rect 15560 1115 15565 1135
rect 15565 1115 15585 1135
rect 15585 1115 15590 1135
rect 15560 1110 15590 1115
rect 15560 1035 15590 1040
rect 15560 1015 15565 1035
rect 15565 1015 15585 1035
rect 15585 1015 15590 1035
rect 15560 1010 15590 1015
rect 15560 935 15590 940
rect 15560 915 15565 935
rect 15565 915 15585 935
rect 15585 915 15590 935
rect 15560 910 15590 915
rect 14510 835 14540 840
rect 14510 815 14515 835
rect 14515 815 14535 835
rect 14535 815 14540 835
rect 14510 810 14540 815
rect 14810 835 14840 840
rect 14810 815 14815 835
rect 14815 815 14835 835
rect 14835 815 14840 835
rect 14810 810 14840 815
rect 15110 835 15140 840
rect 15110 815 15115 835
rect 15115 815 15135 835
rect 15135 815 15140 835
rect 15110 810 15140 815
rect 15410 835 15440 840
rect 15410 815 15415 835
rect 15415 815 15435 835
rect 15435 815 15440 835
rect 15410 810 15440 815
rect 10910 -865 10940 -860
rect 10910 -885 10915 -865
rect 10915 -885 10935 -865
rect 10935 -885 10940 -865
rect 10910 -890 10940 -885
rect 11210 -865 11240 -860
rect 11210 -885 11215 -865
rect 11215 -885 11235 -865
rect 11235 -885 11240 -865
rect 11210 -890 11240 -885
rect 11510 -865 11540 -860
rect 11510 -885 11515 -865
rect 11515 -885 11535 -865
rect 11535 -885 11540 -865
rect 11510 -890 11540 -885
rect 11810 -865 11840 -860
rect 11810 -885 11815 -865
rect 11815 -885 11835 -865
rect 11835 -885 11840 -865
rect 11810 -890 11840 -885
rect 10760 -965 10790 -960
rect 10760 -985 10765 -965
rect 10765 -985 10785 -965
rect 10785 -985 10790 -965
rect 10760 -990 10790 -985
rect 10760 -1065 10790 -1060
rect 10760 -1085 10765 -1065
rect 10765 -1085 10785 -1065
rect 10785 -1085 10790 -1065
rect 10760 -1090 10790 -1085
rect 10760 -1165 10790 -1160
rect 10760 -1185 10765 -1165
rect 10765 -1185 10785 -1165
rect 10785 -1185 10790 -1165
rect 10760 -1190 10790 -1185
rect 10760 -1265 10790 -1260
rect 10760 -1285 10765 -1265
rect 10765 -1285 10785 -1265
rect 10785 -1285 10790 -1265
rect 10760 -1290 10790 -1285
rect 10760 -1365 10790 -1360
rect 10760 -1385 10765 -1365
rect 10765 -1385 10785 -1365
rect 10785 -1385 10790 -1365
rect 10760 -1390 10790 -1385
rect 10760 -1465 10790 -1460
rect 10760 -1485 10765 -1465
rect 10765 -1485 10785 -1465
rect 10785 -1485 10790 -1465
rect 10760 -1490 10790 -1485
rect 10760 -1565 10790 -1560
rect 10760 -1585 10765 -1565
rect 10765 -1585 10785 -1565
rect 10785 -1585 10790 -1565
rect 10760 -1590 10790 -1585
rect 8360 -1715 8390 -1710
rect 8360 -1735 8365 -1715
rect 8365 -1735 8385 -1715
rect 8385 -1735 8390 -1715
rect 8360 -1740 8390 -1735
rect 12110 -865 12140 -860
rect 12110 -885 12115 -865
rect 12115 -885 12135 -865
rect 12135 -885 12140 -865
rect 12110 -890 12140 -885
rect 12410 -865 12440 -860
rect 12410 -885 12415 -865
rect 12415 -885 12435 -865
rect 12435 -885 12440 -865
rect 12410 -890 12440 -885
rect 12560 -890 12590 -860
rect 12710 -865 12740 -860
rect 12710 -885 12715 -865
rect 12715 -885 12735 -865
rect 12735 -885 12740 -865
rect 12710 -890 12740 -885
rect 13010 -865 13040 -860
rect 13010 -885 13015 -865
rect 13015 -885 13035 -865
rect 13035 -885 13040 -865
rect 13010 -890 13040 -885
rect 13160 -890 13190 -860
rect 13310 -865 13340 -860
rect 13310 -885 13315 -865
rect 13315 -885 13335 -865
rect 13335 -885 13340 -865
rect 13310 -890 13340 -885
rect 13610 -865 13640 -860
rect 13610 -885 13615 -865
rect 13615 -885 13635 -865
rect 13635 -885 13640 -865
rect 13610 -890 13640 -885
rect 13760 -890 13790 -860
rect 13910 -865 13940 -860
rect 13910 -885 13915 -865
rect 13915 -885 13935 -865
rect 13935 -885 13940 -865
rect 13910 -890 13940 -885
rect 14210 -865 14240 -860
rect 14210 -885 14215 -865
rect 14215 -885 14235 -865
rect 14235 -885 14240 -865
rect 14210 -890 14240 -885
rect 15710 835 15740 840
rect 15710 815 15715 835
rect 15715 815 15735 835
rect 15735 815 15740 835
rect 15710 810 15740 815
rect 16010 835 16040 840
rect 16010 815 16015 835
rect 16015 815 16035 835
rect 16035 815 16040 835
rect 16010 810 16040 815
rect 16310 835 16340 840
rect 16310 815 16315 835
rect 16315 815 16335 835
rect 16335 815 16340 835
rect 16310 810 16340 815
rect 16610 835 16640 840
rect 16610 815 16615 835
rect 16615 815 16635 835
rect 16635 815 16640 835
rect 16610 810 16640 815
rect 20360 1685 20390 1690
rect 20360 1665 20365 1685
rect 20365 1665 20385 1685
rect 20385 1665 20390 1685
rect 20360 1660 20390 1665
rect 17960 1535 17990 1540
rect 17960 1515 17965 1535
rect 17965 1515 17985 1535
rect 17985 1515 17990 1535
rect 17960 1510 17990 1515
rect 17960 1435 17990 1440
rect 17960 1415 17965 1435
rect 17965 1415 17985 1435
rect 17985 1415 17990 1435
rect 17960 1410 17990 1415
rect 17960 1335 17990 1340
rect 17960 1315 17965 1335
rect 17965 1315 17985 1335
rect 17985 1315 17990 1335
rect 17960 1310 17990 1315
rect 17960 1235 17990 1240
rect 17960 1215 17965 1235
rect 17965 1215 17985 1235
rect 17985 1215 17990 1235
rect 17960 1210 17990 1215
rect 17960 1135 17990 1140
rect 17960 1115 17965 1135
rect 17965 1115 17985 1135
rect 17985 1115 17990 1135
rect 17960 1110 17990 1115
rect 17960 1035 17990 1040
rect 17960 1015 17965 1035
rect 17965 1015 17985 1035
rect 17985 1015 17990 1035
rect 17960 1010 17990 1015
rect 17960 935 17990 940
rect 17960 915 17965 935
rect 17965 915 17985 935
rect 17985 915 17990 935
rect 17960 910 17990 915
rect 16760 810 16790 840
rect 15560 735 15590 740
rect 15560 715 15565 735
rect 15565 715 15585 735
rect 15585 715 15590 735
rect 15560 710 15590 715
rect 15560 635 15590 640
rect 15560 615 15565 635
rect 15565 615 15585 635
rect 15585 615 15590 635
rect 15560 610 15590 615
rect 15560 535 15590 540
rect 15560 515 15565 535
rect 15565 515 15585 535
rect 15585 515 15590 535
rect 15560 510 15590 515
rect 15560 435 15590 440
rect 15560 415 15565 435
rect 15565 415 15585 435
rect 15585 415 15590 435
rect 15560 410 15590 415
rect 15560 335 15590 340
rect 15560 315 15565 335
rect 15565 315 15585 335
rect 15585 315 15590 335
rect 15560 310 15590 315
rect 15560 235 15590 240
rect 15560 215 15565 235
rect 15565 215 15585 235
rect 15585 215 15590 235
rect 15560 210 15590 215
rect 15560 135 15590 140
rect 15560 115 15565 135
rect 15565 115 15585 135
rect 15585 115 15590 135
rect 15560 110 15590 115
rect 16910 835 16940 840
rect 16910 815 16915 835
rect 16915 815 16935 835
rect 16935 815 16940 835
rect 16910 810 16940 815
rect 17210 835 17240 840
rect 17210 815 17215 835
rect 17215 815 17235 835
rect 17235 815 17240 835
rect 17210 810 17240 815
rect 17510 835 17540 840
rect 17510 815 17515 835
rect 17515 815 17535 835
rect 17535 815 17540 835
rect 17510 810 17540 815
rect 17810 835 17840 840
rect 17810 815 17815 835
rect 17815 815 17835 835
rect 17835 815 17840 835
rect 17810 810 17840 815
rect 18110 835 18140 840
rect 18110 815 18115 835
rect 18115 815 18135 835
rect 18135 815 18140 835
rect 18110 810 18140 815
rect 18410 835 18440 840
rect 18410 815 18415 835
rect 18415 815 18435 835
rect 18435 815 18440 835
rect 18410 810 18440 815
rect 18710 835 18740 840
rect 18710 815 18715 835
rect 18715 815 18735 835
rect 18735 815 18740 835
rect 18710 810 18740 815
rect 19010 835 19040 840
rect 19010 815 19015 835
rect 19015 815 19035 835
rect 19035 815 19040 835
rect 19010 810 19040 815
rect 20360 1535 20390 1540
rect 20360 1515 20365 1535
rect 20365 1515 20385 1535
rect 20385 1515 20390 1535
rect 20360 1510 20390 1515
rect 20360 1435 20390 1440
rect 20360 1415 20365 1435
rect 20365 1415 20385 1435
rect 20385 1415 20390 1435
rect 20360 1410 20390 1415
rect 20360 1335 20390 1340
rect 20360 1315 20365 1335
rect 20365 1315 20385 1335
rect 20385 1315 20390 1335
rect 20360 1310 20390 1315
rect 20360 1235 20390 1240
rect 20360 1215 20365 1235
rect 20365 1215 20385 1235
rect 20385 1215 20390 1235
rect 20360 1210 20390 1215
rect 20360 1135 20390 1140
rect 20360 1115 20365 1135
rect 20365 1115 20385 1135
rect 20385 1115 20390 1135
rect 20360 1110 20390 1115
rect 20360 1035 20390 1040
rect 20360 1015 20365 1035
rect 20365 1015 20385 1035
rect 20385 1015 20390 1035
rect 20360 1010 20390 1015
rect 20360 935 20390 940
rect 20360 915 20365 935
rect 20365 915 20385 935
rect 20385 915 20390 935
rect 20360 910 20390 915
rect 19160 810 19190 840
rect 17960 735 17990 740
rect 17960 715 17965 735
rect 17965 715 17985 735
rect 17985 715 17990 735
rect 17960 710 17990 715
rect 17960 635 17990 640
rect 17960 615 17965 635
rect 17965 615 17985 635
rect 17985 615 17990 635
rect 17960 610 17990 615
rect 17960 535 17990 540
rect 17960 515 17965 535
rect 17965 515 17985 535
rect 17985 515 17990 535
rect 17960 510 17990 515
rect 17960 435 17990 440
rect 17960 415 17965 435
rect 17965 415 17985 435
rect 17985 415 17990 435
rect 17960 410 17990 415
rect 17960 335 17990 340
rect 17960 315 17965 335
rect 17965 315 17985 335
rect 17985 315 17990 335
rect 17960 310 17990 315
rect 17960 235 17990 240
rect 17960 215 17965 235
rect 17965 215 17985 235
rect 17985 215 17990 235
rect 17960 210 17990 215
rect 17960 135 17990 140
rect 17960 115 17965 135
rect 17965 115 17985 135
rect 17985 115 17990 135
rect 17960 110 17990 115
rect 15560 -15 15590 -10
rect 15560 -35 15565 -15
rect 15565 -35 15585 -15
rect 15585 -35 15590 -15
rect 15560 -40 15590 -35
rect 19310 835 19340 840
rect 19310 815 19315 835
rect 19315 815 19335 835
rect 19335 815 19340 835
rect 19310 810 19340 815
rect 19610 835 19640 840
rect 19610 815 19615 835
rect 19615 815 19635 835
rect 19635 815 19640 835
rect 19610 810 19640 815
rect 19910 835 19940 840
rect 19910 815 19915 835
rect 19915 815 19935 835
rect 19935 815 19940 835
rect 19910 810 19940 815
rect 20210 835 20240 840
rect 20210 815 20215 835
rect 20215 815 20235 835
rect 20235 815 20240 835
rect 20210 810 20240 815
rect 20360 735 20390 740
rect 20360 715 20365 735
rect 20365 715 20385 735
rect 20385 715 20390 735
rect 20360 710 20390 715
rect 20360 635 20390 640
rect 20360 615 20365 635
rect 20365 615 20385 635
rect 20385 615 20390 635
rect 20360 610 20390 615
rect 20360 535 20390 540
rect 20360 515 20365 535
rect 20365 515 20385 535
rect 20385 515 20390 535
rect 20360 510 20390 515
rect 20360 435 20390 440
rect 20360 415 20365 435
rect 20365 415 20385 435
rect 20385 415 20390 435
rect 20360 410 20390 415
rect 20360 335 20390 340
rect 20360 315 20365 335
rect 20365 315 20385 335
rect 20385 315 20390 335
rect 20360 310 20390 315
rect 20360 235 20390 240
rect 20360 215 20365 235
rect 20365 215 20385 235
rect 20385 215 20390 235
rect 20360 210 20390 215
rect 20360 135 20390 140
rect 20360 115 20365 135
rect 20365 115 20385 135
rect 20385 115 20390 135
rect 20360 110 20390 115
rect 17960 -15 17990 -10
rect 17960 -35 17965 -15
rect 17965 -35 17985 -15
rect 17985 -35 17990 -15
rect 17960 -40 17990 -35
rect 15560 -165 15590 -160
rect 15560 -185 15565 -165
rect 15565 -185 15585 -165
rect 15585 -185 15590 -165
rect 15560 -190 15590 -185
rect 15560 -265 15590 -260
rect 15560 -285 15565 -265
rect 15565 -285 15585 -265
rect 15585 -285 15590 -265
rect 15560 -290 15590 -285
rect 15560 -365 15590 -360
rect 15560 -385 15565 -365
rect 15565 -385 15585 -365
rect 15585 -385 15590 -365
rect 15560 -390 15590 -385
rect 15560 -465 15590 -460
rect 15560 -485 15565 -465
rect 15565 -485 15585 -465
rect 15585 -485 15590 -465
rect 15560 -490 15590 -485
rect 15560 -565 15590 -560
rect 15560 -585 15565 -565
rect 15565 -585 15585 -565
rect 15585 -585 15590 -565
rect 15560 -590 15590 -585
rect 15560 -665 15590 -660
rect 15560 -685 15565 -665
rect 15565 -685 15585 -665
rect 15585 -685 15590 -665
rect 15560 -690 15590 -685
rect 15560 -765 15590 -760
rect 15560 -785 15565 -765
rect 15565 -785 15585 -765
rect 15585 -785 15590 -765
rect 15560 -790 15590 -785
rect 14510 -865 14540 -860
rect 14510 -885 14515 -865
rect 14515 -885 14535 -865
rect 14535 -885 14540 -865
rect 14510 -890 14540 -885
rect 14810 -865 14840 -860
rect 14810 -885 14815 -865
rect 14815 -885 14835 -865
rect 14835 -885 14840 -865
rect 14810 -890 14840 -885
rect 15110 -865 15140 -860
rect 15110 -885 15115 -865
rect 15115 -885 15135 -865
rect 15135 -885 15140 -865
rect 15110 -890 15140 -885
rect 15410 -865 15440 -860
rect 15410 -885 15415 -865
rect 15415 -885 15435 -865
rect 15435 -885 15440 -865
rect 15410 -890 15440 -885
rect 15710 -865 15740 -860
rect 15710 -885 15715 -865
rect 15715 -885 15735 -865
rect 15735 -885 15740 -865
rect 15710 -890 15740 -885
rect 16010 -865 16040 -860
rect 16010 -885 16015 -865
rect 16015 -885 16035 -865
rect 16035 -885 16040 -865
rect 16010 -890 16040 -885
rect 16310 -865 16340 -860
rect 16310 -885 16315 -865
rect 16315 -885 16335 -865
rect 16335 -885 16340 -865
rect 16310 -890 16340 -885
rect 16610 -865 16640 -860
rect 16610 -885 16615 -865
rect 16615 -885 16635 -865
rect 16635 -885 16640 -865
rect 16610 -890 16640 -885
rect 20360 -15 20390 -10
rect 20360 -35 20365 -15
rect 20365 -35 20385 -15
rect 20385 -35 20390 -15
rect 20360 -40 20390 -35
rect 17960 -165 17990 -160
rect 17960 -185 17965 -165
rect 17965 -185 17985 -165
rect 17985 -185 17990 -165
rect 17960 -190 17990 -185
rect 17960 -265 17990 -260
rect 17960 -285 17965 -265
rect 17965 -285 17985 -265
rect 17985 -285 17990 -265
rect 17960 -290 17990 -285
rect 17960 -365 17990 -360
rect 17960 -385 17965 -365
rect 17965 -385 17985 -365
rect 17985 -385 17990 -365
rect 17960 -390 17990 -385
rect 17960 -465 17990 -460
rect 17960 -485 17965 -465
rect 17965 -485 17985 -465
rect 17985 -485 17990 -465
rect 17960 -490 17990 -485
rect 17960 -565 17990 -560
rect 17960 -585 17965 -565
rect 17965 -585 17985 -565
rect 17985 -585 17990 -565
rect 17960 -590 17990 -585
rect 17960 -665 17990 -660
rect 17960 -685 17965 -665
rect 17965 -685 17985 -665
rect 17985 -685 17990 -665
rect 17960 -690 17990 -685
rect 17960 -765 17990 -760
rect 17960 -785 17965 -765
rect 17965 -785 17985 -765
rect 17985 -785 17990 -765
rect 17960 -790 17990 -785
rect 16760 -890 16790 -860
rect 15560 -965 15590 -960
rect 15560 -985 15565 -965
rect 15565 -985 15585 -965
rect 15585 -985 15590 -965
rect 15560 -990 15590 -985
rect 15560 -1065 15590 -1060
rect 15560 -1085 15565 -1065
rect 15565 -1085 15585 -1065
rect 15585 -1085 15590 -1065
rect 15560 -1090 15590 -1085
rect 15560 -1165 15590 -1160
rect 15560 -1185 15565 -1165
rect 15565 -1185 15585 -1165
rect 15585 -1185 15590 -1165
rect 15560 -1190 15590 -1185
rect 15560 -1265 15590 -1260
rect 15560 -1285 15565 -1265
rect 15565 -1285 15585 -1265
rect 15585 -1285 15590 -1265
rect 15560 -1290 15590 -1285
rect 15560 -1365 15590 -1360
rect 15560 -1385 15565 -1365
rect 15565 -1385 15585 -1365
rect 15585 -1385 15590 -1365
rect 15560 -1390 15590 -1385
rect 15560 -1465 15590 -1460
rect 15560 -1485 15565 -1465
rect 15565 -1485 15585 -1465
rect 15585 -1485 15590 -1465
rect 15560 -1490 15590 -1485
rect 15560 -1565 15590 -1560
rect 15560 -1585 15565 -1565
rect 15565 -1585 15585 -1565
rect 15585 -1585 15590 -1565
rect 15560 -1590 15590 -1585
rect 10760 -1715 10790 -1710
rect 10760 -1735 10765 -1715
rect 10765 -1735 10785 -1715
rect 10785 -1735 10790 -1715
rect 10760 -1740 10790 -1735
rect 16910 -865 16940 -860
rect 16910 -885 16915 -865
rect 16915 -885 16935 -865
rect 16935 -885 16940 -865
rect 16910 -890 16940 -885
rect 17210 -865 17240 -860
rect 17210 -885 17215 -865
rect 17215 -885 17235 -865
rect 17235 -885 17240 -865
rect 17210 -890 17240 -885
rect 17510 -865 17540 -860
rect 17510 -885 17515 -865
rect 17515 -885 17535 -865
rect 17535 -885 17540 -865
rect 17510 -890 17540 -885
rect 17810 -865 17840 -860
rect 17810 -885 17815 -865
rect 17815 -885 17835 -865
rect 17835 -885 17840 -865
rect 17810 -890 17840 -885
rect 18110 -865 18140 -860
rect 18110 -885 18115 -865
rect 18115 -885 18135 -865
rect 18135 -885 18140 -865
rect 18110 -890 18140 -885
rect 18410 -865 18440 -860
rect 18410 -885 18415 -865
rect 18415 -885 18435 -865
rect 18435 -885 18440 -865
rect 18410 -890 18440 -885
rect 18710 -865 18740 -860
rect 18710 -885 18715 -865
rect 18715 -885 18735 -865
rect 18735 -885 18740 -865
rect 18710 -890 18740 -885
rect 19010 -865 19040 -860
rect 19010 -885 19015 -865
rect 19015 -885 19035 -865
rect 19035 -885 19040 -865
rect 19010 -890 19040 -885
rect 20360 -165 20390 -160
rect 20360 -185 20365 -165
rect 20365 -185 20385 -165
rect 20385 -185 20390 -165
rect 20360 -190 20390 -185
rect 20360 -265 20390 -260
rect 20360 -285 20365 -265
rect 20365 -285 20385 -265
rect 20385 -285 20390 -265
rect 20360 -290 20390 -285
rect 20360 -365 20390 -360
rect 20360 -385 20365 -365
rect 20365 -385 20385 -365
rect 20385 -385 20390 -365
rect 20360 -390 20390 -385
rect 20360 -465 20390 -460
rect 20360 -485 20365 -465
rect 20365 -485 20385 -465
rect 20385 -485 20390 -465
rect 20360 -490 20390 -485
rect 20360 -565 20390 -560
rect 20360 -585 20365 -565
rect 20365 -585 20385 -565
rect 20385 -585 20390 -565
rect 20360 -590 20390 -585
rect 20360 -665 20390 -660
rect 20360 -685 20365 -665
rect 20365 -685 20385 -665
rect 20385 -685 20390 -665
rect 20360 -690 20390 -685
rect 20360 -765 20390 -760
rect 20360 -785 20365 -765
rect 20365 -785 20385 -765
rect 20385 -785 20390 -765
rect 20360 -790 20390 -785
rect 19160 -890 19190 -860
rect 17960 -965 17990 -960
rect 17960 -985 17965 -965
rect 17965 -985 17985 -965
rect 17985 -985 17990 -965
rect 17960 -990 17990 -985
rect 17960 -1065 17990 -1060
rect 17960 -1085 17965 -1065
rect 17965 -1085 17985 -1065
rect 17985 -1085 17990 -1065
rect 17960 -1090 17990 -1085
rect 17960 -1165 17990 -1160
rect 17960 -1185 17965 -1165
rect 17965 -1185 17985 -1165
rect 17985 -1185 17990 -1165
rect 17960 -1190 17990 -1185
rect 17960 -1265 17990 -1260
rect 17960 -1285 17965 -1265
rect 17965 -1285 17985 -1265
rect 17985 -1285 17990 -1265
rect 17960 -1290 17990 -1285
rect 17960 -1365 17990 -1360
rect 17960 -1385 17965 -1365
rect 17965 -1385 17985 -1365
rect 17985 -1385 17990 -1365
rect 17960 -1390 17990 -1385
rect 17960 -1465 17990 -1460
rect 17960 -1485 17965 -1465
rect 17965 -1485 17985 -1465
rect 17985 -1485 17990 -1465
rect 17960 -1490 17990 -1485
rect 17960 -1565 17990 -1560
rect 17960 -1585 17965 -1565
rect 17965 -1585 17985 -1565
rect 17985 -1585 17990 -1565
rect 17960 -1590 17990 -1585
rect 15560 -1715 15590 -1710
rect 15560 -1735 15565 -1715
rect 15565 -1735 15585 -1715
rect 15585 -1735 15590 -1715
rect 15560 -1740 15590 -1735
rect 19310 -865 19340 -860
rect 19310 -885 19315 -865
rect 19315 -885 19335 -865
rect 19335 -885 19340 -865
rect 19310 -890 19340 -885
rect 19610 -865 19640 -860
rect 19610 -885 19615 -865
rect 19615 -885 19635 -865
rect 19635 -885 19640 -865
rect 19610 -890 19640 -885
rect 19910 -865 19940 -860
rect 19910 -885 19915 -865
rect 19915 -885 19935 -865
rect 19935 -885 19940 -865
rect 19910 -890 19940 -885
rect 20210 -865 20240 -860
rect 20210 -885 20215 -865
rect 20215 -885 20235 -865
rect 20235 -885 20240 -865
rect 20210 -890 20240 -885
rect 20360 -965 20390 -960
rect 20360 -985 20365 -965
rect 20365 -985 20385 -965
rect 20385 -985 20390 -965
rect 20360 -990 20390 -985
rect 20360 -1065 20390 -1060
rect 20360 -1085 20365 -1065
rect 20365 -1085 20385 -1065
rect 20385 -1085 20390 -1065
rect 20360 -1090 20390 -1085
rect 20360 -1165 20390 -1160
rect 20360 -1185 20365 -1165
rect 20365 -1185 20385 -1165
rect 20385 -1185 20390 -1165
rect 20360 -1190 20390 -1185
rect 20360 -1265 20390 -1260
rect 20360 -1285 20365 -1265
rect 20365 -1285 20385 -1265
rect 20385 -1285 20390 -1265
rect 20360 -1290 20390 -1285
rect 20360 -1365 20390 -1360
rect 20360 -1385 20365 -1365
rect 20365 -1385 20385 -1365
rect 20385 -1385 20390 -1365
rect 20360 -1390 20390 -1385
rect 20360 -1465 20390 -1460
rect 20360 -1485 20365 -1465
rect 20365 -1485 20385 -1465
rect 20385 -1485 20390 -1465
rect 20360 -1490 20390 -1485
rect 20360 -1565 20390 -1560
rect 20360 -1585 20365 -1565
rect 20365 -1585 20385 -1565
rect 20385 -1585 20390 -1565
rect 20360 -1590 20390 -1585
rect 17960 -1715 17990 -1710
rect 17960 -1735 17965 -1715
rect 17965 -1735 17985 -1715
rect 17985 -1735 17990 -1715
rect 17960 -1740 17990 -1735
rect 20360 -1715 20390 -1710
rect 20360 -1735 20365 -1715
rect 20365 -1735 20385 -1715
rect 20385 -1735 20390 -1715
rect 20360 -1740 20390 -1735
<< metal2 >>
rect -650 5190 20400 5200
rect -650 5160 -640 5190
rect -610 5160 -40 5190
rect -10 5160 4160 5190
rect 4190 5160 8360 5190
rect 8390 5160 8660 5190
rect 8690 5160 8960 5190
rect 8990 5160 9260 5190
rect 9290 5160 9560 5190
rect 9590 5160 9860 5190
rect 9890 5160 10160 5190
rect 10190 5160 10460 5190
rect 10490 5160 10760 5190
rect 10790 5160 11960 5190
rect 11990 5160 13160 5190
rect 13190 5160 14360 5190
rect 14390 5160 15560 5190
rect 15590 5160 17960 5190
rect 17990 5160 20360 5190
rect 20390 5160 20400 5190
rect -650 5100 20400 5160
rect -650 5040 20400 5050
rect -650 5010 -640 5040
rect -610 5010 8360 5040
rect 8390 5010 8660 5040
rect 8690 5010 8960 5040
rect 8990 5010 9260 5040
rect 9290 5010 9560 5040
rect 9590 5010 9860 5040
rect 9890 5010 10160 5040
rect 10190 5010 10460 5040
rect 10490 5010 10760 5040
rect 10790 5010 11960 5040
rect 11990 5010 13160 5040
rect 13190 5010 14360 5040
rect 14390 5010 15560 5040
rect 15590 5010 20360 5040
rect 20390 5010 20400 5040
rect -650 5000 20400 5010
rect -650 4940 20400 4950
rect -650 4910 -640 4940
rect -610 4910 8360 4940
rect 8390 4910 8660 4940
rect 8690 4910 8960 4940
rect 8990 4910 9260 4940
rect 9290 4910 9560 4940
rect 9590 4910 9860 4940
rect 9890 4910 10160 4940
rect 10190 4910 10460 4940
rect 10490 4910 10760 4940
rect 10790 4910 11960 4940
rect 11990 4910 13160 4940
rect 13190 4910 14360 4940
rect 14390 4910 15560 4940
rect 15590 4910 17960 4940
rect 17990 4910 20360 4940
rect 20390 4910 20400 4940
rect -650 4900 20400 4910
rect -650 4840 20400 4850
rect -650 4810 -640 4840
rect -610 4810 8360 4840
rect 8390 4810 8660 4840
rect 8690 4810 8960 4840
rect 8990 4810 9260 4840
rect 9290 4810 9560 4840
rect 9590 4810 9860 4840
rect 9890 4810 10160 4840
rect 10190 4810 10460 4840
rect 10490 4810 10760 4840
rect 10790 4810 11960 4840
rect 11990 4810 13160 4840
rect 13190 4810 14360 4840
rect 14390 4810 15560 4840
rect 15590 4810 17960 4840
rect 17990 4810 20360 4840
rect 20390 4810 20400 4840
rect -650 4800 20400 4810
rect -650 4740 20400 4750
rect -650 4710 -640 4740
rect -610 4710 8360 4740
rect 8390 4710 8660 4740
rect 8690 4710 8960 4740
rect 8990 4710 9260 4740
rect 9290 4710 9560 4740
rect 9590 4710 9860 4740
rect 9890 4710 10160 4740
rect 10190 4710 10460 4740
rect 10490 4710 10760 4740
rect 10790 4710 11960 4740
rect 11990 4710 13160 4740
rect 13190 4710 14360 4740
rect 14390 4710 15560 4740
rect 15590 4710 17960 4740
rect 17990 4710 20360 4740
rect 20390 4710 20400 4740
rect -650 4700 20400 4710
rect -650 4640 20400 4650
rect -650 4610 -640 4640
rect -610 4610 8360 4640
rect 8390 4610 8660 4640
rect 8690 4610 8960 4640
rect 8990 4610 9260 4640
rect 9290 4610 9560 4640
rect 9590 4610 9860 4640
rect 9890 4610 10160 4640
rect 10190 4610 10460 4640
rect 10490 4610 10760 4640
rect 10790 4610 11960 4640
rect 11990 4610 13160 4640
rect 13190 4610 14360 4640
rect 14390 4610 15560 4640
rect 15590 4610 17960 4640
rect 17990 4610 20360 4640
rect 20390 4610 20400 4640
rect -650 4600 20400 4610
rect -500 4540 -450 4550
rect -500 4510 -490 4540
rect -460 4510 -450 4540
rect -500 4500 -450 4510
rect -350 4540 -300 4550
rect -350 4510 -340 4540
rect -310 4510 -300 4540
rect -350 4500 -300 4510
rect -200 4540 -150 4550
rect -200 4510 -190 4540
rect -160 4510 -150 4540
rect -200 4500 -150 4510
rect 100 4540 150 4550
rect 100 4510 110 4540
rect 140 4510 150 4540
rect 100 4500 150 4510
rect 400 4540 450 4550
rect 400 4510 410 4540
rect 440 4510 450 4540
rect 400 4500 450 4510
rect 700 4540 750 4550
rect 700 4510 710 4540
rect 740 4510 750 4540
rect 700 4500 750 4510
rect 1000 4540 1050 4550
rect 1000 4510 1010 4540
rect 1040 4510 1050 4540
rect 1000 4500 1050 4510
rect 1150 4540 1200 4550
rect 1150 4510 1160 4540
rect 1190 4510 1200 4540
rect 1150 4500 1200 4510
rect 1300 4540 1350 4550
rect 1300 4510 1310 4540
rect 1340 4510 1350 4540
rect 1300 4500 1350 4510
rect 1600 4540 1650 4550
rect 1600 4510 1610 4540
rect 1640 4510 1650 4540
rect 1600 4500 1650 4510
rect 1900 4540 1950 4550
rect 1900 4510 1910 4540
rect 1940 4510 1950 4540
rect 1900 4500 1950 4510
rect 2050 4540 2100 4550
rect 2050 4510 2060 4540
rect 2090 4510 2100 4540
rect 2050 4500 2100 4510
rect 2200 4540 2250 4550
rect 2200 4510 2210 4540
rect 2240 4510 2250 4540
rect 2200 4500 2250 4510
rect 2500 4540 2550 4550
rect 2500 4510 2510 4540
rect 2540 4510 2550 4540
rect 2500 4500 2550 4510
rect 2800 4540 2850 4550
rect 2800 4510 2810 4540
rect 2840 4510 2850 4540
rect 2800 4500 2850 4510
rect 2950 4540 3000 4550
rect 2950 4510 2960 4540
rect 2990 4510 3000 4540
rect 2950 4500 3000 4510
rect 3100 4540 3150 4550
rect 3100 4510 3110 4540
rect 3140 4510 3150 4540
rect 3100 4500 3150 4510
rect 3400 4540 3450 4550
rect 3400 4510 3410 4540
rect 3440 4510 3450 4540
rect 3400 4500 3450 4510
rect 3700 4540 3750 4550
rect 3700 4510 3710 4540
rect 3740 4510 3750 4540
rect 3700 4500 3750 4510
rect 4000 4540 4050 4550
rect 4000 4510 4010 4540
rect 4040 4510 4050 4540
rect 4000 4500 4050 4510
rect 4300 4540 4350 4550
rect 4300 4510 4310 4540
rect 4340 4510 4350 4540
rect 4300 4500 4350 4510
rect 4600 4540 4650 4550
rect 4600 4510 4610 4540
rect 4640 4510 4650 4540
rect 4600 4500 4650 4510
rect 4900 4540 4950 4550
rect 4900 4510 4910 4540
rect 4940 4510 4950 4540
rect 4900 4500 4950 4510
rect 5200 4540 5250 4550
rect 5200 4510 5210 4540
rect 5240 4510 5250 4540
rect 5200 4500 5250 4510
rect 5350 4540 5400 4550
rect 5350 4510 5360 4540
rect 5390 4510 5400 4540
rect 5350 4500 5400 4510
rect 5500 4540 5550 4550
rect 5500 4510 5510 4540
rect 5540 4510 5550 4540
rect 5500 4500 5550 4510
rect 5800 4540 5850 4550
rect 5800 4510 5810 4540
rect 5840 4510 5850 4540
rect 5800 4500 5850 4510
rect 6100 4540 6150 4550
rect 6100 4510 6110 4540
rect 6140 4510 6150 4540
rect 6100 4500 6150 4510
rect 6250 4540 6300 4550
rect 6250 4510 6260 4540
rect 6290 4510 6300 4540
rect 6250 4500 6300 4510
rect 6400 4540 6450 4550
rect 6400 4510 6410 4540
rect 6440 4510 6450 4540
rect 6400 4500 6450 4510
rect 6700 4540 6750 4550
rect 6700 4510 6710 4540
rect 6740 4510 6750 4540
rect 6700 4500 6750 4510
rect 7000 4540 7050 4550
rect 7000 4510 7010 4540
rect 7040 4510 7050 4540
rect 7000 4500 7050 4510
rect 7150 4540 7200 4550
rect 7150 4510 7160 4540
rect 7190 4510 7200 4540
rect 7150 4500 7200 4510
rect 7300 4540 7350 4550
rect 7300 4510 7310 4540
rect 7340 4510 7350 4540
rect 7300 4500 7350 4510
rect 7600 4540 7650 4550
rect 7600 4510 7610 4540
rect 7640 4510 7650 4540
rect 7600 4500 7650 4510
rect 7900 4540 7950 4550
rect 7900 4510 7910 4540
rect 7940 4510 7950 4540
rect 7900 4500 7950 4510
rect 8200 4540 8250 4550
rect 8200 4510 8210 4540
rect 8240 4510 8250 4540
rect 8200 4500 8250 4510
rect 8500 4540 8550 4550
rect 8500 4510 8510 4540
rect 8540 4510 8550 4540
rect 8500 4500 8550 4510
rect 8800 4540 8850 4550
rect 8800 4510 8810 4540
rect 8840 4510 8850 4540
rect 8800 4500 8850 4510
rect 9100 4540 9150 4550
rect 9100 4510 9110 4540
rect 9140 4510 9150 4540
rect 9100 4500 9150 4510
rect 9400 4540 9450 4550
rect 9400 4510 9410 4540
rect 9440 4510 9450 4540
rect 9400 4500 9450 4510
rect 9700 4540 9750 4550
rect 9700 4510 9710 4540
rect 9740 4510 9750 4540
rect 9700 4500 9750 4510
rect 10000 4540 10050 4550
rect 10000 4510 10010 4540
rect 10040 4510 10050 4540
rect 10000 4500 10050 4510
rect 10300 4540 10350 4550
rect 10300 4510 10310 4540
rect 10340 4510 10350 4540
rect 10300 4500 10350 4510
rect 10600 4540 10650 4550
rect 10600 4510 10610 4540
rect 10640 4510 10650 4540
rect 10600 4500 10650 4510
rect 10900 4540 10950 4550
rect 10900 4510 10910 4540
rect 10940 4510 10950 4540
rect 10900 4500 10950 4510
rect 11200 4540 11250 4550
rect 11200 4510 11210 4540
rect 11240 4510 11250 4540
rect 11200 4500 11250 4510
rect 11350 4540 11400 4550
rect 11350 4510 11360 4540
rect 11390 4510 11400 4540
rect 11350 4500 11400 4510
rect 11500 4540 11550 4550
rect 11500 4510 11510 4540
rect 11540 4510 11550 4540
rect 11500 4500 11550 4510
rect 11800 4540 11850 4550
rect 11800 4510 11810 4540
rect 11840 4510 11850 4540
rect 11800 4500 11850 4510
rect 12100 4540 12150 4550
rect 12100 4510 12110 4540
rect 12140 4510 12150 4540
rect 12100 4500 12150 4510
rect 12400 4540 12450 4550
rect 12400 4510 12410 4540
rect 12440 4510 12450 4540
rect 12400 4500 12450 4510
rect 12550 4540 12600 4550
rect 12550 4510 12560 4540
rect 12590 4510 12600 4540
rect 12550 4500 12600 4510
rect 12700 4540 12750 4550
rect 12700 4510 12710 4540
rect 12740 4510 12750 4540
rect 12700 4500 12750 4510
rect 13000 4540 13050 4550
rect 13000 4510 13010 4540
rect 13040 4510 13050 4540
rect 13000 4500 13050 4510
rect 13300 4540 13350 4550
rect 13300 4510 13310 4540
rect 13340 4510 13350 4540
rect 13300 4500 13350 4510
rect 13600 4540 13650 4550
rect 13600 4510 13610 4540
rect 13640 4510 13650 4540
rect 13600 4500 13650 4510
rect 13750 4540 13800 4550
rect 13750 4510 13760 4540
rect 13790 4510 13800 4540
rect 13750 4500 13800 4510
rect 13900 4540 13950 4550
rect 13900 4510 13910 4540
rect 13940 4510 13950 4540
rect 13900 4500 13950 4510
rect 14200 4540 14250 4550
rect 14200 4510 14210 4540
rect 14240 4510 14250 4540
rect 14200 4500 14250 4510
rect 14500 4540 14550 4550
rect 14500 4510 14510 4540
rect 14540 4510 14550 4540
rect 14500 4500 14550 4510
rect 14800 4540 14850 4550
rect 14800 4510 14810 4540
rect 14840 4510 14850 4540
rect 14800 4500 14850 4510
rect 14950 4540 15000 4550
rect 14950 4510 14960 4540
rect 14990 4510 15000 4540
rect 14950 4500 15000 4510
rect 15100 4540 15150 4550
rect 15100 4510 15110 4540
rect 15140 4510 15150 4540
rect 15100 4500 15150 4510
rect 15400 4540 15450 4550
rect 15400 4510 15410 4540
rect 15440 4510 15450 4540
rect 15400 4500 15450 4510
rect 15700 4540 15750 4550
rect 15700 4510 15710 4540
rect 15740 4510 15750 4540
rect 15700 4500 15750 4510
rect 16000 4540 16050 4550
rect 16000 4510 16010 4540
rect 16040 4510 16050 4540
rect 16000 4500 16050 4510
rect 16300 4540 16350 4550
rect 16300 4510 16310 4540
rect 16340 4510 16350 4540
rect 16300 4500 16350 4510
rect 16600 4540 16650 4550
rect 16600 4510 16610 4540
rect 16640 4510 16650 4540
rect 16600 4500 16650 4510
rect 16750 4540 16800 4550
rect 16750 4510 16760 4540
rect 16790 4510 16800 4540
rect 16750 4500 16800 4510
rect 16900 4540 16950 4550
rect 16900 4510 16910 4540
rect 16940 4510 16950 4540
rect 16900 4500 16950 4510
rect 17200 4540 17250 4550
rect 17200 4510 17210 4540
rect 17240 4510 17250 4540
rect 17200 4500 17250 4510
rect 17500 4540 17550 4550
rect 17500 4510 17510 4540
rect 17540 4510 17550 4540
rect 17500 4500 17550 4510
rect 17800 4540 17850 4550
rect 17800 4510 17810 4540
rect 17840 4510 17850 4540
rect 17800 4500 17850 4510
rect 18100 4540 18150 4550
rect 18100 4510 18110 4540
rect 18140 4510 18150 4540
rect 18100 4500 18150 4510
rect 18400 4540 18450 4550
rect 18400 4510 18410 4540
rect 18440 4510 18450 4540
rect 18400 4500 18450 4510
rect 18700 4540 18750 4550
rect 18700 4510 18710 4540
rect 18740 4510 18750 4540
rect 18700 4500 18750 4510
rect 19000 4540 19050 4550
rect 19000 4510 19010 4540
rect 19040 4510 19050 4540
rect 19000 4500 19050 4510
rect 19150 4540 19200 4550
rect 19150 4510 19160 4540
rect 19190 4510 19200 4540
rect 19150 4500 19200 4510
rect 19300 4540 19350 4550
rect 19300 4510 19310 4540
rect 19340 4510 19350 4540
rect 19300 4500 19350 4510
rect 19600 4540 19650 4550
rect 19600 4510 19610 4540
rect 19640 4510 19650 4540
rect 19600 4500 19650 4510
rect 19900 4540 19950 4550
rect 19900 4510 19910 4540
rect 19940 4510 19950 4540
rect 19900 4500 19950 4510
rect 20200 4540 20250 4550
rect 20200 4510 20210 4540
rect 20240 4510 20250 4540
rect 20200 4500 20250 4510
rect -650 4440 20400 4450
rect -650 4410 -640 4440
rect -610 4410 -40 4440
rect -10 4410 4160 4440
rect 4190 4410 8360 4440
rect 8390 4410 8660 4440
rect 8690 4410 8960 4440
rect 8990 4410 9260 4440
rect 9290 4410 9560 4440
rect 9590 4410 9860 4440
rect 9890 4410 10160 4440
rect 10190 4410 10460 4440
rect 10490 4410 10760 4440
rect 10790 4410 11960 4440
rect 11990 4410 13160 4440
rect 13190 4410 14360 4440
rect 14390 4410 15560 4440
rect 15590 4410 17960 4440
rect 17990 4410 20360 4440
rect 20390 4410 20400 4440
rect -650 4400 20400 4410
rect -650 4340 20400 4350
rect -650 4310 -640 4340
rect -610 4310 -40 4340
rect -10 4310 4160 4340
rect 4190 4310 8360 4340
rect 8390 4310 8660 4340
rect 8690 4310 8960 4340
rect 8990 4310 9260 4340
rect 9290 4310 9560 4340
rect 9590 4310 9860 4340
rect 9890 4310 10160 4340
rect 10190 4310 10460 4340
rect 10490 4310 10760 4340
rect 10790 4310 11960 4340
rect 11990 4310 13160 4340
rect 13190 4310 14360 4340
rect 14390 4310 15560 4340
rect 15590 4310 17960 4340
rect 17990 4310 20360 4340
rect 20390 4310 20400 4340
rect -650 4300 20400 4310
rect -650 4240 20400 4250
rect -650 4210 -640 4240
rect -610 4210 -40 4240
rect -10 4210 4160 4240
rect 4190 4210 8360 4240
rect 8390 4210 8660 4240
rect 8690 4210 8960 4240
rect 8990 4210 9260 4240
rect 9290 4210 9560 4240
rect 9590 4210 9860 4240
rect 9890 4210 10160 4240
rect 10190 4210 10460 4240
rect 10490 4210 10760 4240
rect 10790 4210 11960 4240
rect 11990 4210 13160 4240
rect 13190 4210 14360 4240
rect 14390 4210 15560 4240
rect 15590 4210 17960 4240
rect 17990 4210 20360 4240
rect 20390 4210 20400 4240
rect -650 4200 20400 4210
rect -650 4140 20400 4150
rect -650 4110 -640 4140
rect -610 4110 -40 4140
rect -10 4110 4160 4140
rect 4190 4110 8360 4140
rect 8390 4110 8660 4140
rect 8690 4110 8960 4140
rect 8990 4110 9260 4140
rect 9290 4110 9560 4140
rect 9590 4110 9860 4140
rect 9890 4110 10160 4140
rect 10190 4110 10460 4140
rect 10490 4110 10760 4140
rect 10790 4110 11960 4140
rect 11990 4110 13160 4140
rect 13190 4110 14360 4140
rect 14390 4110 15560 4140
rect 15590 4110 17960 4140
rect 17990 4110 20360 4140
rect 20390 4110 20400 4140
rect -650 4100 20400 4110
rect -650 4040 20400 4050
rect -650 4010 -640 4040
rect -610 4010 -40 4040
rect -10 4010 4160 4040
rect 4190 4010 8360 4040
rect 8390 4010 8660 4040
rect 8690 4010 8960 4040
rect 8990 4010 9260 4040
rect 9290 4010 9560 4040
rect 9590 4010 9860 4040
rect 9890 4010 10160 4040
rect 10190 4010 10460 4040
rect 10490 4010 10760 4040
rect 10790 4010 11960 4040
rect 11990 4010 13160 4040
rect 13190 4010 14360 4040
rect 14390 4010 15560 4040
rect 15590 4010 20360 4040
rect 20390 4010 20400 4040
rect -650 4000 20400 4010
rect -650 3890 20400 3950
rect -650 3860 -640 3890
rect -610 3860 -40 3890
rect -10 3860 4160 3890
rect 4190 3860 8360 3890
rect 8390 3860 8660 3890
rect 8690 3860 8960 3890
rect 8990 3860 9260 3890
rect 9290 3860 9560 3890
rect 9590 3860 9860 3890
rect 9890 3860 10160 3890
rect 10190 3860 10460 3890
rect 10490 3860 10760 3890
rect 10790 3860 11960 3890
rect 11990 3860 13160 3890
rect 13190 3860 14360 3890
rect 14390 3860 15560 3890
rect 15590 3860 20360 3890
rect 20390 3860 20400 3890
rect -650 3800 20400 3860
rect -650 3740 20400 3750
rect -650 3710 -640 3740
rect -610 3710 8360 3740
rect 8390 3710 8660 3740
rect 8690 3710 8960 3740
rect 8990 3710 9260 3740
rect 9290 3710 9560 3740
rect 9590 3710 9860 3740
rect 9890 3710 10160 3740
rect 10190 3710 10460 3740
rect 10490 3710 10760 3740
rect 10790 3710 11960 3740
rect 11990 3710 13160 3740
rect 13190 3710 14360 3740
rect 14390 3710 15560 3740
rect 15590 3710 20360 3740
rect 20390 3710 20400 3740
rect -650 3700 20400 3710
rect -650 3640 20400 3650
rect -650 3610 -640 3640
rect -610 3610 8360 3640
rect 8390 3610 8660 3640
rect 8690 3610 8960 3640
rect 8990 3610 9260 3640
rect 9290 3610 9560 3640
rect 9590 3610 9860 3640
rect 9890 3610 10160 3640
rect 10190 3610 10460 3640
rect 10490 3610 10760 3640
rect 10790 3610 11960 3640
rect 11990 3610 13160 3640
rect 13190 3610 14360 3640
rect 14390 3610 15560 3640
rect 15590 3610 17960 3640
rect 17990 3610 20360 3640
rect 20390 3610 20400 3640
rect -650 3600 20400 3610
rect -650 3540 20400 3550
rect -650 3510 -640 3540
rect -610 3510 8360 3540
rect 8390 3510 8660 3540
rect 8690 3510 8960 3540
rect 8990 3510 9260 3540
rect 9290 3510 9560 3540
rect 9590 3510 9860 3540
rect 9890 3510 10160 3540
rect 10190 3510 10460 3540
rect 10490 3510 10760 3540
rect 10790 3510 11960 3540
rect 11990 3510 13160 3540
rect 13190 3510 14360 3540
rect 14390 3510 15560 3540
rect 15590 3510 17960 3540
rect 17990 3510 20360 3540
rect 20390 3510 20400 3540
rect -650 3500 20400 3510
rect -650 3440 20400 3450
rect -650 3410 -640 3440
rect -610 3410 8360 3440
rect 8390 3410 8660 3440
rect 8690 3410 8960 3440
rect 8990 3410 9260 3440
rect 9290 3410 9560 3440
rect 9590 3410 9860 3440
rect 9890 3410 10160 3440
rect 10190 3410 10460 3440
rect 10490 3410 10760 3440
rect 10790 3410 11960 3440
rect 11990 3410 13160 3440
rect 13190 3410 14360 3440
rect 14390 3410 15560 3440
rect 15590 3410 17960 3440
rect 17990 3410 20360 3440
rect 20390 3410 20400 3440
rect -650 3400 20400 3410
rect -650 3340 20400 3350
rect -650 3310 -640 3340
rect -610 3310 8360 3340
rect 8390 3310 8660 3340
rect 8690 3310 8960 3340
rect 8990 3310 9260 3340
rect 9290 3310 9560 3340
rect 9590 3310 9860 3340
rect 9890 3310 10160 3340
rect 10190 3310 10460 3340
rect 10490 3310 10760 3340
rect 10790 3310 11960 3340
rect 11990 3310 13160 3340
rect 13190 3310 14360 3340
rect 14390 3310 15560 3340
rect 15590 3310 17960 3340
rect 17990 3310 20360 3340
rect 20390 3310 20400 3340
rect -650 3300 20400 3310
rect -500 3240 -450 3250
rect -500 3210 -490 3240
rect -460 3210 -450 3240
rect -500 3200 -450 3210
rect -350 3240 -300 3250
rect -350 3210 -340 3240
rect -310 3210 -300 3240
rect -350 3200 -300 3210
rect -200 3240 -150 3250
rect -200 3210 -190 3240
rect -160 3210 -150 3240
rect -200 3200 -150 3210
rect 100 3240 150 3250
rect 100 3210 110 3240
rect 140 3210 150 3240
rect 100 3200 150 3210
rect 400 3240 450 3250
rect 400 3210 410 3240
rect 440 3210 450 3240
rect 400 3200 450 3210
rect 700 3240 750 3250
rect 700 3210 710 3240
rect 740 3210 750 3240
rect 700 3200 750 3210
rect 1000 3240 1050 3250
rect 1000 3210 1010 3240
rect 1040 3210 1050 3240
rect 1000 3200 1050 3210
rect 1150 3240 1200 3250
rect 1150 3210 1160 3240
rect 1190 3210 1200 3240
rect 1150 3200 1200 3210
rect 1300 3240 1350 3250
rect 1300 3210 1310 3240
rect 1340 3210 1350 3240
rect 1300 3200 1350 3210
rect 1600 3240 1650 3250
rect 1600 3210 1610 3240
rect 1640 3210 1650 3240
rect 1600 3200 1650 3210
rect 1900 3240 1950 3250
rect 1900 3210 1910 3240
rect 1940 3210 1950 3240
rect 1900 3200 1950 3210
rect 2050 3240 2100 3250
rect 2050 3210 2060 3240
rect 2090 3210 2100 3240
rect 2050 3200 2100 3210
rect 2200 3240 2250 3250
rect 2200 3210 2210 3240
rect 2240 3210 2250 3240
rect 2200 3200 2250 3210
rect 2500 3240 2550 3250
rect 2500 3210 2510 3240
rect 2540 3210 2550 3240
rect 2500 3200 2550 3210
rect 2800 3240 2850 3250
rect 2800 3210 2810 3240
rect 2840 3210 2850 3240
rect 2800 3200 2850 3210
rect 2950 3240 3000 3250
rect 2950 3210 2960 3240
rect 2990 3210 3000 3240
rect 2950 3200 3000 3210
rect 3100 3240 3150 3250
rect 3100 3210 3110 3240
rect 3140 3210 3150 3240
rect 3100 3200 3150 3210
rect 3400 3240 3450 3250
rect 3400 3210 3410 3240
rect 3440 3210 3450 3240
rect 3400 3200 3450 3210
rect 3700 3240 3750 3250
rect 3700 3210 3710 3240
rect 3740 3210 3750 3240
rect 3700 3200 3750 3210
rect 4000 3240 4050 3250
rect 4000 3210 4010 3240
rect 4040 3210 4050 3240
rect 4000 3200 4050 3210
rect 4300 3240 4350 3250
rect 4300 3210 4310 3240
rect 4340 3210 4350 3240
rect 4300 3200 4350 3210
rect 4600 3240 4650 3250
rect 4600 3210 4610 3240
rect 4640 3210 4650 3240
rect 4600 3200 4650 3210
rect 4900 3240 4950 3250
rect 4900 3210 4910 3240
rect 4940 3210 4950 3240
rect 4900 3200 4950 3210
rect 5200 3240 5250 3250
rect 5200 3210 5210 3240
rect 5240 3210 5250 3240
rect 5200 3200 5250 3210
rect 5350 3240 5400 3250
rect 5350 3210 5360 3240
rect 5390 3210 5400 3240
rect 5350 3200 5400 3210
rect 5500 3240 5550 3250
rect 5500 3210 5510 3240
rect 5540 3210 5550 3240
rect 5500 3200 5550 3210
rect 5800 3240 5850 3250
rect 5800 3210 5810 3240
rect 5840 3210 5850 3240
rect 5800 3200 5850 3210
rect 6100 3240 6150 3250
rect 6100 3210 6110 3240
rect 6140 3210 6150 3240
rect 6100 3200 6150 3210
rect 6250 3240 6300 3250
rect 6250 3210 6260 3240
rect 6290 3210 6300 3240
rect 6250 3200 6300 3210
rect 6400 3240 6450 3250
rect 6400 3210 6410 3240
rect 6440 3210 6450 3240
rect 6400 3200 6450 3210
rect 6700 3240 6750 3250
rect 6700 3210 6710 3240
rect 6740 3210 6750 3240
rect 6700 3200 6750 3210
rect 7000 3240 7050 3250
rect 7000 3210 7010 3240
rect 7040 3210 7050 3240
rect 7000 3200 7050 3210
rect 7150 3240 7200 3250
rect 7150 3210 7160 3240
rect 7190 3210 7200 3240
rect 7150 3200 7200 3210
rect 7300 3240 7350 3250
rect 7300 3210 7310 3240
rect 7340 3210 7350 3240
rect 7300 3200 7350 3210
rect 7600 3240 7650 3250
rect 7600 3210 7610 3240
rect 7640 3210 7650 3240
rect 7600 3200 7650 3210
rect 7900 3240 7950 3250
rect 7900 3210 7910 3240
rect 7940 3210 7950 3240
rect 7900 3200 7950 3210
rect 8200 3240 8250 3250
rect 8200 3210 8210 3240
rect 8240 3210 8250 3240
rect 8200 3200 8250 3210
rect 8500 3240 8550 3250
rect 8500 3210 8510 3240
rect 8540 3210 8550 3240
rect 8500 3200 8550 3210
rect 8800 3240 8850 3250
rect 8800 3210 8810 3240
rect 8840 3210 8850 3240
rect 8800 3200 8850 3210
rect 9100 3240 9150 3250
rect 9100 3210 9110 3240
rect 9140 3210 9150 3240
rect 9100 3200 9150 3210
rect 9400 3240 9450 3250
rect 9400 3210 9410 3240
rect 9440 3210 9450 3240
rect 9400 3200 9450 3210
rect 9700 3240 9750 3250
rect 9700 3210 9710 3240
rect 9740 3210 9750 3240
rect 9700 3200 9750 3210
rect 10000 3240 10050 3250
rect 10000 3210 10010 3240
rect 10040 3210 10050 3240
rect 10000 3200 10050 3210
rect 10300 3240 10350 3250
rect 10300 3210 10310 3240
rect 10340 3210 10350 3240
rect 10300 3200 10350 3210
rect 10600 3240 10650 3250
rect 10600 3210 10610 3240
rect 10640 3210 10650 3240
rect 10600 3200 10650 3210
rect 10900 3240 10950 3250
rect 10900 3210 10910 3240
rect 10940 3210 10950 3240
rect 10900 3200 10950 3210
rect 11200 3240 11250 3250
rect 11200 3210 11210 3240
rect 11240 3210 11250 3240
rect 11200 3200 11250 3210
rect 11350 3240 11400 3250
rect 11350 3210 11360 3240
rect 11390 3210 11400 3240
rect 11350 3200 11400 3210
rect 11500 3240 11550 3250
rect 11500 3210 11510 3240
rect 11540 3210 11550 3240
rect 11500 3200 11550 3210
rect 11800 3240 11850 3250
rect 11800 3210 11810 3240
rect 11840 3210 11850 3240
rect 11800 3200 11850 3210
rect 12100 3240 12150 3250
rect 12100 3210 12110 3240
rect 12140 3210 12150 3240
rect 12100 3200 12150 3210
rect 12400 3240 12450 3250
rect 12400 3210 12410 3240
rect 12440 3210 12450 3240
rect 12400 3200 12450 3210
rect 12550 3240 12600 3250
rect 12550 3210 12560 3240
rect 12590 3210 12600 3240
rect 12550 3200 12600 3210
rect 12700 3240 12750 3250
rect 12700 3210 12710 3240
rect 12740 3210 12750 3240
rect 12700 3200 12750 3210
rect 13000 3240 13050 3250
rect 13000 3210 13010 3240
rect 13040 3210 13050 3240
rect 13000 3200 13050 3210
rect 13300 3240 13350 3250
rect 13300 3210 13310 3240
rect 13340 3210 13350 3240
rect 13300 3200 13350 3210
rect 13600 3240 13650 3250
rect 13600 3210 13610 3240
rect 13640 3210 13650 3240
rect 13600 3200 13650 3210
rect 13750 3240 13800 3250
rect 13750 3210 13760 3240
rect 13790 3210 13800 3240
rect 13750 3200 13800 3210
rect 13900 3240 13950 3250
rect 13900 3210 13910 3240
rect 13940 3210 13950 3240
rect 13900 3200 13950 3210
rect 14200 3240 14250 3250
rect 14200 3210 14210 3240
rect 14240 3210 14250 3240
rect 14200 3200 14250 3210
rect 14500 3240 14550 3250
rect 14500 3210 14510 3240
rect 14540 3210 14550 3240
rect 14500 3200 14550 3210
rect 14800 3240 14850 3250
rect 14800 3210 14810 3240
rect 14840 3210 14850 3240
rect 14800 3200 14850 3210
rect 14950 3240 15000 3250
rect 14950 3210 14960 3240
rect 14990 3210 15000 3240
rect 14950 3200 15000 3210
rect 15100 3240 15150 3250
rect 15100 3210 15110 3240
rect 15140 3210 15150 3240
rect 15100 3200 15150 3210
rect 15400 3240 15450 3250
rect 15400 3210 15410 3240
rect 15440 3210 15450 3240
rect 15400 3200 15450 3210
rect 15700 3240 15750 3250
rect 15700 3210 15710 3240
rect 15740 3210 15750 3240
rect 15700 3200 15750 3210
rect 16000 3240 16050 3250
rect 16000 3210 16010 3240
rect 16040 3210 16050 3240
rect 16000 3200 16050 3210
rect 16300 3240 16350 3250
rect 16300 3210 16310 3240
rect 16340 3210 16350 3240
rect 16300 3200 16350 3210
rect 16600 3240 16650 3250
rect 16600 3210 16610 3240
rect 16640 3210 16650 3240
rect 16600 3200 16650 3210
rect 16750 3240 16800 3250
rect 16750 3210 16760 3240
rect 16790 3210 16800 3240
rect 16750 3200 16800 3210
rect 16900 3240 16950 3250
rect 16900 3210 16910 3240
rect 16940 3210 16950 3240
rect 16900 3200 16950 3210
rect 17200 3240 17250 3250
rect 17200 3210 17210 3240
rect 17240 3210 17250 3240
rect 17200 3200 17250 3210
rect 17500 3240 17550 3250
rect 17500 3210 17510 3240
rect 17540 3210 17550 3240
rect 17500 3200 17550 3210
rect 17800 3240 17850 3250
rect 17800 3210 17810 3240
rect 17840 3210 17850 3240
rect 17800 3200 17850 3210
rect 18100 3240 18150 3250
rect 18100 3210 18110 3240
rect 18140 3210 18150 3240
rect 18100 3200 18150 3210
rect 18400 3240 18450 3250
rect 18400 3210 18410 3240
rect 18440 3210 18450 3240
rect 18400 3200 18450 3210
rect 18700 3240 18750 3250
rect 18700 3210 18710 3240
rect 18740 3210 18750 3240
rect 18700 3200 18750 3210
rect 19000 3240 19050 3250
rect 19000 3210 19010 3240
rect 19040 3210 19050 3240
rect 19000 3200 19050 3210
rect 19150 3240 19200 3250
rect 19150 3210 19160 3240
rect 19190 3210 19200 3240
rect 19150 3200 19200 3210
rect 19300 3240 19350 3250
rect 19300 3210 19310 3240
rect 19340 3210 19350 3240
rect 19300 3200 19350 3210
rect 19600 3240 19650 3250
rect 19600 3210 19610 3240
rect 19640 3210 19650 3240
rect 19600 3200 19650 3210
rect 19900 3240 19950 3250
rect 19900 3210 19910 3240
rect 19940 3210 19950 3240
rect 19900 3200 19950 3210
rect 20200 3240 20250 3250
rect 20200 3210 20210 3240
rect 20240 3210 20250 3240
rect 20200 3200 20250 3210
rect -650 3140 20400 3150
rect -650 3110 -640 3140
rect -610 3110 -40 3140
rect -10 3110 4160 3140
rect 4190 3110 8360 3140
rect 8390 3110 8660 3140
rect 8690 3110 8960 3140
rect 8990 3110 9260 3140
rect 9290 3110 9560 3140
rect 9590 3110 9860 3140
rect 9890 3110 10160 3140
rect 10190 3110 10460 3140
rect 10490 3110 10760 3140
rect 10790 3110 11960 3140
rect 11990 3110 13160 3140
rect 13190 3110 14360 3140
rect 14390 3110 15560 3140
rect 15590 3110 17960 3140
rect 17990 3110 20360 3140
rect 20390 3110 20400 3140
rect -650 3100 20400 3110
rect -650 3040 20400 3050
rect -650 3010 -640 3040
rect -610 3010 -40 3040
rect -10 3010 4160 3040
rect 4190 3010 8360 3040
rect 8390 3010 8660 3040
rect 8690 3010 8960 3040
rect 8990 3010 9260 3040
rect 9290 3010 9560 3040
rect 9590 3010 9860 3040
rect 9890 3010 10160 3040
rect 10190 3010 10460 3040
rect 10490 3010 10760 3040
rect 10790 3010 11960 3040
rect 11990 3010 13160 3040
rect 13190 3010 14360 3040
rect 14390 3010 15560 3040
rect 15590 3010 17960 3040
rect 17990 3010 20360 3040
rect 20390 3010 20400 3040
rect -650 3000 20400 3010
rect -650 2940 20400 2950
rect -650 2910 -640 2940
rect -610 2910 -40 2940
rect -10 2910 4160 2940
rect 4190 2910 8360 2940
rect 8390 2910 8660 2940
rect 8690 2910 8960 2940
rect 8990 2910 9260 2940
rect 9290 2910 9560 2940
rect 9590 2910 9860 2940
rect 9890 2910 10160 2940
rect 10190 2910 10460 2940
rect 10490 2910 10760 2940
rect 10790 2910 11960 2940
rect 11990 2910 13160 2940
rect 13190 2910 14360 2940
rect 14390 2910 15560 2940
rect 15590 2910 17960 2940
rect 17990 2910 20360 2940
rect 20390 2910 20400 2940
rect -650 2900 20400 2910
rect -650 2840 20400 2850
rect -650 2810 -640 2840
rect -610 2810 -40 2840
rect -10 2810 4160 2840
rect 4190 2810 8360 2840
rect 8390 2810 8660 2840
rect 8690 2810 8960 2840
rect 8990 2810 9260 2840
rect 9290 2810 9560 2840
rect 9590 2810 9860 2840
rect 9890 2810 10160 2840
rect 10190 2810 10460 2840
rect 10490 2810 10760 2840
rect 10790 2810 11960 2840
rect 11990 2810 13160 2840
rect 13190 2810 14360 2840
rect 14390 2810 15560 2840
rect 15590 2810 17960 2840
rect 17990 2810 20360 2840
rect 20390 2810 20400 2840
rect -650 2800 20400 2810
rect -650 2740 20400 2750
rect -650 2710 -640 2740
rect -610 2710 -40 2740
rect -10 2710 4160 2740
rect 4190 2710 8360 2740
rect 8390 2710 8660 2740
rect 8690 2710 8960 2740
rect 8990 2710 9260 2740
rect 9290 2710 9560 2740
rect 9590 2710 9860 2740
rect 9890 2710 10160 2740
rect 10190 2710 10460 2740
rect 10490 2710 10760 2740
rect 10790 2710 11960 2740
rect 11990 2710 13160 2740
rect 13190 2710 14360 2740
rect 14390 2710 15560 2740
rect 15590 2710 20360 2740
rect 20390 2710 20400 2740
rect -650 2700 20400 2710
rect -650 2590 20400 2650
rect -650 2560 -640 2590
rect -610 2560 -40 2590
rect -10 2560 4160 2590
rect 4190 2560 8360 2590
rect 8390 2560 8660 2590
rect 8690 2560 8960 2590
rect 8990 2560 9260 2590
rect 9290 2560 9560 2590
rect 9590 2560 9860 2590
rect 9890 2560 10160 2590
rect 10190 2560 10460 2590
rect 10490 2560 10760 2590
rect 10790 2560 11960 2590
rect 11990 2560 13160 2590
rect 13190 2560 14360 2590
rect 14390 2560 15560 2590
rect 15590 2560 17960 2590
rect 17990 2560 20360 2590
rect 20390 2560 20400 2590
rect -650 2550 20400 2560
rect -900 2400 20400 2450
rect -900 2300 20400 2350
rect -900 2200 20400 2250
rect -900 2100 20400 2150
rect -900 2000 20400 2050
rect -900 1690 20400 1700
rect -900 1660 -640 1690
rect -610 1660 -40 1690
rect -10 1660 8360 1690
rect 8390 1660 10760 1690
rect 10790 1660 15560 1690
rect 15590 1660 17960 1690
rect 17990 1660 20360 1690
rect 20390 1660 20400 1690
rect -900 1640 20400 1660
rect -900 1610 -640 1640
rect -610 1610 -40 1640
rect -10 1610 8360 1640
rect 8390 1610 10760 1640
rect 10790 1610 15560 1640
rect 15590 1610 17960 1640
rect 17990 1610 20360 1640
rect 20390 1610 20400 1640
rect -900 1600 20400 1610
rect -900 1540 20400 1550
rect -900 1510 -640 1540
rect -610 1510 -40 1540
rect -10 1510 8360 1540
rect 8390 1510 10760 1540
rect 10790 1510 15560 1540
rect 15590 1510 17960 1540
rect 17990 1510 20360 1540
rect 20390 1510 20400 1540
rect -900 1500 20400 1510
rect -900 1440 20400 1450
rect -900 1410 -640 1440
rect -610 1410 -40 1440
rect -10 1410 8360 1440
rect 8390 1410 10760 1440
rect 10790 1410 15560 1440
rect 15590 1410 17960 1440
rect 17990 1410 20360 1440
rect 20390 1410 20400 1440
rect -900 1400 20400 1410
rect -900 1340 20400 1350
rect -900 1310 -640 1340
rect -610 1310 -40 1340
rect -10 1310 8360 1340
rect 8390 1310 10760 1340
rect 10790 1310 15560 1340
rect 15590 1310 17960 1340
rect 17990 1310 20360 1340
rect 20390 1310 20400 1340
rect -900 1300 20400 1310
rect -900 1240 20400 1250
rect -900 1210 -640 1240
rect -610 1210 -40 1240
rect -10 1210 8360 1240
rect 8390 1210 10760 1240
rect 10790 1210 15560 1240
rect 15590 1210 17960 1240
rect 17990 1210 20360 1240
rect 20390 1210 20400 1240
rect -900 1200 20400 1210
rect -900 1140 20400 1150
rect -900 1110 -640 1140
rect -610 1110 -40 1140
rect -10 1110 8360 1140
rect 8390 1110 10760 1140
rect 10790 1110 15560 1140
rect 15590 1110 17960 1140
rect 17990 1110 20360 1140
rect 20390 1110 20400 1140
rect -900 1100 20400 1110
rect -900 1040 20400 1050
rect -900 1010 -640 1040
rect -610 1010 -40 1040
rect -10 1010 8360 1040
rect 8390 1010 10760 1040
rect 10790 1010 15560 1040
rect 15590 1010 17960 1040
rect 17990 1010 20360 1040
rect 20390 1010 20400 1040
rect -900 1000 20400 1010
rect -900 940 20400 950
rect -900 910 -640 940
rect -610 910 -40 940
rect -10 910 8360 940
rect 8390 910 10760 940
rect 10790 910 15560 940
rect 15590 910 17960 940
rect 17990 910 20360 940
rect 20390 910 20400 940
rect -900 900 20400 910
rect -500 840 -450 850
rect -500 810 -490 840
rect -460 810 -450 840
rect -500 800 -450 810
rect -350 840 -300 850
rect -350 810 -340 840
rect -310 810 -300 840
rect -350 800 -300 810
rect -200 840 -150 850
rect -200 810 -190 840
rect -160 810 -150 840
rect -200 800 -150 810
rect 100 840 150 850
rect 100 810 110 840
rect 140 810 150 840
rect 100 800 150 810
rect 400 840 450 850
rect 400 810 410 840
rect 440 810 450 840
rect 400 800 450 810
rect 700 840 750 850
rect 700 810 710 840
rect 740 810 750 840
rect 700 800 750 810
rect 1000 840 1050 850
rect 1000 810 1010 840
rect 1040 810 1050 840
rect 1000 800 1050 810
rect 1300 840 1350 850
rect 1300 810 1310 840
rect 1340 810 1350 840
rect 1300 800 1350 810
rect 1600 840 1650 850
rect 1600 810 1610 840
rect 1640 810 1650 840
rect 1600 800 1650 810
rect 1900 840 1950 850
rect 1900 810 1910 840
rect 1940 810 1950 840
rect 1900 800 1950 810
rect 2200 840 2250 850
rect 2200 810 2210 840
rect 2240 810 2250 840
rect 2200 800 2250 810
rect 2350 840 2400 850
rect 2350 810 2360 840
rect 2390 810 2400 840
rect 2350 800 2400 810
rect 2500 840 2550 850
rect 2500 810 2510 840
rect 2540 810 2550 840
rect 2500 800 2550 810
rect 2800 840 2850 850
rect 2800 810 2810 840
rect 2840 810 2850 840
rect 2800 800 2850 810
rect 3100 840 3150 850
rect 3100 810 3110 840
rect 3140 810 3150 840
rect 3100 800 3150 810
rect 3400 840 3450 850
rect 3400 810 3410 840
rect 3440 810 3450 840
rect 3400 800 3450 810
rect 3700 840 3750 850
rect 3700 810 3710 840
rect 3740 810 3750 840
rect 3700 800 3750 810
rect 3850 840 3900 850
rect 3850 810 3860 840
rect 3890 810 3900 840
rect 3850 800 3900 810
rect 4000 840 4050 850
rect 4000 810 4010 840
rect 4040 810 4050 840
rect 4000 800 4050 810
rect 4300 840 4350 850
rect 4300 810 4310 840
rect 4340 810 4350 840
rect 4300 800 4350 810
rect 4450 840 4500 850
rect 4450 810 4460 840
rect 4490 810 4500 840
rect 4450 800 4500 810
rect 4600 840 4650 850
rect 4600 810 4610 840
rect 4640 810 4650 840
rect 4600 800 4650 810
rect 4900 840 4950 850
rect 4900 810 4910 840
rect 4940 810 4950 840
rect 4900 800 4950 810
rect 5200 840 5250 850
rect 5200 810 5210 840
rect 5240 810 5250 840
rect 5200 800 5250 810
rect 5500 840 5550 850
rect 5500 810 5510 840
rect 5540 810 5550 840
rect 5500 800 5550 810
rect 5800 840 5850 850
rect 5800 810 5810 840
rect 5840 810 5850 840
rect 5800 800 5850 810
rect 5950 840 6000 850
rect 5950 810 5960 840
rect 5990 810 6000 840
rect 5950 800 6000 810
rect 6100 840 6150 850
rect 6100 810 6110 840
rect 6140 810 6150 840
rect 6100 800 6150 810
rect 6400 840 6450 850
rect 6400 810 6410 840
rect 6440 810 6450 840
rect 6400 800 6450 810
rect 6700 840 6750 850
rect 6700 810 6710 840
rect 6740 810 6750 840
rect 6700 800 6750 810
rect 7000 840 7050 850
rect 7000 810 7010 840
rect 7040 810 7050 840
rect 7000 800 7050 810
rect 7300 840 7350 850
rect 7300 810 7310 840
rect 7340 810 7350 840
rect 7300 800 7350 810
rect 7600 840 7650 850
rect 7600 810 7610 840
rect 7640 810 7650 840
rect 7600 800 7650 810
rect 7900 840 7950 850
rect 7900 810 7910 840
rect 7940 810 7950 840
rect 7900 800 7950 810
rect 8200 840 8250 850
rect 8200 810 8210 840
rect 8240 810 8250 840
rect 8200 800 8250 810
rect 8500 840 8550 850
rect 8500 810 8510 840
rect 8540 810 8550 840
rect 8500 800 8550 810
rect 8800 840 8850 850
rect 8800 810 8810 840
rect 8840 810 8850 840
rect 8800 800 8850 810
rect 9100 840 9150 850
rect 9100 810 9110 840
rect 9140 810 9150 840
rect 9100 800 9150 810
rect 9400 840 9450 850
rect 9400 810 9410 840
rect 9440 810 9450 840
rect 9400 800 9450 810
rect 9550 840 9600 850
rect 9550 810 9560 840
rect 9590 810 9600 840
rect 9550 800 9600 810
rect 9700 840 9750 850
rect 9700 810 9710 840
rect 9740 810 9750 840
rect 9700 800 9750 810
rect 10000 840 10050 850
rect 10000 810 10010 840
rect 10040 810 10050 840
rect 10000 800 10050 810
rect 10300 840 10350 850
rect 10300 810 10310 840
rect 10340 810 10350 840
rect 10300 800 10350 810
rect 10600 840 10650 850
rect 10600 810 10610 840
rect 10640 810 10650 840
rect 10600 800 10650 810
rect 10900 840 10950 850
rect 10900 810 10910 840
rect 10940 810 10950 840
rect 10900 800 10950 810
rect 11200 840 11250 850
rect 11200 810 11210 840
rect 11240 810 11250 840
rect 11200 800 11250 810
rect 11500 840 11550 850
rect 11500 810 11510 840
rect 11540 810 11550 840
rect 11500 800 11550 810
rect 11800 840 11850 850
rect 11800 810 11810 840
rect 11840 810 11850 840
rect 11800 800 11850 810
rect 12100 840 12150 850
rect 12100 810 12110 840
rect 12140 810 12150 840
rect 12100 800 12150 810
rect 12400 840 12450 850
rect 12400 810 12410 840
rect 12440 810 12450 840
rect 12400 800 12450 810
rect 12550 840 12600 850
rect 12550 810 12560 840
rect 12590 810 12600 840
rect 12550 800 12600 810
rect 12700 840 12750 850
rect 12700 810 12710 840
rect 12740 810 12750 840
rect 12700 800 12750 810
rect 13000 840 13050 850
rect 13000 810 13010 840
rect 13040 810 13050 840
rect 13000 800 13050 810
rect 13150 840 13200 850
rect 13150 810 13160 840
rect 13190 810 13200 840
rect 13150 800 13200 810
rect 13300 840 13350 850
rect 13300 810 13310 840
rect 13340 810 13350 840
rect 13300 800 13350 810
rect 13600 840 13650 850
rect 13600 810 13610 840
rect 13640 810 13650 840
rect 13600 800 13650 810
rect 13750 840 13800 850
rect 13750 810 13760 840
rect 13790 810 13800 840
rect 13750 800 13800 810
rect 13900 840 13950 850
rect 13900 810 13910 840
rect 13940 810 13950 840
rect 13900 800 13950 810
rect 14200 840 14250 850
rect 14200 810 14210 840
rect 14240 810 14250 840
rect 14200 800 14250 810
rect 14500 840 14550 850
rect 14500 810 14510 840
rect 14540 810 14550 840
rect 14500 800 14550 810
rect 14800 840 14850 850
rect 14800 810 14810 840
rect 14840 810 14850 840
rect 14800 800 14850 810
rect 15100 840 15150 850
rect 15100 810 15110 840
rect 15140 810 15150 840
rect 15100 800 15150 810
rect 15400 840 15450 850
rect 15400 810 15410 840
rect 15440 810 15450 840
rect 15400 800 15450 810
rect 15700 840 15750 850
rect 15700 810 15710 840
rect 15740 810 15750 840
rect 15700 800 15750 810
rect 16000 840 16050 850
rect 16000 810 16010 840
rect 16040 810 16050 840
rect 16000 800 16050 810
rect 16300 840 16350 850
rect 16300 810 16310 840
rect 16340 810 16350 840
rect 16300 800 16350 810
rect 16600 840 16650 850
rect 16600 810 16610 840
rect 16640 810 16650 840
rect 16600 800 16650 810
rect 16750 840 16800 850
rect 16750 810 16760 840
rect 16790 810 16800 840
rect 16750 800 16800 810
rect 16900 840 16950 850
rect 16900 810 16910 840
rect 16940 810 16950 840
rect 16900 800 16950 810
rect 17200 840 17250 850
rect 17200 810 17210 840
rect 17240 810 17250 840
rect 17200 800 17250 810
rect 17500 840 17550 850
rect 17500 810 17510 840
rect 17540 810 17550 840
rect 17500 800 17550 810
rect 17800 840 17850 850
rect 17800 810 17810 840
rect 17840 810 17850 840
rect 17800 800 17850 810
rect 18100 840 18150 850
rect 18100 810 18110 840
rect 18140 810 18150 840
rect 18100 800 18150 810
rect 18400 840 18450 850
rect 18400 810 18410 840
rect 18440 810 18450 840
rect 18400 800 18450 810
rect 18700 840 18750 850
rect 18700 810 18710 840
rect 18740 810 18750 840
rect 18700 800 18750 810
rect 19000 840 19050 850
rect 19000 810 19010 840
rect 19040 810 19050 840
rect 19000 800 19050 810
rect 19150 840 19200 850
rect 19150 810 19160 840
rect 19190 810 19200 840
rect 19150 800 19200 810
rect 19300 840 19350 850
rect 19300 810 19310 840
rect 19340 810 19350 840
rect 19300 800 19350 810
rect 19600 840 19650 850
rect 19600 810 19610 840
rect 19640 810 19650 840
rect 19600 800 19650 810
rect 19900 840 19950 850
rect 19900 810 19910 840
rect 19940 810 19950 840
rect 19900 800 19950 810
rect 20200 840 20250 850
rect 20200 810 20210 840
rect 20240 810 20250 840
rect 20200 800 20250 810
rect -900 740 20400 750
rect -900 710 -640 740
rect -610 710 -40 740
rect -10 710 8360 740
rect 8390 710 10760 740
rect 10790 710 15560 740
rect 15590 710 17960 740
rect 17990 710 20360 740
rect 20390 710 20400 740
rect -900 700 20400 710
rect -900 640 20400 650
rect -900 610 -640 640
rect -610 610 -40 640
rect -10 610 8360 640
rect 8390 610 10760 640
rect 10790 610 15560 640
rect 15590 610 17960 640
rect 17990 610 20360 640
rect 20390 610 20400 640
rect -900 600 20400 610
rect -900 540 20400 550
rect -900 510 -640 540
rect -610 510 -40 540
rect -10 510 8360 540
rect 8390 510 10760 540
rect 10790 510 15560 540
rect 15590 510 17960 540
rect 17990 510 20360 540
rect 20390 510 20400 540
rect -900 500 20400 510
rect -900 440 20400 450
rect -900 410 -640 440
rect -610 410 -40 440
rect -10 410 8360 440
rect 8390 410 10760 440
rect 10790 410 15560 440
rect 15590 410 17960 440
rect 17990 410 20360 440
rect 20390 410 20400 440
rect -900 400 20400 410
rect -900 340 20400 350
rect -900 310 -640 340
rect -610 310 -40 340
rect -10 310 8360 340
rect 8390 310 10760 340
rect 10790 310 15560 340
rect 15590 310 17960 340
rect 17990 310 20360 340
rect 20390 310 20400 340
rect -900 300 20400 310
rect -900 240 20400 250
rect -900 210 -640 240
rect -610 210 -40 240
rect -10 210 8360 240
rect 8390 210 10760 240
rect 10790 210 15560 240
rect 15590 210 17960 240
rect 17990 210 20360 240
rect 20390 210 20400 240
rect -900 200 20400 210
rect -900 140 20400 150
rect -900 110 -640 140
rect -610 110 -40 140
rect -10 110 8360 140
rect 8390 110 10760 140
rect 10790 110 15560 140
rect 15590 110 17960 140
rect 17990 110 20360 140
rect 20390 110 20400 140
rect -900 100 20400 110
rect -900 40 20400 50
rect -900 10 -640 40
rect -610 10 -40 40
rect -10 10 8360 40
rect 8390 10 10760 40
rect 10790 10 15560 40
rect 15590 10 17960 40
rect 17990 10 20360 40
rect 20390 10 20400 40
rect -900 -10 20400 10
rect -900 -40 -640 -10
rect -610 -40 -40 -10
rect -10 -40 8360 -10
rect 8390 -40 10760 -10
rect 10790 -40 15560 -10
rect 15590 -40 17960 -10
rect 17990 -40 20360 -10
rect 20390 -40 20400 -10
rect -900 -60 20400 -40
rect -900 -90 -640 -60
rect -610 -90 -40 -60
rect -10 -90 8360 -60
rect 8390 -90 10760 -60
rect 10790 -90 15560 -60
rect 15590 -90 17960 -60
rect 17990 -90 20360 -60
rect 20390 -90 20400 -60
rect -900 -100 20400 -90
rect -900 -160 20400 -150
rect -900 -190 -640 -160
rect -610 -190 -40 -160
rect -10 -190 8360 -160
rect 8390 -190 10760 -160
rect 10790 -190 15560 -160
rect 15590 -190 17960 -160
rect 17990 -190 20360 -160
rect 20390 -190 20400 -160
rect -900 -200 20400 -190
rect -900 -260 20400 -250
rect -900 -290 -640 -260
rect -610 -290 -40 -260
rect -10 -290 8360 -260
rect 8390 -290 10760 -260
rect 10790 -290 15560 -260
rect 15590 -290 17960 -260
rect 17990 -290 20360 -260
rect 20390 -290 20400 -260
rect -900 -300 20400 -290
rect -900 -360 20400 -350
rect -900 -390 -640 -360
rect -610 -390 -40 -360
rect -10 -390 8360 -360
rect 8390 -390 10760 -360
rect 10790 -390 15560 -360
rect 15590 -390 17960 -360
rect 17990 -390 20360 -360
rect 20390 -390 20400 -360
rect -900 -400 20400 -390
rect -900 -460 20400 -450
rect -900 -490 -640 -460
rect -610 -490 -40 -460
rect -10 -490 8360 -460
rect 8390 -490 10760 -460
rect 10790 -490 15560 -460
rect 15590 -490 17960 -460
rect 17990 -490 20360 -460
rect 20390 -490 20400 -460
rect -900 -500 20400 -490
rect -900 -560 20400 -550
rect -900 -590 -640 -560
rect -610 -590 -40 -560
rect -10 -590 8360 -560
rect 8390 -590 10760 -560
rect 10790 -590 15560 -560
rect 15590 -590 17960 -560
rect 17990 -590 20360 -560
rect 20390 -590 20400 -560
rect -900 -600 20400 -590
rect -900 -660 20400 -650
rect -900 -690 -640 -660
rect -610 -690 -40 -660
rect -10 -690 8360 -660
rect 8390 -690 10760 -660
rect 10790 -690 15560 -660
rect 15590 -690 17960 -660
rect 17990 -690 20360 -660
rect 20390 -690 20400 -660
rect -900 -700 20400 -690
rect -900 -760 20400 -750
rect -900 -790 -640 -760
rect -610 -790 -40 -760
rect -10 -790 8360 -760
rect 8390 -790 10760 -760
rect 10790 -790 15560 -760
rect 15590 -790 17960 -760
rect 17990 -790 20360 -760
rect 20390 -790 20400 -760
rect -900 -800 20400 -790
rect -500 -860 -450 -850
rect -500 -890 -490 -860
rect -460 -890 -450 -860
rect -500 -900 -450 -890
rect -350 -860 -300 -850
rect -350 -890 -340 -860
rect -310 -890 -300 -860
rect -350 -900 -300 -890
rect -200 -860 -150 -850
rect -200 -890 -190 -860
rect -160 -890 -150 -860
rect -200 -900 -150 -890
rect 100 -860 150 -850
rect 100 -890 110 -860
rect 140 -890 150 -860
rect 100 -900 150 -890
rect 400 -860 450 -850
rect 400 -890 410 -860
rect 440 -890 450 -860
rect 400 -900 450 -890
rect 700 -860 750 -850
rect 700 -890 710 -860
rect 740 -890 750 -860
rect 700 -900 750 -890
rect 1000 -860 1050 -850
rect 1000 -890 1010 -860
rect 1040 -890 1050 -860
rect 1000 -900 1050 -890
rect 1300 -860 1350 -850
rect 1300 -890 1310 -860
rect 1340 -890 1350 -860
rect 1300 -900 1350 -890
rect 1600 -860 1650 -850
rect 1600 -890 1610 -860
rect 1640 -890 1650 -860
rect 1600 -900 1650 -890
rect 1900 -860 1950 -850
rect 1900 -890 1910 -860
rect 1940 -890 1950 -860
rect 1900 -900 1950 -890
rect 2200 -860 2250 -850
rect 2200 -890 2210 -860
rect 2240 -890 2250 -860
rect 2200 -900 2250 -890
rect 2350 -860 2400 -850
rect 2350 -890 2360 -860
rect 2390 -890 2400 -860
rect 2350 -900 2400 -890
rect 2500 -860 2550 -850
rect 2500 -890 2510 -860
rect 2540 -890 2550 -860
rect 2500 -900 2550 -890
rect 2800 -860 2850 -850
rect 2800 -890 2810 -860
rect 2840 -890 2850 -860
rect 2800 -900 2850 -890
rect 3100 -860 3150 -850
rect 3100 -890 3110 -860
rect 3140 -890 3150 -860
rect 3100 -900 3150 -890
rect 3400 -860 3450 -850
rect 3400 -890 3410 -860
rect 3440 -890 3450 -860
rect 3400 -900 3450 -890
rect 3700 -860 3750 -850
rect 3700 -890 3710 -860
rect 3740 -890 3750 -860
rect 3700 -900 3750 -890
rect 3850 -860 3900 -850
rect 3850 -890 3860 -860
rect 3890 -890 3900 -860
rect 3850 -900 3900 -890
rect 4000 -860 4050 -850
rect 4000 -890 4010 -860
rect 4040 -890 4050 -860
rect 4000 -900 4050 -890
rect 4300 -860 4350 -850
rect 4300 -890 4310 -860
rect 4340 -890 4350 -860
rect 4300 -900 4350 -890
rect 4450 -860 4500 -850
rect 4450 -890 4460 -860
rect 4490 -890 4500 -860
rect 4450 -900 4500 -890
rect 4600 -860 4650 -850
rect 4600 -890 4610 -860
rect 4640 -890 4650 -860
rect 4600 -900 4650 -890
rect 4900 -860 4950 -850
rect 4900 -890 4910 -860
rect 4940 -890 4950 -860
rect 4900 -900 4950 -890
rect 5200 -860 5250 -850
rect 5200 -890 5210 -860
rect 5240 -890 5250 -860
rect 5200 -900 5250 -890
rect 5500 -860 5550 -850
rect 5500 -890 5510 -860
rect 5540 -890 5550 -860
rect 5500 -900 5550 -890
rect 5800 -860 5850 -850
rect 5800 -890 5810 -860
rect 5840 -890 5850 -860
rect 5800 -900 5850 -890
rect 5950 -860 6000 -850
rect 5950 -890 5960 -860
rect 5990 -890 6000 -860
rect 5950 -900 6000 -890
rect 6100 -860 6150 -850
rect 6100 -890 6110 -860
rect 6140 -890 6150 -860
rect 6100 -900 6150 -890
rect 6400 -860 6450 -850
rect 6400 -890 6410 -860
rect 6440 -890 6450 -860
rect 6400 -900 6450 -890
rect 6700 -860 6750 -850
rect 6700 -890 6710 -860
rect 6740 -890 6750 -860
rect 6700 -900 6750 -890
rect 7000 -860 7050 -850
rect 7000 -890 7010 -860
rect 7040 -890 7050 -860
rect 7000 -900 7050 -890
rect 7300 -860 7350 -850
rect 7300 -890 7310 -860
rect 7340 -890 7350 -860
rect 7300 -900 7350 -890
rect 7600 -860 7650 -850
rect 7600 -890 7610 -860
rect 7640 -890 7650 -860
rect 7600 -900 7650 -890
rect 7900 -860 7950 -850
rect 7900 -890 7910 -860
rect 7940 -890 7950 -860
rect 7900 -900 7950 -890
rect 8200 -860 8250 -850
rect 8200 -890 8210 -860
rect 8240 -890 8250 -860
rect 8200 -900 8250 -890
rect 8500 -860 8550 -850
rect 8500 -890 8510 -860
rect 8540 -890 8550 -860
rect 8500 -900 8550 -890
rect 8800 -860 8850 -850
rect 8800 -890 8810 -860
rect 8840 -890 8850 -860
rect 8800 -900 8850 -890
rect 9100 -860 9150 -850
rect 9100 -890 9110 -860
rect 9140 -890 9150 -860
rect 9100 -900 9150 -890
rect 9400 -860 9450 -850
rect 9400 -890 9410 -860
rect 9440 -890 9450 -860
rect 9400 -900 9450 -890
rect 9550 -860 9600 -850
rect 9550 -890 9560 -860
rect 9590 -890 9600 -860
rect 9550 -900 9600 -890
rect 9700 -860 9750 -850
rect 9700 -890 9710 -860
rect 9740 -890 9750 -860
rect 9700 -900 9750 -890
rect 10000 -860 10050 -850
rect 10000 -890 10010 -860
rect 10040 -890 10050 -860
rect 10000 -900 10050 -890
rect 10300 -860 10350 -850
rect 10300 -890 10310 -860
rect 10340 -890 10350 -860
rect 10300 -900 10350 -890
rect 10600 -860 10650 -850
rect 10600 -890 10610 -860
rect 10640 -890 10650 -860
rect 10600 -900 10650 -890
rect 10900 -860 10950 -850
rect 10900 -890 10910 -860
rect 10940 -890 10950 -860
rect 10900 -900 10950 -890
rect 11200 -860 11250 -850
rect 11200 -890 11210 -860
rect 11240 -890 11250 -860
rect 11200 -900 11250 -890
rect 11500 -860 11550 -850
rect 11500 -890 11510 -860
rect 11540 -890 11550 -860
rect 11500 -900 11550 -890
rect 11800 -860 11850 -850
rect 11800 -890 11810 -860
rect 11840 -890 11850 -860
rect 11800 -900 11850 -890
rect 12100 -860 12150 -850
rect 12100 -890 12110 -860
rect 12140 -890 12150 -860
rect 12100 -900 12150 -890
rect 12400 -860 12450 -850
rect 12400 -890 12410 -860
rect 12440 -890 12450 -860
rect 12400 -900 12450 -890
rect 12550 -860 12600 -850
rect 12550 -890 12560 -860
rect 12590 -890 12600 -860
rect 12550 -900 12600 -890
rect 12700 -860 12750 -850
rect 12700 -890 12710 -860
rect 12740 -890 12750 -860
rect 12700 -900 12750 -890
rect 13000 -860 13050 -850
rect 13000 -890 13010 -860
rect 13040 -890 13050 -860
rect 13000 -900 13050 -890
rect 13150 -860 13200 -850
rect 13150 -890 13160 -860
rect 13190 -890 13200 -860
rect 13150 -900 13200 -890
rect 13300 -860 13350 -850
rect 13300 -890 13310 -860
rect 13340 -890 13350 -860
rect 13300 -900 13350 -890
rect 13600 -860 13650 -850
rect 13600 -890 13610 -860
rect 13640 -890 13650 -860
rect 13600 -900 13650 -890
rect 13750 -860 13800 -850
rect 13750 -890 13760 -860
rect 13790 -890 13800 -860
rect 13750 -900 13800 -890
rect 13900 -860 13950 -850
rect 13900 -890 13910 -860
rect 13940 -890 13950 -860
rect 13900 -900 13950 -890
rect 14200 -860 14250 -850
rect 14200 -890 14210 -860
rect 14240 -890 14250 -860
rect 14200 -900 14250 -890
rect 14500 -860 14550 -850
rect 14500 -890 14510 -860
rect 14540 -890 14550 -860
rect 14500 -900 14550 -890
rect 14800 -860 14850 -850
rect 14800 -890 14810 -860
rect 14840 -890 14850 -860
rect 14800 -900 14850 -890
rect 15100 -860 15150 -850
rect 15100 -890 15110 -860
rect 15140 -890 15150 -860
rect 15100 -900 15150 -890
rect 15400 -860 15450 -850
rect 15400 -890 15410 -860
rect 15440 -890 15450 -860
rect 15400 -900 15450 -890
rect 15700 -860 15750 -850
rect 15700 -890 15710 -860
rect 15740 -890 15750 -860
rect 15700 -900 15750 -890
rect 16000 -860 16050 -850
rect 16000 -890 16010 -860
rect 16040 -890 16050 -860
rect 16000 -900 16050 -890
rect 16300 -860 16350 -850
rect 16300 -890 16310 -860
rect 16340 -890 16350 -860
rect 16300 -900 16350 -890
rect 16600 -860 16650 -850
rect 16600 -890 16610 -860
rect 16640 -890 16650 -860
rect 16600 -900 16650 -890
rect 16750 -860 16800 -850
rect 16750 -890 16760 -860
rect 16790 -890 16800 -860
rect 16750 -900 16800 -890
rect 16900 -860 16950 -850
rect 16900 -890 16910 -860
rect 16940 -890 16950 -860
rect 16900 -900 16950 -890
rect 17200 -860 17250 -850
rect 17200 -890 17210 -860
rect 17240 -890 17250 -860
rect 17200 -900 17250 -890
rect 17500 -860 17550 -850
rect 17500 -890 17510 -860
rect 17540 -890 17550 -860
rect 17500 -900 17550 -890
rect 17800 -860 17850 -850
rect 17800 -890 17810 -860
rect 17840 -890 17850 -860
rect 17800 -900 17850 -890
rect 18100 -860 18150 -850
rect 18100 -890 18110 -860
rect 18140 -890 18150 -860
rect 18100 -900 18150 -890
rect 18400 -860 18450 -850
rect 18400 -890 18410 -860
rect 18440 -890 18450 -860
rect 18400 -900 18450 -890
rect 18700 -860 18750 -850
rect 18700 -890 18710 -860
rect 18740 -890 18750 -860
rect 18700 -900 18750 -890
rect 19000 -860 19050 -850
rect 19000 -890 19010 -860
rect 19040 -890 19050 -860
rect 19000 -900 19050 -890
rect 19150 -860 19200 -850
rect 19150 -890 19160 -860
rect 19190 -890 19200 -860
rect 19150 -900 19200 -890
rect 19300 -860 19350 -850
rect 19300 -890 19310 -860
rect 19340 -890 19350 -860
rect 19300 -900 19350 -890
rect 19600 -860 19650 -850
rect 19600 -890 19610 -860
rect 19640 -890 19650 -860
rect 19600 -900 19650 -890
rect 19900 -860 19950 -850
rect 19900 -890 19910 -860
rect 19940 -890 19950 -860
rect 19900 -900 19950 -890
rect 20200 -860 20250 -850
rect 20200 -890 20210 -860
rect 20240 -890 20250 -860
rect 20200 -900 20250 -890
rect -900 -960 20400 -950
rect -900 -990 -640 -960
rect -610 -990 -40 -960
rect -10 -990 8360 -960
rect 8390 -990 10760 -960
rect 10790 -990 15560 -960
rect 15590 -990 17960 -960
rect 17990 -990 20360 -960
rect 20390 -990 20400 -960
rect -900 -1000 20400 -990
rect -900 -1060 20400 -1050
rect -900 -1090 -640 -1060
rect -610 -1090 -40 -1060
rect -10 -1090 8360 -1060
rect 8390 -1090 10760 -1060
rect 10790 -1090 15560 -1060
rect 15590 -1090 17960 -1060
rect 17990 -1090 20360 -1060
rect 20390 -1090 20400 -1060
rect -900 -1100 20400 -1090
rect -900 -1160 20400 -1150
rect -900 -1190 -640 -1160
rect -610 -1190 -40 -1160
rect -10 -1190 8360 -1160
rect 8390 -1190 10760 -1160
rect 10790 -1190 15560 -1160
rect 15590 -1190 17960 -1160
rect 17990 -1190 20360 -1160
rect 20390 -1190 20400 -1160
rect -900 -1200 20400 -1190
rect -900 -1260 20400 -1250
rect -900 -1290 -640 -1260
rect -610 -1290 -40 -1260
rect -10 -1290 8360 -1260
rect 8390 -1290 10760 -1260
rect 10790 -1290 15560 -1260
rect 15590 -1290 17960 -1260
rect 17990 -1290 20360 -1260
rect 20390 -1290 20400 -1260
rect -900 -1300 20400 -1290
rect -900 -1360 20400 -1350
rect -900 -1390 -640 -1360
rect -610 -1390 -40 -1360
rect -10 -1390 8360 -1360
rect 8390 -1390 10760 -1360
rect 10790 -1390 15560 -1360
rect 15590 -1390 17960 -1360
rect 17990 -1390 20360 -1360
rect 20390 -1390 20400 -1360
rect -900 -1400 20400 -1390
rect -900 -1460 20400 -1450
rect -900 -1490 -640 -1460
rect -610 -1490 -40 -1460
rect -10 -1490 8360 -1460
rect 8390 -1490 10760 -1460
rect 10790 -1490 15560 -1460
rect 15590 -1490 17960 -1460
rect 17990 -1490 20360 -1460
rect 20390 -1490 20400 -1460
rect -900 -1500 20400 -1490
rect -900 -1560 20400 -1550
rect -900 -1590 -640 -1560
rect -610 -1590 -40 -1560
rect -10 -1590 8360 -1560
rect 8390 -1590 10760 -1560
rect 10790 -1590 15560 -1560
rect 15590 -1590 17960 -1560
rect 17990 -1590 20360 -1560
rect 20390 -1590 20400 -1560
rect -900 -1600 20400 -1590
rect -900 -1660 20400 -1650
rect -900 -1690 -640 -1660
rect -610 -1690 -40 -1660
rect -10 -1690 8360 -1660
rect 8390 -1690 10760 -1660
rect 10790 -1690 15560 -1660
rect 15590 -1690 17960 -1660
rect 17990 -1690 20360 -1660
rect 20390 -1690 20400 -1660
rect -900 -1710 20400 -1690
rect -900 -1740 -640 -1710
rect -610 -1740 -40 -1710
rect -10 -1740 8360 -1710
rect 8390 -1740 10760 -1710
rect 10790 -1740 15560 -1710
rect 15590 -1740 17960 -1710
rect 17990 -1740 20360 -1710
rect 20390 -1740 20400 -1710
rect -900 -1750 20400 -1740
<< via2 >>
rect -640 5160 -610 5190
rect 8360 5160 8390 5190
rect 8660 5160 8690 5190
rect 8960 5160 8990 5190
rect 9260 5160 9290 5190
rect 9560 5160 9590 5190
rect 9860 5160 9890 5190
rect 10160 5160 10190 5190
rect 10460 5160 10490 5190
rect 10760 5160 10790 5190
rect 11960 5160 11990 5190
rect 13160 5160 13190 5190
rect 14360 5160 14390 5190
rect 15560 5160 15590 5190
rect 17960 5160 17990 5190
rect 20360 5160 20390 5190
rect -490 4510 -460 4540
rect -340 4510 -310 4540
rect -190 4510 -160 4540
rect 110 4510 140 4540
rect 410 4510 440 4540
rect 710 4510 740 4540
rect 1010 4510 1040 4540
rect 1160 4510 1190 4540
rect 1310 4510 1340 4540
rect 1610 4510 1640 4540
rect 1910 4510 1940 4540
rect 2060 4510 2090 4540
rect 2210 4510 2240 4540
rect 2510 4510 2540 4540
rect 2810 4510 2840 4540
rect 2960 4510 2990 4540
rect 3110 4510 3140 4540
rect 3410 4510 3440 4540
rect 3710 4510 3740 4540
rect 4010 4510 4040 4540
rect 4310 4510 4340 4540
rect 4610 4510 4640 4540
rect 4910 4510 4940 4540
rect 5210 4510 5240 4540
rect 5360 4510 5390 4540
rect 5510 4510 5540 4540
rect 5810 4510 5840 4540
rect 6110 4510 6140 4540
rect 6260 4510 6290 4540
rect 6410 4510 6440 4540
rect 6710 4510 6740 4540
rect 7010 4510 7040 4540
rect 7160 4510 7190 4540
rect 7310 4510 7340 4540
rect 7610 4510 7640 4540
rect 7910 4510 7940 4540
rect 8210 4510 8240 4540
rect 8510 4510 8540 4540
rect 8810 4510 8840 4540
rect 9110 4510 9140 4540
rect 9410 4510 9440 4540
rect 9710 4510 9740 4540
rect 10010 4510 10040 4540
rect 10310 4510 10340 4540
rect 10610 4510 10640 4540
rect 10910 4510 10940 4540
rect 11210 4510 11240 4540
rect 11360 4510 11390 4540
rect 11510 4510 11540 4540
rect 11810 4510 11840 4540
rect 12110 4510 12140 4540
rect 12410 4510 12440 4540
rect 12560 4510 12590 4540
rect 12710 4510 12740 4540
rect 13010 4510 13040 4540
rect 13310 4510 13340 4540
rect 13610 4510 13640 4540
rect 13760 4510 13790 4540
rect 13910 4510 13940 4540
rect 14210 4510 14240 4540
rect 14510 4510 14540 4540
rect 14810 4510 14840 4540
rect 14960 4510 14990 4540
rect 15110 4510 15140 4540
rect 15410 4510 15440 4540
rect 15710 4510 15740 4540
rect 16010 4510 16040 4540
rect 16310 4510 16340 4540
rect 16610 4510 16640 4540
rect 16760 4510 16790 4540
rect 16910 4510 16940 4540
rect 17210 4510 17240 4540
rect 17510 4510 17540 4540
rect 17810 4510 17840 4540
rect 18110 4510 18140 4540
rect 18410 4510 18440 4540
rect 18710 4510 18740 4540
rect 19010 4510 19040 4540
rect 19160 4510 19190 4540
rect 19310 4510 19340 4540
rect 19610 4510 19640 4540
rect 19910 4510 19940 4540
rect 20210 4510 20240 4540
rect -640 3860 -610 3890
rect -40 3860 -10 3890
rect 4160 3860 4190 3890
rect 8360 3860 8390 3890
rect 8660 3860 8690 3890
rect 8960 3860 8990 3890
rect 9260 3860 9290 3890
rect 9560 3860 9590 3890
rect 9860 3860 9890 3890
rect 10160 3860 10190 3890
rect 10460 3860 10490 3890
rect 10760 3860 10790 3890
rect 11960 3860 11990 3890
rect 13160 3860 13190 3890
rect 14360 3860 14390 3890
rect 15560 3860 15590 3890
rect 20360 3860 20390 3890
rect -490 3210 -460 3240
rect -340 3210 -310 3240
rect -190 3210 -160 3240
rect 110 3210 140 3240
rect 410 3210 440 3240
rect 710 3210 740 3240
rect 1010 3210 1040 3240
rect 1160 3210 1190 3240
rect 1310 3210 1340 3240
rect 1610 3210 1640 3240
rect 1910 3210 1940 3240
rect 2060 3210 2090 3240
rect 2210 3210 2240 3240
rect 2510 3210 2540 3240
rect 2810 3210 2840 3240
rect 2960 3210 2990 3240
rect 3110 3210 3140 3240
rect 3410 3210 3440 3240
rect 3710 3210 3740 3240
rect 4010 3210 4040 3240
rect 4310 3210 4340 3240
rect 4610 3210 4640 3240
rect 4910 3210 4940 3240
rect 5210 3210 5240 3240
rect 5360 3210 5390 3240
rect 5510 3210 5540 3240
rect 5810 3210 5840 3240
rect 6110 3210 6140 3240
rect 6260 3210 6290 3240
rect 6410 3210 6440 3240
rect 6710 3210 6740 3240
rect 7010 3210 7040 3240
rect 7160 3210 7190 3240
rect 7310 3210 7340 3240
rect 7610 3210 7640 3240
rect 7910 3210 7940 3240
rect 8210 3210 8240 3240
rect 8510 3210 8540 3240
rect 8810 3210 8840 3240
rect 9110 3210 9140 3240
rect 9410 3210 9440 3240
rect 9710 3210 9740 3240
rect 10010 3210 10040 3240
rect 10310 3210 10340 3240
rect 10610 3210 10640 3240
rect 10910 3210 10940 3240
rect 11210 3210 11240 3240
rect 11360 3210 11390 3240
rect 11510 3210 11540 3240
rect 11810 3210 11840 3240
rect 12110 3210 12140 3240
rect 12410 3210 12440 3240
rect 12560 3210 12590 3240
rect 12710 3210 12740 3240
rect 13010 3210 13040 3240
rect 13310 3210 13340 3240
rect 13610 3210 13640 3240
rect 13760 3210 13790 3240
rect 13910 3210 13940 3240
rect 14210 3210 14240 3240
rect 14510 3210 14540 3240
rect 14810 3210 14840 3240
rect 14960 3210 14990 3240
rect 15110 3210 15140 3240
rect 15410 3210 15440 3240
rect 15710 3210 15740 3240
rect 16010 3210 16040 3240
rect 16310 3210 16340 3240
rect 16610 3210 16640 3240
rect 16760 3210 16790 3240
rect 16910 3210 16940 3240
rect 17210 3210 17240 3240
rect 17510 3210 17540 3240
rect 17810 3210 17840 3240
rect 18110 3210 18140 3240
rect 18410 3210 18440 3240
rect 18710 3210 18740 3240
rect 19010 3210 19040 3240
rect 19160 3210 19190 3240
rect 19310 3210 19340 3240
rect 19610 3210 19640 3240
rect 19910 3210 19940 3240
rect 20210 3210 20240 3240
rect -640 2560 -610 2590
rect -40 2560 -10 2590
rect 4160 2560 4190 2590
rect 8360 2560 8390 2590
rect 8660 2560 8690 2590
rect 8960 2560 8990 2590
rect 9260 2560 9290 2590
rect 9560 2560 9590 2590
rect 9860 2560 9890 2590
rect 10160 2560 10190 2590
rect 10460 2560 10490 2590
rect 10760 2560 10790 2590
rect 11960 2560 11990 2590
rect 13160 2560 13190 2590
rect 14360 2560 14390 2590
rect 15560 2560 15590 2590
rect 17960 2560 17990 2590
rect 20360 2560 20390 2590
rect -640 1660 -610 1690
rect -40 1660 -10 1690
rect 8360 1660 8390 1690
rect 10760 1660 10790 1690
rect 15560 1660 15590 1690
rect 17960 1660 17990 1690
rect 20360 1660 20390 1690
rect -640 1610 -610 1640
rect -40 1610 -10 1640
rect 8360 1610 8390 1640
rect 10760 1610 10790 1640
rect 15560 1610 15590 1640
rect 17960 1610 17990 1640
rect 20360 1610 20390 1640
rect -490 810 -460 840
rect -340 810 -310 840
rect -190 810 -160 840
rect 110 810 140 840
rect 410 810 440 840
rect 710 810 740 840
rect 1010 810 1040 840
rect 1310 810 1340 840
rect 1610 810 1640 840
rect 1910 810 1940 840
rect 2210 810 2240 840
rect 2360 810 2390 840
rect 2510 810 2540 840
rect 2810 810 2840 840
rect 3110 810 3140 840
rect 3410 810 3440 840
rect 3710 810 3740 840
rect 3860 810 3890 840
rect 4010 810 4040 840
rect 4310 810 4340 840
rect 4460 810 4490 840
rect 4610 810 4640 840
rect 4910 810 4940 840
rect 5210 810 5240 840
rect 5510 810 5540 840
rect 5810 810 5840 840
rect 5960 810 5990 840
rect 6110 810 6140 840
rect 6410 810 6440 840
rect 6710 810 6740 840
rect 7010 810 7040 840
rect 7310 810 7340 840
rect 7610 810 7640 840
rect 7910 810 7940 840
rect 8210 810 8240 840
rect 8510 810 8540 840
rect 8810 810 8840 840
rect 9110 810 9140 840
rect 9410 810 9440 840
rect 9560 810 9590 840
rect 9710 810 9740 840
rect 10010 810 10040 840
rect 10310 810 10340 840
rect 10610 810 10640 840
rect 10910 810 10940 840
rect 11210 810 11240 840
rect 11510 810 11540 840
rect 11810 810 11840 840
rect 12110 810 12140 840
rect 12410 810 12440 840
rect 12560 810 12590 840
rect 12710 810 12740 840
rect 13010 810 13040 840
rect 13160 810 13190 840
rect 13310 810 13340 840
rect 13610 810 13640 840
rect 13760 810 13790 840
rect 13910 810 13940 840
rect 14210 810 14240 840
rect 14510 810 14540 840
rect 14810 810 14840 840
rect 15110 810 15140 840
rect 15410 810 15440 840
rect 15710 810 15740 840
rect 16010 810 16040 840
rect 16310 810 16340 840
rect 16610 810 16640 840
rect 16760 810 16790 840
rect 16910 810 16940 840
rect 17210 810 17240 840
rect 17510 810 17540 840
rect 17810 810 17840 840
rect 18110 810 18140 840
rect 18410 810 18440 840
rect 18710 810 18740 840
rect 19010 810 19040 840
rect 19160 810 19190 840
rect 19310 810 19340 840
rect 19610 810 19640 840
rect 19910 810 19940 840
rect 20210 810 20240 840
rect -640 10 -610 40
rect -40 10 -10 40
rect 8360 10 8390 40
rect 10760 10 10790 40
rect 15560 10 15590 40
rect 17960 10 17990 40
rect 20360 10 20390 40
rect -640 -40 -610 -10
rect -40 -40 -10 -10
rect 8360 -40 8390 -10
rect 10760 -40 10790 -10
rect 15560 -40 15590 -10
rect 17960 -40 17990 -10
rect 20360 -40 20390 -10
rect -640 -90 -610 -60
rect -40 -90 -10 -60
rect 8360 -90 8390 -60
rect 10760 -90 10790 -60
rect 15560 -90 15590 -60
rect 17960 -90 17990 -60
rect 20360 -90 20390 -60
rect -490 -890 -460 -860
rect -340 -890 -310 -860
rect -190 -890 -160 -860
rect 110 -890 140 -860
rect 410 -890 440 -860
rect 710 -890 740 -860
rect 1010 -890 1040 -860
rect 1310 -890 1340 -860
rect 1610 -890 1640 -860
rect 1910 -890 1940 -860
rect 2210 -890 2240 -860
rect 2360 -890 2390 -860
rect 2510 -890 2540 -860
rect 2810 -890 2840 -860
rect 3110 -890 3140 -860
rect 3410 -890 3440 -860
rect 3710 -890 3740 -860
rect 3860 -890 3890 -860
rect 4010 -890 4040 -860
rect 4310 -890 4340 -860
rect 4460 -890 4490 -860
rect 4610 -890 4640 -860
rect 4910 -890 4940 -860
rect 5210 -890 5240 -860
rect 5510 -890 5540 -860
rect 5810 -890 5840 -860
rect 5960 -890 5990 -860
rect 6110 -890 6140 -860
rect 6410 -890 6440 -860
rect 6710 -890 6740 -860
rect 7010 -890 7040 -860
rect 7310 -890 7340 -860
rect 7610 -890 7640 -860
rect 7910 -890 7940 -860
rect 8210 -890 8240 -860
rect 8510 -890 8540 -860
rect 8810 -890 8840 -860
rect 9110 -890 9140 -860
rect 9410 -890 9440 -860
rect 9560 -890 9590 -860
rect 9710 -890 9740 -860
rect 10010 -890 10040 -860
rect 10310 -890 10340 -860
rect 10610 -890 10640 -860
rect 10910 -890 10940 -860
rect 11210 -890 11240 -860
rect 11510 -890 11540 -860
rect 11810 -890 11840 -860
rect 12110 -890 12140 -860
rect 12410 -890 12440 -860
rect 12560 -890 12590 -860
rect 12710 -890 12740 -860
rect 13010 -890 13040 -860
rect 13160 -890 13190 -860
rect 13310 -890 13340 -860
rect 13610 -890 13640 -860
rect 13760 -890 13790 -860
rect 13910 -890 13940 -860
rect 14210 -890 14240 -860
rect 14510 -890 14540 -860
rect 14810 -890 14840 -860
rect 15110 -890 15140 -860
rect 15410 -890 15440 -860
rect 15710 -890 15740 -860
rect 16010 -890 16040 -860
rect 16310 -890 16340 -860
rect 16610 -890 16640 -860
rect 16760 -890 16790 -860
rect 16910 -890 16940 -860
rect 17210 -890 17240 -860
rect 17510 -890 17540 -860
rect 17810 -890 17840 -860
rect 18110 -890 18140 -860
rect 18410 -890 18440 -860
rect 18710 -890 18740 -860
rect 19010 -890 19040 -860
rect 19160 -890 19190 -860
rect 19310 -890 19340 -860
rect 19610 -890 19640 -860
rect 19910 -890 19940 -860
rect 20210 -890 20240 -860
rect -640 -1690 -610 -1660
rect -40 -1690 -10 -1660
rect 8360 -1690 8390 -1660
rect 10760 -1690 10790 -1660
rect 15560 -1690 15590 -1660
rect 17960 -1690 17990 -1660
rect 20360 -1690 20390 -1660
rect -640 -1740 -610 -1710
rect -40 -1740 -10 -1710
rect 8360 -1740 8390 -1710
rect 10760 -1740 10790 -1710
rect 15560 -1740 15590 -1710
rect 17960 -1740 17990 -1710
rect 20360 -1740 20390 -1710
<< metal3 >>
rect -650 5190 20400 5200
rect -650 5160 -640 5190
rect -610 5160 8360 5190
rect 8390 5160 8660 5190
rect 8690 5160 8960 5190
rect 8990 5160 9260 5190
rect 9290 5160 9560 5190
rect 9590 5160 9860 5190
rect 9890 5160 10160 5190
rect 10190 5160 10460 5190
rect 10490 5160 10760 5190
rect 10790 5160 11960 5190
rect 11990 5160 13160 5190
rect 13190 5160 14360 5190
rect 14390 5160 15560 5190
rect 15590 5160 17960 5190
rect 17990 5160 20360 5190
rect 20390 5160 20400 5190
rect -650 5100 20400 5160
rect -650 5000 20400 5050
rect -650 4900 20400 4950
rect -650 4800 20400 4850
rect -650 4700 20400 4750
rect -650 4600 20400 4650
rect -500 4545 -450 4550
rect -500 4505 -495 4545
rect -455 4505 -450 4545
rect -500 4500 -450 4505
rect -350 4545 -300 4550
rect -350 4505 -345 4545
rect -305 4505 -300 4545
rect -350 4500 -300 4505
rect -200 4545 -150 4550
rect -200 4505 -195 4545
rect -155 4505 -150 4545
rect -200 4500 -150 4505
rect 100 4545 150 4550
rect 100 4505 105 4545
rect 145 4505 150 4545
rect 100 4500 150 4505
rect 400 4545 450 4550
rect 400 4505 405 4545
rect 445 4505 450 4545
rect 400 4500 450 4505
rect 700 4545 750 4550
rect 700 4505 705 4545
rect 745 4505 750 4545
rect 700 4500 750 4505
rect 1000 4545 1050 4550
rect 1000 4505 1005 4545
rect 1045 4505 1050 4545
rect 1000 4500 1050 4505
rect 1150 4545 1200 4550
rect 1150 4505 1155 4545
rect 1195 4505 1200 4545
rect 1150 4500 1200 4505
rect 1300 4545 1350 4550
rect 1300 4505 1305 4545
rect 1345 4505 1350 4545
rect 1300 4500 1350 4505
rect 1600 4545 1650 4550
rect 1600 4505 1605 4545
rect 1645 4505 1650 4545
rect 1600 4500 1650 4505
rect 1900 4545 1950 4550
rect 1900 4505 1905 4545
rect 1945 4505 1950 4545
rect 1900 4500 1950 4505
rect 2050 4545 2100 4550
rect 2050 4505 2055 4545
rect 2095 4505 2100 4545
rect 2050 4500 2100 4505
rect 2200 4545 2250 4550
rect 2200 4505 2205 4545
rect 2245 4505 2250 4545
rect 2200 4500 2250 4505
rect 2500 4545 2550 4550
rect 2500 4505 2505 4545
rect 2545 4505 2550 4545
rect 2500 4500 2550 4505
rect 2800 4545 2850 4550
rect 2800 4505 2805 4545
rect 2845 4505 2850 4545
rect 2800 4500 2850 4505
rect 2950 4545 3000 4550
rect 2950 4505 2955 4545
rect 2995 4505 3000 4545
rect 2950 4500 3000 4505
rect 3100 4545 3150 4550
rect 3100 4505 3105 4545
rect 3145 4505 3150 4545
rect 3100 4500 3150 4505
rect 3400 4545 3450 4550
rect 3400 4505 3405 4545
rect 3445 4505 3450 4545
rect 3400 4500 3450 4505
rect 3700 4545 3750 4550
rect 3700 4505 3705 4545
rect 3745 4505 3750 4545
rect 3700 4500 3750 4505
rect 4000 4545 4050 4550
rect 4000 4505 4005 4545
rect 4045 4505 4050 4545
rect 4000 4500 4050 4505
rect 4300 4545 4350 4550
rect 4300 4505 4305 4545
rect 4345 4505 4350 4545
rect 4300 4500 4350 4505
rect 4600 4545 4650 4550
rect 4600 4505 4605 4545
rect 4645 4505 4650 4545
rect 4600 4500 4650 4505
rect 4900 4545 4950 4550
rect 4900 4505 4905 4545
rect 4945 4505 4950 4545
rect 4900 4500 4950 4505
rect 5200 4545 5250 4550
rect 5200 4505 5205 4545
rect 5245 4505 5250 4545
rect 5200 4500 5250 4505
rect 5350 4545 5400 4550
rect 5350 4505 5355 4545
rect 5395 4505 5400 4545
rect 5350 4500 5400 4505
rect 5500 4545 5550 4550
rect 5500 4505 5505 4545
rect 5545 4505 5550 4545
rect 5500 4500 5550 4505
rect 5800 4545 5850 4550
rect 5800 4505 5805 4545
rect 5845 4505 5850 4545
rect 5800 4500 5850 4505
rect 6100 4545 6150 4550
rect 6100 4505 6105 4545
rect 6145 4505 6150 4545
rect 6100 4500 6150 4505
rect 6250 4545 6300 4550
rect 6250 4505 6255 4545
rect 6295 4505 6300 4545
rect 6250 4500 6300 4505
rect 6400 4545 6450 4550
rect 6400 4505 6405 4545
rect 6445 4505 6450 4545
rect 6400 4500 6450 4505
rect 6700 4545 6750 4550
rect 6700 4505 6705 4545
rect 6745 4505 6750 4545
rect 6700 4500 6750 4505
rect 7000 4545 7050 4550
rect 7000 4505 7005 4545
rect 7045 4505 7050 4545
rect 7000 4500 7050 4505
rect 7150 4545 7200 4550
rect 7150 4505 7155 4545
rect 7195 4505 7200 4545
rect 7150 4500 7200 4505
rect 7300 4545 7350 4550
rect 7300 4505 7305 4545
rect 7345 4505 7350 4545
rect 7300 4500 7350 4505
rect 7600 4545 7650 4550
rect 7600 4505 7605 4545
rect 7645 4505 7650 4545
rect 7600 4500 7650 4505
rect 7900 4545 7950 4550
rect 7900 4505 7905 4545
rect 7945 4505 7950 4545
rect 7900 4500 7950 4505
rect 8200 4545 8250 4550
rect 8200 4505 8205 4545
rect 8245 4505 8250 4545
rect 8200 4500 8250 4505
rect 8500 4545 8550 4550
rect 8500 4505 8505 4545
rect 8545 4505 8550 4545
rect 8500 4500 8550 4505
rect 8800 4545 8850 4550
rect 8800 4505 8805 4545
rect 8845 4505 8850 4545
rect 8800 4500 8850 4505
rect 9100 4545 9150 4550
rect 9100 4505 9105 4545
rect 9145 4505 9150 4545
rect 9100 4500 9150 4505
rect 9400 4545 9450 4550
rect 9400 4505 9405 4545
rect 9445 4505 9450 4545
rect 9400 4500 9450 4505
rect 9700 4545 9750 4550
rect 9700 4505 9705 4545
rect 9745 4505 9750 4545
rect 9700 4500 9750 4505
rect 10000 4545 10050 4550
rect 10000 4505 10005 4545
rect 10045 4505 10050 4545
rect 10000 4500 10050 4505
rect 10300 4545 10350 4550
rect 10300 4505 10305 4545
rect 10345 4505 10350 4545
rect 10300 4500 10350 4505
rect 10600 4545 10650 4550
rect 10600 4505 10605 4545
rect 10645 4505 10650 4545
rect 10600 4500 10650 4505
rect 10900 4545 10950 4550
rect 10900 4505 10905 4545
rect 10945 4505 10950 4545
rect 10900 4500 10950 4505
rect 11200 4545 11250 4550
rect 11200 4505 11205 4545
rect 11245 4505 11250 4545
rect 11200 4500 11250 4505
rect 11350 4545 11400 4550
rect 11350 4505 11355 4545
rect 11395 4505 11400 4545
rect 11350 4500 11400 4505
rect 11500 4545 11550 4550
rect 11500 4505 11505 4545
rect 11545 4505 11550 4545
rect 11500 4500 11550 4505
rect 11800 4545 11850 4550
rect 11800 4505 11805 4545
rect 11845 4505 11850 4545
rect 11800 4500 11850 4505
rect 12100 4545 12150 4550
rect 12100 4505 12105 4545
rect 12145 4505 12150 4545
rect 12100 4500 12150 4505
rect 12400 4545 12450 4550
rect 12400 4505 12405 4545
rect 12445 4505 12450 4545
rect 12400 4500 12450 4505
rect 12550 4545 12600 4550
rect 12550 4505 12555 4545
rect 12595 4505 12600 4545
rect 12550 4500 12600 4505
rect 12700 4545 12750 4550
rect 12700 4505 12705 4545
rect 12745 4505 12750 4545
rect 12700 4500 12750 4505
rect 13000 4545 13050 4550
rect 13000 4505 13005 4545
rect 13045 4505 13050 4545
rect 13000 4500 13050 4505
rect 13300 4545 13350 4550
rect 13300 4505 13305 4545
rect 13345 4505 13350 4545
rect 13300 4500 13350 4505
rect 13600 4545 13650 4550
rect 13600 4505 13605 4545
rect 13645 4505 13650 4545
rect 13600 4500 13650 4505
rect 13750 4545 13800 4550
rect 13750 4505 13755 4545
rect 13795 4505 13800 4545
rect 13750 4500 13800 4505
rect 13900 4545 13950 4550
rect 13900 4505 13905 4545
rect 13945 4505 13950 4545
rect 13900 4500 13950 4505
rect 14200 4545 14250 4550
rect 14200 4505 14205 4545
rect 14245 4505 14250 4545
rect 14200 4500 14250 4505
rect 14500 4545 14550 4550
rect 14500 4505 14505 4545
rect 14545 4505 14550 4545
rect 14500 4500 14550 4505
rect 14800 4545 14850 4550
rect 14800 4505 14805 4545
rect 14845 4505 14850 4545
rect 14800 4500 14850 4505
rect 14950 4545 15000 4550
rect 14950 4505 14955 4545
rect 14995 4505 15000 4545
rect 14950 4500 15000 4505
rect 15100 4545 15150 4550
rect 15100 4505 15105 4545
rect 15145 4505 15150 4545
rect 15100 4500 15150 4505
rect 15400 4545 15450 4550
rect 15400 4505 15405 4545
rect 15445 4505 15450 4545
rect 15400 4500 15450 4505
rect 15700 4545 15750 4550
rect 15700 4505 15705 4545
rect 15745 4505 15750 4545
rect 15700 4500 15750 4505
rect 16000 4545 16050 4550
rect 16000 4505 16005 4545
rect 16045 4505 16050 4545
rect 16000 4500 16050 4505
rect 16300 4545 16350 4550
rect 16300 4505 16305 4545
rect 16345 4505 16350 4545
rect 16300 4500 16350 4505
rect 16600 4545 16650 4550
rect 16600 4505 16605 4545
rect 16645 4505 16650 4545
rect 16600 4500 16650 4505
rect 16750 4545 16800 4550
rect 16750 4505 16755 4545
rect 16795 4505 16800 4545
rect 16750 4500 16800 4505
rect 16900 4545 16950 4550
rect 16900 4505 16905 4545
rect 16945 4505 16950 4545
rect 16900 4500 16950 4505
rect 17200 4545 17250 4550
rect 17200 4505 17205 4545
rect 17245 4505 17250 4545
rect 17200 4500 17250 4505
rect 17500 4545 17550 4550
rect 17500 4505 17505 4545
rect 17545 4505 17550 4545
rect 17500 4500 17550 4505
rect 17800 4545 17850 4550
rect 17800 4505 17805 4545
rect 17845 4505 17850 4545
rect 17800 4500 17850 4505
rect 18100 4545 18150 4550
rect 18100 4505 18105 4545
rect 18145 4505 18150 4545
rect 18100 4500 18150 4505
rect 18400 4545 18450 4550
rect 18400 4505 18405 4545
rect 18445 4505 18450 4545
rect 18400 4500 18450 4505
rect 18700 4545 18750 4550
rect 18700 4505 18705 4545
rect 18745 4505 18750 4545
rect 18700 4500 18750 4505
rect 19000 4545 19050 4550
rect 19000 4505 19005 4545
rect 19045 4505 19050 4545
rect 19000 4500 19050 4505
rect 19150 4545 19200 4550
rect 19150 4505 19155 4545
rect 19195 4505 19200 4545
rect 19150 4500 19200 4505
rect 19300 4545 19350 4550
rect 19300 4505 19305 4545
rect 19345 4505 19350 4545
rect 19300 4500 19350 4505
rect 19600 4545 19650 4550
rect 19600 4505 19605 4545
rect 19645 4505 19650 4545
rect 19600 4500 19650 4505
rect 19900 4545 19950 4550
rect 19900 4505 19905 4545
rect 19945 4505 19950 4545
rect 19900 4500 19950 4505
rect 20200 4545 20250 4550
rect 20200 4505 20205 4545
rect 20245 4505 20250 4545
rect 20200 4500 20250 4505
rect -650 4400 20400 4450
rect -650 4345 20400 4350
rect -650 4305 13755 4345
rect 13795 4305 14955 4345
rect 14995 4305 20400 4345
rect -650 4300 20400 4305
rect -650 4200 20400 4250
rect -650 4145 20400 4150
rect -650 4105 11355 4145
rect 11395 4105 12555 4145
rect 12595 4105 20400 4145
rect -650 4100 20400 4105
rect -650 4000 20400 4050
rect -650 3890 20400 3950
rect -650 3860 -640 3890
rect -610 3860 -40 3890
rect -10 3860 4160 3890
rect 4190 3860 8360 3890
rect 8390 3860 8660 3890
rect 8690 3860 8960 3890
rect 8990 3860 9260 3890
rect 9290 3860 9560 3890
rect 9590 3860 9860 3890
rect 9890 3860 10160 3890
rect 10190 3860 10460 3890
rect 10490 3860 10760 3890
rect 10790 3860 11960 3890
rect 11990 3860 13160 3890
rect 13190 3860 14360 3890
rect 14390 3860 15560 3890
rect 15590 3860 20360 3890
rect 20390 3860 20400 3890
rect -650 3800 20400 3860
rect -650 3700 20400 3750
rect -650 3645 20400 3650
rect -650 3605 13305 3645
rect 13345 3605 13605 3645
rect 13645 3605 13905 3645
rect 13945 3605 14205 3645
rect 14245 3605 14505 3645
rect 14545 3605 14805 3645
rect 14845 3605 15105 3645
rect 15145 3605 15405 3645
rect 15445 3605 20400 3645
rect -650 3600 20400 3605
rect -650 3500 20400 3550
rect -650 3445 20400 3450
rect -650 3405 10905 3445
rect 10945 3405 11205 3445
rect 11245 3405 11505 3445
rect 11545 3405 11805 3445
rect 11845 3405 12105 3445
rect 12145 3405 12405 3445
rect 12445 3405 12705 3445
rect 12745 3405 13005 3445
rect 13045 3405 20400 3445
rect -650 3400 20400 3405
rect -650 3300 20400 3350
rect -500 3245 -450 3250
rect -500 3205 -495 3245
rect -455 3205 -450 3245
rect -500 3200 -450 3205
rect -350 3245 -300 3250
rect -350 3205 -345 3245
rect -305 3205 -300 3245
rect -350 3200 -300 3205
rect -200 3245 -150 3250
rect -200 3205 -195 3245
rect -155 3205 -150 3245
rect -200 3200 -150 3205
rect 100 3245 150 3250
rect 100 3205 105 3245
rect 145 3205 150 3245
rect 100 3200 150 3205
rect 400 3245 450 3250
rect 400 3205 405 3245
rect 445 3205 450 3245
rect 400 3200 450 3205
rect 700 3245 750 3250
rect 700 3205 705 3245
rect 745 3205 750 3245
rect 700 3200 750 3205
rect 1000 3245 1050 3250
rect 1000 3205 1005 3245
rect 1045 3205 1050 3245
rect 1000 3200 1050 3205
rect 1150 3245 1200 3250
rect 1150 3205 1155 3245
rect 1195 3205 1200 3245
rect 1150 3200 1200 3205
rect 1300 3245 1350 3250
rect 1300 3205 1305 3245
rect 1345 3205 1350 3245
rect 1300 3200 1350 3205
rect 1600 3245 1650 3250
rect 1600 3205 1605 3245
rect 1645 3205 1650 3245
rect 1600 3200 1650 3205
rect 1900 3245 1950 3250
rect 1900 3205 1905 3245
rect 1945 3205 1950 3245
rect 1900 3200 1950 3205
rect 2050 3245 2100 3250
rect 2050 3205 2055 3245
rect 2095 3205 2100 3245
rect 2050 3200 2100 3205
rect 2200 3245 2250 3250
rect 2200 3205 2205 3245
rect 2245 3205 2250 3245
rect 2200 3200 2250 3205
rect 2500 3245 2550 3250
rect 2500 3205 2505 3245
rect 2545 3205 2550 3245
rect 2500 3200 2550 3205
rect 2800 3245 2850 3250
rect 2800 3205 2805 3245
rect 2845 3205 2850 3245
rect 2800 3200 2850 3205
rect 2950 3245 3000 3250
rect 2950 3205 2955 3245
rect 2995 3205 3000 3245
rect 2950 3200 3000 3205
rect 3100 3245 3150 3250
rect 3100 3205 3105 3245
rect 3145 3205 3150 3245
rect 3100 3200 3150 3205
rect 3400 3245 3450 3250
rect 3400 3205 3405 3245
rect 3445 3205 3450 3245
rect 3400 3200 3450 3205
rect 3700 3245 3750 3250
rect 3700 3205 3705 3245
rect 3745 3205 3750 3245
rect 3700 3200 3750 3205
rect 4000 3245 4050 3250
rect 4000 3205 4005 3245
rect 4045 3205 4050 3245
rect 4000 3200 4050 3205
rect 4300 3245 4350 3250
rect 4300 3205 4305 3245
rect 4345 3205 4350 3245
rect 4300 3200 4350 3205
rect 4600 3245 4650 3250
rect 4600 3205 4605 3245
rect 4645 3205 4650 3245
rect 4600 3200 4650 3205
rect 4900 3245 4950 3250
rect 4900 3205 4905 3245
rect 4945 3205 4950 3245
rect 4900 3200 4950 3205
rect 5200 3245 5250 3250
rect 5200 3205 5205 3245
rect 5245 3205 5250 3245
rect 5200 3200 5250 3205
rect 5350 3245 5400 3250
rect 5350 3205 5355 3245
rect 5395 3205 5400 3245
rect 5350 3200 5400 3205
rect 5500 3245 5550 3250
rect 5500 3205 5505 3245
rect 5545 3205 5550 3245
rect 5500 3200 5550 3205
rect 5800 3245 5850 3250
rect 5800 3205 5805 3245
rect 5845 3205 5850 3245
rect 5800 3200 5850 3205
rect 6100 3245 6150 3250
rect 6100 3205 6105 3245
rect 6145 3205 6150 3245
rect 6100 3200 6150 3205
rect 6250 3245 6300 3250
rect 6250 3205 6255 3245
rect 6295 3205 6300 3245
rect 6250 3200 6300 3205
rect 6400 3245 6450 3250
rect 6400 3205 6405 3245
rect 6445 3205 6450 3245
rect 6400 3200 6450 3205
rect 6700 3245 6750 3250
rect 6700 3205 6705 3245
rect 6745 3205 6750 3245
rect 6700 3200 6750 3205
rect 7000 3245 7050 3250
rect 7000 3205 7005 3245
rect 7045 3205 7050 3245
rect 7000 3200 7050 3205
rect 7150 3245 7200 3250
rect 7150 3205 7155 3245
rect 7195 3205 7200 3245
rect 7150 3200 7200 3205
rect 7300 3245 7350 3250
rect 7300 3205 7305 3245
rect 7345 3205 7350 3245
rect 7300 3200 7350 3205
rect 7600 3245 7650 3250
rect 7600 3205 7605 3245
rect 7645 3205 7650 3245
rect 7600 3200 7650 3205
rect 7900 3245 7950 3250
rect 7900 3205 7905 3245
rect 7945 3205 7950 3245
rect 7900 3200 7950 3205
rect 8200 3245 8250 3250
rect 8200 3205 8205 3245
rect 8245 3205 8250 3245
rect 8200 3200 8250 3205
rect 8500 3245 8550 3250
rect 8500 3205 8505 3245
rect 8545 3205 8550 3245
rect 8500 3200 8550 3205
rect 8800 3245 8850 3250
rect 8800 3205 8805 3245
rect 8845 3205 8850 3245
rect 8800 3200 8850 3205
rect 9100 3245 9150 3250
rect 9100 3205 9105 3245
rect 9145 3205 9150 3245
rect 9100 3200 9150 3205
rect 9400 3245 9450 3250
rect 9400 3205 9405 3245
rect 9445 3205 9450 3245
rect 9400 3200 9450 3205
rect 9700 3245 9750 3250
rect 9700 3205 9705 3245
rect 9745 3205 9750 3245
rect 9700 3200 9750 3205
rect 10000 3245 10050 3250
rect 10000 3205 10005 3245
rect 10045 3205 10050 3245
rect 10000 3200 10050 3205
rect 10300 3245 10350 3250
rect 10300 3205 10305 3245
rect 10345 3205 10350 3245
rect 10300 3200 10350 3205
rect 10600 3245 10650 3250
rect 10600 3205 10605 3245
rect 10645 3205 10650 3245
rect 10600 3200 10650 3205
rect 10900 3245 10950 3250
rect 10900 3205 10905 3245
rect 10945 3205 10950 3245
rect 10900 3200 10950 3205
rect 11200 3245 11250 3250
rect 11200 3205 11205 3245
rect 11245 3205 11250 3245
rect 11200 3200 11250 3205
rect 11350 3245 11400 3250
rect 11350 3205 11355 3245
rect 11395 3205 11400 3245
rect 11350 3200 11400 3205
rect 11500 3245 11550 3250
rect 11500 3205 11505 3245
rect 11545 3205 11550 3245
rect 11500 3200 11550 3205
rect 11800 3245 11850 3250
rect 11800 3205 11805 3245
rect 11845 3205 11850 3245
rect 11800 3200 11850 3205
rect 12100 3245 12150 3250
rect 12100 3205 12105 3245
rect 12145 3205 12150 3245
rect 12100 3200 12150 3205
rect 12400 3245 12450 3250
rect 12400 3205 12405 3245
rect 12445 3205 12450 3245
rect 12400 3200 12450 3205
rect 12550 3245 12600 3250
rect 12550 3205 12555 3245
rect 12595 3205 12600 3245
rect 12550 3200 12600 3205
rect 12700 3245 12750 3250
rect 12700 3205 12705 3245
rect 12745 3205 12750 3245
rect 12700 3200 12750 3205
rect 13000 3245 13050 3250
rect 13000 3205 13005 3245
rect 13045 3205 13050 3245
rect 13000 3200 13050 3205
rect 13300 3245 13350 3250
rect 13300 3205 13305 3245
rect 13345 3205 13350 3245
rect 13300 3200 13350 3205
rect 13600 3245 13650 3250
rect 13600 3205 13605 3245
rect 13645 3205 13650 3245
rect 13600 3200 13650 3205
rect 13750 3245 13800 3250
rect 13750 3205 13755 3245
rect 13795 3205 13800 3245
rect 13750 3200 13800 3205
rect 13900 3245 13950 3250
rect 13900 3205 13905 3245
rect 13945 3205 13950 3245
rect 13900 3200 13950 3205
rect 14200 3245 14250 3250
rect 14200 3205 14205 3245
rect 14245 3205 14250 3245
rect 14200 3200 14250 3205
rect 14500 3245 14550 3250
rect 14500 3205 14505 3245
rect 14545 3205 14550 3245
rect 14500 3200 14550 3205
rect 14800 3245 14850 3250
rect 14800 3205 14805 3245
rect 14845 3205 14850 3245
rect 14800 3200 14850 3205
rect 14950 3245 15000 3250
rect 14950 3205 14955 3245
rect 14995 3205 15000 3245
rect 14950 3200 15000 3205
rect 15100 3245 15150 3250
rect 15100 3205 15105 3245
rect 15145 3205 15150 3245
rect 15100 3200 15150 3205
rect 15400 3245 15450 3250
rect 15400 3205 15405 3245
rect 15445 3205 15450 3245
rect 15400 3200 15450 3205
rect 15700 3245 15750 3250
rect 15700 3205 15705 3245
rect 15745 3205 15750 3245
rect 15700 3200 15750 3205
rect 16000 3245 16050 3250
rect 16000 3205 16005 3245
rect 16045 3205 16050 3245
rect 16000 3200 16050 3205
rect 16300 3245 16350 3250
rect 16300 3205 16305 3245
rect 16345 3205 16350 3245
rect 16300 3200 16350 3205
rect 16600 3245 16650 3250
rect 16600 3205 16605 3245
rect 16645 3205 16650 3245
rect 16600 3200 16650 3205
rect 16750 3245 16800 3250
rect 16750 3205 16755 3245
rect 16795 3205 16800 3245
rect 16750 3200 16800 3205
rect 16900 3245 16950 3250
rect 16900 3205 16905 3245
rect 16945 3205 16950 3245
rect 16900 3200 16950 3205
rect 17200 3245 17250 3250
rect 17200 3205 17205 3245
rect 17245 3205 17250 3245
rect 17200 3200 17250 3205
rect 17500 3245 17550 3250
rect 17500 3205 17505 3245
rect 17545 3205 17550 3245
rect 17500 3200 17550 3205
rect 17800 3245 17850 3250
rect 17800 3205 17805 3245
rect 17845 3205 17850 3245
rect 17800 3200 17850 3205
rect 18100 3245 18150 3250
rect 18100 3205 18105 3245
rect 18145 3205 18150 3245
rect 18100 3200 18150 3205
rect 18400 3245 18450 3250
rect 18400 3205 18405 3245
rect 18445 3205 18450 3245
rect 18400 3200 18450 3205
rect 18700 3245 18750 3250
rect 18700 3205 18705 3245
rect 18745 3205 18750 3245
rect 18700 3200 18750 3205
rect 19000 3245 19050 3250
rect 19000 3205 19005 3245
rect 19045 3205 19050 3245
rect 19000 3200 19050 3205
rect 19150 3245 19200 3250
rect 19150 3205 19155 3245
rect 19195 3205 19200 3245
rect 19150 3200 19200 3205
rect 19300 3245 19350 3250
rect 19300 3205 19305 3245
rect 19345 3205 19350 3245
rect 19300 3200 19350 3205
rect 19600 3245 19650 3250
rect 19600 3205 19605 3245
rect 19645 3205 19650 3245
rect 19600 3200 19650 3205
rect 19900 3245 19950 3250
rect 19900 3205 19905 3245
rect 19945 3205 19950 3245
rect 19900 3200 19950 3205
rect 20200 3245 20250 3250
rect 20200 3205 20205 3245
rect 20245 3205 20250 3245
rect 20200 3200 20250 3205
rect -650 3100 20400 3150
rect -650 3045 20400 3050
rect -650 3005 -345 3045
rect -305 3005 105 3045
rect 145 3005 405 3045
rect 445 3005 2055 3045
rect 2095 3005 3705 3045
rect 3745 3005 4005 3045
rect 4045 3005 4305 3045
rect 4345 3005 4605 3045
rect 4645 3005 6255 3045
rect 6295 3005 7905 3045
rect 7945 3005 8205 3045
rect 8245 3005 20400 3045
rect -650 3000 20400 3005
rect -650 2945 20400 2950
rect -650 2905 705 2945
rect 745 2905 1005 2945
rect 1045 2905 1155 2945
rect 1195 2905 1305 2945
rect 1345 2905 1605 2945
rect 1645 2905 2505 2945
rect 2545 2905 2805 2945
rect 2845 2905 2955 2945
rect 2995 2905 3105 2945
rect 3145 2905 3405 2945
rect 3445 2905 4905 2945
rect 4945 2905 5205 2945
rect 5245 2905 5355 2945
rect 5395 2905 5505 2945
rect 5545 2905 5805 2945
rect 5845 2905 6705 2945
rect 6745 2905 7005 2945
rect 7045 2905 7155 2945
rect 7195 2905 7305 2945
rect 7345 2905 7605 2945
rect 7645 2905 9555 2945
rect 9595 2905 20400 2945
rect -650 2900 20400 2905
rect -650 2845 20400 2850
rect -650 2805 1905 2845
rect 1945 2805 2205 2845
rect 2245 2805 6105 2845
rect 6145 2805 6405 2845
rect 6445 2805 20400 2845
rect -650 2800 20400 2805
rect -650 2745 20400 2750
rect -650 2705 -495 2745
rect -455 2705 -195 2745
rect -155 2705 20400 2745
rect -650 2700 20400 2705
rect -650 2590 20400 2650
rect -650 2560 -640 2590
rect -610 2560 -40 2590
rect -10 2560 4160 2590
rect 4190 2560 8360 2590
rect 8390 2560 8660 2590
rect 8690 2560 8960 2590
rect 8990 2560 9260 2590
rect 9290 2560 9560 2590
rect 9590 2560 9860 2590
rect 9890 2560 10160 2590
rect 10190 2560 10460 2590
rect 10490 2560 10760 2590
rect 10790 2560 11960 2590
rect 11990 2560 13160 2590
rect 13190 2560 14360 2590
rect 14390 2560 15560 2590
rect 15590 2560 17960 2590
rect 17990 2560 20360 2590
rect 20390 2560 20400 2590
rect -650 2550 20400 2560
rect -900 2400 20400 2450
rect -900 2345 20400 2350
rect -900 2305 13305 2345
rect 13345 2305 13605 2345
rect 13645 2305 13905 2345
rect 13945 2305 14205 2345
rect 14245 2305 18705 2345
rect 18745 2305 19005 2345
rect 19045 2305 19305 2345
rect 19345 2305 19605 2345
rect 19645 2305 20400 2345
rect -900 2300 20400 2305
rect -900 2200 20400 2250
rect -900 2145 20400 2150
rect -900 2105 12105 2145
rect 12145 2105 12405 2145
rect 12445 2105 12705 2145
rect 12745 2105 13005 2145
rect 13045 2105 16305 2145
rect 16345 2105 16605 2145
rect 16645 2105 16905 2145
rect 16945 2105 17205 2145
rect 17245 2105 20400 2145
rect -900 2100 20400 2105
rect -900 2000 20400 2050
rect -900 1690 20400 1700
rect -900 1660 -640 1690
rect -610 1660 -40 1690
rect -10 1660 8360 1690
rect 8390 1660 10760 1690
rect 10790 1660 15560 1690
rect 15590 1660 17960 1690
rect 17990 1660 20360 1690
rect 20390 1660 20400 1690
rect -900 1640 20400 1660
rect -900 1610 -640 1640
rect -610 1610 -40 1640
rect -10 1610 8360 1640
rect 8390 1610 10760 1640
rect 10790 1610 15560 1640
rect 15590 1610 17960 1640
rect 17990 1610 20360 1640
rect 20390 1610 20400 1640
rect -900 1600 20400 1610
rect -900 1500 20400 1550
rect -900 1400 20400 1450
rect -900 1345 20400 1350
rect -900 1305 -495 1345
rect -455 1305 -195 1345
rect -155 1305 20400 1345
rect -900 1300 20400 1305
rect -900 1245 20400 1250
rect -900 1205 3705 1245
rect 3745 1205 4005 1245
rect 4045 1205 4305 1245
rect 4345 1205 4605 1245
rect 4645 1205 20400 1245
rect -900 1200 20400 1205
rect -900 1145 20400 1150
rect -900 1105 1305 1145
rect 1345 1105 1605 1145
rect 1645 1105 1905 1145
rect 1945 1105 2205 1145
rect 2245 1105 2355 1145
rect 2395 1105 2505 1145
rect 2545 1105 2805 1145
rect 2845 1105 3105 1145
rect 3145 1105 3405 1145
rect 3445 1105 4905 1145
rect 4945 1105 5205 1145
rect 5245 1105 5505 1145
rect 5545 1105 5805 1145
rect 5845 1105 5955 1145
rect 5995 1105 6105 1145
rect 6145 1105 6405 1145
rect 6445 1105 6705 1145
rect 6745 1105 7005 1145
rect 7045 1105 20400 1145
rect -900 1100 20400 1105
rect -900 1045 20400 1050
rect -900 1005 -345 1045
rect -305 1005 105 1045
rect 145 1005 405 1045
rect 445 1005 705 1045
rect 745 1005 1005 1045
rect 1045 1005 3855 1045
rect 3895 1005 4455 1045
rect 4495 1005 7305 1045
rect 7345 1005 7605 1045
rect 7645 1005 7905 1045
rect 7945 1005 8205 1045
rect 8245 1005 8505 1045
rect 8545 1005 8805 1045
rect 8845 1005 9105 1045
rect 9145 1005 9405 1045
rect 9445 1005 9705 1045
rect 9745 1005 10005 1045
rect 10045 1005 10305 1045
rect 10345 1005 10605 1045
rect 10645 1005 10905 1045
rect 10945 1005 11205 1045
rect 11245 1005 11505 1045
rect 11545 1005 11805 1045
rect 11845 1005 14505 1045
rect 14545 1005 14805 1045
rect 14845 1005 15105 1045
rect 15145 1005 15405 1045
rect 15445 1005 20400 1045
rect -900 1000 20400 1005
rect -900 900 20400 950
rect -500 845 -450 850
rect -500 805 -495 845
rect -455 805 -450 845
rect -500 800 -450 805
rect -350 845 -300 850
rect -350 805 -345 845
rect -305 805 -300 845
rect -350 800 -300 805
rect -200 845 -150 850
rect -200 805 -195 845
rect -155 805 -150 845
rect -200 800 -150 805
rect 100 845 150 850
rect 100 805 105 845
rect 145 805 150 845
rect 100 800 150 805
rect 400 845 450 850
rect 400 805 405 845
rect 445 805 450 845
rect 400 800 450 805
rect 700 845 750 850
rect 700 805 705 845
rect 745 805 750 845
rect 700 800 750 805
rect 1000 845 1050 850
rect 1000 805 1005 845
rect 1045 805 1050 845
rect 1000 800 1050 805
rect 1300 845 1350 850
rect 1300 805 1305 845
rect 1345 805 1350 845
rect 1300 800 1350 805
rect 1600 845 1650 850
rect 1600 805 1605 845
rect 1645 805 1650 845
rect 1600 800 1650 805
rect 1900 845 1950 850
rect 1900 805 1905 845
rect 1945 805 1950 845
rect 1900 800 1950 805
rect 2200 845 2250 850
rect 2200 805 2205 845
rect 2245 805 2250 845
rect 2200 800 2250 805
rect 2350 845 2400 850
rect 2350 805 2355 845
rect 2395 805 2400 845
rect 2350 800 2400 805
rect 2500 845 2550 850
rect 2500 805 2505 845
rect 2545 805 2550 845
rect 2500 800 2550 805
rect 2800 845 2850 850
rect 2800 805 2805 845
rect 2845 805 2850 845
rect 2800 800 2850 805
rect 3100 845 3150 850
rect 3100 805 3105 845
rect 3145 805 3150 845
rect 3100 800 3150 805
rect 3400 845 3450 850
rect 3400 805 3405 845
rect 3445 805 3450 845
rect 3400 800 3450 805
rect 3700 845 3750 850
rect 3700 805 3705 845
rect 3745 805 3750 845
rect 3700 800 3750 805
rect 3850 845 3900 850
rect 3850 805 3855 845
rect 3895 805 3900 845
rect 3850 800 3900 805
rect 4000 845 4050 850
rect 4000 805 4005 845
rect 4045 805 4050 845
rect 4000 800 4050 805
rect 4300 845 4350 850
rect 4300 805 4305 845
rect 4345 805 4350 845
rect 4300 800 4350 805
rect 4450 845 4500 850
rect 4450 805 4455 845
rect 4495 805 4500 845
rect 4450 800 4500 805
rect 4600 845 4650 850
rect 4600 805 4605 845
rect 4645 805 4650 845
rect 4600 800 4650 805
rect 4900 845 4950 850
rect 4900 805 4905 845
rect 4945 805 4950 845
rect 4900 800 4950 805
rect 5200 845 5250 850
rect 5200 805 5205 845
rect 5245 805 5250 845
rect 5200 800 5250 805
rect 5500 845 5550 850
rect 5500 805 5505 845
rect 5545 805 5550 845
rect 5500 800 5550 805
rect 5800 845 5850 850
rect 5800 805 5805 845
rect 5845 805 5850 845
rect 5800 800 5850 805
rect 5950 845 6000 850
rect 5950 805 5955 845
rect 5995 805 6000 845
rect 5950 800 6000 805
rect 6100 845 6150 850
rect 6100 805 6105 845
rect 6145 805 6150 845
rect 6100 800 6150 805
rect 6400 845 6450 850
rect 6400 805 6405 845
rect 6445 805 6450 845
rect 6400 800 6450 805
rect 6700 845 6750 850
rect 6700 805 6705 845
rect 6745 805 6750 845
rect 6700 800 6750 805
rect 7000 845 7050 850
rect 7000 805 7005 845
rect 7045 805 7050 845
rect 7000 800 7050 805
rect 7300 845 7350 850
rect 7300 805 7305 845
rect 7345 805 7350 845
rect 7300 800 7350 805
rect 7600 845 7650 850
rect 7600 805 7605 845
rect 7645 805 7650 845
rect 7600 800 7650 805
rect 7900 845 7950 850
rect 7900 805 7905 845
rect 7945 805 7950 845
rect 7900 800 7950 805
rect 8200 845 8250 850
rect 8200 805 8205 845
rect 8245 805 8250 845
rect 8200 800 8250 805
rect 8500 845 8550 850
rect 8500 805 8505 845
rect 8545 805 8550 845
rect 8500 800 8550 805
rect 8800 845 8850 850
rect 8800 805 8805 845
rect 8845 805 8850 845
rect 8800 800 8850 805
rect 9100 845 9150 850
rect 9100 805 9105 845
rect 9145 805 9150 845
rect 9100 800 9150 805
rect 9400 845 9450 850
rect 9400 805 9405 845
rect 9445 805 9450 845
rect 9400 800 9450 805
rect 9550 845 9600 850
rect 9550 805 9555 845
rect 9595 805 9600 845
rect 9550 800 9600 805
rect 9700 845 9750 850
rect 9700 805 9705 845
rect 9745 805 9750 845
rect 9700 800 9750 805
rect 10000 845 10050 850
rect 10000 805 10005 845
rect 10045 805 10050 845
rect 10000 800 10050 805
rect 10300 845 10350 850
rect 10300 805 10305 845
rect 10345 805 10350 845
rect 10300 800 10350 805
rect 10600 845 10650 850
rect 10600 805 10605 845
rect 10645 805 10650 845
rect 10600 800 10650 805
rect 10900 845 10950 850
rect 10900 805 10905 845
rect 10945 805 10950 845
rect 10900 800 10950 805
rect 11200 845 11250 850
rect 11200 805 11205 845
rect 11245 805 11250 845
rect 11200 800 11250 805
rect 11500 845 11550 850
rect 11500 805 11505 845
rect 11545 805 11550 845
rect 11500 800 11550 805
rect 11800 845 11850 850
rect 11800 805 11805 845
rect 11845 805 11850 845
rect 11800 800 11850 805
rect 12100 845 12150 850
rect 12100 805 12105 845
rect 12145 805 12150 845
rect 12100 800 12150 805
rect 12400 845 12450 850
rect 12400 805 12405 845
rect 12445 805 12450 845
rect 12400 800 12450 805
rect 12550 845 12600 850
rect 12550 805 12555 845
rect 12595 805 12600 845
rect 12550 800 12600 805
rect 12700 845 12750 850
rect 12700 805 12705 845
rect 12745 805 12750 845
rect 12700 800 12750 805
rect 13000 845 13050 850
rect 13000 805 13005 845
rect 13045 805 13050 845
rect 13000 800 13050 805
rect 13150 840 13200 850
rect 13150 810 13160 840
rect 13190 810 13200 840
rect 13150 800 13200 810
rect 13300 845 13350 850
rect 13300 805 13305 845
rect 13345 805 13350 845
rect 13300 800 13350 805
rect 13600 845 13650 850
rect 13600 805 13605 845
rect 13645 805 13650 845
rect 13600 800 13650 805
rect 13750 845 13800 850
rect 13750 805 13755 845
rect 13795 805 13800 845
rect 13750 800 13800 805
rect 13900 845 13950 850
rect 13900 805 13905 845
rect 13945 805 13950 845
rect 13900 800 13950 805
rect 14200 845 14250 850
rect 14200 805 14205 845
rect 14245 805 14250 845
rect 14200 800 14250 805
rect 14500 845 14550 850
rect 14500 805 14505 845
rect 14545 805 14550 845
rect 14500 800 14550 805
rect 14800 845 14850 850
rect 14800 805 14805 845
rect 14845 805 14850 845
rect 14800 800 14850 805
rect 15100 845 15150 850
rect 15100 805 15105 845
rect 15145 805 15150 845
rect 15100 800 15150 805
rect 15400 845 15450 850
rect 15400 805 15405 845
rect 15445 805 15450 845
rect 15400 800 15450 805
rect 15700 845 15750 850
rect 15700 805 15705 845
rect 15745 805 15750 845
rect 15700 800 15750 805
rect 16000 845 16050 850
rect 16000 805 16005 845
rect 16045 805 16050 845
rect 16000 800 16050 805
rect 16300 845 16350 850
rect 16300 805 16305 845
rect 16345 805 16350 845
rect 16300 800 16350 805
rect 16600 845 16650 850
rect 16600 805 16605 845
rect 16645 805 16650 845
rect 16600 800 16650 805
rect 16750 845 16800 850
rect 16750 805 16755 845
rect 16795 805 16800 845
rect 16750 800 16800 805
rect 16900 845 16950 850
rect 16900 805 16905 845
rect 16945 805 16950 845
rect 16900 800 16950 805
rect 17200 845 17250 850
rect 17200 805 17205 845
rect 17245 805 17250 845
rect 17200 800 17250 805
rect 17500 845 17550 850
rect 17500 805 17505 845
rect 17545 805 17550 845
rect 17500 800 17550 805
rect 17800 845 17850 850
rect 17800 805 17805 845
rect 17845 805 17850 845
rect 17800 800 17850 805
rect 18100 845 18150 850
rect 18100 805 18105 845
rect 18145 805 18150 845
rect 18100 800 18150 805
rect 18400 845 18450 850
rect 18400 805 18405 845
rect 18445 805 18450 845
rect 18400 800 18450 805
rect 18700 845 18750 850
rect 18700 805 18705 845
rect 18745 805 18750 845
rect 18700 800 18750 805
rect 19000 845 19050 850
rect 19000 805 19005 845
rect 19045 805 19050 845
rect 19000 800 19050 805
rect 19150 845 19200 850
rect 19150 805 19155 845
rect 19195 805 19200 845
rect 19150 800 19200 805
rect 19300 845 19350 850
rect 19300 805 19305 845
rect 19345 805 19350 845
rect 19300 800 19350 805
rect 19600 845 19650 850
rect 19600 805 19605 845
rect 19645 805 19650 845
rect 19600 800 19650 805
rect 19900 845 19950 850
rect 19900 805 19905 845
rect 19945 805 19950 845
rect 19900 800 19950 805
rect 20200 845 20250 850
rect 20200 805 20205 845
rect 20245 805 20250 845
rect 20200 800 20250 805
rect -900 700 20400 750
rect -900 645 20400 650
rect -900 605 15705 645
rect 15745 605 16005 645
rect 16045 605 16305 645
rect 16345 605 16605 645
rect 16645 605 16905 645
rect 16945 605 17205 645
rect 17245 605 17505 645
rect 17545 605 17805 645
rect 17845 605 20400 645
rect -900 600 20400 605
rect -900 500 20400 550
rect -900 445 20400 450
rect -900 405 18105 445
rect 18145 405 18405 445
rect 18445 405 18705 445
rect 18745 405 19005 445
rect 19045 405 19305 445
rect 19345 405 19605 445
rect 19645 405 19905 445
rect 19945 405 20205 445
rect 20245 405 20400 445
rect -900 400 20400 405
rect -900 300 20400 350
rect -900 200 20400 250
rect -900 100 20400 150
rect -900 40 20400 50
rect -900 10 -640 40
rect -610 10 -40 40
rect -10 10 8360 40
rect 8390 10 10760 40
rect 10790 10 15560 40
rect 15590 10 17960 40
rect 17990 10 20360 40
rect 20390 10 20400 40
rect -900 -10 20400 10
rect -900 -40 -640 -10
rect -610 -40 -40 -10
rect -10 -40 8360 -10
rect 8390 -40 10760 -10
rect 10790 -40 15560 -10
rect 15590 -40 17960 -10
rect 17990 -40 20360 -10
rect 20390 -40 20400 -10
rect -900 -60 20400 -40
rect -900 -90 -640 -60
rect -610 -90 -40 -60
rect -10 -90 8360 -60
rect 8390 -90 10760 -60
rect 10790 -90 15560 -60
rect 15590 -90 17960 -60
rect 17990 -90 20360 -60
rect 20390 -90 20400 -60
rect -900 -100 20400 -90
rect -900 -200 20400 -150
rect -900 -300 20400 -250
rect -900 -400 20400 -350
rect -900 -500 20400 -450
rect -900 -600 20400 -550
rect -900 -700 20400 -650
rect -900 -800 20400 -750
rect -500 -855 -450 -850
rect -500 -895 -495 -855
rect -455 -895 -450 -855
rect -500 -900 -450 -895
rect -350 -855 -300 -850
rect -350 -895 -345 -855
rect -305 -895 -300 -855
rect -350 -900 -300 -895
rect -200 -855 -150 -850
rect -200 -895 -195 -855
rect -155 -895 -150 -855
rect -200 -900 -150 -895
rect 100 -855 150 -850
rect 100 -895 105 -855
rect 145 -895 150 -855
rect 100 -900 150 -895
rect 400 -855 450 -850
rect 400 -895 405 -855
rect 445 -895 450 -855
rect 400 -900 450 -895
rect 700 -855 750 -850
rect 700 -895 705 -855
rect 745 -895 750 -855
rect 700 -900 750 -895
rect 1000 -855 1050 -850
rect 1000 -895 1005 -855
rect 1045 -895 1050 -855
rect 1000 -900 1050 -895
rect 1300 -855 1350 -850
rect 1300 -895 1305 -855
rect 1345 -895 1350 -855
rect 1300 -900 1350 -895
rect 1600 -855 1650 -850
rect 1600 -895 1605 -855
rect 1645 -895 1650 -855
rect 1600 -900 1650 -895
rect 1900 -855 1950 -850
rect 1900 -895 1905 -855
rect 1945 -895 1950 -855
rect 1900 -900 1950 -895
rect 2200 -855 2250 -850
rect 2200 -895 2205 -855
rect 2245 -895 2250 -855
rect 2200 -900 2250 -895
rect 2350 -855 2400 -850
rect 2350 -895 2355 -855
rect 2395 -895 2400 -855
rect 2350 -900 2400 -895
rect 2500 -855 2550 -850
rect 2500 -895 2505 -855
rect 2545 -895 2550 -855
rect 2500 -900 2550 -895
rect 2800 -855 2850 -850
rect 2800 -895 2805 -855
rect 2845 -895 2850 -855
rect 2800 -900 2850 -895
rect 3100 -855 3150 -850
rect 3100 -895 3105 -855
rect 3145 -895 3150 -855
rect 3100 -900 3150 -895
rect 3400 -855 3450 -850
rect 3400 -895 3405 -855
rect 3445 -895 3450 -855
rect 3400 -900 3450 -895
rect 3700 -855 3750 -850
rect 3700 -895 3705 -855
rect 3745 -895 3750 -855
rect 3700 -900 3750 -895
rect 3850 -855 3900 -850
rect 3850 -895 3855 -855
rect 3895 -895 3900 -855
rect 3850 -900 3900 -895
rect 4000 -855 4050 -850
rect 4000 -895 4005 -855
rect 4045 -895 4050 -855
rect 4000 -900 4050 -895
rect 4300 -855 4350 -850
rect 4300 -895 4305 -855
rect 4345 -895 4350 -855
rect 4300 -900 4350 -895
rect 4450 -855 4500 -850
rect 4450 -895 4455 -855
rect 4495 -895 4500 -855
rect 4450 -900 4500 -895
rect 4600 -855 4650 -850
rect 4600 -895 4605 -855
rect 4645 -895 4650 -855
rect 4600 -900 4650 -895
rect 4900 -855 4950 -850
rect 4900 -895 4905 -855
rect 4945 -895 4950 -855
rect 4900 -900 4950 -895
rect 5200 -855 5250 -850
rect 5200 -895 5205 -855
rect 5245 -895 5250 -855
rect 5200 -900 5250 -895
rect 5500 -855 5550 -850
rect 5500 -895 5505 -855
rect 5545 -895 5550 -855
rect 5500 -900 5550 -895
rect 5800 -855 5850 -850
rect 5800 -895 5805 -855
rect 5845 -895 5850 -855
rect 5800 -900 5850 -895
rect 5950 -855 6000 -850
rect 5950 -895 5955 -855
rect 5995 -895 6000 -855
rect 5950 -900 6000 -895
rect 6100 -855 6150 -850
rect 6100 -895 6105 -855
rect 6145 -895 6150 -855
rect 6100 -900 6150 -895
rect 6400 -855 6450 -850
rect 6400 -895 6405 -855
rect 6445 -895 6450 -855
rect 6400 -900 6450 -895
rect 6700 -855 6750 -850
rect 6700 -895 6705 -855
rect 6745 -895 6750 -855
rect 6700 -900 6750 -895
rect 7000 -855 7050 -850
rect 7000 -895 7005 -855
rect 7045 -895 7050 -855
rect 7000 -900 7050 -895
rect 7300 -855 7350 -850
rect 7300 -895 7305 -855
rect 7345 -895 7350 -855
rect 7300 -900 7350 -895
rect 7600 -855 7650 -850
rect 7600 -895 7605 -855
rect 7645 -895 7650 -855
rect 7600 -900 7650 -895
rect 7900 -855 7950 -850
rect 7900 -895 7905 -855
rect 7945 -895 7950 -855
rect 7900 -900 7950 -895
rect 8200 -855 8250 -850
rect 8200 -895 8205 -855
rect 8245 -895 8250 -855
rect 8200 -900 8250 -895
rect 8500 -855 8550 -850
rect 8500 -895 8505 -855
rect 8545 -895 8550 -855
rect 8500 -900 8550 -895
rect 8800 -855 8850 -850
rect 8800 -895 8805 -855
rect 8845 -895 8850 -855
rect 8800 -900 8850 -895
rect 9100 -855 9150 -850
rect 9100 -895 9105 -855
rect 9145 -895 9150 -855
rect 9100 -900 9150 -895
rect 9400 -855 9450 -850
rect 9400 -895 9405 -855
rect 9445 -895 9450 -855
rect 9400 -900 9450 -895
rect 9550 -855 9600 -850
rect 9550 -895 9555 -855
rect 9595 -895 9600 -855
rect 9550 -900 9600 -895
rect 9700 -855 9750 -850
rect 9700 -895 9705 -855
rect 9745 -895 9750 -855
rect 9700 -900 9750 -895
rect 10000 -855 10050 -850
rect 10000 -895 10005 -855
rect 10045 -895 10050 -855
rect 10000 -900 10050 -895
rect 10300 -855 10350 -850
rect 10300 -895 10305 -855
rect 10345 -895 10350 -855
rect 10300 -900 10350 -895
rect 10600 -855 10650 -850
rect 10600 -895 10605 -855
rect 10645 -895 10650 -855
rect 10600 -900 10650 -895
rect 10900 -855 10950 -850
rect 10900 -895 10905 -855
rect 10945 -895 10950 -855
rect 10900 -900 10950 -895
rect 11200 -855 11250 -850
rect 11200 -895 11205 -855
rect 11245 -895 11250 -855
rect 11200 -900 11250 -895
rect 11500 -855 11550 -850
rect 11500 -895 11505 -855
rect 11545 -895 11550 -855
rect 11500 -900 11550 -895
rect 11800 -855 11850 -850
rect 11800 -895 11805 -855
rect 11845 -895 11850 -855
rect 11800 -900 11850 -895
rect 12100 -855 12150 -850
rect 12100 -895 12105 -855
rect 12145 -895 12150 -855
rect 12100 -900 12150 -895
rect 12400 -855 12450 -850
rect 12400 -895 12405 -855
rect 12445 -895 12450 -855
rect 12400 -900 12450 -895
rect 12550 -855 12600 -850
rect 12550 -895 12555 -855
rect 12595 -895 12600 -855
rect 12550 -900 12600 -895
rect 12700 -855 12750 -850
rect 12700 -895 12705 -855
rect 12745 -895 12750 -855
rect 12700 -900 12750 -895
rect 13000 -855 13050 -850
rect 13000 -895 13005 -855
rect 13045 -895 13050 -855
rect 13000 -900 13050 -895
rect 13150 -860 13200 -850
rect 13150 -890 13160 -860
rect 13190 -890 13200 -860
rect 13150 -900 13200 -890
rect 13300 -855 13350 -850
rect 13300 -895 13305 -855
rect 13345 -895 13350 -855
rect 13300 -900 13350 -895
rect 13600 -855 13650 -850
rect 13600 -895 13605 -855
rect 13645 -895 13650 -855
rect 13600 -900 13650 -895
rect 13750 -855 13800 -850
rect 13750 -895 13755 -855
rect 13795 -895 13800 -855
rect 13750 -900 13800 -895
rect 13900 -855 13950 -850
rect 13900 -895 13905 -855
rect 13945 -895 13950 -855
rect 13900 -900 13950 -895
rect 14200 -855 14250 -850
rect 14200 -895 14205 -855
rect 14245 -895 14250 -855
rect 14200 -900 14250 -895
rect 14500 -855 14550 -850
rect 14500 -895 14505 -855
rect 14545 -895 14550 -855
rect 14500 -900 14550 -895
rect 14800 -855 14850 -850
rect 14800 -895 14805 -855
rect 14845 -895 14850 -855
rect 14800 -900 14850 -895
rect 15100 -855 15150 -850
rect 15100 -895 15105 -855
rect 15145 -895 15150 -855
rect 15100 -900 15150 -895
rect 15400 -855 15450 -850
rect 15400 -895 15405 -855
rect 15445 -895 15450 -855
rect 15400 -900 15450 -895
rect 15700 -855 15750 -850
rect 15700 -895 15705 -855
rect 15745 -895 15750 -855
rect 15700 -900 15750 -895
rect 16000 -855 16050 -850
rect 16000 -895 16005 -855
rect 16045 -895 16050 -855
rect 16000 -900 16050 -895
rect 16300 -855 16350 -850
rect 16300 -895 16305 -855
rect 16345 -895 16350 -855
rect 16300 -900 16350 -895
rect 16600 -855 16650 -850
rect 16600 -895 16605 -855
rect 16645 -895 16650 -855
rect 16600 -900 16650 -895
rect 16750 -855 16800 -850
rect 16750 -895 16755 -855
rect 16795 -895 16800 -855
rect 16750 -900 16800 -895
rect 16900 -855 16950 -850
rect 16900 -895 16905 -855
rect 16945 -895 16950 -855
rect 16900 -900 16950 -895
rect 17200 -855 17250 -850
rect 17200 -895 17205 -855
rect 17245 -895 17250 -855
rect 17200 -900 17250 -895
rect 17500 -855 17550 -850
rect 17500 -895 17505 -855
rect 17545 -895 17550 -855
rect 17500 -900 17550 -895
rect 17800 -855 17850 -850
rect 17800 -895 17805 -855
rect 17845 -895 17850 -855
rect 17800 -900 17850 -895
rect 18100 -855 18150 -850
rect 18100 -895 18105 -855
rect 18145 -895 18150 -855
rect 18100 -900 18150 -895
rect 18400 -855 18450 -850
rect 18400 -895 18405 -855
rect 18445 -895 18450 -855
rect 18400 -900 18450 -895
rect 18700 -855 18750 -850
rect 18700 -895 18705 -855
rect 18745 -895 18750 -855
rect 18700 -900 18750 -895
rect 19000 -855 19050 -850
rect 19000 -895 19005 -855
rect 19045 -895 19050 -855
rect 19000 -900 19050 -895
rect 19150 -855 19200 -850
rect 19150 -895 19155 -855
rect 19195 -895 19200 -855
rect 19150 -900 19200 -895
rect 19300 -855 19350 -850
rect 19300 -895 19305 -855
rect 19345 -895 19350 -855
rect 19300 -900 19350 -895
rect 19600 -855 19650 -850
rect 19600 -895 19605 -855
rect 19645 -895 19650 -855
rect 19600 -900 19650 -895
rect 19900 -855 19950 -850
rect 19900 -895 19905 -855
rect 19945 -895 19950 -855
rect 19900 -900 19950 -895
rect 20200 -855 20250 -850
rect 20200 -895 20205 -855
rect 20245 -895 20250 -855
rect 20200 -900 20250 -895
rect -900 -1000 20400 -950
rect -900 -1100 20400 -1050
rect -900 -1200 20400 -1150
rect -900 -1300 20400 -1250
rect -900 -1400 20400 -1350
rect -900 -1500 20400 -1450
rect -900 -1600 20400 -1550
rect -900 -1660 20400 -1650
rect -900 -1690 -640 -1660
rect -610 -1690 -40 -1660
rect -10 -1690 8360 -1660
rect 8390 -1690 10760 -1660
rect 10790 -1690 15560 -1660
rect 15590 -1690 17960 -1660
rect 17990 -1690 20360 -1660
rect 20390 -1690 20400 -1660
rect -900 -1710 20400 -1690
rect -900 -1740 -640 -1710
rect -610 -1740 -40 -1710
rect -10 -1740 8360 -1710
rect 8390 -1740 10760 -1710
rect 10790 -1740 15560 -1710
rect 15590 -1740 17960 -1710
rect 17990 -1740 20360 -1710
rect 20390 -1740 20400 -1710
rect -900 -1750 20400 -1740
<< via3 >>
rect -495 4540 -455 4545
rect -495 4510 -490 4540
rect -490 4510 -460 4540
rect -460 4510 -455 4540
rect -495 4505 -455 4510
rect -345 4540 -305 4545
rect -345 4510 -340 4540
rect -340 4510 -310 4540
rect -310 4510 -305 4540
rect -345 4505 -305 4510
rect -195 4540 -155 4545
rect -195 4510 -190 4540
rect -190 4510 -160 4540
rect -160 4510 -155 4540
rect -195 4505 -155 4510
rect 105 4540 145 4545
rect 105 4510 110 4540
rect 110 4510 140 4540
rect 140 4510 145 4540
rect 105 4505 145 4510
rect 405 4540 445 4545
rect 405 4510 410 4540
rect 410 4510 440 4540
rect 440 4510 445 4540
rect 405 4505 445 4510
rect 705 4540 745 4545
rect 705 4510 710 4540
rect 710 4510 740 4540
rect 740 4510 745 4540
rect 705 4505 745 4510
rect 1005 4540 1045 4545
rect 1005 4510 1010 4540
rect 1010 4510 1040 4540
rect 1040 4510 1045 4540
rect 1005 4505 1045 4510
rect 1155 4540 1195 4545
rect 1155 4510 1160 4540
rect 1160 4510 1190 4540
rect 1190 4510 1195 4540
rect 1155 4505 1195 4510
rect 1305 4540 1345 4545
rect 1305 4510 1310 4540
rect 1310 4510 1340 4540
rect 1340 4510 1345 4540
rect 1305 4505 1345 4510
rect 1605 4540 1645 4545
rect 1605 4510 1610 4540
rect 1610 4510 1640 4540
rect 1640 4510 1645 4540
rect 1605 4505 1645 4510
rect 1905 4540 1945 4545
rect 1905 4510 1910 4540
rect 1910 4510 1940 4540
rect 1940 4510 1945 4540
rect 1905 4505 1945 4510
rect 2055 4540 2095 4545
rect 2055 4510 2060 4540
rect 2060 4510 2090 4540
rect 2090 4510 2095 4540
rect 2055 4505 2095 4510
rect 2205 4540 2245 4545
rect 2205 4510 2210 4540
rect 2210 4510 2240 4540
rect 2240 4510 2245 4540
rect 2205 4505 2245 4510
rect 2505 4540 2545 4545
rect 2505 4510 2510 4540
rect 2510 4510 2540 4540
rect 2540 4510 2545 4540
rect 2505 4505 2545 4510
rect 2805 4540 2845 4545
rect 2805 4510 2810 4540
rect 2810 4510 2840 4540
rect 2840 4510 2845 4540
rect 2805 4505 2845 4510
rect 2955 4540 2995 4545
rect 2955 4510 2960 4540
rect 2960 4510 2990 4540
rect 2990 4510 2995 4540
rect 2955 4505 2995 4510
rect 3105 4540 3145 4545
rect 3105 4510 3110 4540
rect 3110 4510 3140 4540
rect 3140 4510 3145 4540
rect 3105 4505 3145 4510
rect 3405 4540 3445 4545
rect 3405 4510 3410 4540
rect 3410 4510 3440 4540
rect 3440 4510 3445 4540
rect 3405 4505 3445 4510
rect 3705 4540 3745 4545
rect 3705 4510 3710 4540
rect 3710 4510 3740 4540
rect 3740 4510 3745 4540
rect 3705 4505 3745 4510
rect 4005 4540 4045 4545
rect 4005 4510 4010 4540
rect 4010 4510 4040 4540
rect 4040 4510 4045 4540
rect 4005 4505 4045 4510
rect 4305 4540 4345 4545
rect 4305 4510 4310 4540
rect 4310 4510 4340 4540
rect 4340 4510 4345 4540
rect 4305 4505 4345 4510
rect 4605 4540 4645 4545
rect 4605 4510 4610 4540
rect 4610 4510 4640 4540
rect 4640 4510 4645 4540
rect 4605 4505 4645 4510
rect 4905 4540 4945 4545
rect 4905 4510 4910 4540
rect 4910 4510 4940 4540
rect 4940 4510 4945 4540
rect 4905 4505 4945 4510
rect 5205 4540 5245 4545
rect 5205 4510 5210 4540
rect 5210 4510 5240 4540
rect 5240 4510 5245 4540
rect 5205 4505 5245 4510
rect 5355 4540 5395 4545
rect 5355 4510 5360 4540
rect 5360 4510 5390 4540
rect 5390 4510 5395 4540
rect 5355 4505 5395 4510
rect 5505 4540 5545 4545
rect 5505 4510 5510 4540
rect 5510 4510 5540 4540
rect 5540 4510 5545 4540
rect 5505 4505 5545 4510
rect 5805 4540 5845 4545
rect 5805 4510 5810 4540
rect 5810 4510 5840 4540
rect 5840 4510 5845 4540
rect 5805 4505 5845 4510
rect 6105 4540 6145 4545
rect 6105 4510 6110 4540
rect 6110 4510 6140 4540
rect 6140 4510 6145 4540
rect 6105 4505 6145 4510
rect 6255 4540 6295 4545
rect 6255 4510 6260 4540
rect 6260 4510 6290 4540
rect 6290 4510 6295 4540
rect 6255 4505 6295 4510
rect 6405 4540 6445 4545
rect 6405 4510 6410 4540
rect 6410 4510 6440 4540
rect 6440 4510 6445 4540
rect 6405 4505 6445 4510
rect 6705 4540 6745 4545
rect 6705 4510 6710 4540
rect 6710 4510 6740 4540
rect 6740 4510 6745 4540
rect 6705 4505 6745 4510
rect 7005 4540 7045 4545
rect 7005 4510 7010 4540
rect 7010 4510 7040 4540
rect 7040 4510 7045 4540
rect 7005 4505 7045 4510
rect 7155 4540 7195 4545
rect 7155 4510 7160 4540
rect 7160 4510 7190 4540
rect 7190 4510 7195 4540
rect 7155 4505 7195 4510
rect 7305 4540 7345 4545
rect 7305 4510 7310 4540
rect 7310 4510 7340 4540
rect 7340 4510 7345 4540
rect 7305 4505 7345 4510
rect 7605 4540 7645 4545
rect 7605 4510 7610 4540
rect 7610 4510 7640 4540
rect 7640 4510 7645 4540
rect 7605 4505 7645 4510
rect 7905 4540 7945 4545
rect 7905 4510 7910 4540
rect 7910 4510 7940 4540
rect 7940 4510 7945 4540
rect 7905 4505 7945 4510
rect 8205 4540 8245 4545
rect 8205 4510 8210 4540
rect 8210 4510 8240 4540
rect 8240 4510 8245 4540
rect 8205 4505 8245 4510
rect 8505 4540 8545 4545
rect 8505 4510 8510 4540
rect 8510 4510 8540 4540
rect 8540 4510 8545 4540
rect 8505 4505 8545 4510
rect 8805 4540 8845 4545
rect 8805 4510 8810 4540
rect 8810 4510 8840 4540
rect 8840 4510 8845 4540
rect 8805 4505 8845 4510
rect 9105 4540 9145 4545
rect 9105 4510 9110 4540
rect 9110 4510 9140 4540
rect 9140 4510 9145 4540
rect 9105 4505 9145 4510
rect 9405 4540 9445 4545
rect 9405 4510 9410 4540
rect 9410 4510 9440 4540
rect 9440 4510 9445 4540
rect 9405 4505 9445 4510
rect 9705 4540 9745 4545
rect 9705 4510 9710 4540
rect 9710 4510 9740 4540
rect 9740 4510 9745 4540
rect 9705 4505 9745 4510
rect 10005 4540 10045 4545
rect 10005 4510 10010 4540
rect 10010 4510 10040 4540
rect 10040 4510 10045 4540
rect 10005 4505 10045 4510
rect 10305 4540 10345 4545
rect 10305 4510 10310 4540
rect 10310 4510 10340 4540
rect 10340 4510 10345 4540
rect 10305 4505 10345 4510
rect 10605 4540 10645 4545
rect 10605 4510 10610 4540
rect 10610 4510 10640 4540
rect 10640 4510 10645 4540
rect 10605 4505 10645 4510
rect 10905 4540 10945 4545
rect 10905 4510 10910 4540
rect 10910 4510 10940 4540
rect 10940 4510 10945 4540
rect 10905 4505 10945 4510
rect 11205 4540 11245 4545
rect 11205 4510 11210 4540
rect 11210 4510 11240 4540
rect 11240 4510 11245 4540
rect 11205 4505 11245 4510
rect 11355 4540 11395 4545
rect 11355 4510 11360 4540
rect 11360 4510 11390 4540
rect 11390 4510 11395 4540
rect 11355 4505 11395 4510
rect 11505 4540 11545 4545
rect 11505 4510 11510 4540
rect 11510 4510 11540 4540
rect 11540 4510 11545 4540
rect 11505 4505 11545 4510
rect 11805 4540 11845 4545
rect 11805 4510 11810 4540
rect 11810 4510 11840 4540
rect 11840 4510 11845 4540
rect 11805 4505 11845 4510
rect 12105 4540 12145 4545
rect 12105 4510 12110 4540
rect 12110 4510 12140 4540
rect 12140 4510 12145 4540
rect 12105 4505 12145 4510
rect 12405 4540 12445 4545
rect 12405 4510 12410 4540
rect 12410 4510 12440 4540
rect 12440 4510 12445 4540
rect 12405 4505 12445 4510
rect 12555 4540 12595 4545
rect 12555 4510 12560 4540
rect 12560 4510 12590 4540
rect 12590 4510 12595 4540
rect 12555 4505 12595 4510
rect 12705 4540 12745 4545
rect 12705 4510 12710 4540
rect 12710 4510 12740 4540
rect 12740 4510 12745 4540
rect 12705 4505 12745 4510
rect 13005 4540 13045 4545
rect 13005 4510 13010 4540
rect 13010 4510 13040 4540
rect 13040 4510 13045 4540
rect 13005 4505 13045 4510
rect 13305 4540 13345 4545
rect 13305 4510 13310 4540
rect 13310 4510 13340 4540
rect 13340 4510 13345 4540
rect 13305 4505 13345 4510
rect 13605 4540 13645 4545
rect 13605 4510 13610 4540
rect 13610 4510 13640 4540
rect 13640 4510 13645 4540
rect 13605 4505 13645 4510
rect 13755 4540 13795 4545
rect 13755 4510 13760 4540
rect 13760 4510 13790 4540
rect 13790 4510 13795 4540
rect 13755 4505 13795 4510
rect 13905 4540 13945 4545
rect 13905 4510 13910 4540
rect 13910 4510 13940 4540
rect 13940 4510 13945 4540
rect 13905 4505 13945 4510
rect 14205 4540 14245 4545
rect 14205 4510 14210 4540
rect 14210 4510 14240 4540
rect 14240 4510 14245 4540
rect 14205 4505 14245 4510
rect 14505 4540 14545 4545
rect 14505 4510 14510 4540
rect 14510 4510 14540 4540
rect 14540 4510 14545 4540
rect 14505 4505 14545 4510
rect 14805 4540 14845 4545
rect 14805 4510 14810 4540
rect 14810 4510 14840 4540
rect 14840 4510 14845 4540
rect 14805 4505 14845 4510
rect 14955 4540 14995 4545
rect 14955 4510 14960 4540
rect 14960 4510 14990 4540
rect 14990 4510 14995 4540
rect 14955 4505 14995 4510
rect 15105 4540 15145 4545
rect 15105 4510 15110 4540
rect 15110 4510 15140 4540
rect 15140 4510 15145 4540
rect 15105 4505 15145 4510
rect 15405 4540 15445 4545
rect 15405 4510 15410 4540
rect 15410 4510 15440 4540
rect 15440 4510 15445 4540
rect 15405 4505 15445 4510
rect 15705 4540 15745 4545
rect 15705 4510 15710 4540
rect 15710 4510 15740 4540
rect 15740 4510 15745 4540
rect 15705 4505 15745 4510
rect 16005 4540 16045 4545
rect 16005 4510 16010 4540
rect 16010 4510 16040 4540
rect 16040 4510 16045 4540
rect 16005 4505 16045 4510
rect 16305 4540 16345 4545
rect 16305 4510 16310 4540
rect 16310 4510 16340 4540
rect 16340 4510 16345 4540
rect 16305 4505 16345 4510
rect 16605 4540 16645 4545
rect 16605 4510 16610 4540
rect 16610 4510 16640 4540
rect 16640 4510 16645 4540
rect 16605 4505 16645 4510
rect 16755 4540 16795 4545
rect 16755 4510 16760 4540
rect 16760 4510 16790 4540
rect 16790 4510 16795 4540
rect 16755 4505 16795 4510
rect 16905 4540 16945 4545
rect 16905 4510 16910 4540
rect 16910 4510 16940 4540
rect 16940 4510 16945 4540
rect 16905 4505 16945 4510
rect 17205 4540 17245 4545
rect 17205 4510 17210 4540
rect 17210 4510 17240 4540
rect 17240 4510 17245 4540
rect 17205 4505 17245 4510
rect 17505 4540 17545 4545
rect 17505 4510 17510 4540
rect 17510 4510 17540 4540
rect 17540 4510 17545 4540
rect 17505 4505 17545 4510
rect 17805 4540 17845 4545
rect 17805 4510 17810 4540
rect 17810 4510 17840 4540
rect 17840 4510 17845 4540
rect 17805 4505 17845 4510
rect 18105 4540 18145 4545
rect 18105 4510 18110 4540
rect 18110 4510 18140 4540
rect 18140 4510 18145 4540
rect 18105 4505 18145 4510
rect 18405 4540 18445 4545
rect 18405 4510 18410 4540
rect 18410 4510 18440 4540
rect 18440 4510 18445 4540
rect 18405 4505 18445 4510
rect 18705 4540 18745 4545
rect 18705 4510 18710 4540
rect 18710 4510 18740 4540
rect 18740 4510 18745 4540
rect 18705 4505 18745 4510
rect 19005 4540 19045 4545
rect 19005 4510 19010 4540
rect 19010 4510 19040 4540
rect 19040 4510 19045 4540
rect 19005 4505 19045 4510
rect 19155 4540 19195 4545
rect 19155 4510 19160 4540
rect 19160 4510 19190 4540
rect 19190 4510 19195 4540
rect 19155 4505 19195 4510
rect 19305 4540 19345 4545
rect 19305 4510 19310 4540
rect 19310 4510 19340 4540
rect 19340 4510 19345 4540
rect 19305 4505 19345 4510
rect 19605 4540 19645 4545
rect 19605 4510 19610 4540
rect 19610 4510 19640 4540
rect 19640 4510 19645 4540
rect 19605 4505 19645 4510
rect 19905 4540 19945 4545
rect 19905 4510 19910 4540
rect 19910 4510 19940 4540
rect 19940 4510 19945 4540
rect 19905 4505 19945 4510
rect 20205 4540 20245 4545
rect 20205 4510 20210 4540
rect 20210 4510 20240 4540
rect 20240 4510 20245 4540
rect 20205 4505 20245 4510
rect 13755 4305 13795 4345
rect 14955 4305 14995 4345
rect 11355 4105 11395 4145
rect 12555 4105 12595 4145
rect 13305 3605 13345 3645
rect 13605 3605 13645 3645
rect 13905 3605 13945 3645
rect 14205 3605 14245 3645
rect 14505 3605 14545 3645
rect 14805 3605 14845 3645
rect 15105 3605 15145 3645
rect 15405 3605 15445 3645
rect 10905 3405 10945 3445
rect 11205 3405 11245 3445
rect 11505 3405 11545 3445
rect 11805 3405 11845 3445
rect 12105 3405 12145 3445
rect 12405 3405 12445 3445
rect 12705 3405 12745 3445
rect 13005 3405 13045 3445
rect -495 3240 -455 3245
rect -495 3210 -490 3240
rect -490 3210 -460 3240
rect -460 3210 -455 3240
rect -495 3205 -455 3210
rect -345 3240 -305 3245
rect -345 3210 -340 3240
rect -340 3210 -310 3240
rect -310 3210 -305 3240
rect -345 3205 -305 3210
rect -195 3240 -155 3245
rect -195 3210 -190 3240
rect -190 3210 -160 3240
rect -160 3210 -155 3240
rect -195 3205 -155 3210
rect 105 3240 145 3245
rect 105 3210 110 3240
rect 110 3210 140 3240
rect 140 3210 145 3240
rect 105 3205 145 3210
rect 405 3240 445 3245
rect 405 3210 410 3240
rect 410 3210 440 3240
rect 440 3210 445 3240
rect 405 3205 445 3210
rect 705 3240 745 3245
rect 705 3210 710 3240
rect 710 3210 740 3240
rect 740 3210 745 3240
rect 705 3205 745 3210
rect 1005 3240 1045 3245
rect 1005 3210 1010 3240
rect 1010 3210 1040 3240
rect 1040 3210 1045 3240
rect 1005 3205 1045 3210
rect 1155 3240 1195 3245
rect 1155 3210 1160 3240
rect 1160 3210 1190 3240
rect 1190 3210 1195 3240
rect 1155 3205 1195 3210
rect 1305 3240 1345 3245
rect 1305 3210 1310 3240
rect 1310 3210 1340 3240
rect 1340 3210 1345 3240
rect 1305 3205 1345 3210
rect 1605 3240 1645 3245
rect 1605 3210 1610 3240
rect 1610 3210 1640 3240
rect 1640 3210 1645 3240
rect 1605 3205 1645 3210
rect 1905 3240 1945 3245
rect 1905 3210 1910 3240
rect 1910 3210 1940 3240
rect 1940 3210 1945 3240
rect 1905 3205 1945 3210
rect 2055 3240 2095 3245
rect 2055 3210 2060 3240
rect 2060 3210 2090 3240
rect 2090 3210 2095 3240
rect 2055 3205 2095 3210
rect 2205 3240 2245 3245
rect 2205 3210 2210 3240
rect 2210 3210 2240 3240
rect 2240 3210 2245 3240
rect 2205 3205 2245 3210
rect 2505 3240 2545 3245
rect 2505 3210 2510 3240
rect 2510 3210 2540 3240
rect 2540 3210 2545 3240
rect 2505 3205 2545 3210
rect 2805 3240 2845 3245
rect 2805 3210 2810 3240
rect 2810 3210 2840 3240
rect 2840 3210 2845 3240
rect 2805 3205 2845 3210
rect 2955 3240 2995 3245
rect 2955 3210 2960 3240
rect 2960 3210 2990 3240
rect 2990 3210 2995 3240
rect 2955 3205 2995 3210
rect 3105 3240 3145 3245
rect 3105 3210 3110 3240
rect 3110 3210 3140 3240
rect 3140 3210 3145 3240
rect 3105 3205 3145 3210
rect 3405 3240 3445 3245
rect 3405 3210 3410 3240
rect 3410 3210 3440 3240
rect 3440 3210 3445 3240
rect 3405 3205 3445 3210
rect 3705 3240 3745 3245
rect 3705 3210 3710 3240
rect 3710 3210 3740 3240
rect 3740 3210 3745 3240
rect 3705 3205 3745 3210
rect 4005 3240 4045 3245
rect 4005 3210 4010 3240
rect 4010 3210 4040 3240
rect 4040 3210 4045 3240
rect 4005 3205 4045 3210
rect 4305 3240 4345 3245
rect 4305 3210 4310 3240
rect 4310 3210 4340 3240
rect 4340 3210 4345 3240
rect 4305 3205 4345 3210
rect 4605 3240 4645 3245
rect 4605 3210 4610 3240
rect 4610 3210 4640 3240
rect 4640 3210 4645 3240
rect 4605 3205 4645 3210
rect 4905 3240 4945 3245
rect 4905 3210 4910 3240
rect 4910 3210 4940 3240
rect 4940 3210 4945 3240
rect 4905 3205 4945 3210
rect 5205 3240 5245 3245
rect 5205 3210 5210 3240
rect 5210 3210 5240 3240
rect 5240 3210 5245 3240
rect 5205 3205 5245 3210
rect 5355 3240 5395 3245
rect 5355 3210 5360 3240
rect 5360 3210 5390 3240
rect 5390 3210 5395 3240
rect 5355 3205 5395 3210
rect 5505 3240 5545 3245
rect 5505 3210 5510 3240
rect 5510 3210 5540 3240
rect 5540 3210 5545 3240
rect 5505 3205 5545 3210
rect 5805 3240 5845 3245
rect 5805 3210 5810 3240
rect 5810 3210 5840 3240
rect 5840 3210 5845 3240
rect 5805 3205 5845 3210
rect 6105 3240 6145 3245
rect 6105 3210 6110 3240
rect 6110 3210 6140 3240
rect 6140 3210 6145 3240
rect 6105 3205 6145 3210
rect 6255 3240 6295 3245
rect 6255 3210 6260 3240
rect 6260 3210 6290 3240
rect 6290 3210 6295 3240
rect 6255 3205 6295 3210
rect 6405 3240 6445 3245
rect 6405 3210 6410 3240
rect 6410 3210 6440 3240
rect 6440 3210 6445 3240
rect 6405 3205 6445 3210
rect 6705 3240 6745 3245
rect 6705 3210 6710 3240
rect 6710 3210 6740 3240
rect 6740 3210 6745 3240
rect 6705 3205 6745 3210
rect 7005 3240 7045 3245
rect 7005 3210 7010 3240
rect 7010 3210 7040 3240
rect 7040 3210 7045 3240
rect 7005 3205 7045 3210
rect 7155 3240 7195 3245
rect 7155 3210 7160 3240
rect 7160 3210 7190 3240
rect 7190 3210 7195 3240
rect 7155 3205 7195 3210
rect 7305 3240 7345 3245
rect 7305 3210 7310 3240
rect 7310 3210 7340 3240
rect 7340 3210 7345 3240
rect 7305 3205 7345 3210
rect 7605 3240 7645 3245
rect 7605 3210 7610 3240
rect 7610 3210 7640 3240
rect 7640 3210 7645 3240
rect 7605 3205 7645 3210
rect 7905 3240 7945 3245
rect 7905 3210 7910 3240
rect 7910 3210 7940 3240
rect 7940 3210 7945 3240
rect 7905 3205 7945 3210
rect 8205 3240 8245 3245
rect 8205 3210 8210 3240
rect 8210 3210 8240 3240
rect 8240 3210 8245 3240
rect 8205 3205 8245 3210
rect 8505 3240 8545 3245
rect 8505 3210 8510 3240
rect 8510 3210 8540 3240
rect 8540 3210 8545 3240
rect 8505 3205 8545 3210
rect 8805 3240 8845 3245
rect 8805 3210 8810 3240
rect 8810 3210 8840 3240
rect 8840 3210 8845 3240
rect 8805 3205 8845 3210
rect 9105 3240 9145 3245
rect 9105 3210 9110 3240
rect 9110 3210 9140 3240
rect 9140 3210 9145 3240
rect 9105 3205 9145 3210
rect 9405 3240 9445 3245
rect 9405 3210 9410 3240
rect 9410 3210 9440 3240
rect 9440 3210 9445 3240
rect 9405 3205 9445 3210
rect 9705 3240 9745 3245
rect 9705 3210 9710 3240
rect 9710 3210 9740 3240
rect 9740 3210 9745 3240
rect 9705 3205 9745 3210
rect 10005 3240 10045 3245
rect 10005 3210 10010 3240
rect 10010 3210 10040 3240
rect 10040 3210 10045 3240
rect 10005 3205 10045 3210
rect 10305 3240 10345 3245
rect 10305 3210 10310 3240
rect 10310 3210 10340 3240
rect 10340 3210 10345 3240
rect 10305 3205 10345 3210
rect 10605 3240 10645 3245
rect 10605 3210 10610 3240
rect 10610 3210 10640 3240
rect 10640 3210 10645 3240
rect 10605 3205 10645 3210
rect 10905 3240 10945 3245
rect 10905 3210 10910 3240
rect 10910 3210 10940 3240
rect 10940 3210 10945 3240
rect 10905 3205 10945 3210
rect 11205 3240 11245 3245
rect 11205 3210 11210 3240
rect 11210 3210 11240 3240
rect 11240 3210 11245 3240
rect 11205 3205 11245 3210
rect 11355 3240 11395 3245
rect 11355 3210 11360 3240
rect 11360 3210 11390 3240
rect 11390 3210 11395 3240
rect 11355 3205 11395 3210
rect 11505 3240 11545 3245
rect 11505 3210 11510 3240
rect 11510 3210 11540 3240
rect 11540 3210 11545 3240
rect 11505 3205 11545 3210
rect 11805 3240 11845 3245
rect 11805 3210 11810 3240
rect 11810 3210 11840 3240
rect 11840 3210 11845 3240
rect 11805 3205 11845 3210
rect 12105 3240 12145 3245
rect 12105 3210 12110 3240
rect 12110 3210 12140 3240
rect 12140 3210 12145 3240
rect 12105 3205 12145 3210
rect 12405 3240 12445 3245
rect 12405 3210 12410 3240
rect 12410 3210 12440 3240
rect 12440 3210 12445 3240
rect 12405 3205 12445 3210
rect 12555 3240 12595 3245
rect 12555 3210 12560 3240
rect 12560 3210 12590 3240
rect 12590 3210 12595 3240
rect 12555 3205 12595 3210
rect 12705 3240 12745 3245
rect 12705 3210 12710 3240
rect 12710 3210 12740 3240
rect 12740 3210 12745 3240
rect 12705 3205 12745 3210
rect 13005 3240 13045 3245
rect 13005 3210 13010 3240
rect 13010 3210 13040 3240
rect 13040 3210 13045 3240
rect 13005 3205 13045 3210
rect 13305 3240 13345 3245
rect 13305 3210 13310 3240
rect 13310 3210 13340 3240
rect 13340 3210 13345 3240
rect 13305 3205 13345 3210
rect 13605 3240 13645 3245
rect 13605 3210 13610 3240
rect 13610 3210 13640 3240
rect 13640 3210 13645 3240
rect 13605 3205 13645 3210
rect 13755 3240 13795 3245
rect 13755 3210 13760 3240
rect 13760 3210 13790 3240
rect 13790 3210 13795 3240
rect 13755 3205 13795 3210
rect 13905 3240 13945 3245
rect 13905 3210 13910 3240
rect 13910 3210 13940 3240
rect 13940 3210 13945 3240
rect 13905 3205 13945 3210
rect 14205 3240 14245 3245
rect 14205 3210 14210 3240
rect 14210 3210 14240 3240
rect 14240 3210 14245 3240
rect 14205 3205 14245 3210
rect 14505 3240 14545 3245
rect 14505 3210 14510 3240
rect 14510 3210 14540 3240
rect 14540 3210 14545 3240
rect 14505 3205 14545 3210
rect 14805 3240 14845 3245
rect 14805 3210 14810 3240
rect 14810 3210 14840 3240
rect 14840 3210 14845 3240
rect 14805 3205 14845 3210
rect 14955 3240 14995 3245
rect 14955 3210 14960 3240
rect 14960 3210 14990 3240
rect 14990 3210 14995 3240
rect 14955 3205 14995 3210
rect 15105 3240 15145 3245
rect 15105 3210 15110 3240
rect 15110 3210 15140 3240
rect 15140 3210 15145 3240
rect 15105 3205 15145 3210
rect 15405 3240 15445 3245
rect 15405 3210 15410 3240
rect 15410 3210 15440 3240
rect 15440 3210 15445 3240
rect 15405 3205 15445 3210
rect 15705 3240 15745 3245
rect 15705 3210 15710 3240
rect 15710 3210 15740 3240
rect 15740 3210 15745 3240
rect 15705 3205 15745 3210
rect 16005 3240 16045 3245
rect 16005 3210 16010 3240
rect 16010 3210 16040 3240
rect 16040 3210 16045 3240
rect 16005 3205 16045 3210
rect 16305 3240 16345 3245
rect 16305 3210 16310 3240
rect 16310 3210 16340 3240
rect 16340 3210 16345 3240
rect 16305 3205 16345 3210
rect 16605 3240 16645 3245
rect 16605 3210 16610 3240
rect 16610 3210 16640 3240
rect 16640 3210 16645 3240
rect 16605 3205 16645 3210
rect 16755 3240 16795 3245
rect 16755 3210 16760 3240
rect 16760 3210 16790 3240
rect 16790 3210 16795 3240
rect 16755 3205 16795 3210
rect 16905 3240 16945 3245
rect 16905 3210 16910 3240
rect 16910 3210 16940 3240
rect 16940 3210 16945 3240
rect 16905 3205 16945 3210
rect 17205 3240 17245 3245
rect 17205 3210 17210 3240
rect 17210 3210 17240 3240
rect 17240 3210 17245 3240
rect 17205 3205 17245 3210
rect 17505 3240 17545 3245
rect 17505 3210 17510 3240
rect 17510 3210 17540 3240
rect 17540 3210 17545 3240
rect 17505 3205 17545 3210
rect 17805 3240 17845 3245
rect 17805 3210 17810 3240
rect 17810 3210 17840 3240
rect 17840 3210 17845 3240
rect 17805 3205 17845 3210
rect 18105 3240 18145 3245
rect 18105 3210 18110 3240
rect 18110 3210 18140 3240
rect 18140 3210 18145 3240
rect 18105 3205 18145 3210
rect 18405 3240 18445 3245
rect 18405 3210 18410 3240
rect 18410 3210 18440 3240
rect 18440 3210 18445 3240
rect 18405 3205 18445 3210
rect 18705 3240 18745 3245
rect 18705 3210 18710 3240
rect 18710 3210 18740 3240
rect 18740 3210 18745 3240
rect 18705 3205 18745 3210
rect 19005 3240 19045 3245
rect 19005 3210 19010 3240
rect 19010 3210 19040 3240
rect 19040 3210 19045 3240
rect 19005 3205 19045 3210
rect 19155 3240 19195 3245
rect 19155 3210 19160 3240
rect 19160 3210 19190 3240
rect 19190 3210 19195 3240
rect 19155 3205 19195 3210
rect 19305 3240 19345 3245
rect 19305 3210 19310 3240
rect 19310 3210 19340 3240
rect 19340 3210 19345 3240
rect 19305 3205 19345 3210
rect 19605 3240 19645 3245
rect 19605 3210 19610 3240
rect 19610 3210 19640 3240
rect 19640 3210 19645 3240
rect 19605 3205 19645 3210
rect 19905 3240 19945 3245
rect 19905 3210 19910 3240
rect 19910 3210 19940 3240
rect 19940 3210 19945 3240
rect 19905 3205 19945 3210
rect 20205 3240 20245 3245
rect 20205 3210 20210 3240
rect 20210 3210 20240 3240
rect 20240 3210 20245 3240
rect 20205 3205 20245 3210
rect -345 3005 -305 3045
rect 105 3005 145 3045
rect 405 3005 445 3045
rect 2055 3005 2095 3045
rect 3705 3005 3745 3045
rect 4005 3005 4045 3045
rect 4305 3005 4345 3045
rect 4605 3005 4645 3045
rect 6255 3005 6295 3045
rect 7905 3005 7945 3045
rect 8205 3005 8245 3045
rect 705 2905 745 2945
rect 1005 2905 1045 2945
rect 1155 2905 1195 2945
rect 1305 2905 1345 2945
rect 1605 2905 1645 2945
rect 2505 2905 2545 2945
rect 2805 2905 2845 2945
rect 2955 2905 2995 2945
rect 3105 2905 3145 2945
rect 3405 2905 3445 2945
rect 4905 2905 4945 2945
rect 5205 2905 5245 2945
rect 5355 2905 5395 2945
rect 5505 2905 5545 2945
rect 5805 2905 5845 2945
rect 6705 2905 6745 2945
rect 7005 2905 7045 2945
rect 7155 2905 7195 2945
rect 7305 2905 7345 2945
rect 7605 2905 7645 2945
rect 9555 2905 9595 2945
rect 1905 2805 1945 2845
rect 2205 2805 2245 2845
rect 6105 2805 6145 2845
rect 6405 2805 6445 2845
rect -495 2705 -455 2745
rect -195 2705 -155 2745
rect 13305 2305 13345 2345
rect 13605 2305 13645 2345
rect 13905 2305 13945 2345
rect 14205 2305 14245 2345
rect 18705 2305 18745 2345
rect 19005 2305 19045 2345
rect 19305 2305 19345 2345
rect 19605 2305 19645 2345
rect 12105 2105 12145 2145
rect 12405 2105 12445 2145
rect 12705 2105 12745 2145
rect 13005 2105 13045 2145
rect 16305 2105 16345 2145
rect 16605 2105 16645 2145
rect 16905 2105 16945 2145
rect 17205 2105 17245 2145
rect -495 1305 -455 1345
rect -195 1305 -155 1345
rect 3705 1205 3745 1245
rect 4005 1205 4045 1245
rect 4305 1205 4345 1245
rect 4605 1205 4645 1245
rect 1305 1105 1345 1145
rect 1605 1105 1645 1145
rect 1905 1105 1945 1145
rect 2205 1105 2245 1145
rect 2355 1105 2395 1145
rect 2505 1105 2545 1145
rect 2805 1105 2845 1145
rect 3105 1105 3145 1145
rect 3405 1105 3445 1145
rect 4905 1105 4945 1145
rect 5205 1105 5245 1145
rect 5505 1105 5545 1145
rect 5805 1105 5845 1145
rect 5955 1105 5995 1145
rect 6105 1105 6145 1145
rect 6405 1105 6445 1145
rect 6705 1105 6745 1145
rect 7005 1105 7045 1145
rect -345 1005 -305 1045
rect 105 1005 145 1045
rect 405 1005 445 1045
rect 705 1005 745 1045
rect 1005 1005 1045 1045
rect 3855 1005 3895 1045
rect 4455 1005 4495 1045
rect 7305 1005 7345 1045
rect 7605 1005 7645 1045
rect 7905 1005 7945 1045
rect 8205 1005 8245 1045
rect 8505 1005 8545 1045
rect 8805 1005 8845 1045
rect 9105 1005 9145 1045
rect 9405 1005 9445 1045
rect 9705 1005 9745 1045
rect 10005 1005 10045 1045
rect 10305 1005 10345 1045
rect 10605 1005 10645 1045
rect 10905 1005 10945 1045
rect 11205 1005 11245 1045
rect 11505 1005 11545 1045
rect 11805 1005 11845 1045
rect 14505 1005 14545 1045
rect 14805 1005 14845 1045
rect 15105 1005 15145 1045
rect 15405 1005 15445 1045
rect -495 840 -455 845
rect -495 810 -490 840
rect -490 810 -460 840
rect -460 810 -455 840
rect -495 805 -455 810
rect -345 840 -305 845
rect -345 810 -340 840
rect -340 810 -310 840
rect -310 810 -305 840
rect -345 805 -305 810
rect -195 840 -155 845
rect -195 810 -190 840
rect -190 810 -160 840
rect -160 810 -155 840
rect -195 805 -155 810
rect 105 840 145 845
rect 105 810 110 840
rect 110 810 140 840
rect 140 810 145 840
rect 105 805 145 810
rect 405 840 445 845
rect 405 810 410 840
rect 410 810 440 840
rect 440 810 445 840
rect 405 805 445 810
rect 705 840 745 845
rect 705 810 710 840
rect 710 810 740 840
rect 740 810 745 840
rect 705 805 745 810
rect 1005 840 1045 845
rect 1005 810 1010 840
rect 1010 810 1040 840
rect 1040 810 1045 840
rect 1005 805 1045 810
rect 1305 840 1345 845
rect 1305 810 1310 840
rect 1310 810 1340 840
rect 1340 810 1345 840
rect 1305 805 1345 810
rect 1605 840 1645 845
rect 1605 810 1610 840
rect 1610 810 1640 840
rect 1640 810 1645 840
rect 1605 805 1645 810
rect 1905 840 1945 845
rect 1905 810 1910 840
rect 1910 810 1940 840
rect 1940 810 1945 840
rect 1905 805 1945 810
rect 2205 840 2245 845
rect 2205 810 2210 840
rect 2210 810 2240 840
rect 2240 810 2245 840
rect 2205 805 2245 810
rect 2355 840 2395 845
rect 2355 810 2360 840
rect 2360 810 2390 840
rect 2390 810 2395 840
rect 2355 805 2395 810
rect 2505 840 2545 845
rect 2505 810 2510 840
rect 2510 810 2540 840
rect 2540 810 2545 840
rect 2505 805 2545 810
rect 2805 840 2845 845
rect 2805 810 2810 840
rect 2810 810 2840 840
rect 2840 810 2845 840
rect 2805 805 2845 810
rect 3105 840 3145 845
rect 3105 810 3110 840
rect 3110 810 3140 840
rect 3140 810 3145 840
rect 3105 805 3145 810
rect 3405 840 3445 845
rect 3405 810 3410 840
rect 3410 810 3440 840
rect 3440 810 3445 840
rect 3405 805 3445 810
rect 3705 840 3745 845
rect 3705 810 3710 840
rect 3710 810 3740 840
rect 3740 810 3745 840
rect 3705 805 3745 810
rect 3855 840 3895 845
rect 3855 810 3860 840
rect 3860 810 3890 840
rect 3890 810 3895 840
rect 3855 805 3895 810
rect 4005 840 4045 845
rect 4005 810 4010 840
rect 4010 810 4040 840
rect 4040 810 4045 840
rect 4005 805 4045 810
rect 4305 840 4345 845
rect 4305 810 4310 840
rect 4310 810 4340 840
rect 4340 810 4345 840
rect 4305 805 4345 810
rect 4455 840 4495 845
rect 4455 810 4460 840
rect 4460 810 4490 840
rect 4490 810 4495 840
rect 4455 805 4495 810
rect 4605 840 4645 845
rect 4605 810 4610 840
rect 4610 810 4640 840
rect 4640 810 4645 840
rect 4605 805 4645 810
rect 4905 840 4945 845
rect 4905 810 4910 840
rect 4910 810 4940 840
rect 4940 810 4945 840
rect 4905 805 4945 810
rect 5205 840 5245 845
rect 5205 810 5210 840
rect 5210 810 5240 840
rect 5240 810 5245 840
rect 5205 805 5245 810
rect 5505 840 5545 845
rect 5505 810 5510 840
rect 5510 810 5540 840
rect 5540 810 5545 840
rect 5505 805 5545 810
rect 5805 840 5845 845
rect 5805 810 5810 840
rect 5810 810 5840 840
rect 5840 810 5845 840
rect 5805 805 5845 810
rect 5955 840 5995 845
rect 5955 810 5960 840
rect 5960 810 5990 840
rect 5990 810 5995 840
rect 5955 805 5995 810
rect 6105 840 6145 845
rect 6105 810 6110 840
rect 6110 810 6140 840
rect 6140 810 6145 840
rect 6105 805 6145 810
rect 6405 840 6445 845
rect 6405 810 6410 840
rect 6410 810 6440 840
rect 6440 810 6445 840
rect 6405 805 6445 810
rect 6705 840 6745 845
rect 6705 810 6710 840
rect 6710 810 6740 840
rect 6740 810 6745 840
rect 6705 805 6745 810
rect 7005 840 7045 845
rect 7005 810 7010 840
rect 7010 810 7040 840
rect 7040 810 7045 840
rect 7005 805 7045 810
rect 7305 840 7345 845
rect 7305 810 7310 840
rect 7310 810 7340 840
rect 7340 810 7345 840
rect 7305 805 7345 810
rect 7605 840 7645 845
rect 7605 810 7610 840
rect 7610 810 7640 840
rect 7640 810 7645 840
rect 7605 805 7645 810
rect 7905 840 7945 845
rect 7905 810 7910 840
rect 7910 810 7940 840
rect 7940 810 7945 840
rect 7905 805 7945 810
rect 8205 840 8245 845
rect 8205 810 8210 840
rect 8210 810 8240 840
rect 8240 810 8245 840
rect 8205 805 8245 810
rect 8505 840 8545 845
rect 8505 810 8510 840
rect 8510 810 8540 840
rect 8540 810 8545 840
rect 8505 805 8545 810
rect 8805 840 8845 845
rect 8805 810 8810 840
rect 8810 810 8840 840
rect 8840 810 8845 840
rect 8805 805 8845 810
rect 9105 840 9145 845
rect 9105 810 9110 840
rect 9110 810 9140 840
rect 9140 810 9145 840
rect 9105 805 9145 810
rect 9405 840 9445 845
rect 9405 810 9410 840
rect 9410 810 9440 840
rect 9440 810 9445 840
rect 9405 805 9445 810
rect 9555 840 9595 845
rect 9555 810 9560 840
rect 9560 810 9590 840
rect 9590 810 9595 840
rect 9555 805 9595 810
rect 9705 840 9745 845
rect 9705 810 9710 840
rect 9710 810 9740 840
rect 9740 810 9745 840
rect 9705 805 9745 810
rect 10005 840 10045 845
rect 10005 810 10010 840
rect 10010 810 10040 840
rect 10040 810 10045 840
rect 10005 805 10045 810
rect 10305 840 10345 845
rect 10305 810 10310 840
rect 10310 810 10340 840
rect 10340 810 10345 840
rect 10305 805 10345 810
rect 10605 840 10645 845
rect 10605 810 10610 840
rect 10610 810 10640 840
rect 10640 810 10645 840
rect 10605 805 10645 810
rect 10905 840 10945 845
rect 10905 810 10910 840
rect 10910 810 10940 840
rect 10940 810 10945 840
rect 10905 805 10945 810
rect 11205 840 11245 845
rect 11205 810 11210 840
rect 11210 810 11240 840
rect 11240 810 11245 840
rect 11205 805 11245 810
rect 11505 840 11545 845
rect 11505 810 11510 840
rect 11510 810 11540 840
rect 11540 810 11545 840
rect 11505 805 11545 810
rect 11805 840 11845 845
rect 11805 810 11810 840
rect 11810 810 11840 840
rect 11840 810 11845 840
rect 11805 805 11845 810
rect 12105 840 12145 845
rect 12105 810 12110 840
rect 12110 810 12140 840
rect 12140 810 12145 840
rect 12105 805 12145 810
rect 12405 840 12445 845
rect 12405 810 12410 840
rect 12410 810 12440 840
rect 12440 810 12445 840
rect 12405 805 12445 810
rect 12555 840 12595 845
rect 12555 810 12560 840
rect 12560 810 12590 840
rect 12590 810 12595 840
rect 12555 805 12595 810
rect 12705 840 12745 845
rect 12705 810 12710 840
rect 12710 810 12740 840
rect 12740 810 12745 840
rect 12705 805 12745 810
rect 13005 840 13045 845
rect 13005 810 13010 840
rect 13010 810 13040 840
rect 13040 810 13045 840
rect 13005 805 13045 810
rect 13305 840 13345 845
rect 13305 810 13310 840
rect 13310 810 13340 840
rect 13340 810 13345 840
rect 13305 805 13345 810
rect 13605 840 13645 845
rect 13605 810 13610 840
rect 13610 810 13640 840
rect 13640 810 13645 840
rect 13605 805 13645 810
rect 13755 840 13795 845
rect 13755 810 13760 840
rect 13760 810 13790 840
rect 13790 810 13795 840
rect 13755 805 13795 810
rect 13905 840 13945 845
rect 13905 810 13910 840
rect 13910 810 13940 840
rect 13940 810 13945 840
rect 13905 805 13945 810
rect 14205 840 14245 845
rect 14205 810 14210 840
rect 14210 810 14240 840
rect 14240 810 14245 840
rect 14205 805 14245 810
rect 14505 840 14545 845
rect 14505 810 14510 840
rect 14510 810 14540 840
rect 14540 810 14545 840
rect 14505 805 14545 810
rect 14805 840 14845 845
rect 14805 810 14810 840
rect 14810 810 14840 840
rect 14840 810 14845 840
rect 14805 805 14845 810
rect 15105 840 15145 845
rect 15105 810 15110 840
rect 15110 810 15140 840
rect 15140 810 15145 840
rect 15105 805 15145 810
rect 15405 840 15445 845
rect 15405 810 15410 840
rect 15410 810 15440 840
rect 15440 810 15445 840
rect 15405 805 15445 810
rect 15705 840 15745 845
rect 15705 810 15710 840
rect 15710 810 15740 840
rect 15740 810 15745 840
rect 15705 805 15745 810
rect 16005 840 16045 845
rect 16005 810 16010 840
rect 16010 810 16040 840
rect 16040 810 16045 840
rect 16005 805 16045 810
rect 16305 840 16345 845
rect 16305 810 16310 840
rect 16310 810 16340 840
rect 16340 810 16345 840
rect 16305 805 16345 810
rect 16605 840 16645 845
rect 16605 810 16610 840
rect 16610 810 16640 840
rect 16640 810 16645 840
rect 16605 805 16645 810
rect 16755 840 16795 845
rect 16755 810 16760 840
rect 16760 810 16790 840
rect 16790 810 16795 840
rect 16755 805 16795 810
rect 16905 840 16945 845
rect 16905 810 16910 840
rect 16910 810 16940 840
rect 16940 810 16945 840
rect 16905 805 16945 810
rect 17205 840 17245 845
rect 17205 810 17210 840
rect 17210 810 17240 840
rect 17240 810 17245 840
rect 17205 805 17245 810
rect 17505 840 17545 845
rect 17505 810 17510 840
rect 17510 810 17540 840
rect 17540 810 17545 840
rect 17505 805 17545 810
rect 17805 840 17845 845
rect 17805 810 17810 840
rect 17810 810 17840 840
rect 17840 810 17845 840
rect 17805 805 17845 810
rect 18105 840 18145 845
rect 18105 810 18110 840
rect 18110 810 18140 840
rect 18140 810 18145 840
rect 18105 805 18145 810
rect 18405 840 18445 845
rect 18405 810 18410 840
rect 18410 810 18440 840
rect 18440 810 18445 840
rect 18405 805 18445 810
rect 18705 840 18745 845
rect 18705 810 18710 840
rect 18710 810 18740 840
rect 18740 810 18745 840
rect 18705 805 18745 810
rect 19005 840 19045 845
rect 19005 810 19010 840
rect 19010 810 19040 840
rect 19040 810 19045 840
rect 19005 805 19045 810
rect 19155 840 19195 845
rect 19155 810 19160 840
rect 19160 810 19190 840
rect 19190 810 19195 840
rect 19155 805 19195 810
rect 19305 840 19345 845
rect 19305 810 19310 840
rect 19310 810 19340 840
rect 19340 810 19345 840
rect 19305 805 19345 810
rect 19605 840 19645 845
rect 19605 810 19610 840
rect 19610 810 19640 840
rect 19640 810 19645 840
rect 19605 805 19645 810
rect 19905 840 19945 845
rect 19905 810 19910 840
rect 19910 810 19940 840
rect 19940 810 19945 840
rect 19905 805 19945 810
rect 20205 840 20245 845
rect 20205 810 20210 840
rect 20210 810 20240 840
rect 20240 810 20245 840
rect 20205 805 20245 810
rect 15705 605 15745 645
rect 16005 605 16045 645
rect 16305 605 16345 645
rect 16605 605 16645 645
rect 16905 605 16945 645
rect 17205 605 17245 645
rect 17505 605 17545 645
rect 17805 605 17845 645
rect 18105 405 18145 445
rect 18405 405 18445 445
rect 18705 405 18745 445
rect 19005 405 19045 445
rect 19305 405 19345 445
rect 19605 405 19645 445
rect 19905 405 19945 445
rect 20205 405 20245 445
rect -495 -860 -455 -855
rect -495 -890 -490 -860
rect -490 -890 -460 -860
rect -460 -890 -455 -860
rect -495 -895 -455 -890
rect -345 -860 -305 -855
rect -345 -890 -340 -860
rect -340 -890 -310 -860
rect -310 -890 -305 -860
rect -345 -895 -305 -890
rect -195 -860 -155 -855
rect -195 -890 -190 -860
rect -190 -890 -160 -860
rect -160 -890 -155 -860
rect -195 -895 -155 -890
rect 105 -860 145 -855
rect 105 -890 110 -860
rect 110 -890 140 -860
rect 140 -890 145 -860
rect 105 -895 145 -890
rect 405 -860 445 -855
rect 405 -890 410 -860
rect 410 -890 440 -860
rect 440 -890 445 -860
rect 405 -895 445 -890
rect 705 -860 745 -855
rect 705 -890 710 -860
rect 710 -890 740 -860
rect 740 -890 745 -860
rect 705 -895 745 -890
rect 1005 -860 1045 -855
rect 1005 -890 1010 -860
rect 1010 -890 1040 -860
rect 1040 -890 1045 -860
rect 1005 -895 1045 -890
rect 1305 -860 1345 -855
rect 1305 -890 1310 -860
rect 1310 -890 1340 -860
rect 1340 -890 1345 -860
rect 1305 -895 1345 -890
rect 1605 -860 1645 -855
rect 1605 -890 1610 -860
rect 1610 -890 1640 -860
rect 1640 -890 1645 -860
rect 1605 -895 1645 -890
rect 1905 -860 1945 -855
rect 1905 -890 1910 -860
rect 1910 -890 1940 -860
rect 1940 -890 1945 -860
rect 1905 -895 1945 -890
rect 2205 -860 2245 -855
rect 2205 -890 2210 -860
rect 2210 -890 2240 -860
rect 2240 -890 2245 -860
rect 2205 -895 2245 -890
rect 2355 -860 2395 -855
rect 2355 -890 2360 -860
rect 2360 -890 2390 -860
rect 2390 -890 2395 -860
rect 2355 -895 2395 -890
rect 2505 -860 2545 -855
rect 2505 -890 2510 -860
rect 2510 -890 2540 -860
rect 2540 -890 2545 -860
rect 2505 -895 2545 -890
rect 2805 -860 2845 -855
rect 2805 -890 2810 -860
rect 2810 -890 2840 -860
rect 2840 -890 2845 -860
rect 2805 -895 2845 -890
rect 3105 -860 3145 -855
rect 3105 -890 3110 -860
rect 3110 -890 3140 -860
rect 3140 -890 3145 -860
rect 3105 -895 3145 -890
rect 3405 -860 3445 -855
rect 3405 -890 3410 -860
rect 3410 -890 3440 -860
rect 3440 -890 3445 -860
rect 3405 -895 3445 -890
rect 3705 -860 3745 -855
rect 3705 -890 3710 -860
rect 3710 -890 3740 -860
rect 3740 -890 3745 -860
rect 3705 -895 3745 -890
rect 3855 -860 3895 -855
rect 3855 -890 3860 -860
rect 3860 -890 3890 -860
rect 3890 -890 3895 -860
rect 3855 -895 3895 -890
rect 4005 -860 4045 -855
rect 4005 -890 4010 -860
rect 4010 -890 4040 -860
rect 4040 -890 4045 -860
rect 4005 -895 4045 -890
rect 4305 -860 4345 -855
rect 4305 -890 4310 -860
rect 4310 -890 4340 -860
rect 4340 -890 4345 -860
rect 4305 -895 4345 -890
rect 4455 -860 4495 -855
rect 4455 -890 4460 -860
rect 4460 -890 4490 -860
rect 4490 -890 4495 -860
rect 4455 -895 4495 -890
rect 4605 -860 4645 -855
rect 4605 -890 4610 -860
rect 4610 -890 4640 -860
rect 4640 -890 4645 -860
rect 4605 -895 4645 -890
rect 4905 -860 4945 -855
rect 4905 -890 4910 -860
rect 4910 -890 4940 -860
rect 4940 -890 4945 -860
rect 4905 -895 4945 -890
rect 5205 -860 5245 -855
rect 5205 -890 5210 -860
rect 5210 -890 5240 -860
rect 5240 -890 5245 -860
rect 5205 -895 5245 -890
rect 5505 -860 5545 -855
rect 5505 -890 5510 -860
rect 5510 -890 5540 -860
rect 5540 -890 5545 -860
rect 5505 -895 5545 -890
rect 5805 -860 5845 -855
rect 5805 -890 5810 -860
rect 5810 -890 5840 -860
rect 5840 -890 5845 -860
rect 5805 -895 5845 -890
rect 5955 -860 5995 -855
rect 5955 -890 5960 -860
rect 5960 -890 5990 -860
rect 5990 -890 5995 -860
rect 5955 -895 5995 -890
rect 6105 -860 6145 -855
rect 6105 -890 6110 -860
rect 6110 -890 6140 -860
rect 6140 -890 6145 -860
rect 6105 -895 6145 -890
rect 6405 -860 6445 -855
rect 6405 -890 6410 -860
rect 6410 -890 6440 -860
rect 6440 -890 6445 -860
rect 6405 -895 6445 -890
rect 6705 -860 6745 -855
rect 6705 -890 6710 -860
rect 6710 -890 6740 -860
rect 6740 -890 6745 -860
rect 6705 -895 6745 -890
rect 7005 -860 7045 -855
rect 7005 -890 7010 -860
rect 7010 -890 7040 -860
rect 7040 -890 7045 -860
rect 7005 -895 7045 -890
rect 7305 -860 7345 -855
rect 7305 -890 7310 -860
rect 7310 -890 7340 -860
rect 7340 -890 7345 -860
rect 7305 -895 7345 -890
rect 7605 -860 7645 -855
rect 7605 -890 7610 -860
rect 7610 -890 7640 -860
rect 7640 -890 7645 -860
rect 7605 -895 7645 -890
rect 7905 -860 7945 -855
rect 7905 -890 7910 -860
rect 7910 -890 7940 -860
rect 7940 -890 7945 -860
rect 7905 -895 7945 -890
rect 8205 -860 8245 -855
rect 8205 -890 8210 -860
rect 8210 -890 8240 -860
rect 8240 -890 8245 -860
rect 8205 -895 8245 -890
rect 8505 -860 8545 -855
rect 8505 -890 8510 -860
rect 8510 -890 8540 -860
rect 8540 -890 8545 -860
rect 8505 -895 8545 -890
rect 8805 -860 8845 -855
rect 8805 -890 8810 -860
rect 8810 -890 8840 -860
rect 8840 -890 8845 -860
rect 8805 -895 8845 -890
rect 9105 -860 9145 -855
rect 9105 -890 9110 -860
rect 9110 -890 9140 -860
rect 9140 -890 9145 -860
rect 9105 -895 9145 -890
rect 9405 -860 9445 -855
rect 9405 -890 9410 -860
rect 9410 -890 9440 -860
rect 9440 -890 9445 -860
rect 9405 -895 9445 -890
rect 9555 -860 9595 -855
rect 9555 -890 9560 -860
rect 9560 -890 9590 -860
rect 9590 -890 9595 -860
rect 9555 -895 9595 -890
rect 9705 -860 9745 -855
rect 9705 -890 9710 -860
rect 9710 -890 9740 -860
rect 9740 -890 9745 -860
rect 9705 -895 9745 -890
rect 10005 -860 10045 -855
rect 10005 -890 10010 -860
rect 10010 -890 10040 -860
rect 10040 -890 10045 -860
rect 10005 -895 10045 -890
rect 10305 -860 10345 -855
rect 10305 -890 10310 -860
rect 10310 -890 10340 -860
rect 10340 -890 10345 -860
rect 10305 -895 10345 -890
rect 10605 -860 10645 -855
rect 10605 -890 10610 -860
rect 10610 -890 10640 -860
rect 10640 -890 10645 -860
rect 10605 -895 10645 -890
rect 10905 -860 10945 -855
rect 10905 -890 10910 -860
rect 10910 -890 10940 -860
rect 10940 -890 10945 -860
rect 10905 -895 10945 -890
rect 11205 -860 11245 -855
rect 11205 -890 11210 -860
rect 11210 -890 11240 -860
rect 11240 -890 11245 -860
rect 11205 -895 11245 -890
rect 11505 -860 11545 -855
rect 11505 -890 11510 -860
rect 11510 -890 11540 -860
rect 11540 -890 11545 -860
rect 11505 -895 11545 -890
rect 11805 -860 11845 -855
rect 11805 -890 11810 -860
rect 11810 -890 11840 -860
rect 11840 -890 11845 -860
rect 11805 -895 11845 -890
rect 12105 -860 12145 -855
rect 12105 -890 12110 -860
rect 12110 -890 12140 -860
rect 12140 -890 12145 -860
rect 12105 -895 12145 -890
rect 12405 -860 12445 -855
rect 12405 -890 12410 -860
rect 12410 -890 12440 -860
rect 12440 -890 12445 -860
rect 12405 -895 12445 -890
rect 12555 -860 12595 -855
rect 12555 -890 12560 -860
rect 12560 -890 12590 -860
rect 12590 -890 12595 -860
rect 12555 -895 12595 -890
rect 12705 -860 12745 -855
rect 12705 -890 12710 -860
rect 12710 -890 12740 -860
rect 12740 -890 12745 -860
rect 12705 -895 12745 -890
rect 13005 -860 13045 -855
rect 13005 -890 13010 -860
rect 13010 -890 13040 -860
rect 13040 -890 13045 -860
rect 13005 -895 13045 -890
rect 13305 -860 13345 -855
rect 13305 -890 13310 -860
rect 13310 -890 13340 -860
rect 13340 -890 13345 -860
rect 13305 -895 13345 -890
rect 13605 -860 13645 -855
rect 13605 -890 13610 -860
rect 13610 -890 13640 -860
rect 13640 -890 13645 -860
rect 13605 -895 13645 -890
rect 13755 -860 13795 -855
rect 13755 -890 13760 -860
rect 13760 -890 13790 -860
rect 13790 -890 13795 -860
rect 13755 -895 13795 -890
rect 13905 -860 13945 -855
rect 13905 -890 13910 -860
rect 13910 -890 13940 -860
rect 13940 -890 13945 -860
rect 13905 -895 13945 -890
rect 14205 -860 14245 -855
rect 14205 -890 14210 -860
rect 14210 -890 14240 -860
rect 14240 -890 14245 -860
rect 14205 -895 14245 -890
rect 14505 -860 14545 -855
rect 14505 -890 14510 -860
rect 14510 -890 14540 -860
rect 14540 -890 14545 -860
rect 14505 -895 14545 -890
rect 14805 -860 14845 -855
rect 14805 -890 14810 -860
rect 14810 -890 14840 -860
rect 14840 -890 14845 -860
rect 14805 -895 14845 -890
rect 15105 -860 15145 -855
rect 15105 -890 15110 -860
rect 15110 -890 15140 -860
rect 15140 -890 15145 -860
rect 15105 -895 15145 -890
rect 15405 -860 15445 -855
rect 15405 -890 15410 -860
rect 15410 -890 15440 -860
rect 15440 -890 15445 -860
rect 15405 -895 15445 -890
rect 15705 -860 15745 -855
rect 15705 -890 15710 -860
rect 15710 -890 15740 -860
rect 15740 -890 15745 -860
rect 15705 -895 15745 -890
rect 16005 -860 16045 -855
rect 16005 -890 16010 -860
rect 16010 -890 16040 -860
rect 16040 -890 16045 -860
rect 16005 -895 16045 -890
rect 16305 -860 16345 -855
rect 16305 -890 16310 -860
rect 16310 -890 16340 -860
rect 16340 -890 16345 -860
rect 16305 -895 16345 -890
rect 16605 -860 16645 -855
rect 16605 -890 16610 -860
rect 16610 -890 16640 -860
rect 16640 -890 16645 -860
rect 16605 -895 16645 -890
rect 16755 -860 16795 -855
rect 16755 -890 16760 -860
rect 16760 -890 16790 -860
rect 16790 -890 16795 -860
rect 16755 -895 16795 -890
rect 16905 -860 16945 -855
rect 16905 -890 16910 -860
rect 16910 -890 16940 -860
rect 16940 -890 16945 -860
rect 16905 -895 16945 -890
rect 17205 -860 17245 -855
rect 17205 -890 17210 -860
rect 17210 -890 17240 -860
rect 17240 -890 17245 -860
rect 17205 -895 17245 -890
rect 17505 -860 17545 -855
rect 17505 -890 17510 -860
rect 17510 -890 17540 -860
rect 17540 -890 17545 -860
rect 17505 -895 17545 -890
rect 17805 -860 17845 -855
rect 17805 -890 17810 -860
rect 17810 -890 17840 -860
rect 17840 -890 17845 -860
rect 17805 -895 17845 -890
rect 18105 -860 18145 -855
rect 18105 -890 18110 -860
rect 18110 -890 18140 -860
rect 18140 -890 18145 -860
rect 18105 -895 18145 -890
rect 18405 -860 18445 -855
rect 18405 -890 18410 -860
rect 18410 -890 18440 -860
rect 18440 -890 18445 -860
rect 18405 -895 18445 -890
rect 18705 -860 18745 -855
rect 18705 -890 18710 -860
rect 18710 -890 18740 -860
rect 18740 -890 18745 -860
rect 18705 -895 18745 -890
rect 19005 -860 19045 -855
rect 19005 -890 19010 -860
rect 19010 -890 19040 -860
rect 19040 -890 19045 -860
rect 19005 -895 19045 -890
rect 19155 -860 19195 -855
rect 19155 -890 19160 -860
rect 19160 -890 19190 -860
rect 19190 -890 19195 -860
rect 19155 -895 19195 -890
rect 19305 -860 19345 -855
rect 19305 -890 19310 -860
rect 19310 -890 19340 -860
rect 19340 -890 19345 -860
rect 19305 -895 19345 -890
rect 19605 -860 19645 -855
rect 19605 -890 19610 -860
rect 19610 -890 19640 -860
rect 19640 -890 19645 -860
rect 19605 -895 19645 -890
rect 19905 -860 19945 -855
rect 19905 -890 19910 -860
rect 19910 -890 19940 -860
rect 19940 -890 19945 -860
rect 19905 -895 19945 -890
rect 20205 -860 20245 -855
rect 20205 -890 20210 -860
rect 20210 -890 20240 -860
rect 20240 -890 20245 -860
rect 20205 -895 20245 -890
<< metal4 >>
rect -500 4545 -450 4550
rect -500 4505 -495 4545
rect -455 4505 -450 4545
rect -500 3245 -450 4505
rect -500 3205 -495 3245
rect -455 3205 -450 3245
rect -500 2745 -450 3205
rect -350 4545 -300 4600
rect -350 4505 -345 4545
rect -305 4505 -300 4545
rect -350 3245 -300 4505
rect -350 3205 -345 3245
rect -305 3205 -300 3245
rect -350 3045 -300 3205
rect -350 3005 -345 3045
rect -305 3005 -300 3045
rect -350 3000 -300 3005
rect -200 4545 -150 4550
rect -200 4505 -195 4545
rect -155 4505 -150 4545
rect -200 3245 -150 4505
rect -200 3205 -195 3245
rect -155 3205 -150 3245
rect -500 2705 -495 2745
rect -455 2705 -450 2745
rect -500 2700 -450 2705
rect -200 2745 -150 3205
rect 100 4545 150 4550
rect 100 4505 105 4545
rect 145 4505 150 4545
rect 100 3245 150 4505
rect 100 3205 105 3245
rect 145 3205 150 3245
rect 100 3045 150 3205
rect 100 3005 105 3045
rect 145 3005 150 3045
rect 100 3000 150 3005
rect 400 4545 450 4550
rect 400 4505 405 4545
rect 445 4505 450 4545
rect 400 3245 450 4505
rect 400 3205 405 3245
rect 445 3205 450 3245
rect 400 3045 450 3205
rect 400 3005 405 3045
rect 445 3005 450 3045
rect 400 3000 450 3005
rect 700 4545 750 4550
rect 700 4505 705 4545
rect 745 4505 750 4545
rect 700 3245 750 4505
rect 700 3205 705 3245
rect 745 3205 750 3245
rect 700 2945 750 3205
rect 700 2905 705 2945
rect 745 2905 750 2945
rect 700 2900 750 2905
rect 1000 4545 1050 4550
rect 1000 4505 1005 4545
rect 1045 4505 1050 4545
rect 1000 3245 1050 4505
rect 1000 3205 1005 3245
rect 1045 3205 1050 3245
rect 1000 2945 1050 3205
rect 1000 2905 1005 2945
rect 1045 2905 1050 2945
rect 1000 2900 1050 2905
rect 1150 4545 1200 4550
rect 1150 4505 1155 4545
rect 1195 4505 1200 4545
rect 1150 3245 1200 4505
rect 1150 3205 1155 3245
rect 1195 3205 1200 3245
rect 1150 2945 1200 3205
rect 1150 2905 1155 2945
rect 1195 2905 1200 2945
rect 1150 2900 1200 2905
rect 1300 4545 1350 4550
rect 1300 4505 1305 4545
rect 1345 4505 1350 4545
rect 1300 3245 1350 4505
rect 1300 3205 1305 3245
rect 1345 3205 1350 3245
rect 1300 2945 1350 3205
rect 1300 2905 1305 2945
rect 1345 2905 1350 2945
rect 1300 2900 1350 2905
rect 1600 4545 1650 4550
rect 1600 4505 1605 4545
rect 1645 4505 1650 4545
rect 1600 3245 1650 4505
rect 1600 3205 1605 3245
rect 1645 3205 1650 3245
rect 1600 2945 1650 3205
rect 1600 2905 1605 2945
rect 1645 2905 1650 2945
rect 1600 2900 1650 2905
rect 1900 4545 1950 4550
rect 1900 4505 1905 4545
rect 1945 4505 1950 4545
rect 1900 3245 1950 4505
rect 1900 3205 1905 3245
rect 1945 3205 1950 3245
rect 1900 2845 1950 3205
rect 2050 4545 2100 4550
rect 2050 4505 2055 4545
rect 2095 4505 2100 4545
rect 2050 3245 2100 4505
rect 2050 3205 2055 3245
rect 2095 3205 2100 3245
rect 2050 3045 2100 3205
rect 2050 3005 2055 3045
rect 2095 3005 2100 3045
rect 2050 3000 2100 3005
rect 2200 4545 2250 4550
rect 2200 4505 2205 4545
rect 2245 4505 2250 4545
rect 2200 3245 2250 4505
rect 2200 3205 2205 3245
rect 2245 3205 2250 3245
rect 1900 2805 1905 2845
rect 1945 2805 1950 2845
rect 1900 2800 1950 2805
rect 2200 2845 2250 3205
rect 2500 4545 2550 4550
rect 2500 4505 2505 4545
rect 2545 4505 2550 4545
rect 2500 3245 2550 4505
rect 2500 3205 2505 3245
rect 2545 3205 2550 3245
rect 2500 2945 2550 3205
rect 2500 2905 2505 2945
rect 2545 2905 2550 2945
rect 2500 2900 2550 2905
rect 2800 4545 2850 4550
rect 2800 4505 2805 4545
rect 2845 4505 2850 4545
rect 2800 3245 2850 4505
rect 2800 3205 2805 3245
rect 2845 3205 2850 3245
rect 2800 2945 2850 3205
rect 2800 2905 2805 2945
rect 2845 2905 2850 2945
rect 2800 2900 2850 2905
rect 2950 4545 3000 4550
rect 2950 4505 2955 4545
rect 2995 4505 3000 4545
rect 2950 3245 3000 4505
rect 2950 3205 2955 3245
rect 2995 3205 3000 3245
rect 2950 2945 3000 3205
rect 2950 2905 2955 2945
rect 2995 2905 3000 2945
rect 2950 2900 3000 2905
rect 3100 4545 3150 4550
rect 3100 4505 3105 4545
rect 3145 4505 3150 4545
rect 3100 3245 3150 4505
rect 3100 3205 3105 3245
rect 3145 3205 3150 3245
rect 3100 2945 3150 3205
rect 3100 2905 3105 2945
rect 3145 2905 3150 2945
rect 3100 2900 3150 2905
rect 3400 4545 3450 4550
rect 3400 4505 3405 4545
rect 3445 4505 3450 4545
rect 3400 3245 3450 4505
rect 3400 3205 3405 3245
rect 3445 3205 3450 3245
rect 3400 2945 3450 3205
rect 3700 4545 3750 4550
rect 3700 4505 3705 4545
rect 3745 4505 3750 4545
rect 3700 3245 3750 4505
rect 3700 3205 3705 3245
rect 3745 3205 3750 3245
rect 3700 3045 3750 3205
rect 3700 3005 3705 3045
rect 3745 3005 3750 3045
rect 3700 3000 3750 3005
rect 4000 4545 4050 4550
rect 4000 4505 4005 4545
rect 4045 4505 4050 4545
rect 4000 3245 4050 4505
rect 4000 3205 4005 3245
rect 4045 3205 4050 3245
rect 4000 3045 4050 3205
rect 4000 3005 4005 3045
rect 4045 3005 4050 3045
rect 4000 3000 4050 3005
rect 4300 4545 4350 4550
rect 4300 4505 4305 4545
rect 4345 4505 4350 4545
rect 4300 3245 4350 4505
rect 4300 3205 4305 3245
rect 4345 3205 4350 3245
rect 4300 3045 4350 3205
rect 4300 3005 4305 3045
rect 4345 3005 4350 3045
rect 4300 3000 4350 3005
rect 4600 4545 4650 4550
rect 4600 4505 4605 4545
rect 4645 4505 4650 4545
rect 4600 3245 4650 4505
rect 4600 3205 4605 3245
rect 4645 3205 4650 3245
rect 4600 3045 4650 3205
rect 4600 3005 4605 3045
rect 4645 3005 4650 3045
rect 4600 3000 4650 3005
rect 4900 4545 4950 4550
rect 4900 4505 4905 4545
rect 4945 4505 4950 4545
rect 4900 3245 4950 4505
rect 4900 3205 4905 3245
rect 4945 3205 4950 3245
rect 3400 2905 3405 2945
rect 3445 2905 3450 2945
rect 3400 2900 3450 2905
rect 4900 2945 4950 3205
rect 4900 2905 4905 2945
rect 4945 2905 4950 2945
rect 4900 2900 4950 2905
rect 5200 4545 5250 4550
rect 5200 4505 5205 4545
rect 5245 4505 5250 4545
rect 5200 3245 5250 4505
rect 5200 3205 5205 3245
rect 5245 3205 5250 3245
rect 5200 2945 5250 3205
rect 5200 2905 5205 2945
rect 5245 2905 5250 2945
rect 5200 2900 5250 2905
rect 5350 4545 5400 4550
rect 5350 4505 5355 4545
rect 5395 4505 5400 4545
rect 5350 3245 5400 4505
rect 5350 3205 5355 3245
rect 5395 3205 5400 3245
rect 5350 2945 5400 3205
rect 5350 2905 5355 2945
rect 5395 2905 5400 2945
rect 5350 2900 5400 2905
rect 5500 4545 5550 4550
rect 5500 4505 5505 4545
rect 5545 4505 5550 4545
rect 5500 3245 5550 4505
rect 5500 3205 5505 3245
rect 5545 3205 5550 3245
rect 5500 2945 5550 3205
rect 5500 2905 5505 2945
rect 5545 2905 5550 2945
rect 5500 2900 5550 2905
rect 5800 4545 5850 4550
rect 5800 4505 5805 4545
rect 5845 4505 5850 4545
rect 5800 3245 5850 4505
rect 5800 3205 5805 3245
rect 5845 3205 5850 3245
rect 5800 2945 5850 3205
rect 5800 2905 5805 2945
rect 5845 2905 5850 2945
rect 5800 2900 5850 2905
rect 6100 4545 6150 4550
rect 6100 4505 6105 4545
rect 6145 4505 6150 4545
rect 6100 3245 6150 4505
rect 6100 3205 6105 3245
rect 6145 3205 6150 3245
rect 2200 2805 2205 2845
rect 2245 2805 2250 2845
rect 2200 2800 2250 2805
rect 6100 2845 6150 3205
rect 6250 4545 6300 4550
rect 6250 4505 6255 4545
rect 6295 4505 6300 4545
rect 6250 3245 6300 4505
rect 6250 3205 6255 3245
rect 6295 3205 6300 3245
rect 6250 3045 6300 3205
rect 6250 3005 6255 3045
rect 6295 3005 6300 3045
rect 6250 3000 6300 3005
rect 6400 4545 6450 4550
rect 6400 4505 6405 4545
rect 6445 4505 6450 4545
rect 6400 3245 6450 4505
rect 6400 3205 6405 3245
rect 6445 3205 6450 3245
rect 6100 2805 6105 2845
rect 6145 2805 6150 2845
rect 6100 2800 6150 2805
rect 6400 2845 6450 3205
rect 6700 4545 6750 4550
rect 6700 4505 6705 4545
rect 6745 4505 6750 4545
rect 6700 3245 6750 4505
rect 6700 3205 6705 3245
rect 6745 3205 6750 3245
rect 6700 2945 6750 3205
rect 6700 2905 6705 2945
rect 6745 2905 6750 2945
rect 6700 2900 6750 2905
rect 7000 4545 7050 4550
rect 7000 4505 7005 4545
rect 7045 4505 7050 4545
rect 7000 3245 7050 4505
rect 7000 3205 7005 3245
rect 7045 3205 7050 3245
rect 7000 2945 7050 3205
rect 7000 2905 7005 2945
rect 7045 2905 7050 2945
rect 7000 2900 7050 2905
rect 7150 4545 7200 4550
rect 7150 4505 7155 4545
rect 7195 4505 7200 4545
rect 7150 3245 7200 4505
rect 7150 3205 7155 3245
rect 7195 3205 7200 3245
rect 7150 2945 7200 3205
rect 7150 2905 7155 2945
rect 7195 2905 7200 2945
rect 7150 2900 7200 2905
rect 7300 4545 7350 4550
rect 7300 4505 7305 4545
rect 7345 4505 7350 4545
rect 7300 3245 7350 4505
rect 7300 3205 7305 3245
rect 7345 3205 7350 3245
rect 7300 2945 7350 3205
rect 7300 2905 7305 2945
rect 7345 2905 7350 2945
rect 7300 2900 7350 2905
rect 7600 4545 7650 4550
rect 7600 4505 7605 4545
rect 7645 4505 7650 4545
rect 7600 3245 7650 4505
rect 7600 3205 7605 3245
rect 7645 3205 7650 3245
rect 7600 2945 7650 3205
rect 7900 4545 7950 4550
rect 7900 4505 7905 4545
rect 7945 4505 7950 4545
rect 7900 3245 7950 4505
rect 7900 3205 7905 3245
rect 7945 3205 7950 3245
rect 7900 3045 7950 3205
rect 7900 3005 7905 3045
rect 7945 3005 7950 3045
rect 7900 3000 7950 3005
rect 8200 4545 8250 4550
rect 8200 4505 8205 4545
rect 8245 4505 8250 4545
rect 8200 3245 8250 4505
rect 8200 3205 8205 3245
rect 8245 3205 8250 3245
rect 8200 3045 8250 3205
rect 8500 4545 8550 4550
rect 8500 4505 8505 4545
rect 8545 4505 8550 4545
rect 8500 3245 8550 4505
rect 8500 3205 8505 3245
rect 8545 3205 8550 3245
rect 8500 3200 8550 3205
rect 8800 4545 8850 4550
rect 8800 4505 8805 4545
rect 8845 4505 8850 4545
rect 8800 3245 8850 4505
rect 8800 3205 8805 3245
rect 8845 3205 8850 3245
rect 8800 3200 8850 3205
rect 9100 4545 9150 4550
rect 9100 4505 9105 4545
rect 9145 4505 9150 4545
rect 9100 3245 9150 4505
rect 9100 3205 9105 3245
rect 9145 3205 9150 3245
rect 9100 3200 9150 3205
rect 9400 4545 9450 4550
rect 9400 4505 9405 4545
rect 9445 4505 9450 4545
rect 9400 3245 9450 4505
rect 9400 3205 9405 3245
rect 9445 3205 9450 3245
rect 9400 3200 9450 3205
rect 9700 4545 9750 4550
rect 9700 4505 9705 4545
rect 9745 4505 9750 4545
rect 9700 3245 9750 4505
rect 9700 3205 9705 3245
rect 9745 3205 9750 3245
rect 9700 3200 9750 3205
rect 10000 4545 10050 4550
rect 10000 4505 10005 4545
rect 10045 4505 10050 4545
rect 10000 3245 10050 4505
rect 10000 3205 10005 3245
rect 10045 3205 10050 3245
rect 10000 3200 10050 3205
rect 10300 4545 10350 4550
rect 10300 4505 10305 4545
rect 10345 4505 10350 4545
rect 10300 3245 10350 4505
rect 10300 3205 10305 3245
rect 10345 3205 10350 3245
rect 10300 3200 10350 3205
rect 10600 4545 10650 4550
rect 10600 4505 10605 4545
rect 10645 4505 10650 4545
rect 10600 3245 10650 4505
rect 10600 3205 10605 3245
rect 10645 3205 10650 3245
rect 10600 3200 10650 3205
rect 10900 4545 10950 4550
rect 10900 4505 10905 4545
rect 10945 4505 10950 4545
rect 10900 3445 10950 4505
rect 10900 3405 10905 3445
rect 10945 3405 10950 3445
rect 10900 3245 10950 3405
rect 10900 3205 10905 3245
rect 10945 3205 10950 3245
rect 10900 3200 10950 3205
rect 11200 4545 11250 4550
rect 11200 4505 11205 4545
rect 11245 4505 11250 4545
rect 11200 3445 11250 4505
rect 11200 3405 11205 3445
rect 11245 3405 11250 3445
rect 11200 3245 11250 3405
rect 11200 3205 11205 3245
rect 11245 3205 11250 3245
rect 11200 3200 11250 3205
rect 11350 4545 11400 4550
rect 11350 4505 11355 4545
rect 11395 4505 11400 4545
rect 11350 4145 11400 4505
rect 11350 4105 11355 4145
rect 11395 4105 11400 4145
rect 11350 3245 11400 4105
rect 11350 3205 11355 3245
rect 11395 3205 11400 3245
rect 11350 3200 11400 3205
rect 11500 4545 11550 4550
rect 11500 4505 11505 4545
rect 11545 4505 11550 4545
rect 11500 3445 11550 4505
rect 11500 3405 11505 3445
rect 11545 3405 11550 3445
rect 11500 3245 11550 3405
rect 11500 3205 11505 3245
rect 11545 3205 11550 3245
rect 11500 3200 11550 3205
rect 11800 4545 11850 4550
rect 11800 4505 11805 4545
rect 11845 4505 11850 4545
rect 11800 3445 11850 4505
rect 11800 3405 11805 3445
rect 11845 3405 11850 3445
rect 11800 3245 11850 3405
rect 11800 3205 11805 3245
rect 11845 3205 11850 3245
rect 11800 3200 11850 3205
rect 12100 4545 12150 4550
rect 12100 4505 12105 4545
rect 12145 4505 12150 4545
rect 12100 3445 12150 4505
rect 12100 3405 12105 3445
rect 12145 3405 12150 3445
rect 12100 3245 12150 3405
rect 12100 3205 12105 3245
rect 12145 3205 12150 3245
rect 12100 3200 12150 3205
rect 12400 4545 12450 4550
rect 12400 4505 12405 4545
rect 12445 4505 12450 4545
rect 12400 3445 12450 4505
rect 12550 4545 12600 4550
rect 12550 4505 12555 4545
rect 12595 4505 12600 4545
rect 12550 4500 12600 4505
rect 12700 4545 12750 4550
rect 12700 4505 12705 4545
rect 12745 4505 12750 4545
rect 12400 3405 12405 3445
rect 12445 3405 12450 3445
rect 12400 3245 12450 3405
rect 12400 3205 12405 3245
rect 12445 3205 12450 3245
rect 12400 3200 12450 3205
rect 12550 4145 12600 4150
rect 12550 4105 12555 4145
rect 12595 4105 12600 4145
rect 12550 3245 12600 4105
rect 12550 3205 12555 3245
rect 12595 3205 12600 3245
rect 8200 3005 8205 3045
rect 8245 3005 8250 3045
rect 8200 3000 8250 3005
rect 7600 2905 7605 2945
rect 7645 2905 7650 2945
rect 7600 2900 7650 2905
rect 9550 2945 9600 2950
rect 9550 2905 9555 2945
rect 9595 2905 9600 2945
rect 6400 2805 6405 2845
rect 6445 2805 6450 2845
rect 6400 2800 6450 2805
rect -200 2705 -195 2745
rect -155 2705 -150 2745
rect -200 2700 -150 2705
rect -500 1345 -450 1350
rect -500 1305 -495 1345
rect -455 1305 -450 1345
rect -500 845 -450 1305
rect -200 1345 -150 1350
rect -200 1305 -195 1345
rect -155 1305 -150 1345
rect -500 805 -495 845
rect -455 805 -450 845
rect -500 -855 -450 805
rect -500 -895 -495 -855
rect -455 -895 -450 -855
rect -500 -900 -450 -895
rect -350 1045 -300 1050
rect -350 1005 -345 1045
rect -305 1005 -300 1045
rect -350 845 -300 1005
rect -350 805 -345 845
rect -305 805 -300 845
rect -350 -855 -300 805
rect -350 -895 -345 -855
rect -305 -895 -300 -855
rect -350 -950 -300 -895
rect -200 845 -150 1305
rect 3700 1245 3750 1250
rect 3700 1205 3705 1245
rect 3745 1205 3750 1245
rect 1300 1145 1350 1150
rect 1300 1105 1305 1145
rect 1345 1105 1350 1145
rect -200 805 -195 845
rect -155 805 -150 845
rect -200 -855 -150 805
rect -200 -895 -195 -855
rect -155 -895 -150 -855
rect -200 -900 -150 -895
rect 100 1045 150 1050
rect 100 1005 105 1045
rect 145 1005 150 1045
rect 100 845 150 1005
rect 100 805 105 845
rect 145 805 150 845
rect 100 -855 150 805
rect 100 -895 105 -855
rect 145 -895 150 -855
rect 100 -900 150 -895
rect 400 1045 450 1050
rect 400 1005 405 1045
rect 445 1005 450 1045
rect 400 845 450 1005
rect 400 805 405 845
rect 445 805 450 845
rect 400 -855 450 805
rect 400 -895 405 -855
rect 445 -895 450 -855
rect 400 -900 450 -895
rect 700 1045 750 1050
rect 700 1005 705 1045
rect 745 1005 750 1045
rect 700 845 750 1005
rect 700 805 705 845
rect 745 805 750 845
rect 700 -855 750 805
rect 700 -895 705 -855
rect 745 -895 750 -855
rect 700 -900 750 -895
rect 1000 1045 1050 1050
rect 1000 1005 1005 1045
rect 1045 1005 1050 1045
rect 1000 845 1050 1005
rect 1000 805 1005 845
rect 1045 805 1050 845
rect 1000 -855 1050 805
rect 1000 -895 1005 -855
rect 1045 -895 1050 -855
rect 1000 -900 1050 -895
rect 1300 845 1350 1105
rect 1300 805 1305 845
rect 1345 805 1350 845
rect 1300 -855 1350 805
rect 1300 -895 1305 -855
rect 1345 -895 1350 -855
rect 1300 -900 1350 -895
rect 1600 1145 1650 1150
rect 1600 1105 1605 1145
rect 1645 1105 1650 1145
rect 1600 845 1650 1105
rect 1600 805 1605 845
rect 1645 805 1650 845
rect 1600 -855 1650 805
rect 1600 -895 1605 -855
rect 1645 -895 1650 -855
rect 1600 -900 1650 -895
rect 1900 1145 1950 1150
rect 1900 1105 1905 1145
rect 1945 1105 1950 1145
rect 1900 845 1950 1105
rect 1900 805 1905 845
rect 1945 805 1950 845
rect 1900 -855 1950 805
rect 1900 -895 1905 -855
rect 1945 -895 1950 -855
rect 1900 -900 1950 -895
rect 2200 1145 2250 1150
rect 2200 1105 2205 1145
rect 2245 1105 2250 1145
rect 2200 845 2250 1105
rect 2200 805 2205 845
rect 2245 805 2250 845
rect 2200 -855 2250 805
rect 2200 -895 2205 -855
rect 2245 -895 2250 -855
rect 2200 -900 2250 -895
rect 2350 1145 2400 1150
rect 2350 1105 2355 1145
rect 2395 1105 2400 1145
rect 2350 845 2400 1105
rect 2350 805 2355 845
rect 2395 805 2400 845
rect 2350 -855 2400 805
rect 2350 -895 2355 -855
rect 2395 -895 2400 -855
rect 2350 -900 2400 -895
rect 2500 1145 2550 1150
rect 2500 1105 2505 1145
rect 2545 1105 2550 1145
rect 2500 845 2550 1105
rect 2500 805 2505 845
rect 2545 805 2550 845
rect 2500 -855 2550 805
rect 2500 -895 2505 -855
rect 2545 -895 2550 -855
rect 2500 -900 2550 -895
rect 2800 1145 2850 1150
rect 2800 1105 2805 1145
rect 2845 1105 2850 1145
rect 2800 845 2850 1105
rect 2800 805 2805 845
rect 2845 805 2850 845
rect 2800 -855 2850 805
rect 2800 -895 2805 -855
rect 2845 -895 2850 -855
rect 2800 -900 2850 -895
rect 3100 1145 3150 1150
rect 3100 1105 3105 1145
rect 3145 1105 3150 1145
rect 3100 845 3150 1105
rect 3100 805 3105 845
rect 3145 805 3150 845
rect 3100 -855 3150 805
rect 3100 -895 3105 -855
rect 3145 -895 3150 -855
rect 3100 -900 3150 -895
rect 3400 1145 3450 1150
rect 3400 1105 3405 1145
rect 3445 1105 3450 1145
rect 3400 845 3450 1105
rect 3400 805 3405 845
rect 3445 805 3450 845
rect 3400 -855 3450 805
rect 3400 -895 3405 -855
rect 3445 -895 3450 -855
rect 3400 -900 3450 -895
rect 3700 845 3750 1205
rect 4000 1245 4050 1250
rect 4000 1205 4005 1245
rect 4045 1205 4050 1245
rect 3700 805 3705 845
rect 3745 805 3750 845
rect 3700 -855 3750 805
rect 3700 -895 3705 -855
rect 3745 -895 3750 -855
rect 3700 -900 3750 -895
rect 3850 1045 3900 1050
rect 3850 1005 3855 1045
rect 3895 1005 3900 1045
rect 3850 845 3900 1005
rect 3850 805 3855 845
rect 3895 805 3900 845
rect 3850 -855 3900 805
rect 3850 -895 3855 -855
rect 3895 -895 3900 -855
rect 3850 -900 3900 -895
rect 4000 845 4050 1205
rect 4000 805 4005 845
rect 4045 805 4050 845
rect 4000 -855 4050 805
rect 4000 -895 4005 -855
rect 4045 -895 4050 -855
rect 4000 -900 4050 -895
rect 4300 1245 4350 1250
rect 4300 1205 4305 1245
rect 4345 1205 4350 1245
rect 4300 845 4350 1205
rect 4600 1245 4650 1250
rect 4600 1205 4605 1245
rect 4645 1205 4650 1245
rect 4300 805 4305 845
rect 4345 805 4350 845
rect 4300 -855 4350 805
rect 4300 -895 4305 -855
rect 4345 -895 4350 -855
rect 4300 -900 4350 -895
rect 4450 1045 4500 1050
rect 4450 1005 4455 1045
rect 4495 1005 4500 1045
rect 4450 845 4500 1005
rect 4450 805 4455 845
rect 4495 805 4500 845
rect 4450 -855 4500 805
rect 4450 -895 4455 -855
rect 4495 -895 4500 -855
rect 4450 -900 4500 -895
rect 4600 845 4650 1205
rect 4600 805 4605 845
rect 4645 805 4650 845
rect 4600 -855 4650 805
rect 4600 -895 4605 -855
rect 4645 -895 4650 -855
rect 4600 -900 4650 -895
rect 4900 1145 4950 1150
rect 4900 1105 4905 1145
rect 4945 1105 4950 1145
rect 4900 845 4950 1105
rect 4900 805 4905 845
rect 4945 805 4950 845
rect 4900 -855 4950 805
rect 4900 -895 4905 -855
rect 4945 -895 4950 -855
rect 4900 -900 4950 -895
rect 5200 1145 5250 1150
rect 5200 1105 5205 1145
rect 5245 1105 5250 1145
rect 5200 845 5250 1105
rect 5200 805 5205 845
rect 5245 805 5250 845
rect 5200 -855 5250 805
rect 5200 -895 5205 -855
rect 5245 -895 5250 -855
rect 5200 -900 5250 -895
rect 5500 1145 5550 1150
rect 5500 1105 5505 1145
rect 5545 1105 5550 1145
rect 5500 845 5550 1105
rect 5500 805 5505 845
rect 5545 805 5550 845
rect 5500 -855 5550 805
rect 5500 -895 5505 -855
rect 5545 -895 5550 -855
rect 5500 -900 5550 -895
rect 5800 1145 5850 1150
rect 5800 1105 5805 1145
rect 5845 1105 5850 1145
rect 5800 845 5850 1105
rect 5800 805 5805 845
rect 5845 805 5850 845
rect 5800 -855 5850 805
rect 5800 -895 5805 -855
rect 5845 -895 5850 -855
rect 5800 -900 5850 -895
rect 5950 1145 6000 1150
rect 5950 1105 5955 1145
rect 5995 1105 6000 1145
rect 5950 845 6000 1105
rect 5950 805 5955 845
rect 5995 805 6000 845
rect 5950 -855 6000 805
rect 5950 -895 5955 -855
rect 5995 -895 6000 -855
rect 5950 -900 6000 -895
rect 6100 1145 6150 1150
rect 6100 1105 6105 1145
rect 6145 1105 6150 1145
rect 6100 845 6150 1105
rect 6100 805 6105 845
rect 6145 805 6150 845
rect 6100 -855 6150 805
rect 6100 -895 6105 -855
rect 6145 -895 6150 -855
rect 6100 -900 6150 -895
rect 6400 1145 6450 1150
rect 6400 1105 6405 1145
rect 6445 1105 6450 1145
rect 6400 845 6450 1105
rect 6400 805 6405 845
rect 6445 805 6450 845
rect 6400 -855 6450 805
rect 6400 -895 6405 -855
rect 6445 -895 6450 -855
rect 6400 -900 6450 -895
rect 6700 1145 6750 1150
rect 6700 1105 6705 1145
rect 6745 1105 6750 1145
rect 6700 845 6750 1105
rect 6700 805 6705 845
rect 6745 805 6750 845
rect 6700 -855 6750 805
rect 6700 -895 6705 -855
rect 6745 -895 6750 -855
rect 6700 -900 6750 -895
rect 7000 1145 7050 1150
rect 7000 1105 7005 1145
rect 7045 1105 7050 1145
rect 7000 845 7050 1105
rect 7000 805 7005 845
rect 7045 805 7050 845
rect 7000 -855 7050 805
rect 7000 -895 7005 -855
rect 7045 -895 7050 -855
rect 7000 -900 7050 -895
rect 7300 1045 7350 1050
rect 7300 1005 7305 1045
rect 7345 1005 7350 1045
rect 7300 845 7350 1005
rect 7300 805 7305 845
rect 7345 805 7350 845
rect 7300 -855 7350 805
rect 7300 -895 7305 -855
rect 7345 -895 7350 -855
rect 7300 -900 7350 -895
rect 7600 1045 7650 1050
rect 7600 1005 7605 1045
rect 7645 1005 7650 1045
rect 7600 845 7650 1005
rect 7600 805 7605 845
rect 7645 805 7650 845
rect 7600 -855 7650 805
rect 7600 -895 7605 -855
rect 7645 -895 7650 -855
rect 7600 -900 7650 -895
rect 7900 1045 7950 1050
rect 7900 1005 7905 1045
rect 7945 1005 7950 1045
rect 7900 845 7950 1005
rect 7900 805 7905 845
rect 7945 805 7950 845
rect 7900 -855 7950 805
rect 7900 -895 7905 -855
rect 7945 -895 7950 -855
rect 7900 -900 7950 -895
rect 8200 1045 8250 1050
rect 8200 1005 8205 1045
rect 8245 1005 8250 1045
rect 8200 845 8250 1005
rect 8200 805 8205 845
rect 8245 805 8250 845
rect 8200 -855 8250 805
rect 8200 -895 8205 -855
rect 8245 -895 8250 -855
rect 8200 -900 8250 -895
rect 8500 1045 8550 1050
rect 8500 1005 8505 1045
rect 8545 1005 8550 1045
rect 8500 845 8550 1005
rect 8500 805 8505 845
rect 8545 805 8550 845
rect 8500 -855 8550 805
rect 8500 -895 8505 -855
rect 8545 -895 8550 -855
rect 8500 -900 8550 -895
rect 8800 1045 8850 1050
rect 8800 1005 8805 1045
rect 8845 1005 8850 1045
rect 8800 845 8850 1005
rect 8800 805 8805 845
rect 8845 805 8850 845
rect 8800 -855 8850 805
rect 8800 -895 8805 -855
rect 8845 -895 8850 -855
rect 8800 -900 8850 -895
rect 9100 1045 9150 1050
rect 9100 1005 9105 1045
rect 9145 1005 9150 1045
rect 9100 845 9150 1005
rect 9100 805 9105 845
rect 9145 805 9150 845
rect 9100 -855 9150 805
rect 9100 -895 9105 -855
rect 9145 -895 9150 -855
rect 9100 -900 9150 -895
rect 9400 1045 9450 1050
rect 9400 1005 9405 1045
rect 9445 1005 9450 1045
rect 9400 845 9450 1005
rect 9400 805 9405 845
rect 9445 805 9450 845
rect 9400 -855 9450 805
rect 9400 -895 9405 -855
rect 9445 -895 9450 -855
rect 9400 -900 9450 -895
rect 9550 845 9600 2905
rect 12100 2145 12150 2150
rect 12100 2105 12105 2145
rect 12145 2105 12150 2145
rect 9550 805 9555 845
rect 9595 805 9600 845
rect 9550 -855 9600 805
rect 9550 -895 9555 -855
rect 9595 -895 9600 -855
rect 9550 -900 9600 -895
rect 9700 1045 9750 1050
rect 9700 1005 9705 1045
rect 9745 1005 9750 1045
rect 9700 845 9750 1005
rect 9700 805 9705 845
rect 9745 805 9750 845
rect 9700 -855 9750 805
rect 9700 -895 9705 -855
rect 9745 -895 9750 -855
rect 9700 -900 9750 -895
rect 10000 1045 10050 1050
rect 10000 1005 10005 1045
rect 10045 1005 10050 1045
rect 10000 845 10050 1005
rect 10000 805 10005 845
rect 10045 805 10050 845
rect 10000 -855 10050 805
rect 10000 -895 10005 -855
rect 10045 -895 10050 -855
rect 10000 -900 10050 -895
rect 10300 1045 10350 1050
rect 10300 1005 10305 1045
rect 10345 1005 10350 1045
rect 10300 845 10350 1005
rect 10300 805 10305 845
rect 10345 805 10350 845
rect 10300 -855 10350 805
rect 10300 -895 10305 -855
rect 10345 -895 10350 -855
rect 10300 -900 10350 -895
rect 10600 1045 10650 1050
rect 10600 1005 10605 1045
rect 10645 1005 10650 1045
rect 10600 845 10650 1005
rect 10600 805 10605 845
rect 10645 805 10650 845
rect 10600 -855 10650 805
rect 10600 -895 10605 -855
rect 10645 -895 10650 -855
rect 10600 -900 10650 -895
rect 10900 1045 10950 1050
rect 10900 1005 10905 1045
rect 10945 1005 10950 1045
rect 10900 845 10950 1005
rect 10900 805 10905 845
rect 10945 805 10950 845
rect 10900 -855 10950 805
rect 10900 -895 10905 -855
rect 10945 -895 10950 -855
rect 10900 -900 10950 -895
rect 11200 1045 11250 1050
rect 11200 1005 11205 1045
rect 11245 1005 11250 1045
rect 11200 845 11250 1005
rect 11200 805 11205 845
rect 11245 805 11250 845
rect 11200 -855 11250 805
rect 11200 -895 11205 -855
rect 11245 -895 11250 -855
rect 11200 -900 11250 -895
rect 11500 1045 11550 1050
rect 11500 1005 11505 1045
rect 11545 1005 11550 1045
rect 11500 845 11550 1005
rect 11500 805 11505 845
rect 11545 805 11550 845
rect 11500 -855 11550 805
rect 11500 -895 11505 -855
rect 11545 -895 11550 -855
rect 11500 -900 11550 -895
rect 11800 1045 11850 1050
rect 11800 1005 11805 1045
rect 11845 1005 11850 1045
rect 11800 845 11850 1005
rect 11800 805 11805 845
rect 11845 805 11850 845
rect 11800 -855 11850 805
rect 11800 -895 11805 -855
rect 11845 -895 11850 -855
rect 11800 -900 11850 -895
rect 12100 845 12150 2105
rect 12100 805 12105 845
rect 12145 805 12150 845
rect 12100 -855 12150 805
rect 12100 -895 12105 -855
rect 12145 -895 12150 -855
rect 12100 -900 12150 -895
rect 12400 2145 12450 2150
rect 12400 2105 12405 2145
rect 12445 2105 12450 2145
rect 12400 845 12450 2105
rect 12400 805 12405 845
rect 12445 805 12450 845
rect 12400 -855 12450 805
rect 12400 -895 12405 -855
rect 12445 -895 12450 -855
rect 12400 -900 12450 -895
rect 12550 845 12600 3205
rect 12700 3445 12750 4505
rect 12700 3405 12705 3445
rect 12745 3405 12750 3445
rect 12700 3245 12750 3405
rect 12700 3205 12705 3245
rect 12745 3205 12750 3245
rect 12700 3200 12750 3205
rect 13000 4545 13050 4550
rect 13000 4505 13005 4545
rect 13045 4505 13050 4545
rect 13000 3445 13050 4505
rect 13000 3405 13005 3445
rect 13045 3405 13050 3445
rect 13000 3245 13050 3405
rect 13000 3205 13005 3245
rect 13045 3205 13050 3245
rect 13000 3200 13050 3205
rect 13300 4545 13350 4550
rect 13300 4505 13305 4545
rect 13345 4505 13350 4545
rect 13300 3645 13350 4505
rect 13300 3605 13305 3645
rect 13345 3605 13350 3645
rect 13300 3245 13350 3605
rect 13300 3205 13305 3245
rect 13345 3205 13350 3245
rect 13300 3200 13350 3205
rect 13600 4545 13650 4550
rect 13600 4505 13605 4545
rect 13645 4505 13650 4545
rect 13600 3645 13650 4505
rect 13750 4545 13800 4550
rect 13750 4505 13755 4545
rect 13795 4505 13800 4545
rect 13750 4500 13800 4505
rect 13900 4545 13950 4550
rect 13900 4505 13905 4545
rect 13945 4505 13950 4545
rect 13600 3605 13605 3645
rect 13645 3605 13650 3645
rect 13600 3245 13650 3605
rect 13600 3205 13605 3245
rect 13645 3205 13650 3245
rect 13600 3200 13650 3205
rect 13750 4345 13800 4350
rect 13750 4305 13755 4345
rect 13795 4305 13800 4345
rect 13750 3245 13800 4305
rect 13750 3205 13755 3245
rect 13795 3205 13800 3245
rect 13300 2345 13350 2350
rect 13300 2305 13305 2345
rect 13345 2305 13350 2345
rect 12550 805 12555 845
rect 12595 805 12600 845
rect 12550 -855 12600 805
rect 12550 -895 12555 -855
rect 12595 -895 12600 -855
rect 12550 -900 12600 -895
rect 12700 2145 12750 2150
rect 12700 2105 12705 2145
rect 12745 2105 12750 2145
rect 12700 845 12750 2105
rect 12700 805 12705 845
rect 12745 805 12750 845
rect 12700 -855 12750 805
rect 12700 -895 12705 -855
rect 12745 -895 12750 -855
rect 12700 -900 12750 -895
rect 13000 2145 13050 2150
rect 13000 2105 13005 2145
rect 13045 2105 13050 2145
rect 13000 845 13050 2105
rect 13000 805 13005 845
rect 13045 805 13050 845
rect 13000 -855 13050 805
rect 13000 -895 13005 -855
rect 13045 -895 13050 -855
rect 13000 -900 13050 -895
rect 13300 845 13350 2305
rect 13300 805 13305 845
rect 13345 805 13350 845
rect 13300 -855 13350 805
rect 13300 -895 13305 -855
rect 13345 -895 13350 -855
rect 13300 -900 13350 -895
rect 13600 2345 13650 2350
rect 13600 2305 13605 2345
rect 13645 2305 13650 2345
rect 13600 845 13650 2305
rect 13600 805 13605 845
rect 13645 805 13650 845
rect 13600 -855 13650 805
rect 13600 -895 13605 -855
rect 13645 -895 13650 -855
rect 13600 -900 13650 -895
rect 13750 845 13800 3205
rect 13900 3645 13950 4505
rect 13900 3605 13905 3645
rect 13945 3605 13950 3645
rect 13900 3245 13950 3605
rect 13900 3205 13905 3245
rect 13945 3205 13950 3245
rect 13900 3200 13950 3205
rect 14200 4545 14250 4550
rect 14200 4505 14205 4545
rect 14245 4505 14250 4545
rect 14200 3645 14250 4505
rect 14200 3605 14205 3645
rect 14245 3605 14250 3645
rect 14200 3245 14250 3605
rect 14200 3205 14205 3245
rect 14245 3205 14250 3245
rect 14200 3200 14250 3205
rect 14500 4545 14550 4550
rect 14500 4505 14505 4545
rect 14545 4505 14550 4545
rect 14500 3645 14550 4505
rect 14500 3605 14505 3645
rect 14545 3605 14550 3645
rect 14500 3245 14550 3605
rect 14500 3205 14505 3245
rect 14545 3205 14550 3245
rect 14500 3200 14550 3205
rect 14800 4545 14850 4550
rect 14800 4505 14805 4545
rect 14845 4505 14850 4545
rect 14800 3645 14850 4505
rect 14800 3605 14805 3645
rect 14845 3605 14850 3645
rect 14800 3245 14850 3605
rect 14800 3205 14805 3245
rect 14845 3205 14850 3245
rect 14800 3200 14850 3205
rect 14950 4545 15000 4550
rect 14950 4505 14955 4545
rect 14995 4505 15000 4545
rect 14950 4345 15000 4505
rect 14950 4305 14955 4345
rect 14995 4305 15000 4345
rect 14950 3245 15000 4305
rect 14950 3205 14955 3245
rect 14995 3205 15000 3245
rect 14950 3200 15000 3205
rect 15100 4545 15150 4550
rect 15100 4505 15105 4545
rect 15145 4505 15150 4545
rect 15100 3645 15150 4505
rect 15100 3605 15105 3645
rect 15145 3605 15150 3645
rect 15100 3245 15150 3605
rect 15100 3205 15105 3245
rect 15145 3205 15150 3245
rect 15100 3200 15150 3205
rect 15400 4545 15450 4550
rect 15400 4505 15405 4545
rect 15445 4505 15450 4545
rect 15400 3645 15450 4505
rect 15400 3605 15405 3645
rect 15445 3605 15450 3645
rect 15400 3245 15450 3605
rect 15400 3205 15405 3245
rect 15445 3205 15450 3245
rect 15400 3200 15450 3205
rect 15700 4545 15750 4550
rect 15700 4505 15705 4545
rect 15745 4505 15750 4545
rect 15700 3245 15750 4505
rect 15700 3205 15705 3245
rect 15745 3205 15750 3245
rect 15700 3200 15750 3205
rect 16000 4545 16050 4550
rect 16000 4505 16005 4545
rect 16045 4505 16050 4545
rect 16000 3245 16050 4505
rect 16000 3205 16005 3245
rect 16045 3205 16050 3245
rect 16000 3200 16050 3205
rect 16300 4545 16350 5100
rect 16300 4505 16305 4545
rect 16345 4505 16350 4545
rect 16300 3245 16350 4505
rect 16300 3205 16305 3245
rect 16345 3205 16350 3245
rect 13750 805 13755 845
rect 13795 805 13800 845
rect 13750 -855 13800 805
rect 13750 -895 13755 -855
rect 13795 -895 13800 -855
rect 13750 -900 13800 -895
rect 13900 2345 13950 2350
rect 13900 2305 13905 2345
rect 13945 2305 13950 2345
rect 13900 845 13950 2305
rect 13900 805 13905 845
rect 13945 805 13950 845
rect 13900 -855 13950 805
rect 13900 -895 13905 -855
rect 13945 -895 13950 -855
rect 13900 -900 13950 -895
rect 14200 2345 14250 2350
rect 14200 2305 14205 2345
rect 14245 2305 14250 2345
rect 14200 845 14250 2305
rect 16300 2145 16350 3205
rect 16300 2105 16305 2145
rect 16345 2105 16350 2145
rect 16300 2100 16350 2105
rect 16600 4545 16650 5100
rect 16600 4505 16605 4545
rect 16645 4505 16650 4545
rect 16600 3245 16650 4505
rect 16600 3205 16605 3245
rect 16645 3205 16650 3245
rect 16600 2145 16650 3205
rect 16600 2105 16605 2145
rect 16645 2105 16650 2145
rect 16600 2100 16650 2105
rect 16750 4545 16800 4550
rect 16750 4505 16755 4545
rect 16795 4505 16800 4545
rect 16750 3245 16800 4505
rect 16750 3205 16755 3245
rect 16795 3205 16800 3245
rect 14200 805 14205 845
rect 14245 805 14250 845
rect 14200 -855 14250 805
rect 14200 -895 14205 -855
rect 14245 -895 14250 -855
rect 14200 -900 14250 -895
rect 14500 1045 14550 1050
rect 14500 1005 14505 1045
rect 14545 1005 14550 1045
rect 14500 845 14550 1005
rect 14500 805 14505 845
rect 14545 805 14550 845
rect 14500 -855 14550 805
rect 14500 -895 14505 -855
rect 14545 -895 14550 -855
rect 14500 -900 14550 -895
rect 14800 1045 14850 1050
rect 14800 1005 14805 1045
rect 14845 1005 14850 1045
rect 14800 845 14850 1005
rect 14800 805 14805 845
rect 14845 805 14850 845
rect 14800 -855 14850 805
rect 14800 -895 14805 -855
rect 14845 -895 14850 -855
rect 14800 -900 14850 -895
rect 15100 1045 15150 1050
rect 15100 1005 15105 1045
rect 15145 1005 15150 1045
rect 15100 845 15150 1005
rect 15100 805 15105 845
rect 15145 805 15150 845
rect 15100 -855 15150 805
rect 15100 -895 15105 -855
rect 15145 -895 15150 -855
rect 15100 -900 15150 -895
rect 15400 1045 15450 1050
rect 15400 1005 15405 1045
rect 15445 1005 15450 1045
rect 15400 845 15450 1005
rect 15400 805 15405 845
rect 15445 805 15450 845
rect 15400 -855 15450 805
rect 15400 -895 15405 -855
rect 15445 -895 15450 -855
rect 15400 -900 15450 -895
rect 15700 845 15750 850
rect 15700 805 15705 845
rect 15745 805 15750 845
rect 15700 645 15750 805
rect 15700 605 15705 645
rect 15745 605 15750 645
rect 15700 -855 15750 605
rect 15700 -895 15705 -855
rect 15745 -895 15750 -855
rect 15700 -900 15750 -895
rect 16000 845 16050 850
rect 16000 805 16005 845
rect 16045 805 16050 845
rect 16000 645 16050 805
rect 16000 605 16005 645
rect 16045 605 16050 645
rect 16000 -855 16050 605
rect 16000 -895 16005 -855
rect 16045 -895 16050 -855
rect 16000 -900 16050 -895
rect 16300 845 16350 850
rect 16300 805 16305 845
rect 16345 805 16350 845
rect 16300 645 16350 805
rect 16300 605 16305 645
rect 16345 605 16350 645
rect 16300 -855 16350 605
rect 16300 -895 16305 -855
rect 16345 -895 16350 -855
rect 16300 -900 16350 -895
rect 16600 845 16650 850
rect 16600 805 16605 845
rect 16645 805 16650 845
rect 16600 645 16650 805
rect 16600 605 16605 645
rect 16645 605 16650 645
rect 16600 -855 16650 605
rect 16600 -895 16605 -855
rect 16645 -895 16650 -855
rect 16600 -900 16650 -895
rect 16750 845 16800 3205
rect 16900 4545 16950 5100
rect 16900 4505 16905 4545
rect 16945 4505 16950 4545
rect 16900 3245 16950 4505
rect 16900 3205 16905 3245
rect 16945 3205 16950 3245
rect 16900 2145 16950 3205
rect 16900 2105 16905 2145
rect 16945 2105 16950 2145
rect 16900 2100 16950 2105
rect 17200 4545 17250 5100
rect 17200 4505 17205 4545
rect 17245 4505 17250 4545
rect 17200 3245 17250 4505
rect 17200 3205 17205 3245
rect 17245 3205 17250 3245
rect 17200 2145 17250 3205
rect 17500 4545 17550 4550
rect 17500 4505 17505 4545
rect 17545 4505 17550 4545
rect 17500 3245 17550 4505
rect 17500 3205 17505 3245
rect 17545 3205 17550 3245
rect 17500 3200 17550 3205
rect 17800 4545 17850 4550
rect 17800 4505 17805 4545
rect 17845 4505 17850 4545
rect 17800 3245 17850 4505
rect 17800 3205 17805 3245
rect 17845 3205 17850 3245
rect 17800 3200 17850 3205
rect 18100 4545 18150 4550
rect 18100 4505 18105 4545
rect 18145 4505 18150 4545
rect 18100 3245 18150 4505
rect 18100 3205 18105 3245
rect 18145 3205 18150 3245
rect 18100 3200 18150 3205
rect 18400 4545 18450 4550
rect 18400 4505 18405 4545
rect 18445 4505 18450 4545
rect 18400 3245 18450 4505
rect 18400 3205 18405 3245
rect 18445 3205 18450 3245
rect 18400 3200 18450 3205
rect 18700 4545 18750 5100
rect 18700 4505 18705 4545
rect 18745 4505 18750 4545
rect 18700 3245 18750 4505
rect 18700 3205 18705 3245
rect 18745 3205 18750 3245
rect 18700 2345 18750 3205
rect 18700 2305 18705 2345
rect 18745 2305 18750 2345
rect 18700 2300 18750 2305
rect 19000 4545 19050 5100
rect 19000 4505 19005 4545
rect 19045 4505 19050 4545
rect 19000 3245 19050 4505
rect 19000 3205 19005 3245
rect 19045 3205 19050 3245
rect 19000 2345 19050 3205
rect 19000 2305 19005 2345
rect 19045 2305 19050 2345
rect 19000 2300 19050 2305
rect 19150 4545 19200 4550
rect 19150 4505 19155 4545
rect 19195 4505 19200 4545
rect 19150 3245 19200 4505
rect 19150 3205 19155 3245
rect 19195 3205 19200 3245
rect 17200 2105 17205 2145
rect 17245 2105 17250 2145
rect 17200 2100 17250 2105
rect 16750 805 16755 845
rect 16795 805 16800 845
rect 16750 -855 16800 805
rect 16750 -895 16755 -855
rect 16795 -895 16800 -855
rect 16750 -900 16800 -895
rect 16900 845 16950 850
rect 16900 805 16905 845
rect 16945 805 16950 845
rect 16900 645 16950 805
rect 16900 605 16905 645
rect 16945 605 16950 645
rect 16900 -855 16950 605
rect 16900 -895 16905 -855
rect 16945 -895 16950 -855
rect 16900 -900 16950 -895
rect 17200 845 17250 850
rect 17200 805 17205 845
rect 17245 805 17250 845
rect 17200 645 17250 805
rect 17200 605 17205 645
rect 17245 605 17250 645
rect 17200 -855 17250 605
rect 17200 -895 17205 -855
rect 17245 -895 17250 -855
rect 17200 -900 17250 -895
rect 17500 845 17550 850
rect 17500 805 17505 845
rect 17545 805 17550 845
rect 17500 645 17550 805
rect 17500 605 17505 645
rect 17545 605 17550 645
rect 17500 -855 17550 605
rect 17500 -895 17505 -855
rect 17545 -895 17550 -855
rect 17500 -900 17550 -895
rect 17800 845 17850 850
rect 17800 805 17805 845
rect 17845 805 17850 845
rect 17800 645 17850 805
rect 17800 605 17805 645
rect 17845 605 17850 645
rect 17800 -855 17850 605
rect 17800 -895 17805 -855
rect 17845 -895 17850 -855
rect 17800 -900 17850 -895
rect 18100 845 18150 850
rect 18100 805 18105 845
rect 18145 805 18150 845
rect 18100 445 18150 805
rect 18100 405 18105 445
rect 18145 405 18150 445
rect 18100 -855 18150 405
rect 18100 -895 18105 -855
rect 18145 -895 18150 -855
rect 18100 -900 18150 -895
rect 18400 845 18450 850
rect 18400 805 18405 845
rect 18445 805 18450 845
rect 18400 445 18450 805
rect 18400 405 18405 445
rect 18445 405 18450 445
rect 18400 -855 18450 405
rect 18400 -895 18405 -855
rect 18445 -895 18450 -855
rect 18400 -900 18450 -895
rect 18700 845 18750 850
rect 18700 805 18705 845
rect 18745 805 18750 845
rect 18700 445 18750 805
rect 18700 405 18705 445
rect 18745 405 18750 445
rect 18700 -855 18750 405
rect 18700 -895 18705 -855
rect 18745 -895 18750 -855
rect 18700 -900 18750 -895
rect 19000 845 19050 850
rect 19000 805 19005 845
rect 19045 805 19050 845
rect 19000 445 19050 805
rect 19000 405 19005 445
rect 19045 405 19050 445
rect 19000 -855 19050 405
rect 19000 -895 19005 -855
rect 19045 -895 19050 -855
rect 19000 -900 19050 -895
rect 19150 845 19200 3205
rect 19300 4545 19350 5100
rect 19300 4505 19305 4545
rect 19345 4505 19350 4545
rect 19300 3245 19350 4505
rect 19300 3205 19305 3245
rect 19345 3205 19350 3245
rect 19300 2345 19350 3205
rect 19300 2305 19305 2345
rect 19345 2305 19350 2345
rect 19300 2300 19350 2305
rect 19600 4545 19650 5100
rect 19600 4505 19605 4545
rect 19645 4505 19650 4545
rect 19600 3245 19650 4505
rect 19600 3205 19605 3245
rect 19645 3205 19650 3245
rect 19600 2345 19650 3205
rect 19900 4545 19950 4550
rect 19900 4505 19905 4545
rect 19945 4505 19950 4545
rect 19900 3245 19950 4505
rect 19900 3205 19905 3245
rect 19945 3205 19950 3245
rect 19900 3200 19950 3205
rect 20200 4545 20250 4550
rect 20200 4505 20205 4545
rect 20245 4505 20250 4545
rect 20200 3245 20250 4505
rect 20200 3205 20205 3245
rect 20245 3205 20250 3245
rect 20200 3200 20250 3205
rect 19600 2305 19605 2345
rect 19645 2305 19650 2345
rect 19600 2300 19650 2305
rect 19150 805 19155 845
rect 19195 805 19200 845
rect 19150 -855 19200 805
rect 19150 -895 19155 -855
rect 19195 -895 19200 -855
rect 19150 -900 19200 -895
rect 19300 845 19350 850
rect 19300 805 19305 845
rect 19345 805 19350 845
rect 19300 445 19350 805
rect 19300 405 19305 445
rect 19345 405 19350 445
rect 19300 -855 19350 405
rect 19300 -895 19305 -855
rect 19345 -895 19350 -855
rect 19300 -900 19350 -895
rect 19600 845 19650 850
rect 19600 805 19605 845
rect 19645 805 19650 845
rect 19600 445 19650 805
rect 19600 405 19605 445
rect 19645 405 19650 445
rect 19600 -855 19650 405
rect 19600 -895 19605 -855
rect 19645 -895 19650 -855
rect 19600 -900 19650 -895
rect 19900 845 19950 850
rect 19900 805 19905 845
rect 19945 805 19950 845
rect 19900 445 19950 805
rect 19900 405 19905 445
rect 19945 405 19950 445
rect 19900 -855 19950 405
rect 19900 -895 19905 -855
rect 19945 -895 19950 -855
rect 19900 -900 19950 -895
rect 20200 845 20250 850
rect 20200 805 20205 845
rect 20245 805 20250 845
rect 20200 445 20250 805
rect 20200 405 20205 445
rect 20245 405 20250 445
rect 20200 -855 20250 405
rect 20200 -895 20205 -855
rect 20245 -895 20250 -855
rect 20200 -900 20250 -895
<< end >>
