magic
tech sky130A
timestamp 1713037678
<< locali >>
rect 0 0 50 50
<< metal1 >>
rect 39800 11340 39850 11350
rect 39800 11310 39810 11340
rect 39840 11310 39850 11340
rect 39800 11300 39850 11310
rect 39900 11240 40900 11250
rect 39900 11210 39910 11240
rect 39940 11210 39960 11240
rect 39990 11210 40010 11240
rect 40040 11210 40060 11240
rect 40090 11210 40110 11240
rect 40140 11210 40160 11240
rect 40190 11210 40210 11240
rect 40240 11210 40260 11240
rect 40290 11210 40310 11240
rect 40340 11210 40360 11240
rect 40390 11210 40410 11240
rect 40440 11210 40460 11240
rect 40490 11210 40510 11240
rect 40540 11210 40560 11240
rect 40590 11210 40610 11240
rect 40640 11210 40660 11240
rect 40690 11210 40710 11240
rect 40740 11210 40760 11240
rect 40790 11210 40810 11240
rect 40840 11210 40860 11240
rect 40890 11210 40900 11240
rect 39900 11190 40900 11210
rect 39900 11160 39910 11190
rect 39940 11160 39960 11190
rect 39990 11160 40010 11190
rect 40040 11160 40060 11190
rect 40090 11160 40110 11190
rect 40140 11160 40160 11190
rect 40190 11160 40210 11190
rect 40240 11160 40260 11190
rect 40290 11160 40310 11190
rect 40340 11160 40360 11190
rect 40390 11160 40410 11190
rect 40440 11160 40460 11190
rect 40490 11160 40510 11190
rect 40540 11160 40560 11190
rect 40590 11160 40610 11190
rect 40640 11160 40660 11190
rect 40690 11160 40710 11190
rect 40740 11160 40760 11190
rect 40790 11160 40810 11190
rect 40840 11160 40860 11190
rect 40890 11160 40900 11190
rect 39900 11140 40900 11160
rect 39900 11110 39910 11140
rect 39940 11110 39960 11140
rect 39990 11110 40010 11140
rect 40040 11110 40060 11140
rect 40090 11110 40110 11140
rect 40140 11110 40160 11140
rect 40190 11110 40210 11140
rect 40240 11110 40260 11140
rect 40290 11110 40310 11140
rect 40340 11110 40360 11140
rect 40390 11110 40410 11140
rect 40440 11110 40460 11140
rect 40490 11110 40510 11140
rect 40540 11110 40560 11140
rect 40590 11110 40610 11140
rect 40640 11110 40660 11140
rect 40690 11110 40710 11140
rect 40740 11110 40760 11140
rect 40790 11110 40810 11140
rect 40840 11110 40860 11140
rect 40890 11110 40900 11140
rect 39900 11090 40900 11110
rect 39900 11060 39910 11090
rect 39940 11060 39960 11090
rect 39990 11060 40010 11090
rect 40040 11060 40060 11090
rect 40090 11060 40110 11090
rect 40140 11060 40160 11090
rect 40190 11060 40210 11090
rect 40240 11060 40260 11090
rect 40290 11060 40310 11090
rect 40340 11060 40360 11090
rect 40390 11060 40410 11090
rect 40440 11060 40460 11090
rect 40490 11060 40510 11090
rect 40540 11060 40560 11090
rect 40590 11060 40610 11090
rect 40640 11060 40660 11090
rect 40690 11060 40710 11090
rect 40740 11060 40760 11090
rect 40790 11060 40810 11090
rect 40840 11060 40860 11090
rect 40890 11060 40900 11090
rect 39900 11040 40900 11060
rect 39900 11010 39910 11040
rect 39940 11010 39960 11040
rect 39990 11010 40010 11040
rect 40040 11010 40060 11040
rect 40090 11010 40110 11040
rect 40140 11010 40160 11040
rect 40190 11010 40210 11040
rect 40240 11010 40260 11040
rect 40290 11010 40310 11040
rect 40340 11010 40360 11040
rect 40390 11010 40410 11040
rect 40440 11010 40460 11040
rect 40490 11010 40510 11040
rect 40540 11010 40560 11040
rect 40590 11010 40610 11040
rect 40640 11010 40660 11040
rect 40690 11010 40710 11040
rect 40740 11010 40760 11040
rect 40790 11010 40810 11040
rect 40840 11010 40860 11040
rect 40890 11010 40900 11040
rect 39900 11000 40900 11010
rect 39800 10940 39850 10950
rect 39800 10910 39810 10940
rect 39840 10910 39850 10940
rect 39800 10900 39850 10910
rect 39800 4740 39850 4750
rect 39800 4710 39810 4740
rect 39840 4710 39850 4740
rect 39800 4700 39850 4710
rect 39900 4640 40900 4650
rect 39900 4610 39910 4640
rect 39940 4610 39960 4640
rect 39990 4610 40010 4640
rect 40040 4610 40060 4640
rect 40090 4610 40110 4640
rect 40140 4610 40160 4640
rect 40190 4610 40210 4640
rect 40240 4610 40260 4640
rect 40290 4610 40310 4640
rect 40340 4610 40360 4640
rect 40390 4610 40410 4640
rect 40440 4610 40460 4640
rect 40490 4610 40510 4640
rect 40540 4610 40560 4640
rect 40590 4610 40610 4640
rect 40640 4610 40660 4640
rect 40690 4610 40710 4640
rect 40740 4610 40760 4640
rect 40790 4610 40810 4640
rect 40840 4610 40860 4640
rect 40890 4610 40900 4640
rect 39900 4590 40900 4610
rect 39900 4560 39910 4590
rect 39940 4560 39960 4590
rect 39990 4560 40010 4590
rect 40040 4560 40060 4590
rect 40090 4560 40110 4590
rect 40140 4560 40160 4590
rect 40190 4560 40210 4590
rect 40240 4560 40260 4590
rect 40290 4560 40310 4590
rect 40340 4560 40360 4590
rect 40390 4560 40410 4590
rect 40440 4560 40460 4590
rect 40490 4560 40510 4590
rect 40540 4560 40560 4590
rect 40590 4560 40610 4590
rect 40640 4560 40660 4590
rect 40690 4560 40710 4590
rect 40740 4560 40760 4590
rect 40790 4560 40810 4590
rect 40840 4560 40860 4590
rect 40890 4560 40900 4590
rect 39900 4540 40900 4560
rect 39900 4510 39910 4540
rect 39940 4510 39960 4540
rect 39990 4510 40010 4540
rect 40040 4510 40060 4540
rect 40090 4510 40110 4540
rect 40140 4510 40160 4540
rect 40190 4510 40210 4540
rect 40240 4510 40260 4540
rect 40290 4510 40310 4540
rect 40340 4510 40360 4540
rect 40390 4510 40410 4540
rect 40440 4510 40460 4540
rect 40490 4510 40510 4540
rect 40540 4510 40560 4540
rect 40590 4510 40610 4540
rect 40640 4510 40660 4540
rect 40690 4510 40710 4540
rect 40740 4510 40760 4540
rect 40790 4510 40810 4540
rect 40840 4510 40860 4540
rect 40890 4510 40900 4540
rect 39900 4490 40900 4510
rect 39900 4460 39910 4490
rect 39940 4460 39960 4490
rect 39990 4460 40010 4490
rect 40040 4460 40060 4490
rect 40090 4460 40110 4490
rect 40140 4460 40160 4490
rect 40190 4460 40210 4490
rect 40240 4460 40260 4490
rect 40290 4460 40310 4490
rect 40340 4460 40360 4490
rect 40390 4460 40410 4490
rect 40440 4460 40460 4490
rect 40490 4460 40510 4490
rect 40540 4460 40560 4490
rect 40590 4460 40610 4490
rect 40640 4460 40660 4490
rect 40690 4460 40710 4490
rect 40740 4460 40760 4490
rect 40790 4460 40810 4490
rect 40840 4460 40860 4490
rect 40890 4460 40900 4490
rect 39900 4440 40900 4460
rect 39900 4410 39910 4440
rect 39940 4410 39960 4440
rect 39990 4410 40010 4440
rect 40040 4410 40060 4440
rect 40090 4410 40110 4440
rect 40140 4410 40160 4440
rect 40190 4410 40210 4440
rect 40240 4410 40260 4440
rect 40290 4410 40310 4440
rect 40340 4410 40360 4440
rect 40390 4410 40410 4440
rect 40440 4410 40460 4440
rect 40490 4410 40510 4440
rect 40540 4410 40560 4440
rect 40590 4410 40610 4440
rect 40640 4410 40660 4440
rect 40690 4410 40710 4440
rect 40740 4410 40760 4440
rect 40790 4410 40810 4440
rect 40840 4410 40860 4440
rect 40890 4410 40900 4440
rect 39900 4400 40900 4410
rect 39800 4340 39850 4350
rect 39800 4310 39810 4340
rect 39840 4310 39850 4340
rect 39800 4300 39850 4310
<< via1 >>
rect 39810 11310 39840 11340
rect 39910 11210 39940 11240
rect 39960 11210 39990 11240
rect 40010 11210 40040 11240
rect 40060 11210 40090 11240
rect 40110 11210 40140 11240
rect 40160 11210 40190 11240
rect 40210 11210 40240 11240
rect 40260 11210 40290 11240
rect 40310 11210 40340 11240
rect 40360 11210 40390 11240
rect 40410 11210 40440 11240
rect 40460 11210 40490 11240
rect 40510 11210 40540 11240
rect 40560 11210 40590 11240
rect 40610 11210 40640 11240
rect 40660 11210 40690 11240
rect 40710 11210 40740 11240
rect 40760 11210 40790 11240
rect 40810 11210 40840 11240
rect 40860 11210 40890 11240
rect 39910 11160 39940 11190
rect 39960 11160 39990 11190
rect 40010 11160 40040 11190
rect 40060 11160 40090 11190
rect 40110 11160 40140 11190
rect 40160 11160 40190 11190
rect 40210 11160 40240 11190
rect 40260 11160 40290 11190
rect 40310 11160 40340 11190
rect 40360 11160 40390 11190
rect 40410 11160 40440 11190
rect 40460 11160 40490 11190
rect 40510 11160 40540 11190
rect 40560 11160 40590 11190
rect 40610 11160 40640 11190
rect 40660 11160 40690 11190
rect 40710 11160 40740 11190
rect 40760 11160 40790 11190
rect 40810 11160 40840 11190
rect 40860 11160 40890 11190
rect 39910 11110 39940 11140
rect 39960 11110 39990 11140
rect 40010 11110 40040 11140
rect 40060 11110 40090 11140
rect 40110 11110 40140 11140
rect 40160 11110 40190 11140
rect 40210 11110 40240 11140
rect 40260 11110 40290 11140
rect 40310 11110 40340 11140
rect 40360 11110 40390 11140
rect 40410 11110 40440 11140
rect 40460 11110 40490 11140
rect 40510 11110 40540 11140
rect 40560 11110 40590 11140
rect 40610 11110 40640 11140
rect 40660 11110 40690 11140
rect 40710 11110 40740 11140
rect 40760 11110 40790 11140
rect 40810 11110 40840 11140
rect 40860 11110 40890 11140
rect 39910 11060 39940 11090
rect 39960 11060 39990 11090
rect 40010 11060 40040 11090
rect 40060 11060 40090 11090
rect 40110 11060 40140 11090
rect 40160 11060 40190 11090
rect 40210 11060 40240 11090
rect 40260 11060 40290 11090
rect 40310 11060 40340 11090
rect 40360 11060 40390 11090
rect 40410 11060 40440 11090
rect 40460 11060 40490 11090
rect 40510 11060 40540 11090
rect 40560 11060 40590 11090
rect 40610 11060 40640 11090
rect 40660 11060 40690 11090
rect 40710 11060 40740 11090
rect 40760 11060 40790 11090
rect 40810 11060 40840 11090
rect 40860 11060 40890 11090
rect 39910 11010 39940 11040
rect 39960 11010 39990 11040
rect 40010 11010 40040 11040
rect 40060 11010 40090 11040
rect 40110 11010 40140 11040
rect 40160 11010 40190 11040
rect 40210 11010 40240 11040
rect 40260 11010 40290 11040
rect 40310 11010 40340 11040
rect 40360 11010 40390 11040
rect 40410 11010 40440 11040
rect 40460 11010 40490 11040
rect 40510 11010 40540 11040
rect 40560 11010 40590 11040
rect 40610 11010 40640 11040
rect 40660 11010 40690 11040
rect 40710 11010 40740 11040
rect 40760 11010 40790 11040
rect 40810 11010 40840 11040
rect 40860 11010 40890 11040
rect 39810 10910 39840 10940
rect 39810 4710 39840 4740
rect 39910 4610 39940 4640
rect 39960 4610 39990 4640
rect 40010 4610 40040 4640
rect 40060 4610 40090 4640
rect 40110 4610 40140 4640
rect 40160 4610 40190 4640
rect 40210 4610 40240 4640
rect 40260 4610 40290 4640
rect 40310 4610 40340 4640
rect 40360 4610 40390 4640
rect 40410 4610 40440 4640
rect 40460 4610 40490 4640
rect 40510 4610 40540 4640
rect 40560 4610 40590 4640
rect 40610 4610 40640 4640
rect 40660 4610 40690 4640
rect 40710 4610 40740 4640
rect 40760 4610 40790 4640
rect 40810 4610 40840 4640
rect 40860 4610 40890 4640
rect 39910 4560 39940 4590
rect 39960 4560 39990 4590
rect 40010 4560 40040 4590
rect 40060 4560 40090 4590
rect 40110 4560 40140 4590
rect 40160 4560 40190 4590
rect 40210 4560 40240 4590
rect 40260 4560 40290 4590
rect 40310 4560 40340 4590
rect 40360 4560 40390 4590
rect 40410 4560 40440 4590
rect 40460 4560 40490 4590
rect 40510 4560 40540 4590
rect 40560 4560 40590 4590
rect 40610 4560 40640 4590
rect 40660 4560 40690 4590
rect 40710 4560 40740 4590
rect 40760 4560 40790 4590
rect 40810 4560 40840 4590
rect 40860 4560 40890 4590
rect 39910 4510 39940 4540
rect 39960 4510 39990 4540
rect 40010 4510 40040 4540
rect 40060 4510 40090 4540
rect 40110 4510 40140 4540
rect 40160 4510 40190 4540
rect 40210 4510 40240 4540
rect 40260 4510 40290 4540
rect 40310 4510 40340 4540
rect 40360 4510 40390 4540
rect 40410 4510 40440 4540
rect 40460 4510 40490 4540
rect 40510 4510 40540 4540
rect 40560 4510 40590 4540
rect 40610 4510 40640 4540
rect 40660 4510 40690 4540
rect 40710 4510 40740 4540
rect 40760 4510 40790 4540
rect 40810 4510 40840 4540
rect 40860 4510 40890 4540
rect 39910 4460 39940 4490
rect 39960 4460 39990 4490
rect 40010 4460 40040 4490
rect 40060 4460 40090 4490
rect 40110 4460 40140 4490
rect 40160 4460 40190 4490
rect 40210 4460 40240 4490
rect 40260 4460 40290 4490
rect 40310 4460 40340 4490
rect 40360 4460 40390 4490
rect 40410 4460 40440 4490
rect 40460 4460 40490 4490
rect 40510 4460 40540 4490
rect 40560 4460 40590 4490
rect 40610 4460 40640 4490
rect 40660 4460 40690 4490
rect 40710 4460 40740 4490
rect 40760 4460 40790 4490
rect 40810 4460 40840 4490
rect 40860 4460 40890 4490
rect 39910 4410 39940 4440
rect 39960 4410 39990 4440
rect 40010 4410 40040 4440
rect 40060 4410 40090 4440
rect 40110 4410 40140 4440
rect 40160 4410 40190 4440
rect 40210 4410 40240 4440
rect 40260 4410 40290 4440
rect 40310 4410 40340 4440
rect 40360 4410 40390 4440
rect 40410 4410 40440 4440
rect 40460 4410 40490 4440
rect 40510 4410 40540 4440
rect 40560 4410 40590 4440
rect 40610 4410 40640 4440
rect 40660 4410 40690 4440
rect 40710 4410 40740 4440
rect 40760 4410 40790 4440
rect 40810 4410 40840 4440
rect 40860 4410 40890 4440
rect 39810 4310 39840 4340
<< metal2 >>
rect -3500 16940 -50 16950
rect -3500 16910 -3490 16940
rect -3460 16910 -3290 16940
rect -3260 16910 -3090 16940
rect -3060 16910 -1590 16940
rect -1560 16910 -1190 16940
rect -1160 16910 -1090 16940
rect -1060 16910 -990 16940
rect -960 16910 -890 16940
rect -860 16910 -790 16940
rect -760 16910 -690 16940
rect -660 16910 -590 16940
rect -560 16910 -490 16940
rect -460 16910 -390 16940
rect -360 16910 -290 16940
rect -260 16910 -190 16940
rect -160 16910 -90 16940
rect -60 16910 -50 16940
rect -3500 16900 -50 16910
rect -3500 15740 -50 15750
rect -3500 15710 -3490 15740
rect -3460 15710 -3290 15740
rect -3260 15710 -3090 15740
rect -3060 15710 -1590 15740
rect -1560 15710 -1190 15740
rect -1160 15710 -1090 15740
rect -1060 15710 -990 15740
rect -960 15710 -890 15740
rect -860 15710 -690 15740
rect -660 15710 -590 15740
rect -560 15710 -490 15740
rect -460 15710 -290 15740
rect -260 15710 -190 15740
rect -160 15710 -90 15740
rect -60 15710 -50 15740
rect -3500 15700 -50 15710
rect -3500 15340 0 15350
rect -3500 15310 -3490 15340
rect -3460 15310 -3290 15340
rect -3260 15310 -3090 15340
rect -3060 15310 -1590 15340
rect -1560 15310 -1090 15340
rect -1060 15310 -890 15340
rect -860 15310 -690 15340
rect -660 15310 -490 15340
rect -460 15310 -290 15340
rect -260 15310 -90 15340
rect -60 15310 0 15340
rect -3500 15290 0 15310
rect -3500 15260 -3490 15290
rect -3460 15260 -3290 15290
rect -3260 15260 -3090 15290
rect -3060 15260 -1590 15290
rect -1560 15260 -1090 15290
rect -1060 15260 -890 15290
rect -860 15260 -690 15290
rect -660 15260 -490 15290
rect -460 15260 -290 15290
rect -260 15260 -90 15290
rect -60 15260 0 15290
rect -3500 15240 0 15260
rect -3500 15210 -3490 15240
rect -3460 15210 -3290 15240
rect -3260 15210 -3090 15240
rect -3060 15210 -1590 15240
rect -1560 15210 -1090 15240
rect -1060 15210 -890 15240
rect -860 15210 -690 15240
rect -660 15210 -490 15240
rect -460 15210 -290 15240
rect -260 15210 -90 15240
rect -60 15210 0 15240
rect -3500 15200 0 15210
rect -3500 13640 0 13650
rect -3500 13610 -3490 13640
rect -3460 13610 -3290 13640
rect -3260 13610 -3090 13640
rect -3060 13610 -1590 13640
rect -1560 13610 -1090 13640
rect -1060 13610 -890 13640
rect -860 13610 -690 13640
rect -660 13610 -490 13640
rect -460 13610 -290 13640
rect -260 13610 -90 13640
rect -60 13610 0 13640
rect -3500 13590 0 13610
rect -3500 13560 -3490 13590
rect -3460 13560 -3290 13590
rect -3260 13560 -3090 13590
rect -3060 13560 -1590 13590
rect -1560 13560 -1090 13590
rect -1060 13560 -890 13590
rect -860 13560 -690 13590
rect -660 13560 -490 13590
rect -460 13560 -290 13590
rect -260 13560 -90 13590
rect -60 13560 0 13590
rect -3500 13540 0 13560
rect -3500 13510 -3490 13540
rect -3460 13510 -3290 13540
rect -3260 13510 -3090 13540
rect -3060 13510 -1590 13540
rect -1560 13510 -1090 13540
rect -1060 13510 -890 13540
rect -860 13510 -690 13540
rect -660 13510 -490 13540
rect -460 13510 -290 13540
rect -260 13510 -90 13540
rect -60 13510 0 13540
rect -3500 13500 0 13510
rect -3500 11940 0 11950
rect -3500 11910 -3490 11940
rect -3460 11910 -3290 11940
rect -3260 11910 -3090 11940
rect -3060 11910 -1590 11940
rect -1560 11910 -1090 11940
rect -1060 11910 -890 11940
rect -860 11910 -690 11940
rect -660 11910 -490 11940
rect -460 11910 -290 11940
rect -260 11910 -90 11940
rect -60 11910 0 11940
rect -3500 11890 0 11910
rect -3500 11860 -3490 11890
rect -3460 11860 -3290 11890
rect -3260 11860 -3090 11890
rect -3060 11860 -1590 11890
rect -1560 11860 -1090 11890
rect -1060 11860 -890 11890
rect -860 11860 -690 11890
rect -660 11860 -490 11890
rect -460 11860 -290 11890
rect -260 11860 -90 11890
rect -60 11860 0 11890
rect -3500 11840 0 11860
rect -3500 11810 -3490 11840
rect -3460 11810 -3290 11840
rect -3260 11810 -3090 11840
rect -3060 11810 -1590 11840
rect -1560 11810 -1090 11840
rect -1060 11810 -890 11840
rect -860 11810 -690 11840
rect -660 11810 -490 11840
rect -460 11810 -290 11840
rect -260 11810 -90 11840
rect -60 11810 0 11840
rect -3500 11800 0 11810
rect 39750 11340 39900 11350
rect 39750 11310 39810 11340
rect 39840 11310 39900 11340
rect 39750 11300 39900 11310
rect 39750 11240 40900 11250
rect 39750 11210 39910 11240
rect 39940 11210 39960 11240
rect 39990 11210 40010 11240
rect 40040 11210 40060 11240
rect 40090 11210 40110 11240
rect 40140 11210 40160 11240
rect 40190 11210 40210 11240
rect 40240 11210 40260 11240
rect 40290 11210 40310 11240
rect 40340 11210 40360 11240
rect 40390 11210 40410 11240
rect 40440 11210 40460 11240
rect 40490 11210 40510 11240
rect 40540 11210 40560 11240
rect 40590 11210 40610 11240
rect 40640 11210 40660 11240
rect 40690 11210 40710 11240
rect 40740 11210 40760 11240
rect 40790 11210 40810 11240
rect 40840 11210 40860 11240
rect 40890 11210 40900 11240
rect 39750 11190 40900 11210
rect 39750 11160 39910 11190
rect 39940 11160 39960 11190
rect 39990 11160 40010 11190
rect 40040 11160 40060 11190
rect 40090 11160 40110 11190
rect 40140 11160 40160 11190
rect 40190 11160 40210 11190
rect 40240 11160 40260 11190
rect 40290 11160 40310 11190
rect 40340 11160 40360 11190
rect 40390 11160 40410 11190
rect 40440 11160 40460 11190
rect 40490 11160 40510 11190
rect 40540 11160 40560 11190
rect 40590 11160 40610 11190
rect 40640 11160 40660 11190
rect 40690 11160 40710 11190
rect 40740 11160 40760 11190
rect 40790 11160 40810 11190
rect 40840 11160 40860 11190
rect 40890 11160 40900 11190
rect 39750 11140 40900 11160
rect 39750 11110 39910 11140
rect 39940 11110 39960 11140
rect 39990 11110 40010 11140
rect 40040 11110 40060 11140
rect 40090 11110 40110 11140
rect 40140 11110 40160 11140
rect 40190 11110 40210 11140
rect 40240 11110 40260 11140
rect 40290 11110 40310 11140
rect 40340 11110 40360 11140
rect 40390 11110 40410 11140
rect 40440 11110 40460 11140
rect 40490 11110 40510 11140
rect 40540 11110 40560 11140
rect 40590 11110 40610 11140
rect 40640 11110 40660 11140
rect 40690 11110 40710 11140
rect 40740 11110 40760 11140
rect 40790 11110 40810 11140
rect 40840 11110 40860 11140
rect 40890 11110 40900 11140
rect 39750 11090 40900 11110
rect 39750 11060 39910 11090
rect 39940 11060 39960 11090
rect 39990 11060 40010 11090
rect 40040 11060 40060 11090
rect 40090 11060 40110 11090
rect 40140 11060 40160 11090
rect 40190 11060 40210 11090
rect 40240 11060 40260 11090
rect 40290 11060 40310 11090
rect 40340 11060 40360 11090
rect 40390 11060 40410 11090
rect 40440 11060 40460 11090
rect 40490 11060 40510 11090
rect 40540 11060 40560 11090
rect 40590 11060 40610 11090
rect 40640 11060 40660 11090
rect 40690 11060 40710 11090
rect 40740 11060 40760 11090
rect 40790 11060 40810 11090
rect 40840 11060 40860 11090
rect 40890 11060 40900 11090
rect 39750 11040 40900 11060
rect 39750 11010 39910 11040
rect 39940 11010 39960 11040
rect 39990 11010 40010 11040
rect 40040 11010 40060 11040
rect 40090 11010 40110 11040
rect 40140 11010 40160 11040
rect 40190 11010 40210 11040
rect 40240 11010 40260 11040
rect 40290 11010 40310 11040
rect 40340 11010 40360 11040
rect 40390 11010 40410 11040
rect 40440 11010 40460 11040
rect 40490 11010 40510 11040
rect 40540 11010 40560 11040
rect 40590 11010 40610 11040
rect 40640 11010 40660 11040
rect 40690 11010 40710 11040
rect 40740 11010 40760 11040
rect 40790 11010 40810 11040
rect 40840 11010 40860 11040
rect 40890 11010 40900 11040
rect 39750 11000 40900 11010
rect 39750 10940 39900 10950
rect 39750 10910 39810 10940
rect 39840 10910 39900 10940
rect 39750 10900 39900 10910
rect -3100 10640 0 10650
rect -3100 10610 -2990 10640
rect -2960 10610 -2790 10640
rect -2760 10610 -2590 10640
rect -2560 10610 -2390 10640
rect -2360 10610 -2190 10640
rect -2160 10610 -1990 10640
rect -1960 10610 -1690 10640
rect -1660 10610 0 10640
rect -3100 10590 0 10610
rect -3100 10560 -2990 10590
rect -2960 10560 -2790 10590
rect -2760 10560 -2590 10590
rect -2560 10560 -2390 10590
rect -2360 10560 -2190 10590
rect -2160 10560 -1990 10590
rect -1960 10560 -1690 10590
rect -1660 10560 0 10590
rect -3100 10540 0 10560
rect -3100 10510 -2990 10540
rect -2960 10510 -2790 10540
rect -2760 10510 -2590 10540
rect -2560 10510 -2390 10540
rect -2360 10510 -2190 10540
rect -2160 10510 -1990 10540
rect -1960 10510 -1690 10540
rect -1660 10510 0 10540
rect -3100 10500 0 10510
rect -3100 9340 0 9350
rect -3100 9310 -2990 9340
rect -2960 9310 -2790 9340
rect -2760 9310 -2590 9340
rect -2560 9310 -2390 9340
rect -2360 9310 -2190 9340
rect -2160 9310 -1990 9340
rect -1960 9310 -1690 9340
rect -1660 9310 0 9340
rect -3100 9290 0 9310
rect -3100 9260 -2990 9290
rect -2960 9260 -2790 9290
rect -2760 9260 -2590 9290
rect -2560 9260 -2390 9290
rect -2360 9260 -2190 9290
rect -2160 9260 -1990 9290
rect -1960 9260 -1690 9290
rect -1660 9260 0 9290
rect -3100 9240 0 9260
rect -3100 9210 -2990 9240
rect -2960 9210 -2790 9240
rect -2760 9210 -2590 9240
rect -2560 9210 -2390 9240
rect -2360 9210 -2190 9240
rect -2160 9210 -1990 9240
rect -1960 9210 -1690 9240
rect -1660 9210 0 9240
rect -3100 9200 0 9210
rect -3100 8040 0 8050
rect -3100 8010 -2990 8040
rect -2960 8010 -2790 8040
rect -2760 8010 -2590 8040
rect -2560 8010 -2390 8040
rect -2360 8010 -2190 8040
rect -2160 8010 -1990 8040
rect -1960 8010 -1690 8040
rect -1660 8010 0 8040
rect -3100 7990 0 8010
rect -3100 7960 -2990 7990
rect -2960 7960 -2790 7990
rect -2760 7960 -2590 7990
rect -2560 7960 -2390 7990
rect -2360 7960 -2190 7990
rect -2160 7960 -1990 7990
rect -1960 7960 -1690 7990
rect -1660 7960 0 7990
rect -3100 7940 0 7960
rect -3100 7910 -2990 7940
rect -2960 7910 -2790 7940
rect -2760 7910 -2590 7940
rect -2560 7910 -2390 7940
rect -2360 7910 -2190 7940
rect -2160 7910 -1990 7940
rect -1960 7910 -1690 7940
rect -1660 7910 0 7940
rect -3100 7900 0 7910
rect -3100 7740 0 7750
rect -3100 7710 -2990 7740
rect -2960 7710 -2790 7740
rect -2760 7710 -2590 7740
rect -2560 7710 -2390 7740
rect -2360 7710 -2190 7740
rect -2160 7710 -1990 7740
rect -1960 7710 -1690 7740
rect -1660 7710 0 7740
rect -3100 7690 0 7710
rect -3100 7660 -2990 7690
rect -2960 7660 -2790 7690
rect -2760 7660 -2590 7690
rect -2560 7660 -2390 7690
rect -2360 7660 -2190 7690
rect -2160 7660 -1990 7690
rect -1960 7660 -1690 7690
rect -1660 7660 0 7690
rect -3100 7640 0 7660
rect -3100 7610 -2990 7640
rect -2960 7610 -2790 7640
rect -2760 7610 -2590 7640
rect -2560 7610 -2390 7640
rect -2360 7610 -2190 7640
rect -2160 7610 -1990 7640
rect -1960 7610 -1690 7640
rect -1660 7610 0 7640
rect -3100 7600 0 7610
rect -3100 6440 0 6450
rect -3100 6410 -2990 6440
rect -2960 6410 -2790 6440
rect -2760 6410 -2590 6440
rect -2560 6410 -2390 6440
rect -2360 6410 -2190 6440
rect -2160 6410 -1990 6440
rect -1960 6410 -1690 6440
rect -1660 6410 0 6440
rect -3100 6390 0 6410
rect -3100 6360 -2990 6390
rect -2960 6360 -2790 6390
rect -2760 6360 -2590 6390
rect -2560 6360 -2390 6390
rect -2360 6360 -2190 6390
rect -2160 6360 -1990 6390
rect -1960 6360 -1690 6390
rect -1660 6360 0 6390
rect -3100 6340 0 6360
rect -3100 6310 -2990 6340
rect -2960 6310 -2790 6340
rect -2760 6310 -2590 6340
rect -2560 6310 -2390 6340
rect -2360 6310 -2190 6340
rect -2160 6310 -1990 6340
rect -1960 6310 -1690 6340
rect -1660 6310 0 6340
rect -3100 6300 0 6310
rect -3100 5140 0 5150
rect -3100 5110 -2990 5140
rect -2960 5110 -2790 5140
rect -2760 5110 -2590 5140
rect -2560 5110 -2390 5140
rect -2360 5110 -2190 5140
rect -2160 5110 -1990 5140
rect -1960 5110 -1690 5140
rect -1660 5110 0 5140
rect -3100 5090 0 5110
rect -3100 5060 -2990 5090
rect -2960 5060 -2790 5090
rect -2760 5060 -2590 5090
rect -2560 5060 -2390 5090
rect -2360 5060 -2190 5090
rect -2160 5060 -1990 5090
rect -1960 5060 -1690 5090
rect -1660 5060 0 5090
rect -3100 5040 0 5060
rect -3100 5010 -2990 5040
rect -2960 5010 -2790 5040
rect -2760 5010 -2590 5040
rect -2560 5010 -2390 5040
rect -2360 5010 -2190 5040
rect -2160 5010 -1990 5040
rect -1960 5010 -1690 5040
rect -1660 5010 0 5040
rect -3100 5000 0 5010
rect 39750 4740 39900 4750
rect 39750 4710 39810 4740
rect 39840 4710 39900 4740
rect 39750 4700 39900 4710
rect 39750 4640 40900 4650
rect 39750 4610 39910 4640
rect 39940 4610 39960 4640
rect 39990 4610 40010 4640
rect 40040 4610 40060 4640
rect 40090 4610 40110 4640
rect 40140 4610 40160 4640
rect 40190 4610 40210 4640
rect 40240 4610 40260 4640
rect 40290 4610 40310 4640
rect 40340 4610 40360 4640
rect 40390 4610 40410 4640
rect 40440 4610 40460 4640
rect 40490 4610 40510 4640
rect 40540 4610 40560 4640
rect 40590 4610 40610 4640
rect 40640 4610 40660 4640
rect 40690 4610 40710 4640
rect 40740 4610 40760 4640
rect 40790 4610 40810 4640
rect 40840 4610 40860 4640
rect 40890 4610 40900 4640
rect 39750 4590 40900 4610
rect 39750 4560 39910 4590
rect 39940 4560 39960 4590
rect 39990 4560 40010 4590
rect 40040 4560 40060 4590
rect 40090 4560 40110 4590
rect 40140 4560 40160 4590
rect 40190 4560 40210 4590
rect 40240 4560 40260 4590
rect 40290 4560 40310 4590
rect 40340 4560 40360 4590
rect 40390 4560 40410 4590
rect 40440 4560 40460 4590
rect 40490 4560 40510 4590
rect 40540 4560 40560 4590
rect 40590 4560 40610 4590
rect 40640 4560 40660 4590
rect 40690 4560 40710 4590
rect 40740 4560 40760 4590
rect 40790 4560 40810 4590
rect 40840 4560 40860 4590
rect 40890 4560 40900 4590
rect 39750 4540 40900 4560
rect 39750 4510 39910 4540
rect 39940 4510 39960 4540
rect 39990 4510 40010 4540
rect 40040 4510 40060 4540
rect 40090 4510 40110 4540
rect 40140 4510 40160 4540
rect 40190 4510 40210 4540
rect 40240 4510 40260 4540
rect 40290 4510 40310 4540
rect 40340 4510 40360 4540
rect 40390 4510 40410 4540
rect 40440 4510 40460 4540
rect 40490 4510 40510 4540
rect 40540 4510 40560 4540
rect 40590 4510 40610 4540
rect 40640 4510 40660 4540
rect 40690 4510 40710 4540
rect 40740 4510 40760 4540
rect 40790 4510 40810 4540
rect 40840 4510 40860 4540
rect 40890 4510 40900 4540
rect 39750 4490 40900 4510
rect 39750 4460 39910 4490
rect 39940 4460 39960 4490
rect 39990 4460 40010 4490
rect 40040 4460 40060 4490
rect 40090 4460 40110 4490
rect 40140 4460 40160 4490
rect 40190 4460 40210 4490
rect 40240 4460 40260 4490
rect 40290 4460 40310 4490
rect 40340 4460 40360 4490
rect 40390 4460 40410 4490
rect 40440 4460 40460 4490
rect 40490 4460 40510 4490
rect 40540 4460 40560 4490
rect 40590 4460 40610 4490
rect 40640 4460 40660 4490
rect 40690 4460 40710 4490
rect 40740 4460 40760 4490
rect 40790 4460 40810 4490
rect 40840 4460 40860 4490
rect 40890 4460 40900 4490
rect 39750 4440 40900 4460
rect 39750 4410 39910 4440
rect 39940 4410 39960 4440
rect 39990 4410 40010 4440
rect 40040 4410 40060 4440
rect 40090 4410 40110 4440
rect 40140 4410 40160 4440
rect 40190 4410 40210 4440
rect 40240 4410 40260 4440
rect 40290 4410 40310 4440
rect 40340 4410 40360 4440
rect 40390 4410 40410 4440
rect 40440 4410 40460 4440
rect 40490 4410 40510 4440
rect 40540 4410 40560 4440
rect 40590 4410 40610 4440
rect 40640 4410 40660 4440
rect 40690 4410 40710 4440
rect 40740 4410 40760 4440
rect 40790 4410 40810 4440
rect 40840 4410 40860 4440
rect 40890 4410 40900 4440
rect 39750 4400 40900 4410
rect 39750 4340 39900 4350
rect 39750 4310 39810 4340
rect 39840 4310 39900 4340
rect 39750 4300 39900 4310
rect -3500 3840 0 3850
rect -3500 3810 -3490 3840
rect -3460 3810 -3290 3840
rect -3260 3810 -3090 3840
rect -3060 3810 -1590 3840
rect -1560 3810 -1090 3840
rect -1060 3810 -890 3840
rect -860 3810 -690 3840
rect -660 3810 -490 3840
rect -460 3810 -290 3840
rect -260 3810 -90 3840
rect -60 3810 0 3840
rect -3500 3790 0 3810
rect -3500 3760 -3490 3790
rect -3460 3760 -3290 3790
rect -3260 3760 -3090 3790
rect -3060 3760 -1590 3790
rect -1560 3760 -1090 3790
rect -1060 3760 -890 3790
rect -860 3760 -690 3790
rect -660 3760 -490 3790
rect -460 3760 -290 3790
rect -260 3760 -90 3790
rect -60 3760 0 3790
rect -3500 3740 0 3760
rect -3500 3710 -3490 3740
rect -3460 3710 -3290 3740
rect -3260 3710 -3090 3740
rect -3060 3710 -1590 3740
rect -1560 3710 -1090 3740
rect -1060 3710 -890 3740
rect -860 3710 -690 3740
rect -660 3710 -490 3740
rect -460 3710 -290 3740
rect -260 3710 -90 3740
rect -60 3710 0 3740
rect -3500 3700 0 3710
rect -3500 2140 0 2150
rect -3500 2110 -3490 2140
rect -3460 2110 -3290 2140
rect -3260 2110 -3090 2140
rect -3060 2110 -1590 2140
rect -1560 2110 -1090 2140
rect -1060 2110 -890 2140
rect -860 2110 -690 2140
rect -660 2110 -490 2140
rect -460 2110 -290 2140
rect -260 2110 -90 2140
rect -60 2110 0 2140
rect -3500 2090 0 2110
rect -3500 2060 -3490 2090
rect -3460 2060 -3290 2090
rect -3260 2060 -3090 2090
rect -3060 2060 -1590 2090
rect -1560 2060 -1090 2090
rect -1060 2060 -890 2090
rect -860 2060 -690 2090
rect -660 2060 -490 2090
rect -460 2060 -290 2090
rect -260 2060 -90 2090
rect -60 2060 0 2090
rect -3500 2040 0 2060
rect -3500 2010 -3490 2040
rect -3460 2010 -3290 2040
rect -3260 2010 -3090 2040
rect -3060 2010 -1590 2040
rect -1560 2010 -1090 2040
rect -1060 2010 -890 2040
rect -860 2010 -690 2040
rect -660 2010 -490 2040
rect -460 2010 -290 2040
rect -260 2010 -90 2040
rect -60 2010 0 2040
rect -3500 2000 0 2010
rect -3500 440 0 450
rect -3500 410 -3490 440
rect -3460 410 -3290 440
rect -3260 410 -3090 440
rect -3060 410 -1590 440
rect -1560 410 -1090 440
rect -1060 410 -890 440
rect -860 410 -690 440
rect -660 410 -490 440
rect -460 410 -290 440
rect -260 410 -90 440
rect -60 410 0 440
rect -3500 390 0 410
rect -3500 360 -3490 390
rect -3460 360 -3290 390
rect -3260 360 -3090 390
rect -3060 360 -1590 390
rect -1560 360 -1090 390
rect -1060 360 -890 390
rect -860 360 -690 390
rect -660 360 -490 390
rect -460 360 -290 390
rect -260 360 -90 390
rect -60 360 0 390
rect -3500 340 0 360
rect -3500 310 -3490 340
rect -3460 310 -3290 340
rect -3260 310 -3090 340
rect -3060 310 -1590 340
rect -1560 310 -1090 340
rect -1060 310 -890 340
rect -860 310 -690 340
rect -660 310 -490 340
rect -460 310 -290 340
rect -260 310 -90 340
rect -60 310 0 340
rect -3500 300 0 310
<< via2 >>
rect -3490 16910 -3460 16940
rect -3290 16910 -3260 16940
rect -3090 16910 -3060 16940
rect -1590 16910 -1560 16940
rect -1190 16910 -1160 16940
rect -1090 16910 -1060 16940
rect -990 16910 -960 16940
rect -890 16910 -860 16940
rect -790 16910 -760 16940
rect -690 16910 -660 16940
rect -590 16910 -560 16940
rect -490 16910 -460 16940
rect -390 16910 -360 16940
rect -290 16910 -260 16940
rect -190 16910 -160 16940
rect -90 16910 -60 16940
rect -3490 15710 -3460 15740
rect -3290 15710 -3260 15740
rect -3090 15710 -3060 15740
rect -1590 15710 -1560 15740
rect -1190 15710 -1160 15740
rect -1090 15710 -1060 15740
rect -990 15710 -960 15740
rect -890 15710 -860 15740
rect -690 15710 -660 15740
rect -590 15710 -560 15740
rect -490 15710 -460 15740
rect -290 15710 -260 15740
rect -190 15710 -160 15740
rect -90 15710 -60 15740
rect -3490 15310 -3460 15340
rect -3290 15310 -3260 15340
rect -3090 15310 -3060 15340
rect -1590 15310 -1560 15340
rect -1090 15310 -1060 15340
rect -890 15310 -860 15340
rect -690 15310 -660 15340
rect -490 15310 -460 15340
rect -290 15310 -260 15340
rect -90 15310 -60 15340
rect -3490 15260 -3460 15290
rect -3290 15260 -3260 15290
rect -3090 15260 -3060 15290
rect -1590 15260 -1560 15290
rect -1090 15260 -1060 15290
rect -890 15260 -860 15290
rect -690 15260 -660 15290
rect -490 15260 -460 15290
rect -290 15260 -260 15290
rect -90 15260 -60 15290
rect -3490 15210 -3460 15240
rect -3290 15210 -3260 15240
rect -3090 15210 -3060 15240
rect -1590 15210 -1560 15240
rect -1090 15210 -1060 15240
rect -890 15210 -860 15240
rect -690 15210 -660 15240
rect -490 15210 -460 15240
rect -290 15210 -260 15240
rect -90 15210 -60 15240
rect -3490 13610 -3460 13640
rect -3290 13610 -3260 13640
rect -3090 13610 -3060 13640
rect -1590 13610 -1560 13640
rect -1090 13610 -1060 13640
rect -890 13610 -860 13640
rect -690 13610 -660 13640
rect -490 13610 -460 13640
rect -290 13610 -260 13640
rect -90 13610 -60 13640
rect -3490 13560 -3460 13590
rect -3290 13560 -3260 13590
rect -3090 13560 -3060 13590
rect -1590 13560 -1560 13590
rect -1090 13560 -1060 13590
rect -890 13560 -860 13590
rect -690 13560 -660 13590
rect -490 13560 -460 13590
rect -290 13560 -260 13590
rect -90 13560 -60 13590
rect -3490 13510 -3460 13540
rect -3290 13510 -3260 13540
rect -3090 13510 -3060 13540
rect -1590 13510 -1560 13540
rect -1090 13510 -1060 13540
rect -890 13510 -860 13540
rect -690 13510 -660 13540
rect -490 13510 -460 13540
rect -290 13510 -260 13540
rect -90 13510 -60 13540
rect -3490 11910 -3460 11940
rect -3290 11910 -3260 11940
rect -3090 11910 -3060 11940
rect -1590 11910 -1560 11940
rect -1090 11910 -1060 11940
rect -890 11910 -860 11940
rect -690 11910 -660 11940
rect -490 11910 -460 11940
rect -290 11910 -260 11940
rect -90 11910 -60 11940
rect -3490 11860 -3460 11890
rect -3290 11860 -3260 11890
rect -3090 11860 -3060 11890
rect -1590 11860 -1560 11890
rect -1090 11860 -1060 11890
rect -890 11860 -860 11890
rect -690 11860 -660 11890
rect -490 11860 -460 11890
rect -290 11860 -260 11890
rect -90 11860 -60 11890
rect -3490 11810 -3460 11840
rect -3290 11810 -3260 11840
rect -3090 11810 -3060 11840
rect -1590 11810 -1560 11840
rect -1090 11810 -1060 11840
rect -890 11810 -860 11840
rect -690 11810 -660 11840
rect -490 11810 -460 11840
rect -290 11810 -260 11840
rect -90 11810 -60 11840
rect 39810 11310 39840 11340
rect 39910 11210 39940 11240
rect 39960 11210 39990 11240
rect 40010 11210 40040 11240
rect 40060 11210 40090 11240
rect 40110 11210 40140 11240
rect 40160 11210 40190 11240
rect 40210 11210 40240 11240
rect 40260 11210 40290 11240
rect 40310 11210 40340 11240
rect 40360 11210 40390 11240
rect 40410 11210 40440 11240
rect 40460 11210 40490 11240
rect 40510 11210 40540 11240
rect 40560 11210 40590 11240
rect 40610 11210 40640 11240
rect 40660 11210 40690 11240
rect 40710 11210 40740 11240
rect 40760 11210 40790 11240
rect 40810 11210 40840 11240
rect 40860 11210 40890 11240
rect 39910 11160 39940 11190
rect 39960 11160 39990 11190
rect 40010 11160 40040 11190
rect 40060 11160 40090 11190
rect 40110 11160 40140 11190
rect 40160 11160 40190 11190
rect 40210 11160 40240 11190
rect 40260 11160 40290 11190
rect 40310 11160 40340 11190
rect 40360 11160 40390 11190
rect 40410 11160 40440 11190
rect 40460 11160 40490 11190
rect 40510 11160 40540 11190
rect 40560 11160 40590 11190
rect 40610 11160 40640 11190
rect 40660 11160 40690 11190
rect 40710 11160 40740 11190
rect 40760 11160 40790 11190
rect 40810 11160 40840 11190
rect 40860 11160 40890 11190
rect 39910 11110 39940 11140
rect 39960 11110 39990 11140
rect 40010 11110 40040 11140
rect 40060 11110 40090 11140
rect 40110 11110 40140 11140
rect 40160 11110 40190 11140
rect 40210 11110 40240 11140
rect 40260 11110 40290 11140
rect 40310 11110 40340 11140
rect 40360 11110 40390 11140
rect 40410 11110 40440 11140
rect 40460 11110 40490 11140
rect 40510 11110 40540 11140
rect 40560 11110 40590 11140
rect 40610 11110 40640 11140
rect 40660 11110 40690 11140
rect 40710 11110 40740 11140
rect 40760 11110 40790 11140
rect 40810 11110 40840 11140
rect 40860 11110 40890 11140
rect 39910 11060 39940 11090
rect 39960 11060 39990 11090
rect 40010 11060 40040 11090
rect 40060 11060 40090 11090
rect 40110 11060 40140 11090
rect 40160 11060 40190 11090
rect 40210 11060 40240 11090
rect 40260 11060 40290 11090
rect 40310 11060 40340 11090
rect 40360 11060 40390 11090
rect 40410 11060 40440 11090
rect 40460 11060 40490 11090
rect 40510 11060 40540 11090
rect 40560 11060 40590 11090
rect 40610 11060 40640 11090
rect 40660 11060 40690 11090
rect 40710 11060 40740 11090
rect 40760 11060 40790 11090
rect 40810 11060 40840 11090
rect 40860 11060 40890 11090
rect 39910 11010 39940 11040
rect 39960 11010 39990 11040
rect 40010 11010 40040 11040
rect 40060 11010 40090 11040
rect 40110 11010 40140 11040
rect 40160 11010 40190 11040
rect 40210 11010 40240 11040
rect 40260 11010 40290 11040
rect 40310 11010 40340 11040
rect 40360 11010 40390 11040
rect 40410 11010 40440 11040
rect 40460 11010 40490 11040
rect 40510 11010 40540 11040
rect 40560 11010 40590 11040
rect 40610 11010 40640 11040
rect 40660 11010 40690 11040
rect 40710 11010 40740 11040
rect 40760 11010 40790 11040
rect 40810 11010 40840 11040
rect 40860 11010 40890 11040
rect 39810 10910 39840 10940
rect -2990 10610 -2960 10640
rect -2790 10610 -2760 10640
rect -2590 10610 -2560 10640
rect -2390 10610 -2360 10640
rect -2190 10610 -2160 10640
rect -1990 10610 -1960 10640
rect -1690 10610 -1660 10640
rect -2990 10560 -2960 10590
rect -2790 10560 -2760 10590
rect -2590 10560 -2560 10590
rect -2390 10560 -2360 10590
rect -2190 10560 -2160 10590
rect -1990 10560 -1960 10590
rect -1690 10560 -1660 10590
rect -2990 10510 -2960 10540
rect -2790 10510 -2760 10540
rect -2590 10510 -2560 10540
rect -2390 10510 -2360 10540
rect -2190 10510 -2160 10540
rect -1990 10510 -1960 10540
rect -1690 10510 -1660 10540
rect -2990 9310 -2960 9340
rect -2790 9310 -2760 9340
rect -2590 9310 -2560 9340
rect -2390 9310 -2360 9340
rect -2190 9310 -2160 9340
rect -1990 9310 -1960 9340
rect -1690 9310 -1660 9340
rect -2990 9260 -2960 9290
rect -2790 9260 -2760 9290
rect -2590 9260 -2560 9290
rect -2390 9260 -2360 9290
rect -2190 9260 -2160 9290
rect -1990 9260 -1960 9290
rect -1690 9260 -1660 9290
rect -2990 9210 -2960 9240
rect -2790 9210 -2760 9240
rect -2590 9210 -2560 9240
rect -2390 9210 -2360 9240
rect -2190 9210 -2160 9240
rect -1990 9210 -1960 9240
rect -1690 9210 -1660 9240
rect -2990 8010 -2960 8040
rect -2790 8010 -2760 8040
rect -2590 8010 -2560 8040
rect -2390 8010 -2360 8040
rect -2190 8010 -2160 8040
rect -1990 8010 -1960 8040
rect -1690 8010 -1660 8040
rect -2990 7960 -2960 7990
rect -2790 7960 -2760 7990
rect -2590 7960 -2560 7990
rect -2390 7960 -2360 7990
rect -2190 7960 -2160 7990
rect -1990 7960 -1960 7990
rect -1690 7960 -1660 7990
rect -2990 7910 -2960 7940
rect -2790 7910 -2760 7940
rect -2590 7910 -2560 7940
rect -2390 7910 -2360 7940
rect -2190 7910 -2160 7940
rect -1990 7910 -1960 7940
rect -1690 7910 -1660 7940
rect -2990 7710 -2960 7740
rect -2790 7710 -2760 7740
rect -2590 7710 -2560 7740
rect -2390 7710 -2360 7740
rect -2190 7710 -2160 7740
rect -1990 7710 -1960 7740
rect -1690 7710 -1660 7740
rect -2990 7660 -2960 7690
rect -2790 7660 -2760 7690
rect -2590 7660 -2560 7690
rect -2390 7660 -2360 7690
rect -2190 7660 -2160 7690
rect -1990 7660 -1960 7690
rect -1690 7660 -1660 7690
rect -2990 7610 -2960 7640
rect -2790 7610 -2760 7640
rect -2590 7610 -2560 7640
rect -2390 7610 -2360 7640
rect -2190 7610 -2160 7640
rect -1990 7610 -1960 7640
rect -1690 7610 -1660 7640
rect -2990 6410 -2960 6440
rect -2790 6410 -2760 6440
rect -2590 6410 -2560 6440
rect -2390 6410 -2360 6440
rect -2190 6410 -2160 6440
rect -1990 6410 -1960 6440
rect -1690 6410 -1660 6440
rect -2990 6360 -2960 6390
rect -2790 6360 -2760 6390
rect -2590 6360 -2560 6390
rect -2390 6360 -2360 6390
rect -2190 6360 -2160 6390
rect -1990 6360 -1960 6390
rect -1690 6360 -1660 6390
rect -2990 6310 -2960 6340
rect -2790 6310 -2760 6340
rect -2590 6310 -2560 6340
rect -2390 6310 -2360 6340
rect -2190 6310 -2160 6340
rect -1990 6310 -1960 6340
rect -1690 6310 -1660 6340
rect -2990 5110 -2960 5140
rect -2790 5110 -2760 5140
rect -2590 5110 -2560 5140
rect -2390 5110 -2360 5140
rect -2190 5110 -2160 5140
rect -1990 5110 -1960 5140
rect -1690 5110 -1660 5140
rect -2990 5060 -2960 5090
rect -2790 5060 -2760 5090
rect -2590 5060 -2560 5090
rect -2390 5060 -2360 5090
rect -2190 5060 -2160 5090
rect -1990 5060 -1960 5090
rect -1690 5060 -1660 5090
rect -2990 5010 -2960 5040
rect -2790 5010 -2760 5040
rect -2590 5010 -2560 5040
rect -2390 5010 -2360 5040
rect -2190 5010 -2160 5040
rect -1990 5010 -1960 5040
rect -1690 5010 -1660 5040
rect 39810 4710 39840 4740
rect 39910 4610 39940 4640
rect 39960 4610 39990 4640
rect 40010 4610 40040 4640
rect 40060 4610 40090 4640
rect 40110 4610 40140 4640
rect 40160 4610 40190 4640
rect 40210 4610 40240 4640
rect 40260 4610 40290 4640
rect 40310 4610 40340 4640
rect 40360 4610 40390 4640
rect 40410 4610 40440 4640
rect 40460 4610 40490 4640
rect 40510 4610 40540 4640
rect 40560 4610 40590 4640
rect 40610 4610 40640 4640
rect 40660 4610 40690 4640
rect 40710 4610 40740 4640
rect 40760 4610 40790 4640
rect 40810 4610 40840 4640
rect 40860 4610 40890 4640
rect 39910 4560 39940 4590
rect 39960 4560 39990 4590
rect 40010 4560 40040 4590
rect 40060 4560 40090 4590
rect 40110 4560 40140 4590
rect 40160 4560 40190 4590
rect 40210 4560 40240 4590
rect 40260 4560 40290 4590
rect 40310 4560 40340 4590
rect 40360 4560 40390 4590
rect 40410 4560 40440 4590
rect 40460 4560 40490 4590
rect 40510 4560 40540 4590
rect 40560 4560 40590 4590
rect 40610 4560 40640 4590
rect 40660 4560 40690 4590
rect 40710 4560 40740 4590
rect 40760 4560 40790 4590
rect 40810 4560 40840 4590
rect 40860 4560 40890 4590
rect 39910 4510 39940 4540
rect 39960 4510 39990 4540
rect 40010 4510 40040 4540
rect 40060 4510 40090 4540
rect 40110 4510 40140 4540
rect 40160 4510 40190 4540
rect 40210 4510 40240 4540
rect 40260 4510 40290 4540
rect 40310 4510 40340 4540
rect 40360 4510 40390 4540
rect 40410 4510 40440 4540
rect 40460 4510 40490 4540
rect 40510 4510 40540 4540
rect 40560 4510 40590 4540
rect 40610 4510 40640 4540
rect 40660 4510 40690 4540
rect 40710 4510 40740 4540
rect 40760 4510 40790 4540
rect 40810 4510 40840 4540
rect 40860 4510 40890 4540
rect 39910 4460 39940 4490
rect 39960 4460 39990 4490
rect 40010 4460 40040 4490
rect 40060 4460 40090 4490
rect 40110 4460 40140 4490
rect 40160 4460 40190 4490
rect 40210 4460 40240 4490
rect 40260 4460 40290 4490
rect 40310 4460 40340 4490
rect 40360 4460 40390 4490
rect 40410 4460 40440 4490
rect 40460 4460 40490 4490
rect 40510 4460 40540 4490
rect 40560 4460 40590 4490
rect 40610 4460 40640 4490
rect 40660 4460 40690 4490
rect 40710 4460 40740 4490
rect 40760 4460 40790 4490
rect 40810 4460 40840 4490
rect 40860 4460 40890 4490
rect 39910 4410 39940 4440
rect 39960 4410 39990 4440
rect 40010 4410 40040 4440
rect 40060 4410 40090 4440
rect 40110 4410 40140 4440
rect 40160 4410 40190 4440
rect 40210 4410 40240 4440
rect 40260 4410 40290 4440
rect 40310 4410 40340 4440
rect 40360 4410 40390 4440
rect 40410 4410 40440 4440
rect 40460 4410 40490 4440
rect 40510 4410 40540 4440
rect 40560 4410 40590 4440
rect 40610 4410 40640 4440
rect 40660 4410 40690 4440
rect 40710 4410 40740 4440
rect 40760 4410 40790 4440
rect 40810 4410 40840 4440
rect 40860 4410 40890 4440
rect 39810 4310 39840 4340
rect -3490 3810 -3460 3840
rect -3290 3810 -3260 3840
rect -3090 3810 -3060 3840
rect -1590 3810 -1560 3840
rect -1090 3810 -1060 3840
rect -890 3810 -860 3840
rect -690 3810 -660 3840
rect -490 3810 -460 3840
rect -290 3810 -260 3840
rect -90 3810 -60 3840
rect -3490 3760 -3460 3790
rect -3290 3760 -3260 3790
rect -3090 3760 -3060 3790
rect -1590 3760 -1560 3790
rect -1090 3760 -1060 3790
rect -890 3760 -860 3790
rect -690 3760 -660 3790
rect -490 3760 -460 3790
rect -290 3760 -260 3790
rect -90 3760 -60 3790
rect -3490 3710 -3460 3740
rect -3290 3710 -3260 3740
rect -3090 3710 -3060 3740
rect -1590 3710 -1560 3740
rect -1090 3710 -1060 3740
rect -890 3710 -860 3740
rect -690 3710 -660 3740
rect -490 3710 -460 3740
rect -290 3710 -260 3740
rect -90 3710 -60 3740
rect -3490 2110 -3460 2140
rect -3290 2110 -3260 2140
rect -3090 2110 -3060 2140
rect -1590 2110 -1560 2140
rect -1090 2110 -1060 2140
rect -890 2110 -860 2140
rect -690 2110 -660 2140
rect -490 2110 -460 2140
rect -290 2110 -260 2140
rect -90 2110 -60 2140
rect -3490 2060 -3460 2090
rect -3290 2060 -3260 2090
rect -3090 2060 -3060 2090
rect -1590 2060 -1560 2090
rect -1090 2060 -1060 2090
rect -890 2060 -860 2090
rect -690 2060 -660 2090
rect -490 2060 -460 2090
rect -290 2060 -260 2090
rect -90 2060 -60 2090
rect -3490 2010 -3460 2040
rect -3290 2010 -3260 2040
rect -3090 2010 -3060 2040
rect -1590 2010 -1560 2040
rect -1090 2010 -1060 2040
rect -890 2010 -860 2040
rect -690 2010 -660 2040
rect -490 2010 -460 2040
rect -290 2010 -260 2040
rect -90 2010 -60 2040
rect -3490 410 -3460 440
rect -3290 410 -3260 440
rect -3090 410 -3060 440
rect -1590 410 -1560 440
rect -1090 410 -1060 440
rect -890 410 -860 440
rect -690 410 -660 440
rect -490 410 -460 440
rect -290 410 -260 440
rect -90 410 -60 440
rect -3490 360 -3460 390
rect -3290 360 -3260 390
rect -3090 360 -3060 390
rect -1590 360 -1560 390
rect -1090 360 -1060 390
rect -890 360 -860 390
rect -690 360 -660 390
rect -490 360 -460 390
rect -290 360 -260 390
rect -90 360 -60 390
rect -3490 310 -3460 340
rect -3290 310 -3260 340
rect -3090 310 -3060 340
rect -1590 310 -1560 340
rect -1090 310 -1060 340
rect -890 310 -860 340
rect -690 310 -660 340
rect -490 310 -460 340
rect -290 310 -260 340
rect -90 310 -60 340
<< metal3 >>
rect 0 18145 40900 18150
rect 0 18105 5 18145
rect 45 18105 55 18145
rect 95 18105 105 18145
rect 145 18105 155 18145
rect 195 18105 205 18145
rect 245 18105 255 18145
rect 295 18105 305 18145
rect 345 18105 355 18145
rect 395 18105 405 18145
rect 445 18105 455 18145
rect 495 18105 505 18145
rect 545 18105 555 18145
rect 595 18105 605 18145
rect 645 18105 655 18145
rect 695 18105 705 18145
rect 745 18105 755 18145
rect 795 18105 805 18145
rect 845 18105 855 18145
rect 895 18105 905 18145
rect 945 18105 955 18145
rect 995 18105 1005 18145
rect 1045 18105 1055 18145
rect 1095 18105 1105 18145
rect 1145 18105 1155 18145
rect 1195 18105 1205 18145
rect 1245 18105 1255 18145
rect 1295 18105 1305 18145
rect 1345 18105 1355 18145
rect 1395 18105 1405 18145
rect 1445 18105 1455 18145
rect 1495 18105 1505 18145
rect 1545 18105 1555 18145
rect 1595 18105 1605 18145
rect 1645 18105 1655 18145
rect 1695 18105 1705 18145
rect 1745 18105 1755 18145
rect 1795 18105 1805 18145
rect 1845 18105 1855 18145
rect 1895 18105 1905 18145
rect 1945 18105 1955 18145
rect 1995 18105 2005 18145
rect 2045 18105 2055 18145
rect 2095 18105 2105 18145
rect 2145 18105 2155 18145
rect 2195 18105 2205 18145
rect 2245 18105 2255 18145
rect 2295 18105 2305 18145
rect 2345 18105 2355 18145
rect 2395 18105 2405 18145
rect 2445 18105 2455 18145
rect 2495 18105 2505 18145
rect 2545 18105 2555 18145
rect 2595 18105 2605 18145
rect 2645 18105 2655 18145
rect 2695 18105 2705 18145
rect 2745 18105 2755 18145
rect 2795 18105 2805 18145
rect 2845 18105 2855 18145
rect 2895 18105 2905 18145
rect 2945 18105 2955 18145
rect 2995 18105 3005 18145
rect 3045 18105 3055 18145
rect 3095 18105 3105 18145
rect 3145 18105 3155 18145
rect 3195 18105 3205 18145
rect 3245 18105 3255 18145
rect 3295 18105 3305 18145
rect 3345 18105 3355 18145
rect 3395 18105 3405 18145
rect 3445 18105 3455 18145
rect 3495 18105 3505 18145
rect 3545 18105 3555 18145
rect 3595 18105 3605 18145
rect 3645 18105 3655 18145
rect 3695 18105 3705 18145
rect 3745 18105 3755 18145
rect 3795 18105 3805 18145
rect 3845 18105 3855 18145
rect 3895 18105 3905 18145
rect 3945 18105 3955 18145
rect 3995 18105 4005 18145
rect 4045 18105 4055 18145
rect 4095 18105 4105 18145
rect 4145 18105 4155 18145
rect 4195 18105 4205 18145
rect 4245 18105 4255 18145
rect 4295 18105 4305 18145
rect 4345 18105 4355 18145
rect 4395 18105 4405 18145
rect 4445 18105 4455 18145
rect 4495 18105 4505 18145
rect 4545 18105 4555 18145
rect 4595 18105 4605 18145
rect 4645 18105 4655 18145
rect 4695 18105 4705 18145
rect 4745 18105 4755 18145
rect 4795 18105 4805 18145
rect 4845 18105 4855 18145
rect 4895 18105 4905 18145
rect 4945 18105 4955 18145
rect 4995 18105 5005 18145
rect 5045 18105 5055 18145
rect 5095 18105 5105 18145
rect 5145 18105 5155 18145
rect 5195 18105 5205 18145
rect 5245 18105 5255 18145
rect 5295 18105 5305 18145
rect 5345 18105 5355 18145
rect 5395 18105 5405 18145
rect 5445 18105 5455 18145
rect 5495 18105 5505 18145
rect 5545 18105 5555 18145
rect 5595 18105 5605 18145
rect 5645 18105 5655 18145
rect 5695 18105 5705 18145
rect 5745 18105 5755 18145
rect 5795 18105 5805 18145
rect 5845 18105 5855 18145
rect 5895 18105 5905 18145
rect 5945 18105 5955 18145
rect 5995 18105 6005 18145
rect 6045 18105 6055 18145
rect 6095 18105 6105 18145
rect 6145 18105 6155 18145
rect 6195 18105 6205 18145
rect 6245 18105 6255 18145
rect 6295 18105 6305 18145
rect 6345 18105 6355 18145
rect 6395 18105 6405 18145
rect 6445 18105 6455 18145
rect 6495 18105 6505 18145
rect 6545 18105 6555 18145
rect 6595 18105 6605 18145
rect 6645 18105 6655 18145
rect 6695 18105 6705 18145
rect 6745 18105 6755 18145
rect 6795 18105 6805 18145
rect 6845 18105 6855 18145
rect 6895 18105 6905 18145
rect 6945 18105 6955 18145
rect 6995 18105 7005 18145
rect 7045 18105 7055 18145
rect 7095 18105 7105 18145
rect 7145 18105 7155 18145
rect 7195 18105 7205 18145
rect 7245 18105 7255 18145
rect 7295 18105 7305 18145
rect 7345 18105 7355 18145
rect 7395 18105 7405 18145
rect 7445 18105 7455 18145
rect 7495 18105 7505 18145
rect 7545 18105 7555 18145
rect 7595 18105 7605 18145
rect 7645 18105 7655 18145
rect 7695 18105 7705 18145
rect 7745 18105 7755 18145
rect 7795 18105 7805 18145
rect 7845 18105 7855 18145
rect 7895 18105 7905 18145
rect 7945 18105 7955 18145
rect 7995 18105 8005 18145
rect 8045 18105 8055 18145
rect 8095 18105 8105 18145
rect 8145 18105 8155 18145
rect 8195 18105 8205 18145
rect 8245 18105 8255 18145
rect 8295 18105 8305 18145
rect 8345 18105 8355 18145
rect 8395 18105 8405 18145
rect 8445 18105 8455 18145
rect 8495 18105 8505 18145
rect 8545 18105 8555 18145
rect 8595 18105 8605 18145
rect 8645 18105 8655 18145
rect 8695 18105 8705 18145
rect 8745 18105 8755 18145
rect 8795 18105 8805 18145
rect 8845 18105 8855 18145
rect 8895 18105 8905 18145
rect 8945 18105 8955 18145
rect 8995 18105 9005 18145
rect 9045 18105 9055 18145
rect 9095 18105 9105 18145
rect 9145 18105 9155 18145
rect 9195 18105 9205 18145
rect 9245 18105 9255 18145
rect 9295 18105 9305 18145
rect 9345 18105 9355 18145
rect 9395 18105 9405 18145
rect 9445 18105 9455 18145
rect 9495 18105 9505 18145
rect 9545 18105 9555 18145
rect 9595 18105 9605 18145
rect 9645 18105 9655 18145
rect 9695 18105 9705 18145
rect 9745 18105 9755 18145
rect 9795 18105 9805 18145
rect 9845 18105 9855 18145
rect 9895 18105 9905 18145
rect 9945 18105 9955 18145
rect 9995 18105 10005 18145
rect 10045 18105 10055 18145
rect 10095 18105 10105 18145
rect 10145 18105 10155 18145
rect 10195 18105 10205 18145
rect 10245 18105 10255 18145
rect 10295 18105 10305 18145
rect 10345 18105 10355 18145
rect 10395 18105 10405 18145
rect 10445 18105 10455 18145
rect 10495 18105 10505 18145
rect 10545 18105 10555 18145
rect 10595 18105 10605 18145
rect 10645 18105 10655 18145
rect 10695 18105 10705 18145
rect 10745 18105 10755 18145
rect 10795 18105 10805 18145
rect 10845 18105 10855 18145
rect 10895 18105 10905 18145
rect 10945 18105 10955 18145
rect 10995 18105 11005 18145
rect 11045 18105 11055 18145
rect 11095 18105 11105 18145
rect 11145 18105 11155 18145
rect 11195 18105 11205 18145
rect 11245 18105 11255 18145
rect 11295 18105 11305 18145
rect 11345 18105 11355 18145
rect 11395 18105 11405 18145
rect 11445 18105 11455 18145
rect 11495 18105 11505 18145
rect 11545 18105 11555 18145
rect 11595 18105 11605 18145
rect 11645 18105 11655 18145
rect 11695 18105 11705 18145
rect 11745 18105 11755 18145
rect 11795 18105 11805 18145
rect 11845 18105 11855 18145
rect 11895 18105 11905 18145
rect 11945 18105 11955 18145
rect 11995 18105 12005 18145
rect 12045 18105 12055 18145
rect 12095 18105 12105 18145
rect 12145 18105 12155 18145
rect 12195 18105 12205 18145
rect 12245 18105 12255 18145
rect 12295 18105 12305 18145
rect 12345 18105 12355 18145
rect 12395 18105 12405 18145
rect 12445 18105 12455 18145
rect 12495 18105 12505 18145
rect 12545 18105 12555 18145
rect 12595 18105 12605 18145
rect 12645 18105 12655 18145
rect 12695 18105 12705 18145
rect 12745 18105 12755 18145
rect 12795 18105 12805 18145
rect 12845 18105 12855 18145
rect 12895 18105 12905 18145
rect 12945 18105 12955 18145
rect 12995 18105 13005 18145
rect 13045 18105 13055 18145
rect 13095 18105 13105 18145
rect 13145 18105 13155 18145
rect 13195 18105 13205 18145
rect 13245 18105 13255 18145
rect 13295 18105 13305 18145
rect 13345 18105 13355 18145
rect 13395 18105 13405 18145
rect 13445 18105 13455 18145
rect 13495 18105 13505 18145
rect 13545 18105 13555 18145
rect 13595 18105 13605 18145
rect 13645 18105 13655 18145
rect 13695 18105 13705 18145
rect 13745 18105 13755 18145
rect 13795 18105 13805 18145
rect 13845 18105 13855 18145
rect 13895 18105 13905 18145
rect 13945 18105 13955 18145
rect 13995 18105 14005 18145
rect 14045 18105 14055 18145
rect 14095 18105 14105 18145
rect 14145 18105 14155 18145
rect 14195 18105 14205 18145
rect 14245 18105 14255 18145
rect 14295 18105 14305 18145
rect 14345 18105 14355 18145
rect 14395 18105 14405 18145
rect 14445 18105 14455 18145
rect 14495 18105 14505 18145
rect 14545 18105 14555 18145
rect 14595 18105 14605 18145
rect 14645 18105 14655 18145
rect 14695 18105 14705 18145
rect 14745 18105 14755 18145
rect 14795 18105 14805 18145
rect 14845 18105 14855 18145
rect 14895 18105 14905 18145
rect 14945 18105 14955 18145
rect 14995 18105 15005 18145
rect 15045 18105 15055 18145
rect 15095 18105 15105 18145
rect 15145 18105 15155 18145
rect 15195 18105 15205 18145
rect 15245 18105 15255 18145
rect 15295 18105 15305 18145
rect 15345 18105 15355 18145
rect 15395 18105 15405 18145
rect 15445 18105 15455 18145
rect 15495 18105 15505 18145
rect 15545 18105 15555 18145
rect 15595 18105 15605 18145
rect 15645 18105 15655 18145
rect 15695 18105 15705 18145
rect 15745 18105 15755 18145
rect 15795 18105 15805 18145
rect 15845 18105 15855 18145
rect 15895 18105 15905 18145
rect 15945 18105 15955 18145
rect 15995 18105 16005 18145
rect 16045 18105 16055 18145
rect 16095 18105 16105 18145
rect 16145 18105 16155 18145
rect 16195 18105 16205 18145
rect 16245 18105 16255 18145
rect 16295 18105 16305 18145
rect 16345 18105 16355 18145
rect 16395 18105 16405 18145
rect 16445 18105 16455 18145
rect 16495 18105 16505 18145
rect 16545 18105 16555 18145
rect 16595 18105 16605 18145
rect 16645 18105 16655 18145
rect 16695 18105 16705 18145
rect 16745 18105 16755 18145
rect 16795 18105 16805 18145
rect 16845 18105 16855 18145
rect 16895 18105 16905 18145
rect 16945 18105 16955 18145
rect 16995 18105 17005 18145
rect 17045 18105 17055 18145
rect 17095 18105 17105 18145
rect 17145 18105 17155 18145
rect 17195 18105 17205 18145
rect 17245 18105 17255 18145
rect 17295 18105 17305 18145
rect 17345 18105 17355 18145
rect 17395 18105 17405 18145
rect 17445 18105 17455 18145
rect 17495 18105 17505 18145
rect 17545 18105 17555 18145
rect 17595 18105 17605 18145
rect 17645 18105 17655 18145
rect 17695 18105 17705 18145
rect 17745 18105 17755 18145
rect 17795 18105 17805 18145
rect 17845 18105 17855 18145
rect 17895 18105 17905 18145
rect 17945 18105 17955 18145
rect 17995 18105 18005 18145
rect 18045 18105 18055 18145
rect 18095 18105 18105 18145
rect 18145 18105 18155 18145
rect 18195 18105 18205 18145
rect 18245 18105 18255 18145
rect 18295 18105 18305 18145
rect 18345 18105 18355 18145
rect 18395 18105 18405 18145
rect 18445 18105 18455 18145
rect 18495 18105 18505 18145
rect 18545 18105 18555 18145
rect 18595 18105 18605 18145
rect 18645 18105 18655 18145
rect 18695 18105 18705 18145
rect 18745 18105 18755 18145
rect 18795 18105 18805 18145
rect 18845 18105 18855 18145
rect 18895 18105 18905 18145
rect 18945 18105 18955 18145
rect 18995 18105 19005 18145
rect 19045 18105 19055 18145
rect 19095 18105 19105 18145
rect 19145 18105 19155 18145
rect 19195 18105 19205 18145
rect 19245 18105 19255 18145
rect 19295 18105 19305 18145
rect 19345 18105 19355 18145
rect 19395 18105 19405 18145
rect 19445 18105 19455 18145
rect 19495 18105 19505 18145
rect 19545 18105 19555 18145
rect 19595 18105 19605 18145
rect 19645 18105 19655 18145
rect 19695 18105 19705 18145
rect 19745 18105 19755 18145
rect 19795 18105 19805 18145
rect 19845 18105 19855 18145
rect 19895 18105 19905 18145
rect 19945 18105 19955 18145
rect 19995 18105 20005 18145
rect 20045 18105 20055 18145
rect 20095 18105 20105 18145
rect 20145 18105 20155 18145
rect 20195 18105 20205 18145
rect 20245 18105 20255 18145
rect 20295 18105 20305 18145
rect 20345 18105 20355 18145
rect 20395 18105 20405 18145
rect 20445 18105 20455 18145
rect 20495 18105 20505 18145
rect 20545 18105 20555 18145
rect 20595 18105 20605 18145
rect 20645 18105 20655 18145
rect 20695 18105 20705 18145
rect 20745 18105 20755 18145
rect 20795 18105 20805 18145
rect 20845 18105 20855 18145
rect 20895 18105 20905 18145
rect 20945 18105 20955 18145
rect 20995 18105 21005 18145
rect 21045 18105 21055 18145
rect 21095 18105 21105 18145
rect 21145 18105 21155 18145
rect 21195 18105 21205 18145
rect 21245 18105 21255 18145
rect 21295 18105 21305 18145
rect 21345 18105 21355 18145
rect 21395 18105 21405 18145
rect 21445 18105 21455 18145
rect 21495 18105 21505 18145
rect 21545 18105 21555 18145
rect 21595 18105 21605 18145
rect 21645 18105 21655 18145
rect 21695 18105 21705 18145
rect 21745 18105 21755 18145
rect 21795 18105 21805 18145
rect 21845 18105 21855 18145
rect 21895 18105 21905 18145
rect 21945 18105 21955 18145
rect 21995 18105 22005 18145
rect 22045 18105 22055 18145
rect 22095 18105 22105 18145
rect 22145 18105 22155 18145
rect 22195 18105 22205 18145
rect 22245 18105 22255 18145
rect 22295 18105 22305 18145
rect 22345 18105 22355 18145
rect 22395 18105 22405 18145
rect 22445 18105 22455 18145
rect 22495 18105 22505 18145
rect 22545 18105 22555 18145
rect 22595 18105 22605 18145
rect 22645 18105 22655 18145
rect 22695 18105 22705 18145
rect 22745 18105 22755 18145
rect 22795 18105 22805 18145
rect 22845 18105 22855 18145
rect 22895 18105 22905 18145
rect 22945 18105 22955 18145
rect 22995 18105 23005 18145
rect 23045 18105 23055 18145
rect 23095 18105 23105 18145
rect 23145 18105 23155 18145
rect 23195 18105 23205 18145
rect 23245 18105 23255 18145
rect 23295 18105 23305 18145
rect 23345 18105 23355 18145
rect 23395 18105 23405 18145
rect 23445 18105 23455 18145
rect 23495 18105 23505 18145
rect 23545 18105 23555 18145
rect 23595 18105 23605 18145
rect 23645 18105 23655 18145
rect 23695 18105 23705 18145
rect 23745 18105 23755 18145
rect 23795 18105 23805 18145
rect 23845 18105 23855 18145
rect 23895 18105 23905 18145
rect 23945 18105 23955 18145
rect 23995 18105 24005 18145
rect 24045 18105 24055 18145
rect 24095 18105 24105 18145
rect 24145 18105 24155 18145
rect 24195 18105 24205 18145
rect 24245 18105 24255 18145
rect 24295 18105 24305 18145
rect 24345 18105 24355 18145
rect 24395 18105 24405 18145
rect 24445 18105 24455 18145
rect 24495 18105 24505 18145
rect 24545 18105 24555 18145
rect 24595 18105 24605 18145
rect 24645 18105 24655 18145
rect 24695 18105 24705 18145
rect 24745 18105 24755 18145
rect 24795 18105 24805 18145
rect 24845 18105 24855 18145
rect 24895 18105 24905 18145
rect 24945 18105 24955 18145
rect 24995 18105 25005 18145
rect 25045 18105 25055 18145
rect 25095 18105 25105 18145
rect 25145 18105 25155 18145
rect 25195 18105 25205 18145
rect 25245 18105 25255 18145
rect 25295 18105 25305 18145
rect 25345 18105 25355 18145
rect 25395 18105 25405 18145
rect 25445 18105 25455 18145
rect 25495 18105 25505 18145
rect 25545 18105 25555 18145
rect 25595 18105 25605 18145
rect 25645 18105 25655 18145
rect 25695 18105 25705 18145
rect 25745 18105 25755 18145
rect 25795 18105 25805 18145
rect 25845 18105 25855 18145
rect 25895 18105 25905 18145
rect 25945 18105 25955 18145
rect 25995 18105 26005 18145
rect 26045 18105 26055 18145
rect 26095 18105 26105 18145
rect 26145 18105 26155 18145
rect 26195 18105 26205 18145
rect 26245 18105 26255 18145
rect 26295 18105 26305 18145
rect 26345 18105 26355 18145
rect 26395 18105 26405 18145
rect 26445 18105 26455 18145
rect 26495 18105 26505 18145
rect 26545 18105 26555 18145
rect 26595 18105 26605 18145
rect 26645 18105 26655 18145
rect 26695 18105 26705 18145
rect 26745 18105 26755 18145
rect 26795 18105 26805 18145
rect 26845 18105 26855 18145
rect 26895 18105 26905 18145
rect 26945 18105 26955 18145
rect 26995 18105 27005 18145
rect 27045 18105 27055 18145
rect 27095 18105 27105 18145
rect 27145 18105 27155 18145
rect 27195 18105 27205 18145
rect 27245 18105 27255 18145
rect 27295 18105 27305 18145
rect 27345 18105 27355 18145
rect 27395 18105 27405 18145
rect 27445 18105 27455 18145
rect 27495 18105 27505 18145
rect 27545 18105 27555 18145
rect 27595 18105 27605 18145
rect 27645 18105 27655 18145
rect 27695 18105 27705 18145
rect 27745 18105 27755 18145
rect 27795 18105 27805 18145
rect 27845 18105 27855 18145
rect 27895 18105 27905 18145
rect 27945 18105 27955 18145
rect 27995 18105 28005 18145
rect 28045 18105 28055 18145
rect 28095 18105 28105 18145
rect 28145 18105 28155 18145
rect 28195 18105 28205 18145
rect 28245 18105 28255 18145
rect 28295 18105 28305 18145
rect 28345 18105 28355 18145
rect 28395 18105 28405 18145
rect 28445 18105 28455 18145
rect 28495 18105 28505 18145
rect 28545 18105 28555 18145
rect 28595 18105 28605 18145
rect 28645 18105 28655 18145
rect 28695 18105 28705 18145
rect 28745 18105 28755 18145
rect 28795 18105 28805 18145
rect 28845 18105 28855 18145
rect 28895 18105 28905 18145
rect 28945 18105 28955 18145
rect 28995 18105 29005 18145
rect 29045 18105 29055 18145
rect 29095 18105 29105 18145
rect 29145 18105 29155 18145
rect 29195 18105 29205 18145
rect 29245 18105 29255 18145
rect 29295 18105 29305 18145
rect 29345 18105 29355 18145
rect 29395 18105 29405 18145
rect 29445 18105 29455 18145
rect 29495 18105 29505 18145
rect 29545 18105 29555 18145
rect 29595 18105 29605 18145
rect 29645 18105 29655 18145
rect 29695 18105 29705 18145
rect 29745 18105 29755 18145
rect 29795 18105 29805 18145
rect 29845 18105 29855 18145
rect 29895 18105 29905 18145
rect 29945 18105 29955 18145
rect 29995 18105 30005 18145
rect 30045 18105 30055 18145
rect 30095 18105 30105 18145
rect 30145 18105 30155 18145
rect 30195 18105 30205 18145
rect 30245 18105 30255 18145
rect 30295 18105 30305 18145
rect 30345 18105 30355 18145
rect 30395 18105 30405 18145
rect 30445 18105 30455 18145
rect 30495 18105 30505 18145
rect 30545 18105 30555 18145
rect 30595 18105 30605 18145
rect 30645 18105 30655 18145
rect 30695 18105 30705 18145
rect 30745 18105 30755 18145
rect 30795 18105 30805 18145
rect 30845 18105 30855 18145
rect 30895 18105 30905 18145
rect 30945 18105 30955 18145
rect 30995 18105 31005 18145
rect 31045 18105 31055 18145
rect 31095 18105 31105 18145
rect 31145 18105 31155 18145
rect 31195 18105 31205 18145
rect 31245 18105 31255 18145
rect 31295 18105 31305 18145
rect 31345 18105 31355 18145
rect 31395 18105 31405 18145
rect 31445 18105 31455 18145
rect 31495 18105 31505 18145
rect 31545 18105 31555 18145
rect 31595 18105 31605 18145
rect 31645 18105 31655 18145
rect 31695 18105 31705 18145
rect 31745 18105 31755 18145
rect 31795 18105 31805 18145
rect 31845 18105 31855 18145
rect 31895 18105 31905 18145
rect 31945 18105 31955 18145
rect 31995 18105 32005 18145
rect 32045 18105 32055 18145
rect 32095 18105 32105 18145
rect 32145 18105 32155 18145
rect 32195 18105 32205 18145
rect 32245 18105 32255 18145
rect 32295 18105 32305 18145
rect 32345 18105 32355 18145
rect 32395 18105 32405 18145
rect 32445 18105 32455 18145
rect 32495 18105 32505 18145
rect 32545 18105 32555 18145
rect 32595 18105 32605 18145
rect 32645 18105 32655 18145
rect 32695 18105 32705 18145
rect 32745 18105 32755 18145
rect 32795 18105 32805 18145
rect 32845 18105 32855 18145
rect 32895 18105 32905 18145
rect 32945 18105 32955 18145
rect 32995 18105 33005 18145
rect 33045 18105 33055 18145
rect 33095 18105 33105 18145
rect 33145 18105 33155 18145
rect 33195 18105 33205 18145
rect 33245 18105 33255 18145
rect 33295 18105 33305 18145
rect 33345 18105 33355 18145
rect 33395 18105 33405 18145
rect 33445 18105 33455 18145
rect 33495 18105 33505 18145
rect 33545 18105 33555 18145
rect 33595 18105 33605 18145
rect 33645 18105 33655 18145
rect 33695 18105 33705 18145
rect 33745 18105 33755 18145
rect 33795 18105 33805 18145
rect 33845 18105 33855 18145
rect 33895 18105 33905 18145
rect 33945 18105 33955 18145
rect 33995 18105 34005 18145
rect 34045 18105 34055 18145
rect 34095 18105 34105 18145
rect 34145 18105 34155 18145
rect 34195 18105 34205 18145
rect 34245 18105 34255 18145
rect 34295 18105 34305 18145
rect 34345 18105 34355 18145
rect 34395 18105 34405 18145
rect 34445 18105 34455 18145
rect 34495 18105 34505 18145
rect 34545 18105 34555 18145
rect 34595 18105 34605 18145
rect 34645 18105 34655 18145
rect 34695 18105 34705 18145
rect 34745 18105 34755 18145
rect 34795 18105 34805 18145
rect 34845 18105 34855 18145
rect 34895 18105 34905 18145
rect 34945 18105 34955 18145
rect 34995 18105 35005 18145
rect 35045 18105 35055 18145
rect 35095 18105 35105 18145
rect 35145 18105 35155 18145
rect 35195 18105 35205 18145
rect 35245 18105 35255 18145
rect 35295 18105 35305 18145
rect 35345 18105 35355 18145
rect 35395 18105 35405 18145
rect 35445 18105 35455 18145
rect 35495 18105 35505 18145
rect 35545 18105 35555 18145
rect 35595 18105 35605 18145
rect 35645 18105 35655 18145
rect 35695 18105 35705 18145
rect 35745 18105 35755 18145
rect 35795 18105 35805 18145
rect 35845 18105 35855 18145
rect 35895 18105 35905 18145
rect 35945 18105 35955 18145
rect 35995 18105 36005 18145
rect 36045 18105 36055 18145
rect 36095 18105 36105 18145
rect 36145 18105 36155 18145
rect 36195 18105 36205 18145
rect 36245 18105 36255 18145
rect 36295 18105 36305 18145
rect 36345 18105 36355 18145
rect 36395 18105 36405 18145
rect 36445 18105 36455 18145
rect 36495 18105 36505 18145
rect 36545 18105 36555 18145
rect 36595 18105 36605 18145
rect 36645 18105 36655 18145
rect 36695 18105 36705 18145
rect 36745 18105 36755 18145
rect 36795 18105 36805 18145
rect 36845 18105 36855 18145
rect 36895 18105 36905 18145
rect 36945 18105 36955 18145
rect 36995 18105 37005 18145
rect 37045 18105 37055 18145
rect 37095 18105 37105 18145
rect 37145 18105 37155 18145
rect 37195 18105 37205 18145
rect 37245 18105 37255 18145
rect 37295 18105 37305 18145
rect 37345 18105 37355 18145
rect 37395 18105 37405 18145
rect 37445 18105 37455 18145
rect 37495 18105 37505 18145
rect 37545 18105 37555 18145
rect 37595 18105 37605 18145
rect 37645 18105 37655 18145
rect 37695 18105 37705 18145
rect 37745 18105 37755 18145
rect 37795 18105 37805 18145
rect 37845 18105 37855 18145
rect 37895 18105 37905 18145
rect 37945 18105 37955 18145
rect 37995 18105 38005 18145
rect 38045 18105 38055 18145
rect 38095 18105 38105 18145
rect 38145 18105 38155 18145
rect 38195 18105 38205 18145
rect 38245 18105 38255 18145
rect 38295 18105 38305 18145
rect 38345 18105 38355 18145
rect 38395 18105 38405 18145
rect 38445 18105 38455 18145
rect 38495 18105 38505 18145
rect 38545 18105 38555 18145
rect 38595 18105 38605 18145
rect 38645 18105 38655 18145
rect 38695 18105 38705 18145
rect 38745 18105 38755 18145
rect 38795 18105 38805 18145
rect 38845 18105 38855 18145
rect 38895 18105 38905 18145
rect 38945 18105 38955 18145
rect 38995 18105 39005 18145
rect 39045 18105 39055 18145
rect 39095 18105 39105 18145
rect 39145 18105 39155 18145
rect 39195 18105 39205 18145
rect 39245 18105 39255 18145
rect 39295 18105 39305 18145
rect 39345 18105 39355 18145
rect 39395 18105 39405 18145
rect 39445 18105 39455 18145
rect 39495 18105 39505 18145
rect 39545 18105 39555 18145
rect 39595 18105 39605 18145
rect 39645 18105 39655 18145
rect 39695 18105 39705 18145
rect 39745 18105 39905 18145
rect 39945 18105 39955 18145
rect 39995 18105 40005 18145
rect 40045 18105 40055 18145
rect 40095 18105 40105 18145
rect 40145 18105 40155 18145
rect 40195 18105 40205 18145
rect 40245 18105 40255 18145
rect 40295 18105 40305 18145
rect 40345 18105 40355 18145
rect 40395 18105 40405 18145
rect 40445 18105 40455 18145
rect 40495 18105 40505 18145
rect 40545 18105 40555 18145
rect 40595 18105 40605 18145
rect 40645 18105 40655 18145
rect 40695 18105 40705 18145
rect 40745 18105 40755 18145
rect 40795 18105 40805 18145
rect 40845 18105 40855 18145
rect 40895 18105 40900 18145
rect 0 18100 40900 18105
rect 0 18045 39750 18050
rect 0 18005 5 18045
rect 45 18005 55 18045
rect 95 18005 105 18045
rect 145 18005 155 18045
rect 195 18005 205 18045
rect 245 18005 255 18045
rect 295 18005 305 18045
rect 345 18005 355 18045
rect 395 18005 405 18045
rect 445 18005 455 18045
rect 495 18005 505 18045
rect 545 18005 555 18045
rect 595 18005 605 18045
rect 645 18005 655 18045
rect 695 18005 705 18045
rect 745 18005 755 18045
rect 795 18005 805 18045
rect 845 18005 855 18045
rect 895 18005 905 18045
rect 945 18005 955 18045
rect 995 18005 1005 18045
rect 1045 18005 1055 18045
rect 1095 18005 1105 18045
rect 1145 18005 1155 18045
rect 1195 18005 1205 18045
rect 1245 18005 1255 18045
rect 1295 18005 1305 18045
rect 1345 18005 1355 18045
rect 1395 18005 1405 18045
rect 1445 18005 1455 18045
rect 1495 18005 1505 18045
rect 1545 18005 1555 18045
rect 1595 18005 1605 18045
rect 1645 18005 1655 18045
rect 1695 18005 1705 18045
rect 1745 18005 1755 18045
rect 1795 18005 1805 18045
rect 1845 18005 1855 18045
rect 1895 18005 1905 18045
rect 1945 18005 1955 18045
rect 1995 18005 2005 18045
rect 2045 18005 2055 18045
rect 2095 18005 2105 18045
rect 2145 18005 2155 18045
rect 2195 18005 2205 18045
rect 2245 18005 2255 18045
rect 2295 18005 2305 18045
rect 2345 18005 2355 18045
rect 2395 18005 2405 18045
rect 2445 18005 2455 18045
rect 2495 18005 2505 18045
rect 2545 18005 2555 18045
rect 2595 18005 2605 18045
rect 2645 18005 2655 18045
rect 2695 18005 2705 18045
rect 2745 18005 2755 18045
rect 2795 18005 2805 18045
rect 2845 18005 2855 18045
rect 2895 18005 2905 18045
rect 2945 18005 2955 18045
rect 2995 18005 3005 18045
rect 3045 18005 3055 18045
rect 3095 18005 3105 18045
rect 3145 18005 3155 18045
rect 3195 18005 3205 18045
rect 3245 18005 3255 18045
rect 3295 18005 3305 18045
rect 3345 18005 3355 18045
rect 3395 18005 3405 18045
rect 3445 18005 3455 18045
rect 3495 18005 3505 18045
rect 3545 18005 3555 18045
rect 3595 18005 3605 18045
rect 3645 18005 3655 18045
rect 3695 18005 3705 18045
rect 3745 18005 3755 18045
rect 3795 18005 3805 18045
rect 3845 18005 3855 18045
rect 3895 18005 3905 18045
rect 3945 18005 3955 18045
rect 3995 18005 4005 18045
rect 4045 18005 4055 18045
rect 4095 18005 4105 18045
rect 4145 18005 4155 18045
rect 4195 18005 4205 18045
rect 4245 18005 4255 18045
rect 4295 18005 4305 18045
rect 4345 18005 4355 18045
rect 4395 18005 4405 18045
rect 4445 18005 4455 18045
rect 4495 18005 4505 18045
rect 4545 18005 4555 18045
rect 4595 18005 4605 18045
rect 4645 18005 4655 18045
rect 4695 18005 4705 18045
rect 4745 18005 4755 18045
rect 4795 18005 4805 18045
rect 4845 18005 4855 18045
rect 4895 18005 4905 18045
rect 4945 18005 4955 18045
rect 4995 18005 5005 18045
rect 5045 18005 5055 18045
rect 5095 18005 5105 18045
rect 5145 18005 5155 18045
rect 5195 18005 5205 18045
rect 5245 18005 5255 18045
rect 5295 18005 5305 18045
rect 5345 18005 5355 18045
rect 5395 18005 5405 18045
rect 5445 18005 5455 18045
rect 5495 18005 5505 18045
rect 5545 18005 5555 18045
rect 5595 18005 5605 18045
rect 5645 18005 5655 18045
rect 5695 18005 5705 18045
rect 5745 18005 5755 18045
rect 5795 18005 5805 18045
rect 5845 18005 5855 18045
rect 5895 18005 5905 18045
rect 5945 18005 5955 18045
rect 5995 18005 6005 18045
rect 6045 18005 6055 18045
rect 6095 18005 6105 18045
rect 6145 18005 6155 18045
rect 6195 18005 6205 18045
rect 6245 18005 6255 18045
rect 6295 18005 6305 18045
rect 6345 18005 6355 18045
rect 6395 18005 6405 18045
rect 6445 18005 6455 18045
rect 6495 18005 6505 18045
rect 6545 18005 6555 18045
rect 6595 18005 6605 18045
rect 6645 18005 6655 18045
rect 6695 18005 6705 18045
rect 6745 18005 6755 18045
rect 6795 18005 6805 18045
rect 6845 18005 6855 18045
rect 6895 18005 6905 18045
rect 6945 18005 6955 18045
rect 6995 18005 7005 18045
rect 7045 18005 7055 18045
rect 7095 18005 7105 18045
rect 7145 18005 7155 18045
rect 7195 18005 7205 18045
rect 7245 18005 7255 18045
rect 7295 18005 7305 18045
rect 7345 18005 7355 18045
rect 7395 18005 7405 18045
rect 7445 18005 7455 18045
rect 7495 18005 7505 18045
rect 7545 18005 7555 18045
rect 7595 18005 7605 18045
rect 7645 18005 7655 18045
rect 7695 18005 7705 18045
rect 7745 18005 7755 18045
rect 7795 18005 7805 18045
rect 7845 18005 7855 18045
rect 7895 18005 7905 18045
rect 7945 18005 7955 18045
rect 7995 18005 8005 18045
rect 8045 18005 8055 18045
rect 8095 18005 8105 18045
rect 8145 18005 8155 18045
rect 8195 18005 8205 18045
rect 8245 18005 8255 18045
rect 8295 18005 8305 18045
rect 8345 18005 8355 18045
rect 8395 18005 8405 18045
rect 8445 18005 8455 18045
rect 8495 18005 8505 18045
rect 8545 18005 8555 18045
rect 8595 18005 8605 18045
rect 8645 18005 8655 18045
rect 8695 18005 8705 18045
rect 8745 18005 8755 18045
rect 8795 18005 8805 18045
rect 8845 18005 8855 18045
rect 8895 18005 8905 18045
rect 8945 18005 8955 18045
rect 8995 18005 9005 18045
rect 9045 18005 9055 18045
rect 9095 18005 9105 18045
rect 9145 18005 9155 18045
rect 9195 18005 9205 18045
rect 9245 18005 9255 18045
rect 9295 18005 9305 18045
rect 9345 18005 9355 18045
rect 9395 18005 9405 18045
rect 9445 18005 9455 18045
rect 9495 18005 9505 18045
rect 9545 18005 9555 18045
rect 9595 18005 9605 18045
rect 9645 18005 9655 18045
rect 9695 18005 9705 18045
rect 9745 18005 9755 18045
rect 9795 18005 9805 18045
rect 9845 18005 9855 18045
rect 9895 18005 9905 18045
rect 9945 18005 9955 18045
rect 9995 18005 10005 18045
rect 10045 18005 10055 18045
rect 10095 18005 10105 18045
rect 10145 18005 10155 18045
rect 10195 18005 10205 18045
rect 10245 18005 10255 18045
rect 10295 18005 10305 18045
rect 10345 18005 10355 18045
rect 10395 18005 10405 18045
rect 10445 18005 10455 18045
rect 10495 18005 10505 18045
rect 10545 18005 10555 18045
rect 10595 18005 10605 18045
rect 10645 18005 10655 18045
rect 10695 18005 10705 18045
rect 10745 18005 10755 18045
rect 10795 18005 10805 18045
rect 10845 18005 10855 18045
rect 10895 18005 10905 18045
rect 10945 18005 10955 18045
rect 10995 18005 11005 18045
rect 11045 18005 11055 18045
rect 11095 18005 11105 18045
rect 11145 18005 11155 18045
rect 11195 18005 11205 18045
rect 11245 18005 11255 18045
rect 11295 18005 11305 18045
rect 11345 18005 11355 18045
rect 11395 18005 11405 18045
rect 11445 18005 11455 18045
rect 11495 18005 11505 18045
rect 11545 18005 11555 18045
rect 11595 18005 11605 18045
rect 11645 18005 11655 18045
rect 11695 18005 11705 18045
rect 11745 18005 11755 18045
rect 11795 18005 11805 18045
rect 11845 18005 11855 18045
rect 11895 18005 11905 18045
rect 11945 18005 11955 18045
rect 11995 18005 12005 18045
rect 12045 18005 12055 18045
rect 12095 18005 12105 18045
rect 12145 18005 12155 18045
rect 12195 18005 12205 18045
rect 12245 18005 12255 18045
rect 12295 18005 12305 18045
rect 12345 18005 12355 18045
rect 12395 18005 12405 18045
rect 12445 18005 12455 18045
rect 12495 18005 12505 18045
rect 12545 18005 12555 18045
rect 12595 18005 12605 18045
rect 12645 18005 12655 18045
rect 12695 18005 12705 18045
rect 12745 18005 12755 18045
rect 12795 18005 12805 18045
rect 12845 18005 12855 18045
rect 12895 18005 12905 18045
rect 12945 18005 12955 18045
rect 12995 18005 13005 18045
rect 13045 18005 13055 18045
rect 13095 18005 13105 18045
rect 13145 18005 13155 18045
rect 13195 18005 13205 18045
rect 13245 18005 13255 18045
rect 13295 18005 13305 18045
rect 13345 18005 13355 18045
rect 13395 18005 13405 18045
rect 13445 18005 13455 18045
rect 13495 18005 13505 18045
rect 13545 18005 13555 18045
rect 13595 18005 13605 18045
rect 13645 18005 13655 18045
rect 13695 18005 13705 18045
rect 13745 18005 13755 18045
rect 13795 18005 13805 18045
rect 13845 18005 13855 18045
rect 13895 18005 13905 18045
rect 13945 18005 13955 18045
rect 13995 18005 14005 18045
rect 14045 18005 14055 18045
rect 14095 18005 14105 18045
rect 14145 18005 14155 18045
rect 14195 18005 14205 18045
rect 14245 18005 14255 18045
rect 14295 18005 14305 18045
rect 14345 18005 14355 18045
rect 14395 18005 14405 18045
rect 14445 18005 14455 18045
rect 14495 18005 14505 18045
rect 14545 18005 14555 18045
rect 14595 18005 14605 18045
rect 14645 18005 14655 18045
rect 14695 18005 14705 18045
rect 14745 18005 14755 18045
rect 14795 18005 14805 18045
rect 14845 18005 14855 18045
rect 14895 18005 14905 18045
rect 14945 18005 14955 18045
rect 14995 18005 15005 18045
rect 15045 18005 15055 18045
rect 15095 18005 15105 18045
rect 15145 18005 15155 18045
rect 15195 18005 15205 18045
rect 15245 18005 15255 18045
rect 15295 18005 15305 18045
rect 15345 18005 15355 18045
rect 15395 18005 15405 18045
rect 15445 18005 15455 18045
rect 15495 18005 15505 18045
rect 15545 18005 15555 18045
rect 15595 18005 15605 18045
rect 15645 18005 15655 18045
rect 15695 18005 15705 18045
rect 15745 18005 15755 18045
rect 15795 18005 15805 18045
rect 15845 18005 15855 18045
rect 15895 18005 15905 18045
rect 15945 18005 15955 18045
rect 15995 18005 16005 18045
rect 16045 18005 16055 18045
rect 16095 18005 16105 18045
rect 16145 18005 16155 18045
rect 16195 18005 16205 18045
rect 16245 18005 16255 18045
rect 16295 18005 16305 18045
rect 16345 18005 16355 18045
rect 16395 18005 16405 18045
rect 16445 18005 16455 18045
rect 16495 18005 16505 18045
rect 16545 18005 16555 18045
rect 16595 18005 16605 18045
rect 16645 18005 16655 18045
rect 16695 18005 16705 18045
rect 16745 18005 16755 18045
rect 16795 18005 16805 18045
rect 16845 18005 16855 18045
rect 16895 18005 16905 18045
rect 16945 18005 16955 18045
rect 16995 18005 17005 18045
rect 17045 18005 17055 18045
rect 17095 18005 17105 18045
rect 17145 18005 17155 18045
rect 17195 18005 17205 18045
rect 17245 18005 17255 18045
rect 17295 18005 17305 18045
rect 17345 18005 17355 18045
rect 17395 18005 17405 18045
rect 17445 18005 17455 18045
rect 17495 18005 17505 18045
rect 17545 18005 17555 18045
rect 17595 18005 17605 18045
rect 17645 18005 17655 18045
rect 17695 18005 17705 18045
rect 17745 18005 17755 18045
rect 17795 18005 17805 18045
rect 17845 18005 17855 18045
rect 17895 18005 17905 18045
rect 17945 18005 17955 18045
rect 17995 18005 18005 18045
rect 18045 18005 18055 18045
rect 18095 18005 18105 18045
rect 18145 18005 18155 18045
rect 18195 18005 18205 18045
rect 18245 18005 18255 18045
rect 18295 18005 18305 18045
rect 18345 18005 18355 18045
rect 18395 18005 18405 18045
rect 18445 18005 18455 18045
rect 18495 18005 18505 18045
rect 18545 18005 18555 18045
rect 18595 18005 18605 18045
rect 18645 18005 18655 18045
rect 18695 18005 18705 18045
rect 18745 18005 18755 18045
rect 18795 18005 18805 18045
rect 18845 18005 18855 18045
rect 18895 18005 18905 18045
rect 18945 18005 18955 18045
rect 18995 18005 19005 18045
rect 19045 18005 19055 18045
rect 19095 18005 19105 18045
rect 19145 18005 19155 18045
rect 19195 18005 19205 18045
rect 19245 18005 19255 18045
rect 19295 18005 19305 18045
rect 19345 18005 19355 18045
rect 19395 18005 19405 18045
rect 19445 18005 19455 18045
rect 19495 18005 19505 18045
rect 19545 18005 19555 18045
rect 19595 18005 19605 18045
rect 19645 18005 19655 18045
rect 19695 18005 19705 18045
rect 19745 18005 19755 18045
rect 19795 18005 19805 18045
rect 19845 18005 19855 18045
rect 19895 18005 19905 18045
rect 19945 18005 19955 18045
rect 19995 18005 20005 18045
rect 20045 18005 20055 18045
rect 20095 18005 20105 18045
rect 20145 18005 20155 18045
rect 20195 18005 20205 18045
rect 20245 18005 20255 18045
rect 20295 18005 20305 18045
rect 20345 18005 20355 18045
rect 20395 18005 20405 18045
rect 20445 18005 20455 18045
rect 20495 18005 20505 18045
rect 20545 18005 20555 18045
rect 20595 18005 20605 18045
rect 20645 18005 20655 18045
rect 20695 18005 20705 18045
rect 20745 18005 20755 18045
rect 20795 18005 20805 18045
rect 20845 18005 20855 18045
rect 20895 18005 20905 18045
rect 20945 18005 20955 18045
rect 20995 18005 21005 18045
rect 21045 18005 21055 18045
rect 21095 18005 21105 18045
rect 21145 18005 21155 18045
rect 21195 18005 21205 18045
rect 21245 18005 21255 18045
rect 21295 18005 21305 18045
rect 21345 18005 21355 18045
rect 21395 18005 21405 18045
rect 21445 18005 21455 18045
rect 21495 18005 21505 18045
rect 21545 18005 21555 18045
rect 21595 18005 21605 18045
rect 21645 18005 21655 18045
rect 21695 18005 21705 18045
rect 21745 18005 21755 18045
rect 21795 18005 21805 18045
rect 21845 18005 21855 18045
rect 21895 18005 21905 18045
rect 21945 18005 21955 18045
rect 21995 18005 22005 18045
rect 22045 18005 22055 18045
rect 22095 18005 22105 18045
rect 22145 18005 22155 18045
rect 22195 18005 22205 18045
rect 22245 18005 22255 18045
rect 22295 18005 22305 18045
rect 22345 18005 22355 18045
rect 22395 18005 22405 18045
rect 22445 18005 22455 18045
rect 22495 18005 22505 18045
rect 22545 18005 22555 18045
rect 22595 18005 22605 18045
rect 22645 18005 22655 18045
rect 22695 18005 22705 18045
rect 22745 18005 22755 18045
rect 22795 18005 22805 18045
rect 22845 18005 22855 18045
rect 22895 18005 22905 18045
rect 22945 18005 22955 18045
rect 22995 18005 23005 18045
rect 23045 18005 23055 18045
rect 23095 18005 23105 18045
rect 23145 18005 23155 18045
rect 23195 18005 23205 18045
rect 23245 18005 23255 18045
rect 23295 18005 23305 18045
rect 23345 18005 23355 18045
rect 23395 18005 23405 18045
rect 23445 18005 23455 18045
rect 23495 18005 23505 18045
rect 23545 18005 23555 18045
rect 23595 18005 23605 18045
rect 23645 18005 23655 18045
rect 23695 18005 23705 18045
rect 23745 18005 23755 18045
rect 23795 18005 23805 18045
rect 23845 18005 23855 18045
rect 23895 18005 23905 18045
rect 23945 18005 23955 18045
rect 23995 18005 24005 18045
rect 24045 18005 24055 18045
rect 24095 18005 24105 18045
rect 24145 18005 24155 18045
rect 24195 18005 24205 18045
rect 24245 18005 24255 18045
rect 24295 18005 24305 18045
rect 24345 18005 24355 18045
rect 24395 18005 24405 18045
rect 24445 18005 24455 18045
rect 24495 18005 24505 18045
rect 24545 18005 24555 18045
rect 24595 18005 24605 18045
rect 24645 18005 24655 18045
rect 24695 18005 24705 18045
rect 24745 18005 24755 18045
rect 24795 18005 24805 18045
rect 24845 18005 24855 18045
rect 24895 18005 24905 18045
rect 24945 18005 24955 18045
rect 24995 18005 25005 18045
rect 25045 18005 25055 18045
rect 25095 18005 25105 18045
rect 25145 18005 25155 18045
rect 25195 18005 25205 18045
rect 25245 18005 25255 18045
rect 25295 18005 25305 18045
rect 25345 18005 25355 18045
rect 25395 18005 25405 18045
rect 25445 18005 25455 18045
rect 25495 18005 25505 18045
rect 25545 18005 25555 18045
rect 25595 18005 25605 18045
rect 25645 18005 25655 18045
rect 25695 18005 25705 18045
rect 25745 18005 25755 18045
rect 25795 18005 25805 18045
rect 25845 18005 25855 18045
rect 25895 18005 25905 18045
rect 25945 18005 25955 18045
rect 25995 18005 26005 18045
rect 26045 18005 26055 18045
rect 26095 18005 26105 18045
rect 26145 18005 26155 18045
rect 26195 18005 26205 18045
rect 26245 18005 26255 18045
rect 26295 18005 26305 18045
rect 26345 18005 26355 18045
rect 26395 18005 26405 18045
rect 26445 18005 26455 18045
rect 26495 18005 26505 18045
rect 26545 18005 26555 18045
rect 26595 18005 26605 18045
rect 26645 18005 26655 18045
rect 26695 18005 26705 18045
rect 26745 18005 26755 18045
rect 26795 18005 26805 18045
rect 26845 18005 26855 18045
rect 26895 18005 26905 18045
rect 26945 18005 26955 18045
rect 26995 18005 27005 18045
rect 27045 18005 27055 18045
rect 27095 18005 27105 18045
rect 27145 18005 27155 18045
rect 27195 18005 27205 18045
rect 27245 18005 27255 18045
rect 27295 18005 27305 18045
rect 27345 18005 27355 18045
rect 27395 18005 27405 18045
rect 27445 18005 27455 18045
rect 27495 18005 27505 18045
rect 27545 18005 27555 18045
rect 27595 18005 27605 18045
rect 27645 18005 27655 18045
rect 27695 18005 27705 18045
rect 27745 18005 27755 18045
rect 27795 18005 27805 18045
rect 27845 18005 27855 18045
rect 27895 18005 27905 18045
rect 27945 18005 27955 18045
rect 27995 18005 28005 18045
rect 28045 18005 28055 18045
rect 28095 18005 28105 18045
rect 28145 18005 28155 18045
rect 28195 18005 28205 18045
rect 28245 18005 28255 18045
rect 28295 18005 28305 18045
rect 28345 18005 28355 18045
rect 28395 18005 28405 18045
rect 28445 18005 28455 18045
rect 28495 18005 28505 18045
rect 28545 18005 28555 18045
rect 28595 18005 28605 18045
rect 28645 18005 28655 18045
rect 28695 18005 28705 18045
rect 28745 18005 28755 18045
rect 28795 18005 28805 18045
rect 28845 18005 28855 18045
rect 28895 18005 28905 18045
rect 28945 18005 28955 18045
rect 28995 18005 29005 18045
rect 29045 18005 29055 18045
rect 29095 18005 29105 18045
rect 29145 18005 29155 18045
rect 29195 18005 29205 18045
rect 29245 18005 29255 18045
rect 29295 18005 29305 18045
rect 29345 18005 29355 18045
rect 29395 18005 29405 18045
rect 29445 18005 29455 18045
rect 29495 18005 29505 18045
rect 29545 18005 29555 18045
rect 29595 18005 29605 18045
rect 29645 18005 29655 18045
rect 29695 18005 29705 18045
rect 29745 18005 29755 18045
rect 29795 18005 29805 18045
rect 29845 18005 29855 18045
rect 29895 18005 29905 18045
rect 29945 18005 29955 18045
rect 29995 18005 30005 18045
rect 30045 18005 30055 18045
rect 30095 18005 30105 18045
rect 30145 18005 30155 18045
rect 30195 18005 30205 18045
rect 30245 18005 30255 18045
rect 30295 18005 30305 18045
rect 30345 18005 30355 18045
rect 30395 18005 30405 18045
rect 30445 18005 30455 18045
rect 30495 18005 30505 18045
rect 30545 18005 30555 18045
rect 30595 18005 30605 18045
rect 30645 18005 30655 18045
rect 30695 18005 30705 18045
rect 30745 18005 30755 18045
rect 30795 18005 30805 18045
rect 30845 18005 30855 18045
rect 30895 18005 30905 18045
rect 30945 18005 30955 18045
rect 30995 18005 31005 18045
rect 31045 18005 31055 18045
rect 31095 18005 31105 18045
rect 31145 18005 31155 18045
rect 31195 18005 31205 18045
rect 31245 18005 31255 18045
rect 31295 18005 31305 18045
rect 31345 18005 31355 18045
rect 31395 18005 31405 18045
rect 31445 18005 31455 18045
rect 31495 18005 31505 18045
rect 31545 18005 31555 18045
rect 31595 18005 31605 18045
rect 31645 18005 31655 18045
rect 31695 18005 31705 18045
rect 31745 18005 31755 18045
rect 31795 18005 31805 18045
rect 31845 18005 31855 18045
rect 31895 18005 31905 18045
rect 31945 18005 31955 18045
rect 31995 18005 32005 18045
rect 32045 18005 32055 18045
rect 32095 18005 32105 18045
rect 32145 18005 32155 18045
rect 32195 18005 32205 18045
rect 32245 18005 32255 18045
rect 32295 18005 32305 18045
rect 32345 18005 32355 18045
rect 32395 18005 32405 18045
rect 32445 18005 32455 18045
rect 32495 18005 32505 18045
rect 32545 18005 32555 18045
rect 32595 18005 32605 18045
rect 32645 18005 32655 18045
rect 32695 18005 32705 18045
rect 32745 18005 32755 18045
rect 32795 18005 32805 18045
rect 32845 18005 32855 18045
rect 32895 18005 32905 18045
rect 32945 18005 32955 18045
rect 32995 18005 33005 18045
rect 33045 18005 33055 18045
rect 33095 18005 33105 18045
rect 33145 18005 33155 18045
rect 33195 18005 33205 18045
rect 33245 18005 33255 18045
rect 33295 18005 33305 18045
rect 33345 18005 33355 18045
rect 33395 18005 33405 18045
rect 33445 18005 33455 18045
rect 33495 18005 33505 18045
rect 33545 18005 33555 18045
rect 33595 18005 33605 18045
rect 33645 18005 33655 18045
rect 33695 18005 33705 18045
rect 33745 18005 33755 18045
rect 33795 18005 33805 18045
rect 33845 18005 33855 18045
rect 33895 18005 33905 18045
rect 33945 18005 33955 18045
rect 33995 18005 34005 18045
rect 34045 18005 34055 18045
rect 34095 18005 34105 18045
rect 34145 18005 34155 18045
rect 34195 18005 34205 18045
rect 34245 18005 34255 18045
rect 34295 18005 34305 18045
rect 34345 18005 34355 18045
rect 34395 18005 34405 18045
rect 34445 18005 34455 18045
rect 34495 18005 34505 18045
rect 34545 18005 34555 18045
rect 34595 18005 34605 18045
rect 34645 18005 34655 18045
rect 34695 18005 34705 18045
rect 34745 18005 34755 18045
rect 34795 18005 34805 18045
rect 34845 18005 34855 18045
rect 34895 18005 34905 18045
rect 34945 18005 34955 18045
rect 34995 18005 35005 18045
rect 35045 18005 35055 18045
rect 35095 18005 35105 18045
rect 35145 18005 35155 18045
rect 35195 18005 35205 18045
rect 35245 18005 35255 18045
rect 35295 18005 35305 18045
rect 35345 18005 35355 18045
rect 35395 18005 35405 18045
rect 35445 18005 35455 18045
rect 35495 18005 35505 18045
rect 35545 18005 35555 18045
rect 35595 18005 35605 18045
rect 35645 18005 35655 18045
rect 35695 18005 35705 18045
rect 35745 18005 35755 18045
rect 35795 18005 35805 18045
rect 35845 18005 35855 18045
rect 35895 18005 35905 18045
rect 35945 18005 35955 18045
rect 35995 18005 36005 18045
rect 36045 18005 36055 18045
rect 36095 18005 36105 18045
rect 36145 18005 36155 18045
rect 36195 18005 36205 18045
rect 36245 18005 36255 18045
rect 36295 18005 36305 18045
rect 36345 18005 36355 18045
rect 36395 18005 36405 18045
rect 36445 18005 36455 18045
rect 36495 18005 36505 18045
rect 36545 18005 36555 18045
rect 36595 18005 36605 18045
rect 36645 18005 36655 18045
rect 36695 18005 36705 18045
rect 36745 18005 36755 18045
rect 36795 18005 36805 18045
rect 36845 18005 36855 18045
rect 36895 18005 36905 18045
rect 36945 18005 36955 18045
rect 36995 18005 37005 18045
rect 37045 18005 37055 18045
rect 37095 18005 37105 18045
rect 37145 18005 37155 18045
rect 37195 18005 37205 18045
rect 37245 18005 37255 18045
rect 37295 18005 37305 18045
rect 37345 18005 37355 18045
rect 37395 18005 37405 18045
rect 37445 18005 37455 18045
rect 37495 18005 37505 18045
rect 37545 18005 37555 18045
rect 37595 18005 37605 18045
rect 37645 18005 37655 18045
rect 37695 18005 37705 18045
rect 37745 18005 37755 18045
rect 37795 18005 37805 18045
rect 37845 18005 37855 18045
rect 37895 18005 37905 18045
rect 37945 18005 37955 18045
rect 37995 18005 38005 18045
rect 38045 18005 38055 18045
rect 38095 18005 38105 18045
rect 38145 18005 38155 18045
rect 38195 18005 38205 18045
rect 38245 18005 38255 18045
rect 38295 18005 38305 18045
rect 38345 18005 38355 18045
rect 38395 18005 38405 18045
rect 38445 18005 38455 18045
rect 38495 18005 38505 18045
rect 38545 18005 38555 18045
rect 38595 18005 38605 18045
rect 38645 18005 38655 18045
rect 38695 18005 38705 18045
rect 38745 18005 38755 18045
rect 38795 18005 38805 18045
rect 38845 18005 38855 18045
rect 38895 18005 38905 18045
rect 38945 18005 38955 18045
rect 38995 18005 39005 18045
rect 39045 18005 39055 18045
rect 39095 18005 39105 18045
rect 39145 18005 39155 18045
rect 39195 18005 39205 18045
rect 39245 18005 39255 18045
rect 39295 18005 39305 18045
rect 39345 18005 39355 18045
rect 39395 18005 39405 18045
rect 39445 18005 39455 18045
rect 39495 18005 39505 18045
rect 39545 18005 39555 18045
rect 39595 18005 39605 18045
rect 39645 18005 39655 18045
rect 39695 18005 39705 18045
rect 39745 18005 39750 18045
rect 0 18000 39750 18005
rect 100 17100 3200 18000
rect 3350 17100 6450 18000
rect 6600 17100 9700 18000
rect 9850 17100 12950 18000
rect 13100 17100 16200 18000
rect 16350 17100 19450 18000
rect 19600 17100 22700 18000
rect 22850 17100 25950 18000
rect 26100 17100 29200 18000
rect 29350 17100 32450 18000
rect 32600 17100 35700 18000
rect 35850 17100 38950 18000
rect 39100 17100 39750 18000
rect -2700 17045 39750 17050
rect -2700 17005 -2695 17045
rect -2655 17005 105 17045
rect 145 17005 155 17045
rect 195 17005 205 17045
rect 245 17005 255 17045
rect 295 17005 305 17045
rect 345 17005 355 17045
rect 395 17005 405 17045
rect 445 17005 455 17045
rect 495 17005 505 17045
rect 545 17005 555 17045
rect 595 17005 605 17045
rect 645 17005 655 17045
rect 695 17005 705 17045
rect 745 17005 755 17045
rect 795 17005 805 17045
rect 845 17005 855 17045
rect 895 17005 905 17045
rect 945 17005 955 17045
rect 995 17005 1005 17045
rect 1045 17005 1055 17045
rect 1095 17005 1105 17045
rect 1145 17005 1155 17045
rect 1195 17005 1205 17045
rect 1245 17005 1255 17045
rect 1295 17005 1305 17045
rect 1345 17005 1355 17045
rect 1395 17005 1405 17045
rect 1445 17005 1455 17045
rect 1495 17005 1505 17045
rect 1545 17005 1555 17045
rect 1595 17005 1605 17045
rect 1645 17005 1655 17045
rect 1695 17005 1705 17045
rect 1745 17005 1755 17045
rect 1795 17005 1805 17045
rect 1845 17005 1855 17045
rect 1895 17005 1905 17045
rect 1945 17005 1955 17045
rect 1995 17005 2005 17045
rect 2045 17005 2055 17045
rect 2095 17005 2105 17045
rect 2145 17005 2155 17045
rect 2195 17005 2205 17045
rect 2245 17005 2255 17045
rect 2295 17005 2305 17045
rect 2345 17005 2355 17045
rect 2395 17005 2405 17045
rect 2445 17005 2455 17045
rect 2495 17005 2505 17045
rect 2545 17005 2555 17045
rect 2595 17005 2605 17045
rect 2645 17005 2655 17045
rect 2695 17005 2705 17045
rect 2745 17005 2755 17045
rect 2795 17005 2805 17045
rect 2845 17005 2855 17045
rect 2895 17005 2905 17045
rect 2945 17005 2955 17045
rect 2995 17005 3005 17045
rect 3045 17005 3055 17045
rect 3095 17005 3105 17045
rect 3145 17005 3155 17045
rect 3195 17005 3205 17045
rect 3245 17005 3255 17045
rect 3295 17005 3305 17045
rect 3345 17005 3355 17045
rect 3395 17005 3405 17045
rect 3445 17005 3455 17045
rect 3495 17005 3505 17045
rect 3545 17005 3555 17045
rect 3595 17005 3605 17045
rect 3645 17005 3655 17045
rect 3695 17005 3705 17045
rect 3745 17005 3755 17045
rect 3795 17005 3805 17045
rect 3845 17005 3855 17045
rect 3895 17005 3905 17045
rect 3945 17005 3955 17045
rect 3995 17005 4005 17045
rect 4045 17005 4055 17045
rect 4095 17005 4105 17045
rect 4145 17005 4155 17045
rect 4195 17005 4205 17045
rect 4245 17005 4255 17045
rect 4295 17005 4305 17045
rect 4345 17005 4355 17045
rect 4395 17005 4405 17045
rect 4445 17005 4455 17045
rect 4495 17005 4505 17045
rect 4545 17005 4555 17045
rect 4595 17005 4605 17045
rect 4645 17005 4655 17045
rect 4695 17005 4705 17045
rect 4745 17005 4755 17045
rect 4795 17005 4805 17045
rect 4845 17005 4855 17045
rect 4895 17005 4905 17045
rect 4945 17005 4955 17045
rect 4995 17005 5005 17045
rect 5045 17005 5055 17045
rect 5095 17005 5105 17045
rect 5145 17005 5155 17045
rect 5195 17005 5205 17045
rect 5245 17005 5255 17045
rect 5295 17005 5305 17045
rect 5345 17005 5355 17045
rect 5395 17005 5405 17045
rect 5445 17005 5455 17045
rect 5495 17005 5505 17045
rect 5545 17005 5555 17045
rect 5595 17005 5605 17045
rect 5645 17005 5655 17045
rect 5695 17005 5705 17045
rect 5745 17005 5755 17045
rect 5795 17005 5805 17045
rect 5845 17005 5855 17045
rect 5895 17005 5905 17045
rect 5945 17005 5955 17045
rect 5995 17005 6005 17045
rect 6045 17005 6055 17045
rect 6095 17005 6105 17045
rect 6145 17005 6155 17045
rect 6195 17005 6205 17045
rect 6245 17005 6255 17045
rect 6295 17005 6305 17045
rect 6345 17005 6355 17045
rect 6395 17005 6405 17045
rect 6445 17005 6455 17045
rect 6495 17005 6505 17045
rect 6545 17005 6555 17045
rect 6595 17005 6605 17045
rect 6645 17005 6655 17045
rect 6695 17005 6705 17045
rect 6745 17005 6755 17045
rect 6795 17005 6805 17045
rect 6845 17005 6855 17045
rect 6895 17005 6905 17045
rect 6945 17005 6955 17045
rect 6995 17005 7005 17045
rect 7045 17005 7055 17045
rect 7095 17005 7105 17045
rect 7145 17005 7155 17045
rect 7195 17005 7205 17045
rect 7245 17005 7255 17045
rect 7295 17005 7305 17045
rect 7345 17005 7355 17045
rect 7395 17005 7405 17045
rect 7445 17005 7455 17045
rect 7495 17005 7505 17045
rect 7545 17005 7555 17045
rect 7595 17005 7605 17045
rect 7645 17005 7655 17045
rect 7695 17005 7705 17045
rect 7745 17005 7755 17045
rect 7795 17005 7805 17045
rect 7845 17005 7855 17045
rect 7895 17005 7905 17045
rect 7945 17005 7955 17045
rect 7995 17005 8005 17045
rect 8045 17005 8055 17045
rect 8095 17005 8105 17045
rect 8145 17005 8155 17045
rect 8195 17005 8205 17045
rect 8245 17005 8255 17045
rect 8295 17005 8305 17045
rect 8345 17005 8355 17045
rect 8395 17005 8405 17045
rect 8445 17005 8455 17045
rect 8495 17005 8505 17045
rect 8545 17005 8555 17045
rect 8595 17005 8605 17045
rect 8645 17005 8655 17045
rect 8695 17005 8705 17045
rect 8745 17005 8755 17045
rect 8795 17005 8805 17045
rect 8845 17005 8855 17045
rect 8895 17005 8905 17045
rect 8945 17005 8955 17045
rect 8995 17005 9005 17045
rect 9045 17005 9055 17045
rect 9095 17005 9105 17045
rect 9145 17005 9155 17045
rect 9195 17005 9205 17045
rect 9245 17005 9255 17045
rect 9295 17005 9305 17045
rect 9345 17005 9355 17045
rect 9395 17005 9405 17045
rect 9445 17005 9455 17045
rect 9495 17005 9505 17045
rect 9545 17005 9555 17045
rect 9595 17005 9605 17045
rect 9645 17005 9655 17045
rect 9695 17005 9705 17045
rect 9745 17005 9755 17045
rect 9795 17005 9805 17045
rect 9845 17005 9855 17045
rect 9895 17005 9905 17045
rect 9945 17005 9955 17045
rect 9995 17005 10005 17045
rect 10045 17005 10055 17045
rect 10095 17005 10105 17045
rect 10145 17005 10155 17045
rect 10195 17005 10205 17045
rect 10245 17005 10255 17045
rect 10295 17005 10305 17045
rect 10345 17005 10355 17045
rect 10395 17005 10405 17045
rect 10445 17005 10455 17045
rect 10495 17005 10505 17045
rect 10545 17005 10555 17045
rect 10595 17005 10605 17045
rect 10645 17005 10655 17045
rect 10695 17005 10705 17045
rect 10745 17005 10755 17045
rect 10795 17005 10805 17045
rect 10845 17005 10855 17045
rect 10895 17005 10905 17045
rect 10945 17005 10955 17045
rect 10995 17005 11005 17045
rect 11045 17005 11055 17045
rect 11095 17005 11105 17045
rect 11145 17005 11155 17045
rect 11195 17005 11205 17045
rect 11245 17005 11255 17045
rect 11295 17005 11305 17045
rect 11345 17005 11355 17045
rect 11395 17005 11405 17045
rect 11445 17005 11455 17045
rect 11495 17005 11505 17045
rect 11545 17005 11555 17045
rect 11595 17005 11605 17045
rect 11645 17005 11655 17045
rect 11695 17005 11705 17045
rect 11745 17005 11755 17045
rect 11795 17005 11805 17045
rect 11845 17005 11855 17045
rect 11895 17005 11905 17045
rect 11945 17005 11955 17045
rect 11995 17005 12005 17045
rect 12045 17005 12055 17045
rect 12095 17005 12105 17045
rect 12145 17005 12155 17045
rect 12195 17005 12205 17045
rect 12245 17005 12255 17045
rect 12295 17005 12305 17045
rect 12345 17005 12355 17045
rect 12395 17005 12405 17045
rect 12445 17005 12455 17045
rect 12495 17005 12505 17045
rect 12545 17005 12555 17045
rect 12595 17005 12605 17045
rect 12645 17005 12655 17045
rect 12695 17005 12705 17045
rect 12745 17005 12755 17045
rect 12795 17005 12805 17045
rect 12845 17005 12855 17045
rect 12895 17005 12905 17045
rect 12945 17005 12955 17045
rect 12995 17005 13005 17045
rect 13045 17005 13055 17045
rect 13095 17005 13105 17045
rect 13145 17005 13155 17045
rect 13195 17005 13205 17045
rect 13245 17005 13255 17045
rect 13295 17005 13305 17045
rect 13345 17005 13355 17045
rect 13395 17005 13405 17045
rect 13445 17005 13455 17045
rect 13495 17005 13505 17045
rect 13545 17005 13555 17045
rect 13595 17005 13605 17045
rect 13645 17005 13655 17045
rect 13695 17005 13705 17045
rect 13745 17005 13755 17045
rect 13795 17005 13805 17045
rect 13845 17005 13855 17045
rect 13895 17005 13905 17045
rect 13945 17005 13955 17045
rect 13995 17005 14005 17045
rect 14045 17005 14055 17045
rect 14095 17005 14105 17045
rect 14145 17005 14155 17045
rect 14195 17005 14205 17045
rect 14245 17005 14255 17045
rect 14295 17005 14305 17045
rect 14345 17005 14355 17045
rect 14395 17005 14405 17045
rect 14445 17005 14455 17045
rect 14495 17005 14505 17045
rect 14545 17005 14555 17045
rect 14595 17005 14605 17045
rect 14645 17005 14655 17045
rect 14695 17005 14705 17045
rect 14745 17005 14755 17045
rect 14795 17005 14805 17045
rect 14845 17005 14855 17045
rect 14895 17005 14905 17045
rect 14945 17005 14955 17045
rect 14995 17005 15005 17045
rect 15045 17005 15055 17045
rect 15095 17005 15105 17045
rect 15145 17005 15155 17045
rect 15195 17005 15205 17045
rect 15245 17005 15255 17045
rect 15295 17005 15305 17045
rect 15345 17005 15355 17045
rect 15395 17005 15405 17045
rect 15445 17005 15455 17045
rect 15495 17005 15505 17045
rect 15545 17005 15555 17045
rect 15595 17005 15605 17045
rect 15645 17005 15655 17045
rect 15695 17005 15705 17045
rect 15745 17005 15755 17045
rect 15795 17005 15805 17045
rect 15845 17005 15855 17045
rect 15895 17005 15905 17045
rect 15945 17005 15955 17045
rect 15995 17005 16005 17045
rect 16045 17005 16055 17045
rect 16095 17005 16105 17045
rect 16145 17005 16155 17045
rect 16195 17005 16205 17045
rect 16245 17005 16255 17045
rect 16295 17005 16305 17045
rect 16345 17005 16355 17045
rect 16395 17005 16405 17045
rect 16445 17005 16455 17045
rect 16495 17005 16505 17045
rect 16545 17005 16555 17045
rect 16595 17005 16605 17045
rect 16645 17005 16655 17045
rect 16695 17005 16705 17045
rect 16745 17005 16755 17045
rect 16795 17005 16805 17045
rect 16845 17005 16855 17045
rect 16895 17005 16905 17045
rect 16945 17005 16955 17045
rect 16995 17005 17005 17045
rect 17045 17005 17055 17045
rect 17095 17005 17105 17045
rect 17145 17005 17155 17045
rect 17195 17005 17205 17045
rect 17245 17005 17255 17045
rect 17295 17005 17305 17045
rect 17345 17005 17355 17045
rect 17395 17005 17405 17045
rect 17445 17005 17455 17045
rect 17495 17005 17505 17045
rect 17545 17005 17555 17045
rect 17595 17005 17605 17045
rect 17645 17005 17655 17045
rect 17695 17005 17705 17045
rect 17745 17005 17755 17045
rect 17795 17005 17805 17045
rect 17845 17005 17855 17045
rect 17895 17005 17905 17045
rect 17945 17005 17955 17045
rect 17995 17005 18005 17045
rect 18045 17005 18055 17045
rect 18095 17005 18105 17045
rect 18145 17005 18155 17045
rect 18195 17005 18205 17045
rect 18245 17005 18255 17045
rect 18295 17005 18305 17045
rect 18345 17005 18355 17045
rect 18395 17005 18405 17045
rect 18445 17005 18455 17045
rect 18495 17005 18505 17045
rect 18545 17005 18555 17045
rect 18595 17005 18605 17045
rect 18645 17005 18655 17045
rect 18695 17005 18705 17045
rect 18745 17005 18755 17045
rect 18795 17005 18805 17045
rect 18845 17005 18855 17045
rect 18895 17005 18905 17045
rect 18945 17005 18955 17045
rect 18995 17005 19005 17045
rect 19045 17005 19055 17045
rect 19095 17005 19105 17045
rect 19145 17005 19155 17045
rect 19195 17005 19205 17045
rect 19245 17005 19255 17045
rect 19295 17005 19305 17045
rect 19345 17005 19355 17045
rect 19395 17005 19405 17045
rect 19445 17005 19455 17045
rect 19495 17005 19505 17045
rect 19545 17005 19555 17045
rect 19595 17005 19605 17045
rect 19645 17005 19655 17045
rect 19695 17005 19705 17045
rect 19745 17005 19755 17045
rect 19795 17005 19805 17045
rect 19845 17005 19855 17045
rect 19895 17005 19905 17045
rect 19945 17005 19955 17045
rect 19995 17005 20005 17045
rect 20045 17005 20055 17045
rect 20095 17005 20105 17045
rect 20145 17005 20155 17045
rect 20195 17005 20205 17045
rect 20245 17005 20255 17045
rect 20295 17005 20305 17045
rect 20345 17005 20355 17045
rect 20395 17005 20405 17045
rect 20445 17005 20455 17045
rect 20495 17005 20505 17045
rect 20545 17005 20555 17045
rect 20595 17005 20605 17045
rect 20645 17005 20655 17045
rect 20695 17005 20705 17045
rect 20745 17005 20755 17045
rect 20795 17005 20805 17045
rect 20845 17005 20855 17045
rect 20895 17005 20905 17045
rect 20945 17005 20955 17045
rect 20995 17005 21005 17045
rect 21045 17005 21055 17045
rect 21095 17005 21105 17045
rect 21145 17005 21155 17045
rect 21195 17005 21205 17045
rect 21245 17005 21255 17045
rect 21295 17005 21305 17045
rect 21345 17005 21355 17045
rect 21395 17005 21405 17045
rect 21445 17005 21455 17045
rect 21495 17005 21505 17045
rect 21545 17005 21555 17045
rect 21595 17005 21605 17045
rect 21645 17005 21655 17045
rect 21695 17005 21705 17045
rect 21745 17005 21755 17045
rect 21795 17005 21805 17045
rect 21845 17005 21855 17045
rect 21895 17005 21905 17045
rect 21945 17005 21955 17045
rect 21995 17005 22005 17045
rect 22045 17005 22055 17045
rect 22095 17005 22105 17045
rect 22145 17005 22155 17045
rect 22195 17005 22205 17045
rect 22245 17005 22255 17045
rect 22295 17005 22305 17045
rect 22345 17005 22355 17045
rect 22395 17005 22405 17045
rect 22445 17005 22455 17045
rect 22495 17005 22505 17045
rect 22545 17005 22555 17045
rect 22595 17005 22605 17045
rect 22645 17005 22655 17045
rect 22695 17005 22705 17045
rect 22745 17005 22755 17045
rect 22795 17005 22805 17045
rect 22845 17005 22855 17045
rect 22895 17005 22905 17045
rect 22945 17005 22955 17045
rect 22995 17005 23005 17045
rect 23045 17005 23055 17045
rect 23095 17005 23105 17045
rect 23145 17005 23155 17045
rect 23195 17005 23205 17045
rect 23245 17005 23255 17045
rect 23295 17005 23305 17045
rect 23345 17005 23355 17045
rect 23395 17005 23405 17045
rect 23445 17005 23455 17045
rect 23495 17005 23505 17045
rect 23545 17005 23555 17045
rect 23595 17005 23605 17045
rect 23645 17005 23655 17045
rect 23695 17005 23705 17045
rect 23745 17005 23755 17045
rect 23795 17005 23805 17045
rect 23845 17005 23855 17045
rect 23895 17005 23905 17045
rect 23945 17005 23955 17045
rect 23995 17005 24005 17045
rect 24045 17005 24055 17045
rect 24095 17005 24105 17045
rect 24145 17005 24155 17045
rect 24195 17005 24205 17045
rect 24245 17005 24255 17045
rect 24295 17005 24305 17045
rect 24345 17005 24355 17045
rect 24395 17005 24405 17045
rect 24445 17005 24455 17045
rect 24495 17005 24505 17045
rect 24545 17005 24555 17045
rect 24595 17005 24605 17045
rect 24645 17005 24655 17045
rect 24695 17005 24705 17045
rect 24745 17005 24755 17045
rect 24795 17005 24805 17045
rect 24845 17005 24855 17045
rect 24895 17005 24905 17045
rect 24945 17005 24955 17045
rect 24995 17005 25005 17045
rect 25045 17005 25055 17045
rect 25095 17005 25105 17045
rect 25145 17005 25155 17045
rect 25195 17005 25205 17045
rect 25245 17005 25255 17045
rect 25295 17005 25305 17045
rect 25345 17005 25355 17045
rect 25395 17005 25405 17045
rect 25445 17005 25455 17045
rect 25495 17005 25505 17045
rect 25545 17005 25555 17045
rect 25595 17005 25605 17045
rect 25645 17005 25655 17045
rect 25695 17005 25705 17045
rect 25745 17005 25755 17045
rect 25795 17005 25805 17045
rect 25845 17005 25855 17045
rect 25895 17005 25905 17045
rect 25945 17005 25955 17045
rect 25995 17005 26005 17045
rect 26045 17005 26055 17045
rect 26095 17005 26105 17045
rect 26145 17005 26155 17045
rect 26195 17005 26205 17045
rect 26245 17005 26255 17045
rect 26295 17005 26305 17045
rect 26345 17005 26355 17045
rect 26395 17005 26405 17045
rect 26445 17005 26455 17045
rect 26495 17005 26505 17045
rect 26545 17005 26555 17045
rect 26595 17005 26605 17045
rect 26645 17005 26655 17045
rect 26695 17005 26705 17045
rect 26745 17005 26755 17045
rect 26795 17005 26805 17045
rect 26845 17005 26855 17045
rect 26895 17005 26905 17045
rect 26945 17005 26955 17045
rect 26995 17005 27005 17045
rect 27045 17005 27055 17045
rect 27095 17005 27105 17045
rect 27145 17005 27155 17045
rect 27195 17005 27205 17045
rect 27245 17005 27255 17045
rect 27295 17005 27305 17045
rect 27345 17005 27355 17045
rect 27395 17005 27405 17045
rect 27445 17005 27455 17045
rect 27495 17005 27505 17045
rect 27545 17005 27555 17045
rect 27595 17005 27605 17045
rect 27645 17005 27655 17045
rect 27695 17005 27705 17045
rect 27745 17005 27755 17045
rect 27795 17005 27805 17045
rect 27845 17005 27855 17045
rect 27895 17005 27905 17045
rect 27945 17005 27955 17045
rect 27995 17005 28005 17045
rect 28045 17005 28055 17045
rect 28095 17005 28105 17045
rect 28145 17005 28155 17045
rect 28195 17005 28205 17045
rect 28245 17005 28255 17045
rect 28295 17005 28305 17045
rect 28345 17005 28355 17045
rect 28395 17005 28405 17045
rect 28445 17005 28455 17045
rect 28495 17005 28505 17045
rect 28545 17005 28555 17045
rect 28595 17005 28605 17045
rect 28645 17005 28655 17045
rect 28695 17005 28705 17045
rect 28745 17005 28755 17045
rect 28795 17005 28805 17045
rect 28845 17005 28855 17045
rect 28895 17005 28905 17045
rect 28945 17005 28955 17045
rect 28995 17005 29005 17045
rect 29045 17005 29055 17045
rect 29095 17005 29105 17045
rect 29145 17005 29155 17045
rect 29195 17005 29205 17045
rect 29245 17005 29255 17045
rect 29295 17005 29305 17045
rect 29345 17005 29355 17045
rect 29395 17005 29405 17045
rect 29445 17005 29455 17045
rect 29495 17005 29505 17045
rect 29545 17005 29555 17045
rect 29595 17005 29605 17045
rect 29645 17005 29655 17045
rect 29695 17005 29705 17045
rect 29745 17005 29755 17045
rect 29795 17005 29805 17045
rect 29845 17005 29855 17045
rect 29895 17005 29905 17045
rect 29945 17005 29955 17045
rect 29995 17005 30005 17045
rect 30045 17005 30055 17045
rect 30095 17005 30105 17045
rect 30145 17005 30155 17045
rect 30195 17005 30205 17045
rect 30245 17005 30255 17045
rect 30295 17005 30305 17045
rect 30345 17005 30355 17045
rect 30395 17005 30405 17045
rect 30445 17005 30455 17045
rect 30495 17005 30505 17045
rect 30545 17005 30555 17045
rect 30595 17005 30605 17045
rect 30645 17005 30655 17045
rect 30695 17005 30705 17045
rect 30745 17005 30755 17045
rect 30795 17005 30805 17045
rect 30845 17005 30855 17045
rect 30895 17005 30905 17045
rect 30945 17005 30955 17045
rect 30995 17005 31005 17045
rect 31045 17005 31055 17045
rect 31095 17005 31105 17045
rect 31145 17005 31155 17045
rect 31195 17005 31205 17045
rect 31245 17005 31255 17045
rect 31295 17005 31305 17045
rect 31345 17005 31355 17045
rect 31395 17005 31405 17045
rect 31445 17005 31455 17045
rect 31495 17005 31505 17045
rect 31545 17005 31555 17045
rect 31595 17005 31605 17045
rect 31645 17005 31655 17045
rect 31695 17005 31705 17045
rect 31745 17005 31755 17045
rect 31795 17005 31805 17045
rect 31845 17005 31855 17045
rect 31895 17005 31905 17045
rect 31945 17005 31955 17045
rect 31995 17005 32005 17045
rect 32045 17005 32055 17045
rect 32095 17005 32105 17045
rect 32145 17005 32155 17045
rect 32195 17005 32205 17045
rect 32245 17005 32255 17045
rect 32295 17005 32305 17045
rect 32345 17005 32355 17045
rect 32395 17005 32405 17045
rect 32445 17005 32455 17045
rect 32495 17005 32505 17045
rect 32545 17005 32555 17045
rect 32595 17005 32605 17045
rect 32645 17005 32655 17045
rect 32695 17005 32705 17045
rect 32745 17005 32755 17045
rect 32795 17005 32805 17045
rect 32845 17005 32855 17045
rect 32895 17005 32905 17045
rect 32945 17005 32955 17045
rect 32995 17005 33005 17045
rect 33045 17005 33055 17045
rect 33095 17005 33105 17045
rect 33145 17005 33155 17045
rect 33195 17005 33205 17045
rect 33245 17005 33255 17045
rect 33295 17005 33305 17045
rect 33345 17005 33355 17045
rect 33395 17005 33405 17045
rect 33445 17005 33455 17045
rect 33495 17005 33505 17045
rect 33545 17005 33555 17045
rect 33595 17005 33605 17045
rect 33645 17005 33655 17045
rect 33695 17005 33705 17045
rect 33745 17005 33755 17045
rect 33795 17005 33805 17045
rect 33845 17005 33855 17045
rect 33895 17005 33905 17045
rect 33945 17005 33955 17045
rect 33995 17005 34005 17045
rect 34045 17005 34055 17045
rect 34095 17005 34105 17045
rect 34145 17005 34155 17045
rect 34195 17005 34205 17045
rect 34245 17005 34255 17045
rect 34295 17005 34305 17045
rect 34345 17005 34355 17045
rect 34395 17005 34405 17045
rect 34445 17005 34455 17045
rect 34495 17005 34505 17045
rect 34545 17005 34555 17045
rect 34595 17005 34605 17045
rect 34645 17005 34655 17045
rect 34695 17005 34705 17045
rect 34745 17005 34755 17045
rect 34795 17005 34805 17045
rect 34845 17005 34855 17045
rect 34895 17005 34905 17045
rect 34945 17005 34955 17045
rect 34995 17005 35005 17045
rect 35045 17005 35055 17045
rect 35095 17005 35105 17045
rect 35145 17005 35155 17045
rect 35195 17005 35205 17045
rect 35245 17005 35255 17045
rect 35295 17005 35305 17045
rect 35345 17005 35355 17045
rect 35395 17005 35405 17045
rect 35445 17005 35455 17045
rect 35495 17005 35505 17045
rect 35545 17005 35555 17045
rect 35595 17005 35605 17045
rect 35645 17005 35655 17045
rect 35695 17005 35705 17045
rect 35745 17005 35755 17045
rect 35795 17005 35805 17045
rect 35845 17005 35855 17045
rect 35895 17005 35905 17045
rect 35945 17005 35955 17045
rect 35995 17005 36005 17045
rect 36045 17005 36055 17045
rect 36095 17005 36105 17045
rect 36145 17005 36155 17045
rect 36195 17005 36205 17045
rect 36245 17005 36255 17045
rect 36295 17005 36305 17045
rect 36345 17005 36355 17045
rect 36395 17005 36405 17045
rect 36445 17005 36455 17045
rect 36495 17005 36505 17045
rect 36545 17005 36555 17045
rect 36595 17005 36605 17045
rect 36645 17005 36655 17045
rect 36695 17005 36705 17045
rect 36745 17005 36755 17045
rect 36795 17005 36805 17045
rect 36845 17005 36855 17045
rect 36895 17005 36905 17045
rect 36945 17005 36955 17045
rect 36995 17005 37005 17045
rect 37045 17005 37055 17045
rect 37095 17005 37105 17045
rect 37145 17005 37155 17045
rect 37195 17005 37205 17045
rect 37245 17005 37255 17045
rect 37295 17005 37305 17045
rect 37345 17005 37355 17045
rect 37395 17005 37405 17045
rect 37445 17005 37455 17045
rect 37495 17005 37505 17045
rect 37545 17005 37555 17045
rect 37595 17005 37605 17045
rect 37645 17005 37655 17045
rect 37695 17005 37705 17045
rect 37745 17005 37755 17045
rect 37795 17005 37805 17045
rect 37845 17005 37855 17045
rect 37895 17005 37905 17045
rect 37945 17005 37955 17045
rect 37995 17005 38005 17045
rect 38045 17005 38055 17045
rect 38095 17005 38105 17045
rect 38145 17005 38155 17045
rect 38195 17005 38205 17045
rect 38245 17005 38255 17045
rect 38295 17005 38305 17045
rect 38345 17005 38355 17045
rect 38395 17005 38405 17045
rect 38445 17005 38455 17045
rect 38495 17005 38505 17045
rect 38545 17005 38555 17045
rect 38595 17005 38605 17045
rect 38645 17005 38655 17045
rect 38695 17005 38705 17045
rect 38745 17005 38755 17045
rect 38795 17005 38805 17045
rect 38845 17005 38855 17045
rect 38895 17005 38905 17045
rect 38945 17005 38955 17045
rect 38995 17005 39005 17045
rect 39045 17005 39055 17045
rect 39095 17005 39105 17045
rect 39145 17005 39155 17045
rect 39195 17005 39205 17045
rect 39245 17005 39255 17045
rect 39295 17005 39305 17045
rect 39345 17005 39355 17045
rect 39395 17005 39405 17045
rect 39445 17005 39455 17045
rect 39495 17005 39505 17045
rect 39545 17005 39555 17045
rect 39595 17005 39605 17045
rect 39645 17005 39655 17045
rect 39695 17005 39705 17045
rect 39745 17005 39750 17045
rect -2700 17000 39750 17005
rect -3500 16945 -50 16950
rect -3500 16905 -3495 16945
rect -3455 16905 -3295 16945
rect -3255 16905 -3095 16945
rect -3055 16905 -1595 16945
rect -1555 16905 -1195 16945
rect -1155 16905 -1095 16945
rect -1055 16905 -995 16945
rect -955 16905 -895 16945
rect -855 16905 -795 16945
rect -755 16905 -695 16945
rect -655 16905 -595 16945
rect -555 16905 -495 16945
rect -455 16905 -395 16945
rect -355 16905 -295 16945
rect -255 16905 -195 16945
rect -155 16905 -95 16945
rect -55 16905 -50 16945
rect -3500 16900 -50 16905
rect 0 16945 40900 16950
rect 0 16905 5 16945
rect 45 16905 55 16945
rect 95 16905 105 16945
rect 145 16905 155 16945
rect 195 16905 205 16945
rect 245 16905 255 16945
rect 295 16905 305 16945
rect 345 16905 355 16945
rect 395 16905 405 16945
rect 445 16905 455 16945
rect 495 16905 505 16945
rect 545 16905 555 16945
rect 595 16905 605 16945
rect 645 16905 655 16945
rect 695 16905 705 16945
rect 745 16905 755 16945
rect 795 16905 805 16945
rect 845 16905 855 16945
rect 895 16905 905 16945
rect 945 16905 955 16945
rect 995 16905 1005 16945
rect 1045 16905 1055 16945
rect 1095 16905 1105 16945
rect 1145 16905 1155 16945
rect 1195 16905 1205 16945
rect 1245 16905 1255 16945
rect 1295 16905 1305 16945
rect 1345 16905 1355 16945
rect 1395 16905 1405 16945
rect 1445 16905 1455 16945
rect 1495 16905 1505 16945
rect 1545 16905 1555 16945
rect 1595 16905 1605 16945
rect 1645 16905 1655 16945
rect 1695 16905 1705 16945
rect 1745 16905 1755 16945
rect 1795 16905 1805 16945
rect 1845 16905 1855 16945
rect 1895 16905 1905 16945
rect 1945 16905 1955 16945
rect 1995 16905 2005 16945
rect 2045 16905 2055 16945
rect 2095 16905 2105 16945
rect 2145 16905 2155 16945
rect 2195 16905 2205 16945
rect 2245 16905 2255 16945
rect 2295 16905 2305 16945
rect 2345 16905 2355 16945
rect 2395 16905 2405 16945
rect 2445 16905 2455 16945
rect 2495 16905 2505 16945
rect 2545 16905 2555 16945
rect 2595 16905 2605 16945
rect 2645 16905 2655 16945
rect 2695 16905 2705 16945
rect 2745 16905 2755 16945
rect 2795 16905 2805 16945
rect 2845 16905 2855 16945
rect 2895 16905 2905 16945
rect 2945 16905 2955 16945
rect 2995 16905 3005 16945
rect 3045 16905 3055 16945
rect 3095 16905 3105 16945
rect 3145 16905 3155 16945
rect 3195 16905 3205 16945
rect 3245 16905 3255 16945
rect 3295 16905 3305 16945
rect 3345 16905 3355 16945
rect 3395 16905 3405 16945
rect 3445 16905 3455 16945
rect 3495 16905 3505 16945
rect 3545 16905 3555 16945
rect 3595 16905 3605 16945
rect 3645 16905 3655 16945
rect 3695 16905 3705 16945
rect 3745 16905 3755 16945
rect 3795 16905 3805 16945
rect 3845 16905 3855 16945
rect 3895 16905 3905 16945
rect 3945 16905 3955 16945
rect 3995 16905 4005 16945
rect 4045 16905 4055 16945
rect 4095 16905 4105 16945
rect 4145 16905 4155 16945
rect 4195 16905 4205 16945
rect 4245 16905 4255 16945
rect 4295 16905 4305 16945
rect 4345 16905 4355 16945
rect 4395 16905 4405 16945
rect 4445 16905 4455 16945
rect 4495 16905 4505 16945
rect 4545 16905 4555 16945
rect 4595 16905 4605 16945
rect 4645 16905 4655 16945
rect 4695 16905 4705 16945
rect 4745 16905 4755 16945
rect 4795 16905 4805 16945
rect 4845 16905 4855 16945
rect 4895 16905 4905 16945
rect 4945 16905 4955 16945
rect 4995 16905 5005 16945
rect 5045 16905 5055 16945
rect 5095 16905 5105 16945
rect 5145 16905 5155 16945
rect 5195 16905 5205 16945
rect 5245 16905 5255 16945
rect 5295 16905 5305 16945
rect 5345 16905 5355 16945
rect 5395 16905 5405 16945
rect 5445 16905 5455 16945
rect 5495 16905 5505 16945
rect 5545 16905 5555 16945
rect 5595 16905 5605 16945
rect 5645 16905 5655 16945
rect 5695 16905 5705 16945
rect 5745 16905 5755 16945
rect 5795 16905 5805 16945
rect 5845 16905 5855 16945
rect 5895 16905 5905 16945
rect 5945 16905 5955 16945
rect 5995 16905 6005 16945
rect 6045 16905 6055 16945
rect 6095 16905 6105 16945
rect 6145 16905 6155 16945
rect 6195 16905 6205 16945
rect 6245 16905 6255 16945
rect 6295 16905 6305 16945
rect 6345 16905 6355 16945
rect 6395 16905 6405 16945
rect 6445 16905 6455 16945
rect 6495 16905 6505 16945
rect 6545 16905 6555 16945
rect 6595 16905 6605 16945
rect 6645 16905 6655 16945
rect 6695 16905 6705 16945
rect 6745 16905 6755 16945
rect 6795 16905 6805 16945
rect 6845 16905 6855 16945
rect 6895 16905 6905 16945
rect 6945 16905 6955 16945
rect 6995 16905 7005 16945
rect 7045 16905 7055 16945
rect 7095 16905 7105 16945
rect 7145 16905 7155 16945
rect 7195 16905 7205 16945
rect 7245 16905 7255 16945
rect 7295 16905 7305 16945
rect 7345 16905 7355 16945
rect 7395 16905 7405 16945
rect 7445 16905 7455 16945
rect 7495 16905 7505 16945
rect 7545 16905 7555 16945
rect 7595 16905 7605 16945
rect 7645 16905 7655 16945
rect 7695 16905 7705 16945
rect 7745 16905 7755 16945
rect 7795 16905 7805 16945
rect 7845 16905 7855 16945
rect 7895 16905 7905 16945
rect 7945 16905 7955 16945
rect 7995 16905 8005 16945
rect 8045 16905 8055 16945
rect 8095 16905 8105 16945
rect 8145 16905 8155 16945
rect 8195 16905 8205 16945
rect 8245 16905 8255 16945
rect 8295 16905 8305 16945
rect 8345 16905 8355 16945
rect 8395 16905 8405 16945
rect 8445 16905 8455 16945
rect 8495 16905 8505 16945
rect 8545 16905 8555 16945
rect 8595 16905 8605 16945
rect 8645 16905 8655 16945
rect 8695 16905 8705 16945
rect 8745 16905 8755 16945
rect 8795 16905 8805 16945
rect 8845 16905 8855 16945
rect 8895 16905 8905 16945
rect 8945 16905 8955 16945
rect 8995 16905 9005 16945
rect 9045 16905 9055 16945
rect 9095 16905 9105 16945
rect 9145 16905 9155 16945
rect 9195 16905 9205 16945
rect 9245 16905 9255 16945
rect 9295 16905 9305 16945
rect 9345 16905 9355 16945
rect 9395 16905 9405 16945
rect 9445 16905 9455 16945
rect 9495 16905 9505 16945
rect 9545 16905 9555 16945
rect 9595 16905 9605 16945
rect 9645 16905 9655 16945
rect 9695 16905 9705 16945
rect 9745 16905 9755 16945
rect 9795 16905 9805 16945
rect 9845 16905 9855 16945
rect 9895 16905 9905 16945
rect 9945 16905 9955 16945
rect 9995 16905 10005 16945
rect 10045 16905 10055 16945
rect 10095 16905 10105 16945
rect 10145 16905 10155 16945
rect 10195 16905 10205 16945
rect 10245 16905 10255 16945
rect 10295 16905 10305 16945
rect 10345 16905 10355 16945
rect 10395 16905 10405 16945
rect 10445 16905 10455 16945
rect 10495 16905 10505 16945
rect 10545 16905 10555 16945
rect 10595 16905 10605 16945
rect 10645 16905 10655 16945
rect 10695 16905 10705 16945
rect 10745 16905 10755 16945
rect 10795 16905 10805 16945
rect 10845 16905 10855 16945
rect 10895 16905 10905 16945
rect 10945 16905 10955 16945
rect 10995 16905 11005 16945
rect 11045 16905 11055 16945
rect 11095 16905 11105 16945
rect 11145 16905 11155 16945
rect 11195 16905 11205 16945
rect 11245 16905 11255 16945
rect 11295 16905 11305 16945
rect 11345 16905 11355 16945
rect 11395 16905 11405 16945
rect 11445 16905 11455 16945
rect 11495 16905 11505 16945
rect 11545 16905 11555 16945
rect 11595 16905 11605 16945
rect 11645 16905 11655 16945
rect 11695 16905 11705 16945
rect 11745 16905 11755 16945
rect 11795 16905 11805 16945
rect 11845 16905 11855 16945
rect 11895 16905 11905 16945
rect 11945 16905 11955 16945
rect 11995 16905 12005 16945
rect 12045 16905 12055 16945
rect 12095 16905 12105 16945
rect 12145 16905 12155 16945
rect 12195 16905 12205 16945
rect 12245 16905 12255 16945
rect 12295 16905 12305 16945
rect 12345 16905 12355 16945
rect 12395 16905 12405 16945
rect 12445 16905 12455 16945
rect 12495 16905 12505 16945
rect 12545 16905 12555 16945
rect 12595 16905 12605 16945
rect 12645 16905 12655 16945
rect 12695 16905 12705 16945
rect 12745 16905 12755 16945
rect 12795 16905 12805 16945
rect 12845 16905 12855 16945
rect 12895 16905 12905 16945
rect 12945 16905 12955 16945
rect 12995 16905 13005 16945
rect 13045 16905 13055 16945
rect 13095 16905 13105 16945
rect 13145 16905 13155 16945
rect 13195 16905 13205 16945
rect 13245 16905 13255 16945
rect 13295 16905 13305 16945
rect 13345 16905 13355 16945
rect 13395 16905 13405 16945
rect 13445 16905 13455 16945
rect 13495 16905 13505 16945
rect 13545 16905 13555 16945
rect 13595 16905 13605 16945
rect 13645 16905 13655 16945
rect 13695 16905 13705 16945
rect 13745 16905 13755 16945
rect 13795 16905 13805 16945
rect 13845 16905 13855 16945
rect 13895 16905 13905 16945
rect 13945 16905 13955 16945
rect 13995 16905 14005 16945
rect 14045 16905 14055 16945
rect 14095 16905 14105 16945
rect 14145 16905 14155 16945
rect 14195 16905 14205 16945
rect 14245 16905 14255 16945
rect 14295 16905 14305 16945
rect 14345 16905 14355 16945
rect 14395 16905 14405 16945
rect 14445 16905 14455 16945
rect 14495 16905 14505 16945
rect 14545 16905 14555 16945
rect 14595 16905 14605 16945
rect 14645 16905 14655 16945
rect 14695 16905 14705 16945
rect 14745 16905 14755 16945
rect 14795 16905 14805 16945
rect 14845 16905 14855 16945
rect 14895 16905 14905 16945
rect 14945 16905 14955 16945
rect 14995 16905 15005 16945
rect 15045 16905 15055 16945
rect 15095 16905 15105 16945
rect 15145 16905 15155 16945
rect 15195 16905 15205 16945
rect 15245 16905 15255 16945
rect 15295 16905 15305 16945
rect 15345 16905 15355 16945
rect 15395 16905 15405 16945
rect 15445 16905 15455 16945
rect 15495 16905 15505 16945
rect 15545 16905 15555 16945
rect 15595 16905 15605 16945
rect 15645 16905 15655 16945
rect 15695 16905 15705 16945
rect 15745 16905 15755 16945
rect 15795 16905 15805 16945
rect 15845 16905 15855 16945
rect 15895 16905 15905 16945
rect 15945 16905 15955 16945
rect 15995 16905 16005 16945
rect 16045 16905 16055 16945
rect 16095 16905 16105 16945
rect 16145 16905 16155 16945
rect 16195 16905 16205 16945
rect 16245 16905 16255 16945
rect 16295 16905 16305 16945
rect 16345 16905 16355 16945
rect 16395 16905 16405 16945
rect 16445 16905 16455 16945
rect 16495 16905 16505 16945
rect 16545 16905 16555 16945
rect 16595 16905 16605 16945
rect 16645 16905 16655 16945
rect 16695 16905 16705 16945
rect 16745 16905 16755 16945
rect 16795 16905 16805 16945
rect 16845 16905 16855 16945
rect 16895 16905 16905 16945
rect 16945 16905 16955 16945
rect 16995 16905 17005 16945
rect 17045 16905 17055 16945
rect 17095 16905 17105 16945
rect 17145 16905 17155 16945
rect 17195 16905 17205 16945
rect 17245 16905 17255 16945
rect 17295 16905 17305 16945
rect 17345 16905 17355 16945
rect 17395 16905 17405 16945
rect 17445 16905 17455 16945
rect 17495 16905 17505 16945
rect 17545 16905 17555 16945
rect 17595 16905 17605 16945
rect 17645 16905 17655 16945
rect 17695 16905 17705 16945
rect 17745 16905 17755 16945
rect 17795 16905 17805 16945
rect 17845 16905 17855 16945
rect 17895 16905 17905 16945
rect 17945 16905 17955 16945
rect 17995 16905 18005 16945
rect 18045 16905 18055 16945
rect 18095 16905 18105 16945
rect 18145 16905 18155 16945
rect 18195 16905 18205 16945
rect 18245 16905 18255 16945
rect 18295 16905 18305 16945
rect 18345 16905 18355 16945
rect 18395 16905 18405 16945
rect 18445 16905 18455 16945
rect 18495 16905 18505 16945
rect 18545 16905 18555 16945
rect 18595 16905 18605 16945
rect 18645 16905 18655 16945
rect 18695 16905 18705 16945
rect 18745 16905 18755 16945
rect 18795 16905 18805 16945
rect 18845 16905 18855 16945
rect 18895 16905 18905 16945
rect 18945 16905 18955 16945
rect 18995 16905 19005 16945
rect 19045 16905 19055 16945
rect 19095 16905 19105 16945
rect 19145 16905 19155 16945
rect 19195 16905 19205 16945
rect 19245 16905 19255 16945
rect 19295 16905 19305 16945
rect 19345 16905 19355 16945
rect 19395 16905 19405 16945
rect 19445 16905 19455 16945
rect 19495 16905 19505 16945
rect 19545 16905 19555 16945
rect 19595 16905 19605 16945
rect 19645 16905 19655 16945
rect 19695 16905 19705 16945
rect 19745 16905 19755 16945
rect 19795 16905 19805 16945
rect 19845 16905 19855 16945
rect 19895 16905 19905 16945
rect 19945 16905 19955 16945
rect 19995 16905 20005 16945
rect 20045 16905 20055 16945
rect 20095 16905 20105 16945
rect 20145 16905 20155 16945
rect 20195 16905 20205 16945
rect 20245 16905 20255 16945
rect 20295 16905 20305 16945
rect 20345 16905 20355 16945
rect 20395 16905 20405 16945
rect 20445 16905 20455 16945
rect 20495 16905 20505 16945
rect 20545 16905 20555 16945
rect 20595 16905 20605 16945
rect 20645 16905 20655 16945
rect 20695 16905 20705 16945
rect 20745 16905 20755 16945
rect 20795 16905 20805 16945
rect 20845 16905 20855 16945
rect 20895 16905 20905 16945
rect 20945 16905 20955 16945
rect 20995 16905 21005 16945
rect 21045 16905 21055 16945
rect 21095 16905 21105 16945
rect 21145 16905 21155 16945
rect 21195 16905 21205 16945
rect 21245 16905 21255 16945
rect 21295 16905 21305 16945
rect 21345 16905 21355 16945
rect 21395 16905 21405 16945
rect 21445 16905 21455 16945
rect 21495 16905 21505 16945
rect 21545 16905 21555 16945
rect 21595 16905 21605 16945
rect 21645 16905 21655 16945
rect 21695 16905 21705 16945
rect 21745 16905 21755 16945
rect 21795 16905 21805 16945
rect 21845 16905 21855 16945
rect 21895 16905 21905 16945
rect 21945 16905 21955 16945
rect 21995 16905 22005 16945
rect 22045 16905 22055 16945
rect 22095 16905 22105 16945
rect 22145 16905 22155 16945
rect 22195 16905 22205 16945
rect 22245 16905 22255 16945
rect 22295 16905 22305 16945
rect 22345 16905 22355 16945
rect 22395 16905 22405 16945
rect 22445 16905 22455 16945
rect 22495 16905 22505 16945
rect 22545 16905 22555 16945
rect 22595 16905 22605 16945
rect 22645 16905 22655 16945
rect 22695 16905 22705 16945
rect 22745 16905 22755 16945
rect 22795 16905 22805 16945
rect 22845 16905 22855 16945
rect 22895 16905 22905 16945
rect 22945 16905 22955 16945
rect 22995 16905 23005 16945
rect 23045 16905 23055 16945
rect 23095 16905 23105 16945
rect 23145 16905 23155 16945
rect 23195 16905 23205 16945
rect 23245 16905 23255 16945
rect 23295 16905 23305 16945
rect 23345 16905 23355 16945
rect 23395 16905 23405 16945
rect 23445 16905 23455 16945
rect 23495 16905 23505 16945
rect 23545 16905 23555 16945
rect 23595 16905 23605 16945
rect 23645 16905 23655 16945
rect 23695 16905 23705 16945
rect 23745 16905 23755 16945
rect 23795 16905 23805 16945
rect 23845 16905 23855 16945
rect 23895 16905 23905 16945
rect 23945 16905 23955 16945
rect 23995 16905 24005 16945
rect 24045 16905 24055 16945
rect 24095 16905 24105 16945
rect 24145 16905 24155 16945
rect 24195 16905 24205 16945
rect 24245 16905 24255 16945
rect 24295 16905 24305 16945
rect 24345 16905 24355 16945
rect 24395 16905 24405 16945
rect 24445 16905 24455 16945
rect 24495 16905 24505 16945
rect 24545 16905 24555 16945
rect 24595 16905 24605 16945
rect 24645 16905 24655 16945
rect 24695 16905 24705 16945
rect 24745 16905 24755 16945
rect 24795 16905 24805 16945
rect 24845 16905 24855 16945
rect 24895 16905 24905 16945
rect 24945 16905 24955 16945
rect 24995 16905 25005 16945
rect 25045 16905 25055 16945
rect 25095 16905 25105 16945
rect 25145 16905 25155 16945
rect 25195 16905 25205 16945
rect 25245 16905 25255 16945
rect 25295 16905 25305 16945
rect 25345 16905 25355 16945
rect 25395 16905 25405 16945
rect 25445 16905 25455 16945
rect 25495 16905 25505 16945
rect 25545 16905 25555 16945
rect 25595 16905 25605 16945
rect 25645 16905 25655 16945
rect 25695 16905 25705 16945
rect 25745 16905 25755 16945
rect 25795 16905 25805 16945
rect 25845 16905 25855 16945
rect 25895 16905 25905 16945
rect 25945 16905 25955 16945
rect 25995 16905 26005 16945
rect 26045 16905 26055 16945
rect 26095 16905 26105 16945
rect 26145 16905 26155 16945
rect 26195 16905 26205 16945
rect 26245 16905 26255 16945
rect 26295 16905 26305 16945
rect 26345 16905 26355 16945
rect 26395 16905 26405 16945
rect 26445 16905 26455 16945
rect 26495 16905 26505 16945
rect 26545 16905 26555 16945
rect 26595 16905 26605 16945
rect 26645 16905 26655 16945
rect 26695 16905 26705 16945
rect 26745 16905 26755 16945
rect 26795 16905 26805 16945
rect 26845 16905 26855 16945
rect 26895 16905 26905 16945
rect 26945 16905 26955 16945
rect 26995 16905 27005 16945
rect 27045 16905 27055 16945
rect 27095 16905 27105 16945
rect 27145 16905 27155 16945
rect 27195 16905 27205 16945
rect 27245 16905 27255 16945
rect 27295 16905 27305 16945
rect 27345 16905 27355 16945
rect 27395 16905 27405 16945
rect 27445 16905 27455 16945
rect 27495 16905 27505 16945
rect 27545 16905 27555 16945
rect 27595 16905 27605 16945
rect 27645 16905 27655 16945
rect 27695 16905 27705 16945
rect 27745 16905 27755 16945
rect 27795 16905 27805 16945
rect 27845 16905 27855 16945
rect 27895 16905 27905 16945
rect 27945 16905 27955 16945
rect 27995 16905 28005 16945
rect 28045 16905 28055 16945
rect 28095 16905 28105 16945
rect 28145 16905 28155 16945
rect 28195 16905 28205 16945
rect 28245 16905 28255 16945
rect 28295 16905 28305 16945
rect 28345 16905 28355 16945
rect 28395 16905 28405 16945
rect 28445 16905 28455 16945
rect 28495 16905 28505 16945
rect 28545 16905 28555 16945
rect 28595 16905 28605 16945
rect 28645 16905 28655 16945
rect 28695 16905 28705 16945
rect 28745 16905 28755 16945
rect 28795 16905 28805 16945
rect 28845 16905 28855 16945
rect 28895 16905 28905 16945
rect 28945 16905 28955 16945
rect 28995 16905 29005 16945
rect 29045 16905 29055 16945
rect 29095 16905 29105 16945
rect 29145 16905 29155 16945
rect 29195 16905 29205 16945
rect 29245 16905 29255 16945
rect 29295 16905 29305 16945
rect 29345 16905 29355 16945
rect 29395 16905 29405 16945
rect 29445 16905 29455 16945
rect 29495 16905 29505 16945
rect 29545 16905 29555 16945
rect 29595 16905 29605 16945
rect 29645 16905 29655 16945
rect 29695 16905 29705 16945
rect 29745 16905 29755 16945
rect 29795 16905 29805 16945
rect 29845 16905 29855 16945
rect 29895 16905 29905 16945
rect 29945 16905 29955 16945
rect 29995 16905 30005 16945
rect 30045 16905 30055 16945
rect 30095 16905 30105 16945
rect 30145 16905 30155 16945
rect 30195 16905 30205 16945
rect 30245 16905 30255 16945
rect 30295 16905 30305 16945
rect 30345 16905 30355 16945
rect 30395 16905 30405 16945
rect 30445 16905 30455 16945
rect 30495 16905 30505 16945
rect 30545 16905 30555 16945
rect 30595 16905 30605 16945
rect 30645 16905 30655 16945
rect 30695 16905 30705 16945
rect 30745 16905 30755 16945
rect 30795 16905 30805 16945
rect 30845 16905 30855 16945
rect 30895 16905 30905 16945
rect 30945 16905 30955 16945
rect 30995 16905 31005 16945
rect 31045 16905 31055 16945
rect 31095 16905 31105 16945
rect 31145 16905 31155 16945
rect 31195 16905 31205 16945
rect 31245 16905 31255 16945
rect 31295 16905 31305 16945
rect 31345 16905 31355 16945
rect 31395 16905 31405 16945
rect 31445 16905 31455 16945
rect 31495 16905 31505 16945
rect 31545 16905 31555 16945
rect 31595 16905 31605 16945
rect 31645 16905 31655 16945
rect 31695 16905 31705 16945
rect 31745 16905 31755 16945
rect 31795 16905 31805 16945
rect 31845 16905 31855 16945
rect 31895 16905 31905 16945
rect 31945 16905 31955 16945
rect 31995 16905 32005 16945
rect 32045 16905 32055 16945
rect 32095 16905 32105 16945
rect 32145 16905 32155 16945
rect 32195 16905 32205 16945
rect 32245 16905 32255 16945
rect 32295 16905 32305 16945
rect 32345 16905 32355 16945
rect 32395 16905 32405 16945
rect 32445 16905 32455 16945
rect 32495 16905 32505 16945
rect 32545 16905 32555 16945
rect 32595 16905 32605 16945
rect 32645 16905 32655 16945
rect 32695 16905 32705 16945
rect 32745 16905 32755 16945
rect 32795 16905 32805 16945
rect 32845 16905 32855 16945
rect 32895 16905 32905 16945
rect 32945 16905 32955 16945
rect 32995 16905 33005 16945
rect 33045 16905 33055 16945
rect 33095 16905 33105 16945
rect 33145 16905 33155 16945
rect 33195 16905 33205 16945
rect 33245 16905 33255 16945
rect 33295 16905 33305 16945
rect 33345 16905 33355 16945
rect 33395 16905 33405 16945
rect 33445 16905 33455 16945
rect 33495 16905 33505 16945
rect 33545 16905 33555 16945
rect 33595 16905 33605 16945
rect 33645 16905 33655 16945
rect 33695 16905 33705 16945
rect 33745 16905 33755 16945
rect 33795 16905 33805 16945
rect 33845 16905 33855 16945
rect 33895 16905 33905 16945
rect 33945 16905 33955 16945
rect 33995 16905 34005 16945
rect 34045 16905 34055 16945
rect 34095 16905 34105 16945
rect 34145 16905 34155 16945
rect 34195 16905 34205 16945
rect 34245 16905 34255 16945
rect 34295 16905 34305 16945
rect 34345 16905 34355 16945
rect 34395 16905 34405 16945
rect 34445 16905 34455 16945
rect 34495 16905 34505 16945
rect 34545 16905 34555 16945
rect 34595 16905 34605 16945
rect 34645 16905 34655 16945
rect 34695 16905 34705 16945
rect 34745 16905 34755 16945
rect 34795 16905 34805 16945
rect 34845 16905 34855 16945
rect 34895 16905 34905 16945
rect 34945 16905 34955 16945
rect 34995 16905 35005 16945
rect 35045 16905 35055 16945
rect 35095 16905 35105 16945
rect 35145 16905 35155 16945
rect 35195 16905 35205 16945
rect 35245 16905 35255 16945
rect 35295 16905 35305 16945
rect 35345 16905 35355 16945
rect 35395 16905 35405 16945
rect 35445 16905 35455 16945
rect 35495 16905 35505 16945
rect 35545 16905 35555 16945
rect 35595 16905 35605 16945
rect 35645 16905 35655 16945
rect 35695 16905 35705 16945
rect 35745 16905 35755 16945
rect 35795 16905 35805 16945
rect 35845 16905 35855 16945
rect 35895 16905 35905 16945
rect 35945 16905 35955 16945
rect 35995 16905 36005 16945
rect 36045 16905 36055 16945
rect 36095 16905 36105 16945
rect 36145 16905 36155 16945
rect 36195 16905 36205 16945
rect 36245 16905 36255 16945
rect 36295 16905 36305 16945
rect 36345 16905 36355 16945
rect 36395 16905 36405 16945
rect 36445 16905 36455 16945
rect 36495 16905 36505 16945
rect 36545 16905 36555 16945
rect 36595 16905 36605 16945
rect 36645 16905 36655 16945
rect 36695 16905 36705 16945
rect 36745 16905 36755 16945
rect 36795 16905 36805 16945
rect 36845 16905 36855 16945
rect 36895 16905 36905 16945
rect 36945 16905 36955 16945
rect 36995 16905 37005 16945
rect 37045 16905 37055 16945
rect 37095 16905 37105 16945
rect 37145 16905 37155 16945
rect 37195 16905 37205 16945
rect 37245 16905 37255 16945
rect 37295 16905 37305 16945
rect 37345 16905 37355 16945
rect 37395 16905 37405 16945
rect 37445 16905 37455 16945
rect 37495 16905 37505 16945
rect 37545 16905 37555 16945
rect 37595 16905 37605 16945
rect 37645 16905 37655 16945
rect 37695 16905 37705 16945
rect 37745 16905 37755 16945
rect 37795 16905 37805 16945
rect 37845 16905 37855 16945
rect 37895 16905 37905 16945
rect 37945 16905 37955 16945
rect 37995 16905 38005 16945
rect 38045 16905 38055 16945
rect 38095 16905 38105 16945
rect 38145 16905 38155 16945
rect 38195 16905 38205 16945
rect 38245 16905 38255 16945
rect 38295 16905 38305 16945
rect 38345 16905 38355 16945
rect 38395 16905 38405 16945
rect 38445 16905 38455 16945
rect 38495 16905 38505 16945
rect 38545 16905 38555 16945
rect 38595 16905 38605 16945
rect 38645 16905 38655 16945
rect 38695 16905 38705 16945
rect 38745 16905 38755 16945
rect 38795 16905 38805 16945
rect 38845 16905 38855 16945
rect 38895 16905 38905 16945
rect 38945 16905 38955 16945
rect 38995 16905 39005 16945
rect 39045 16905 39055 16945
rect 39095 16905 39105 16945
rect 39145 16905 39155 16945
rect 39195 16905 39205 16945
rect 39245 16905 39255 16945
rect 39295 16905 39305 16945
rect 39345 16905 39355 16945
rect 39395 16905 39405 16945
rect 39445 16905 39455 16945
rect 39495 16905 39505 16945
rect 39545 16905 39555 16945
rect 39595 16905 39605 16945
rect 39645 16905 39655 16945
rect 39695 16905 39705 16945
rect 39745 16905 39905 16945
rect 39945 16905 39955 16945
rect 39995 16905 40005 16945
rect 40045 16905 40055 16945
rect 40095 16905 40105 16945
rect 40145 16905 40155 16945
rect 40195 16905 40205 16945
rect 40245 16905 40255 16945
rect 40295 16905 40305 16945
rect 40345 16905 40355 16945
rect 40395 16905 40405 16945
rect 40445 16905 40455 16945
rect 40495 16905 40505 16945
rect 40545 16905 40555 16945
rect 40595 16905 40605 16945
rect 40645 16905 40655 16945
rect 40695 16905 40705 16945
rect 40745 16905 40755 16945
rect 40795 16905 40805 16945
rect 40845 16905 40855 16945
rect 40895 16905 40900 16945
rect 0 16900 40900 16905
rect -400 16845 39750 16850
rect -400 16805 -395 16845
rect -355 16805 105 16845
rect 145 16805 155 16845
rect 195 16805 205 16845
rect 245 16805 255 16845
rect 295 16805 305 16845
rect 345 16805 355 16845
rect 395 16805 405 16845
rect 445 16805 455 16845
rect 495 16805 505 16845
rect 545 16805 555 16845
rect 595 16805 605 16845
rect 645 16805 655 16845
rect 695 16805 705 16845
rect 745 16805 755 16845
rect 795 16805 805 16845
rect 845 16805 855 16845
rect 895 16805 905 16845
rect 945 16805 955 16845
rect 995 16805 1005 16845
rect 1045 16805 1055 16845
rect 1095 16805 1105 16845
rect 1145 16805 1155 16845
rect 1195 16805 1205 16845
rect 1245 16805 1255 16845
rect 1295 16805 1305 16845
rect 1345 16805 1355 16845
rect 1395 16805 1405 16845
rect 1445 16805 1455 16845
rect 1495 16805 1505 16845
rect 1545 16805 1555 16845
rect 1595 16805 1605 16845
rect 1645 16805 1655 16845
rect 1695 16805 1705 16845
rect 1745 16805 1755 16845
rect 1795 16805 1805 16845
rect 1845 16805 1855 16845
rect 1895 16805 1905 16845
rect 1945 16805 1955 16845
rect 1995 16805 2005 16845
rect 2045 16805 2055 16845
rect 2095 16805 2105 16845
rect 2145 16805 2155 16845
rect 2195 16805 2205 16845
rect 2245 16805 2255 16845
rect 2295 16805 2305 16845
rect 2345 16805 2355 16845
rect 2395 16805 2405 16845
rect 2445 16805 2455 16845
rect 2495 16805 2505 16845
rect 2545 16805 2555 16845
rect 2595 16805 2605 16845
rect 2645 16805 2655 16845
rect 2695 16805 2705 16845
rect 2745 16805 2755 16845
rect 2795 16805 2805 16845
rect 2845 16805 2855 16845
rect 2895 16805 2905 16845
rect 2945 16805 2955 16845
rect 2995 16805 3005 16845
rect 3045 16805 3055 16845
rect 3095 16805 3105 16845
rect 3145 16805 3155 16845
rect 3195 16805 3205 16845
rect 3245 16805 3255 16845
rect 3295 16805 3305 16845
rect 3345 16805 3355 16845
rect 3395 16805 3405 16845
rect 3445 16805 3455 16845
rect 3495 16805 3505 16845
rect 3545 16805 3555 16845
rect 3595 16805 3605 16845
rect 3645 16805 3655 16845
rect 3695 16805 3705 16845
rect 3745 16805 3755 16845
rect 3795 16805 3805 16845
rect 3845 16805 3855 16845
rect 3895 16805 3905 16845
rect 3945 16805 3955 16845
rect 3995 16805 4005 16845
rect 4045 16805 4055 16845
rect 4095 16805 4105 16845
rect 4145 16805 4155 16845
rect 4195 16805 4205 16845
rect 4245 16805 4255 16845
rect 4295 16805 4305 16845
rect 4345 16805 4355 16845
rect 4395 16805 4405 16845
rect 4445 16805 4455 16845
rect 4495 16805 4505 16845
rect 4545 16805 4555 16845
rect 4595 16805 4605 16845
rect 4645 16805 4655 16845
rect 4695 16805 4705 16845
rect 4745 16805 4755 16845
rect 4795 16805 4805 16845
rect 4845 16805 4855 16845
rect 4895 16805 4905 16845
rect 4945 16805 4955 16845
rect 4995 16805 5005 16845
rect 5045 16805 5055 16845
rect 5095 16805 5105 16845
rect 5145 16805 5155 16845
rect 5195 16805 5205 16845
rect 5245 16805 5255 16845
rect 5295 16805 5305 16845
rect 5345 16805 5355 16845
rect 5395 16805 5405 16845
rect 5445 16805 5455 16845
rect 5495 16805 5505 16845
rect 5545 16805 5555 16845
rect 5595 16805 5605 16845
rect 5645 16805 5655 16845
rect 5695 16805 5705 16845
rect 5745 16805 5755 16845
rect 5795 16805 5805 16845
rect 5845 16805 5855 16845
rect 5895 16805 5905 16845
rect 5945 16805 5955 16845
rect 5995 16805 6005 16845
rect 6045 16805 6055 16845
rect 6095 16805 6105 16845
rect 6145 16805 6155 16845
rect 6195 16805 6205 16845
rect 6245 16805 6255 16845
rect 6295 16805 6305 16845
rect 6345 16805 6355 16845
rect 6395 16805 6405 16845
rect 6445 16805 6455 16845
rect 6495 16805 6505 16845
rect 6545 16805 6555 16845
rect 6595 16805 6605 16845
rect 6645 16805 6655 16845
rect 6695 16805 6705 16845
rect 6745 16805 6755 16845
rect 6795 16805 6805 16845
rect 6845 16805 6855 16845
rect 6895 16805 6905 16845
rect 6945 16805 6955 16845
rect 6995 16805 7005 16845
rect 7045 16805 7055 16845
rect 7095 16805 7105 16845
rect 7145 16805 7155 16845
rect 7195 16805 7205 16845
rect 7245 16805 7255 16845
rect 7295 16805 7305 16845
rect 7345 16805 7355 16845
rect 7395 16805 7405 16845
rect 7445 16805 7455 16845
rect 7495 16805 7505 16845
rect 7545 16805 7555 16845
rect 7595 16805 7605 16845
rect 7645 16805 7655 16845
rect 7695 16805 7705 16845
rect 7745 16805 7755 16845
rect 7795 16805 7805 16845
rect 7845 16805 7855 16845
rect 7895 16805 7905 16845
rect 7945 16805 7955 16845
rect 7995 16805 8005 16845
rect 8045 16805 8055 16845
rect 8095 16805 8105 16845
rect 8145 16805 8155 16845
rect 8195 16805 8205 16845
rect 8245 16805 8255 16845
rect 8295 16805 8305 16845
rect 8345 16805 8355 16845
rect 8395 16805 8405 16845
rect 8445 16805 8455 16845
rect 8495 16805 8505 16845
rect 8545 16805 8555 16845
rect 8595 16805 8605 16845
rect 8645 16805 8655 16845
rect 8695 16805 8705 16845
rect 8745 16805 8755 16845
rect 8795 16805 8805 16845
rect 8845 16805 8855 16845
rect 8895 16805 8905 16845
rect 8945 16805 8955 16845
rect 8995 16805 9005 16845
rect 9045 16805 9055 16845
rect 9095 16805 9105 16845
rect 9145 16805 9155 16845
rect 9195 16805 9205 16845
rect 9245 16805 9255 16845
rect 9295 16805 9305 16845
rect 9345 16805 9355 16845
rect 9395 16805 9405 16845
rect 9445 16805 9455 16845
rect 9495 16805 9505 16845
rect 9545 16805 9555 16845
rect 9595 16805 9605 16845
rect 9645 16805 9655 16845
rect 9695 16805 9705 16845
rect 9745 16805 9755 16845
rect 9795 16805 9805 16845
rect 9845 16805 9855 16845
rect 9895 16805 9905 16845
rect 9945 16805 9955 16845
rect 9995 16805 10005 16845
rect 10045 16805 10055 16845
rect 10095 16805 10105 16845
rect 10145 16805 10155 16845
rect 10195 16805 10205 16845
rect 10245 16805 10255 16845
rect 10295 16805 10305 16845
rect 10345 16805 10355 16845
rect 10395 16805 10405 16845
rect 10445 16805 10455 16845
rect 10495 16805 10505 16845
rect 10545 16805 10555 16845
rect 10595 16805 10605 16845
rect 10645 16805 10655 16845
rect 10695 16805 10705 16845
rect 10745 16805 10755 16845
rect 10795 16805 10805 16845
rect 10845 16805 10855 16845
rect 10895 16805 10905 16845
rect 10945 16805 10955 16845
rect 10995 16805 11005 16845
rect 11045 16805 11055 16845
rect 11095 16805 11105 16845
rect 11145 16805 11155 16845
rect 11195 16805 11205 16845
rect 11245 16805 11255 16845
rect 11295 16805 11305 16845
rect 11345 16805 11355 16845
rect 11395 16805 11405 16845
rect 11445 16805 11455 16845
rect 11495 16805 11505 16845
rect 11545 16805 11555 16845
rect 11595 16805 11605 16845
rect 11645 16805 11655 16845
rect 11695 16805 11705 16845
rect 11745 16805 11755 16845
rect 11795 16805 11805 16845
rect 11845 16805 11855 16845
rect 11895 16805 11905 16845
rect 11945 16805 11955 16845
rect 11995 16805 12005 16845
rect 12045 16805 12055 16845
rect 12095 16805 12105 16845
rect 12145 16805 12155 16845
rect 12195 16805 12205 16845
rect 12245 16805 12255 16845
rect 12295 16805 12305 16845
rect 12345 16805 12355 16845
rect 12395 16805 12405 16845
rect 12445 16805 12455 16845
rect 12495 16805 12505 16845
rect 12545 16805 12555 16845
rect 12595 16805 12605 16845
rect 12645 16805 12655 16845
rect 12695 16805 12705 16845
rect 12745 16805 12755 16845
rect 12795 16805 12805 16845
rect 12845 16805 12855 16845
rect 12895 16805 12905 16845
rect 12945 16805 12955 16845
rect 12995 16805 13005 16845
rect 13045 16805 13055 16845
rect 13095 16805 13105 16845
rect 13145 16805 13155 16845
rect 13195 16805 13205 16845
rect 13245 16805 13255 16845
rect 13295 16805 13305 16845
rect 13345 16805 13355 16845
rect 13395 16805 13405 16845
rect 13445 16805 13455 16845
rect 13495 16805 13505 16845
rect 13545 16805 13555 16845
rect 13595 16805 13605 16845
rect 13645 16805 13655 16845
rect 13695 16805 13705 16845
rect 13745 16805 13755 16845
rect 13795 16805 13805 16845
rect 13845 16805 13855 16845
rect 13895 16805 13905 16845
rect 13945 16805 13955 16845
rect 13995 16805 14005 16845
rect 14045 16805 14055 16845
rect 14095 16805 14105 16845
rect 14145 16805 14155 16845
rect 14195 16805 14205 16845
rect 14245 16805 14255 16845
rect 14295 16805 14305 16845
rect 14345 16805 14355 16845
rect 14395 16805 14405 16845
rect 14445 16805 14455 16845
rect 14495 16805 14505 16845
rect 14545 16805 14555 16845
rect 14595 16805 14605 16845
rect 14645 16805 14655 16845
rect 14695 16805 14705 16845
rect 14745 16805 14755 16845
rect 14795 16805 14805 16845
rect 14845 16805 14855 16845
rect 14895 16805 14905 16845
rect 14945 16805 14955 16845
rect 14995 16805 15005 16845
rect 15045 16805 15055 16845
rect 15095 16805 15105 16845
rect 15145 16805 15155 16845
rect 15195 16805 15205 16845
rect 15245 16805 15255 16845
rect 15295 16805 15305 16845
rect 15345 16805 15355 16845
rect 15395 16805 15405 16845
rect 15445 16805 15455 16845
rect 15495 16805 15505 16845
rect 15545 16805 15555 16845
rect 15595 16805 15605 16845
rect 15645 16805 15655 16845
rect 15695 16805 15705 16845
rect 15745 16805 15755 16845
rect 15795 16805 15805 16845
rect 15845 16805 15855 16845
rect 15895 16805 15905 16845
rect 15945 16805 15955 16845
rect 15995 16805 16005 16845
rect 16045 16805 16055 16845
rect 16095 16805 16105 16845
rect 16145 16805 16155 16845
rect 16195 16805 16205 16845
rect 16245 16805 16255 16845
rect 16295 16805 16305 16845
rect 16345 16805 16355 16845
rect 16395 16805 16405 16845
rect 16445 16805 16455 16845
rect 16495 16805 16505 16845
rect 16545 16805 16555 16845
rect 16595 16805 16605 16845
rect 16645 16805 16655 16845
rect 16695 16805 16705 16845
rect 16745 16805 16755 16845
rect 16795 16805 16805 16845
rect 16845 16805 16855 16845
rect 16895 16805 16905 16845
rect 16945 16805 16955 16845
rect 16995 16805 17005 16845
rect 17045 16805 17055 16845
rect 17095 16805 17105 16845
rect 17145 16805 17155 16845
rect 17195 16805 17205 16845
rect 17245 16805 17255 16845
rect 17295 16805 17305 16845
rect 17345 16805 17355 16845
rect 17395 16805 17405 16845
rect 17445 16805 17455 16845
rect 17495 16805 17505 16845
rect 17545 16805 17555 16845
rect 17595 16805 17605 16845
rect 17645 16805 17655 16845
rect 17695 16805 17705 16845
rect 17745 16805 17755 16845
rect 17795 16805 17805 16845
rect 17845 16805 17855 16845
rect 17895 16805 17905 16845
rect 17945 16805 17955 16845
rect 17995 16805 18005 16845
rect 18045 16805 18055 16845
rect 18095 16805 18105 16845
rect 18145 16805 18155 16845
rect 18195 16805 18205 16845
rect 18245 16805 18255 16845
rect 18295 16805 18305 16845
rect 18345 16805 18355 16845
rect 18395 16805 18405 16845
rect 18445 16805 18455 16845
rect 18495 16805 18505 16845
rect 18545 16805 18555 16845
rect 18595 16805 18605 16845
rect 18645 16805 18655 16845
rect 18695 16805 18705 16845
rect 18745 16805 18755 16845
rect 18795 16805 18805 16845
rect 18845 16805 18855 16845
rect 18895 16805 18905 16845
rect 18945 16805 18955 16845
rect 18995 16805 19005 16845
rect 19045 16805 19055 16845
rect 19095 16805 19105 16845
rect 19145 16805 19155 16845
rect 19195 16805 19205 16845
rect 19245 16805 19255 16845
rect 19295 16805 19305 16845
rect 19345 16805 19355 16845
rect 19395 16805 19405 16845
rect 19445 16805 19455 16845
rect 19495 16805 19505 16845
rect 19545 16805 19555 16845
rect 19595 16805 19605 16845
rect 19645 16805 19655 16845
rect 19695 16805 19705 16845
rect 19745 16805 19755 16845
rect 19795 16805 19805 16845
rect 19845 16805 19855 16845
rect 19895 16805 19905 16845
rect 19945 16805 19955 16845
rect 19995 16805 20005 16845
rect 20045 16805 20055 16845
rect 20095 16805 20105 16845
rect 20145 16805 20155 16845
rect 20195 16805 20205 16845
rect 20245 16805 20255 16845
rect 20295 16805 20305 16845
rect 20345 16805 20355 16845
rect 20395 16805 20405 16845
rect 20445 16805 20455 16845
rect 20495 16805 20505 16845
rect 20545 16805 20555 16845
rect 20595 16805 20605 16845
rect 20645 16805 20655 16845
rect 20695 16805 20705 16845
rect 20745 16805 20755 16845
rect 20795 16805 20805 16845
rect 20845 16805 20855 16845
rect 20895 16805 20905 16845
rect 20945 16805 20955 16845
rect 20995 16805 21005 16845
rect 21045 16805 21055 16845
rect 21095 16805 21105 16845
rect 21145 16805 21155 16845
rect 21195 16805 21205 16845
rect 21245 16805 21255 16845
rect 21295 16805 21305 16845
rect 21345 16805 21355 16845
rect 21395 16805 21405 16845
rect 21445 16805 21455 16845
rect 21495 16805 21505 16845
rect 21545 16805 21555 16845
rect 21595 16805 21605 16845
rect 21645 16805 21655 16845
rect 21695 16805 21705 16845
rect 21745 16805 21755 16845
rect 21795 16805 21805 16845
rect 21845 16805 21855 16845
rect 21895 16805 21905 16845
rect 21945 16805 21955 16845
rect 21995 16805 22005 16845
rect 22045 16805 22055 16845
rect 22095 16805 22105 16845
rect 22145 16805 22155 16845
rect 22195 16805 22205 16845
rect 22245 16805 22255 16845
rect 22295 16805 22305 16845
rect 22345 16805 22355 16845
rect 22395 16805 22405 16845
rect 22445 16805 22455 16845
rect 22495 16805 22505 16845
rect 22545 16805 22555 16845
rect 22595 16805 22605 16845
rect 22645 16805 22655 16845
rect 22695 16805 22705 16845
rect 22745 16805 22755 16845
rect 22795 16805 22805 16845
rect 22845 16805 22855 16845
rect 22895 16805 22905 16845
rect 22945 16805 22955 16845
rect 22995 16805 23005 16845
rect 23045 16805 23055 16845
rect 23095 16805 23105 16845
rect 23145 16805 23155 16845
rect 23195 16805 23205 16845
rect 23245 16805 23255 16845
rect 23295 16805 23305 16845
rect 23345 16805 23355 16845
rect 23395 16805 23405 16845
rect 23445 16805 23455 16845
rect 23495 16805 23505 16845
rect 23545 16805 23555 16845
rect 23595 16805 23605 16845
rect 23645 16805 23655 16845
rect 23695 16805 23705 16845
rect 23745 16805 23755 16845
rect 23795 16805 23805 16845
rect 23845 16805 23855 16845
rect 23895 16805 23905 16845
rect 23945 16805 23955 16845
rect 23995 16805 24005 16845
rect 24045 16805 24055 16845
rect 24095 16805 24105 16845
rect 24145 16805 24155 16845
rect 24195 16805 24205 16845
rect 24245 16805 24255 16845
rect 24295 16805 24305 16845
rect 24345 16805 24355 16845
rect 24395 16805 24405 16845
rect 24445 16805 24455 16845
rect 24495 16805 24505 16845
rect 24545 16805 24555 16845
rect 24595 16805 24605 16845
rect 24645 16805 24655 16845
rect 24695 16805 24705 16845
rect 24745 16805 24755 16845
rect 24795 16805 24805 16845
rect 24845 16805 24855 16845
rect 24895 16805 24905 16845
rect 24945 16805 24955 16845
rect 24995 16805 25005 16845
rect 25045 16805 25055 16845
rect 25095 16805 25105 16845
rect 25145 16805 25155 16845
rect 25195 16805 25205 16845
rect 25245 16805 25255 16845
rect 25295 16805 25305 16845
rect 25345 16805 25355 16845
rect 25395 16805 25405 16845
rect 25445 16805 25455 16845
rect 25495 16805 25505 16845
rect 25545 16805 25555 16845
rect 25595 16805 25605 16845
rect 25645 16805 25655 16845
rect 25695 16805 25705 16845
rect 25745 16805 25755 16845
rect 25795 16805 25805 16845
rect 25845 16805 25855 16845
rect 25895 16805 25905 16845
rect 25945 16805 25955 16845
rect 25995 16805 26005 16845
rect 26045 16805 26055 16845
rect 26095 16805 26105 16845
rect 26145 16805 26155 16845
rect 26195 16805 26205 16845
rect 26245 16805 26255 16845
rect 26295 16805 26305 16845
rect 26345 16805 26355 16845
rect 26395 16805 26405 16845
rect 26445 16805 26455 16845
rect 26495 16805 26505 16845
rect 26545 16805 26555 16845
rect 26595 16805 26605 16845
rect 26645 16805 26655 16845
rect 26695 16805 26705 16845
rect 26745 16805 26755 16845
rect 26795 16805 26805 16845
rect 26845 16805 26855 16845
rect 26895 16805 26905 16845
rect 26945 16805 26955 16845
rect 26995 16805 27005 16845
rect 27045 16805 27055 16845
rect 27095 16805 27105 16845
rect 27145 16805 27155 16845
rect 27195 16805 27205 16845
rect 27245 16805 27255 16845
rect 27295 16805 27305 16845
rect 27345 16805 27355 16845
rect 27395 16805 27405 16845
rect 27445 16805 27455 16845
rect 27495 16805 27505 16845
rect 27545 16805 27555 16845
rect 27595 16805 27605 16845
rect 27645 16805 27655 16845
rect 27695 16805 27705 16845
rect 27745 16805 27755 16845
rect 27795 16805 27805 16845
rect 27845 16805 27855 16845
rect 27895 16805 27905 16845
rect 27945 16805 27955 16845
rect 27995 16805 28005 16845
rect 28045 16805 28055 16845
rect 28095 16805 28105 16845
rect 28145 16805 28155 16845
rect 28195 16805 28205 16845
rect 28245 16805 28255 16845
rect 28295 16805 28305 16845
rect 28345 16805 28355 16845
rect 28395 16805 28405 16845
rect 28445 16805 28455 16845
rect 28495 16805 28505 16845
rect 28545 16805 28555 16845
rect 28595 16805 28605 16845
rect 28645 16805 28655 16845
rect 28695 16805 28705 16845
rect 28745 16805 28755 16845
rect 28795 16805 28805 16845
rect 28845 16805 28855 16845
rect 28895 16805 28905 16845
rect 28945 16805 28955 16845
rect 28995 16805 29005 16845
rect 29045 16805 29055 16845
rect 29095 16805 29105 16845
rect 29145 16805 29155 16845
rect 29195 16805 29205 16845
rect 29245 16805 29255 16845
rect 29295 16805 29305 16845
rect 29345 16805 29355 16845
rect 29395 16805 29405 16845
rect 29445 16805 29455 16845
rect 29495 16805 29505 16845
rect 29545 16805 29555 16845
rect 29595 16805 29605 16845
rect 29645 16805 29655 16845
rect 29695 16805 29705 16845
rect 29745 16805 29755 16845
rect 29795 16805 29805 16845
rect 29845 16805 29855 16845
rect 29895 16805 29905 16845
rect 29945 16805 29955 16845
rect 29995 16805 30005 16845
rect 30045 16805 30055 16845
rect 30095 16805 30105 16845
rect 30145 16805 30155 16845
rect 30195 16805 30205 16845
rect 30245 16805 30255 16845
rect 30295 16805 30305 16845
rect 30345 16805 30355 16845
rect 30395 16805 30405 16845
rect 30445 16805 30455 16845
rect 30495 16805 30505 16845
rect 30545 16805 30555 16845
rect 30595 16805 30605 16845
rect 30645 16805 30655 16845
rect 30695 16805 30705 16845
rect 30745 16805 30755 16845
rect 30795 16805 30805 16845
rect 30845 16805 30855 16845
rect 30895 16805 30905 16845
rect 30945 16805 30955 16845
rect 30995 16805 31005 16845
rect 31045 16805 31055 16845
rect 31095 16805 31105 16845
rect 31145 16805 31155 16845
rect 31195 16805 31205 16845
rect 31245 16805 31255 16845
rect 31295 16805 31305 16845
rect 31345 16805 31355 16845
rect 31395 16805 31405 16845
rect 31445 16805 31455 16845
rect 31495 16805 31505 16845
rect 31545 16805 31555 16845
rect 31595 16805 31605 16845
rect 31645 16805 31655 16845
rect 31695 16805 31705 16845
rect 31745 16805 31755 16845
rect 31795 16805 31805 16845
rect 31845 16805 31855 16845
rect 31895 16805 31905 16845
rect 31945 16805 31955 16845
rect 31995 16805 32005 16845
rect 32045 16805 32055 16845
rect 32095 16805 32105 16845
rect 32145 16805 32155 16845
rect 32195 16805 32205 16845
rect 32245 16805 32255 16845
rect 32295 16805 32305 16845
rect 32345 16805 32355 16845
rect 32395 16805 32405 16845
rect 32445 16805 32455 16845
rect 32495 16805 32505 16845
rect 32545 16805 32555 16845
rect 32595 16805 32605 16845
rect 32645 16805 32655 16845
rect 32695 16805 32705 16845
rect 32745 16805 32755 16845
rect 32795 16805 32805 16845
rect 32845 16805 32855 16845
rect 32895 16805 32905 16845
rect 32945 16805 32955 16845
rect 32995 16805 33005 16845
rect 33045 16805 33055 16845
rect 33095 16805 33105 16845
rect 33145 16805 33155 16845
rect 33195 16805 33205 16845
rect 33245 16805 33255 16845
rect 33295 16805 33305 16845
rect 33345 16805 33355 16845
rect 33395 16805 33405 16845
rect 33445 16805 33455 16845
rect 33495 16805 33505 16845
rect 33545 16805 33555 16845
rect 33595 16805 33605 16845
rect 33645 16805 33655 16845
rect 33695 16805 33705 16845
rect 33745 16805 33755 16845
rect 33795 16805 33805 16845
rect 33845 16805 33855 16845
rect 33895 16805 33905 16845
rect 33945 16805 33955 16845
rect 33995 16805 34005 16845
rect 34045 16805 34055 16845
rect 34095 16805 34105 16845
rect 34145 16805 34155 16845
rect 34195 16805 34205 16845
rect 34245 16805 34255 16845
rect 34295 16805 34305 16845
rect 34345 16805 34355 16845
rect 34395 16805 34405 16845
rect 34445 16805 34455 16845
rect 34495 16805 34505 16845
rect 34545 16805 34555 16845
rect 34595 16805 34605 16845
rect 34645 16805 34655 16845
rect 34695 16805 34705 16845
rect 34745 16805 34755 16845
rect 34795 16805 34805 16845
rect 34845 16805 34855 16845
rect 34895 16805 34905 16845
rect 34945 16805 34955 16845
rect 34995 16805 35005 16845
rect 35045 16805 35055 16845
rect 35095 16805 35105 16845
rect 35145 16805 35155 16845
rect 35195 16805 35205 16845
rect 35245 16805 35255 16845
rect 35295 16805 35305 16845
rect 35345 16805 35355 16845
rect 35395 16805 35405 16845
rect 35445 16805 35455 16845
rect 35495 16805 35505 16845
rect 35545 16805 35555 16845
rect 35595 16805 35605 16845
rect 35645 16805 35655 16845
rect 35695 16805 35705 16845
rect 35745 16805 35755 16845
rect 35795 16805 35805 16845
rect 35845 16805 35855 16845
rect 35895 16805 35905 16845
rect 35945 16805 35955 16845
rect 35995 16805 36005 16845
rect 36045 16805 36055 16845
rect 36095 16805 36105 16845
rect 36145 16805 36155 16845
rect 36195 16805 36205 16845
rect 36245 16805 36255 16845
rect 36295 16805 36305 16845
rect 36345 16805 36355 16845
rect 36395 16805 36405 16845
rect 36445 16805 36455 16845
rect 36495 16805 36505 16845
rect 36545 16805 36555 16845
rect 36595 16805 36605 16845
rect 36645 16805 36655 16845
rect 36695 16805 36705 16845
rect 36745 16805 36755 16845
rect 36795 16805 36805 16845
rect 36845 16805 36855 16845
rect 36895 16805 36905 16845
rect 36945 16805 36955 16845
rect 36995 16805 37005 16845
rect 37045 16805 37055 16845
rect 37095 16805 37105 16845
rect 37145 16805 37155 16845
rect 37195 16805 37205 16845
rect 37245 16805 37255 16845
rect 37295 16805 37305 16845
rect 37345 16805 37355 16845
rect 37395 16805 37405 16845
rect 37445 16805 37455 16845
rect 37495 16805 37505 16845
rect 37545 16805 37555 16845
rect 37595 16805 37605 16845
rect 37645 16805 37655 16845
rect 37695 16805 37705 16845
rect 37745 16805 37755 16845
rect 37795 16805 37805 16845
rect 37845 16805 37855 16845
rect 37895 16805 37905 16845
rect 37945 16805 37955 16845
rect 37995 16805 38005 16845
rect 38045 16805 38055 16845
rect 38095 16805 38105 16845
rect 38145 16805 38155 16845
rect 38195 16805 38205 16845
rect 38245 16805 38255 16845
rect 38295 16805 38305 16845
rect 38345 16805 38355 16845
rect 38395 16805 38405 16845
rect 38445 16805 38455 16845
rect 38495 16805 38505 16845
rect 38545 16805 38555 16845
rect 38595 16805 38605 16845
rect 38645 16805 38655 16845
rect 38695 16805 38705 16845
rect 38745 16805 38755 16845
rect 38795 16805 38805 16845
rect 38845 16805 38855 16845
rect 38895 16805 38905 16845
rect 38945 16805 38955 16845
rect 38995 16805 39005 16845
rect 39045 16805 39055 16845
rect 39095 16805 39105 16845
rect 39145 16805 39155 16845
rect 39195 16805 39205 16845
rect 39245 16805 39255 16845
rect 39295 16805 39305 16845
rect 39345 16805 39355 16845
rect 39395 16805 39405 16845
rect 39445 16805 39455 16845
rect 39495 16805 39505 16845
rect 39545 16805 39555 16845
rect 39595 16805 39605 16845
rect 39645 16805 39655 16845
rect 39695 16805 39705 16845
rect 39745 16805 39750 16845
rect -400 16800 39750 16805
rect 100 15850 3200 16750
rect 3350 15850 6450 16750
rect 6600 15850 9700 16750
rect 9850 15850 12950 16750
rect 13100 15850 16200 16750
rect 16350 15850 19450 16750
rect 19600 15850 22700 16750
rect 22850 15850 25950 16750
rect 26100 15850 29200 16750
rect 29350 15850 32450 16750
rect 32600 15850 35700 16750
rect 35850 15850 38950 16750
rect 39100 15850 39750 16750
rect 0 15845 39750 15850
rect 0 15805 5 15845
rect 45 15805 55 15845
rect 95 15805 105 15845
rect 145 15805 155 15845
rect 195 15805 205 15845
rect 245 15805 255 15845
rect 295 15805 305 15845
rect 345 15805 355 15845
rect 395 15805 405 15845
rect 445 15805 455 15845
rect 495 15805 505 15845
rect 545 15805 555 15845
rect 595 15805 605 15845
rect 645 15805 655 15845
rect 695 15805 705 15845
rect 745 15805 755 15845
rect 795 15805 805 15845
rect 845 15805 855 15845
rect 895 15805 905 15845
rect 945 15805 955 15845
rect 995 15805 1005 15845
rect 1045 15805 1055 15845
rect 1095 15805 1105 15845
rect 1145 15805 1155 15845
rect 1195 15805 1205 15845
rect 1245 15805 1255 15845
rect 1295 15805 1305 15845
rect 1345 15805 1355 15845
rect 1395 15805 1405 15845
rect 1445 15805 1455 15845
rect 1495 15805 1505 15845
rect 1545 15805 1555 15845
rect 1595 15805 1605 15845
rect 1645 15805 1655 15845
rect 1695 15805 1705 15845
rect 1745 15805 1755 15845
rect 1795 15805 1805 15845
rect 1845 15805 1855 15845
rect 1895 15805 1905 15845
rect 1945 15805 1955 15845
rect 1995 15805 2005 15845
rect 2045 15805 2055 15845
rect 2095 15805 2105 15845
rect 2145 15805 2155 15845
rect 2195 15805 2205 15845
rect 2245 15805 2255 15845
rect 2295 15805 2305 15845
rect 2345 15805 2355 15845
rect 2395 15805 2405 15845
rect 2445 15805 2455 15845
rect 2495 15805 2505 15845
rect 2545 15805 2555 15845
rect 2595 15805 2605 15845
rect 2645 15805 2655 15845
rect 2695 15805 2705 15845
rect 2745 15805 2755 15845
rect 2795 15805 2805 15845
rect 2845 15805 2855 15845
rect 2895 15805 2905 15845
rect 2945 15805 2955 15845
rect 2995 15805 3005 15845
rect 3045 15805 3055 15845
rect 3095 15805 3105 15845
rect 3145 15805 3155 15845
rect 3195 15805 3205 15845
rect 3245 15805 3255 15845
rect 3295 15805 3305 15845
rect 3345 15805 3355 15845
rect 3395 15805 3405 15845
rect 3445 15805 3455 15845
rect 3495 15805 3505 15845
rect 3545 15805 3555 15845
rect 3595 15805 3605 15845
rect 3645 15805 3655 15845
rect 3695 15805 3705 15845
rect 3745 15805 3755 15845
rect 3795 15805 3805 15845
rect 3845 15805 3855 15845
rect 3895 15805 3905 15845
rect 3945 15805 3955 15845
rect 3995 15805 4005 15845
rect 4045 15805 4055 15845
rect 4095 15805 4105 15845
rect 4145 15805 4155 15845
rect 4195 15805 4205 15845
rect 4245 15805 4255 15845
rect 4295 15805 4305 15845
rect 4345 15805 4355 15845
rect 4395 15805 4405 15845
rect 4445 15805 4455 15845
rect 4495 15805 4505 15845
rect 4545 15805 4555 15845
rect 4595 15805 4605 15845
rect 4645 15805 4655 15845
rect 4695 15805 4705 15845
rect 4745 15805 4755 15845
rect 4795 15805 4805 15845
rect 4845 15805 4855 15845
rect 4895 15805 4905 15845
rect 4945 15805 4955 15845
rect 4995 15805 5005 15845
rect 5045 15805 5055 15845
rect 5095 15805 5105 15845
rect 5145 15805 5155 15845
rect 5195 15805 5205 15845
rect 5245 15805 5255 15845
rect 5295 15805 5305 15845
rect 5345 15805 5355 15845
rect 5395 15805 5405 15845
rect 5445 15805 5455 15845
rect 5495 15805 5505 15845
rect 5545 15805 5555 15845
rect 5595 15805 5605 15845
rect 5645 15805 5655 15845
rect 5695 15805 5705 15845
rect 5745 15805 5755 15845
rect 5795 15805 5805 15845
rect 5845 15805 5855 15845
rect 5895 15805 5905 15845
rect 5945 15805 5955 15845
rect 5995 15805 6005 15845
rect 6045 15805 6055 15845
rect 6095 15805 6105 15845
rect 6145 15805 6155 15845
rect 6195 15805 6205 15845
rect 6245 15805 6255 15845
rect 6295 15805 6305 15845
rect 6345 15805 6355 15845
rect 6395 15805 6405 15845
rect 6445 15805 6455 15845
rect 6495 15805 6505 15845
rect 6545 15805 6555 15845
rect 6595 15805 6605 15845
rect 6645 15805 6655 15845
rect 6695 15805 6705 15845
rect 6745 15805 6755 15845
rect 6795 15805 6805 15845
rect 6845 15805 6855 15845
rect 6895 15805 6905 15845
rect 6945 15805 6955 15845
rect 6995 15805 7005 15845
rect 7045 15805 7055 15845
rect 7095 15805 7105 15845
rect 7145 15805 7155 15845
rect 7195 15805 7205 15845
rect 7245 15805 7255 15845
rect 7295 15805 7305 15845
rect 7345 15805 7355 15845
rect 7395 15805 7405 15845
rect 7445 15805 7455 15845
rect 7495 15805 7505 15845
rect 7545 15805 7555 15845
rect 7595 15805 7605 15845
rect 7645 15805 7655 15845
rect 7695 15805 7705 15845
rect 7745 15805 7755 15845
rect 7795 15805 7805 15845
rect 7845 15805 7855 15845
rect 7895 15805 7905 15845
rect 7945 15805 7955 15845
rect 7995 15805 8005 15845
rect 8045 15805 8055 15845
rect 8095 15805 8105 15845
rect 8145 15805 8155 15845
rect 8195 15805 8205 15845
rect 8245 15805 8255 15845
rect 8295 15805 8305 15845
rect 8345 15805 8355 15845
rect 8395 15805 8405 15845
rect 8445 15805 8455 15845
rect 8495 15805 8505 15845
rect 8545 15805 8555 15845
rect 8595 15805 8605 15845
rect 8645 15805 8655 15845
rect 8695 15805 8705 15845
rect 8745 15805 8755 15845
rect 8795 15805 8805 15845
rect 8845 15805 8855 15845
rect 8895 15805 8905 15845
rect 8945 15805 8955 15845
rect 8995 15805 9005 15845
rect 9045 15805 9055 15845
rect 9095 15805 9105 15845
rect 9145 15805 9155 15845
rect 9195 15805 9205 15845
rect 9245 15805 9255 15845
rect 9295 15805 9305 15845
rect 9345 15805 9355 15845
rect 9395 15805 9405 15845
rect 9445 15805 9455 15845
rect 9495 15805 9505 15845
rect 9545 15805 9555 15845
rect 9595 15805 9605 15845
rect 9645 15805 9655 15845
rect 9695 15805 9705 15845
rect 9745 15805 9755 15845
rect 9795 15805 9805 15845
rect 9845 15805 9855 15845
rect 9895 15805 9905 15845
rect 9945 15805 9955 15845
rect 9995 15805 10005 15845
rect 10045 15805 10055 15845
rect 10095 15805 10105 15845
rect 10145 15805 10155 15845
rect 10195 15805 10205 15845
rect 10245 15805 10255 15845
rect 10295 15805 10305 15845
rect 10345 15805 10355 15845
rect 10395 15805 10405 15845
rect 10445 15805 10455 15845
rect 10495 15805 10505 15845
rect 10545 15805 10555 15845
rect 10595 15805 10605 15845
rect 10645 15805 10655 15845
rect 10695 15805 10705 15845
rect 10745 15805 10755 15845
rect 10795 15805 10805 15845
rect 10845 15805 10855 15845
rect 10895 15805 10905 15845
rect 10945 15805 10955 15845
rect 10995 15805 11005 15845
rect 11045 15805 11055 15845
rect 11095 15805 11105 15845
rect 11145 15805 11155 15845
rect 11195 15805 11205 15845
rect 11245 15805 11255 15845
rect 11295 15805 11305 15845
rect 11345 15805 11355 15845
rect 11395 15805 11405 15845
rect 11445 15805 11455 15845
rect 11495 15805 11505 15845
rect 11545 15805 11555 15845
rect 11595 15805 11605 15845
rect 11645 15805 11655 15845
rect 11695 15805 11705 15845
rect 11745 15805 11755 15845
rect 11795 15805 11805 15845
rect 11845 15805 11855 15845
rect 11895 15805 11905 15845
rect 11945 15805 11955 15845
rect 11995 15805 12005 15845
rect 12045 15805 12055 15845
rect 12095 15805 12105 15845
rect 12145 15805 12155 15845
rect 12195 15805 12205 15845
rect 12245 15805 12255 15845
rect 12295 15805 12305 15845
rect 12345 15805 12355 15845
rect 12395 15805 12405 15845
rect 12445 15805 12455 15845
rect 12495 15805 12505 15845
rect 12545 15805 12555 15845
rect 12595 15805 12605 15845
rect 12645 15805 12655 15845
rect 12695 15805 12705 15845
rect 12745 15805 12755 15845
rect 12795 15805 12805 15845
rect 12845 15805 12855 15845
rect 12895 15805 12905 15845
rect 12945 15805 12955 15845
rect 12995 15805 13005 15845
rect 13045 15805 13055 15845
rect 13095 15805 13105 15845
rect 13145 15805 13155 15845
rect 13195 15805 13205 15845
rect 13245 15805 13255 15845
rect 13295 15805 13305 15845
rect 13345 15805 13355 15845
rect 13395 15805 13405 15845
rect 13445 15805 13455 15845
rect 13495 15805 13505 15845
rect 13545 15805 13555 15845
rect 13595 15805 13605 15845
rect 13645 15805 13655 15845
rect 13695 15805 13705 15845
rect 13745 15805 13755 15845
rect 13795 15805 13805 15845
rect 13845 15805 13855 15845
rect 13895 15805 13905 15845
rect 13945 15805 13955 15845
rect 13995 15805 14005 15845
rect 14045 15805 14055 15845
rect 14095 15805 14105 15845
rect 14145 15805 14155 15845
rect 14195 15805 14205 15845
rect 14245 15805 14255 15845
rect 14295 15805 14305 15845
rect 14345 15805 14355 15845
rect 14395 15805 14405 15845
rect 14445 15805 14455 15845
rect 14495 15805 14505 15845
rect 14545 15805 14555 15845
rect 14595 15805 14605 15845
rect 14645 15805 14655 15845
rect 14695 15805 14705 15845
rect 14745 15805 14755 15845
rect 14795 15805 14805 15845
rect 14845 15805 14855 15845
rect 14895 15805 14905 15845
rect 14945 15805 14955 15845
rect 14995 15805 15005 15845
rect 15045 15805 15055 15845
rect 15095 15805 15105 15845
rect 15145 15805 15155 15845
rect 15195 15805 15205 15845
rect 15245 15805 15255 15845
rect 15295 15805 15305 15845
rect 15345 15805 15355 15845
rect 15395 15805 15405 15845
rect 15445 15805 15455 15845
rect 15495 15805 15505 15845
rect 15545 15805 15555 15845
rect 15595 15805 15605 15845
rect 15645 15805 15655 15845
rect 15695 15805 15705 15845
rect 15745 15805 15755 15845
rect 15795 15805 15805 15845
rect 15845 15805 15855 15845
rect 15895 15805 15905 15845
rect 15945 15805 15955 15845
rect 15995 15805 16005 15845
rect 16045 15805 16055 15845
rect 16095 15805 16105 15845
rect 16145 15805 16155 15845
rect 16195 15805 16205 15845
rect 16245 15805 16255 15845
rect 16295 15805 16305 15845
rect 16345 15805 16355 15845
rect 16395 15805 16405 15845
rect 16445 15805 16455 15845
rect 16495 15805 16505 15845
rect 16545 15805 16555 15845
rect 16595 15805 16605 15845
rect 16645 15805 16655 15845
rect 16695 15805 16705 15845
rect 16745 15805 16755 15845
rect 16795 15805 16805 15845
rect 16845 15805 16855 15845
rect 16895 15805 16905 15845
rect 16945 15805 16955 15845
rect 16995 15805 17005 15845
rect 17045 15805 17055 15845
rect 17095 15805 17105 15845
rect 17145 15805 17155 15845
rect 17195 15805 17205 15845
rect 17245 15805 17255 15845
rect 17295 15805 17305 15845
rect 17345 15805 17355 15845
rect 17395 15805 17405 15845
rect 17445 15805 17455 15845
rect 17495 15805 17505 15845
rect 17545 15805 17555 15845
rect 17595 15805 17605 15845
rect 17645 15805 17655 15845
rect 17695 15805 17705 15845
rect 17745 15805 17755 15845
rect 17795 15805 17805 15845
rect 17845 15805 17855 15845
rect 17895 15805 17905 15845
rect 17945 15805 17955 15845
rect 17995 15805 18005 15845
rect 18045 15805 18055 15845
rect 18095 15805 18105 15845
rect 18145 15805 18155 15845
rect 18195 15805 18205 15845
rect 18245 15805 18255 15845
rect 18295 15805 18305 15845
rect 18345 15805 18355 15845
rect 18395 15805 18405 15845
rect 18445 15805 18455 15845
rect 18495 15805 18505 15845
rect 18545 15805 18555 15845
rect 18595 15805 18605 15845
rect 18645 15805 18655 15845
rect 18695 15805 18705 15845
rect 18745 15805 18755 15845
rect 18795 15805 18805 15845
rect 18845 15805 18855 15845
rect 18895 15805 18905 15845
rect 18945 15805 18955 15845
rect 18995 15805 19005 15845
rect 19045 15805 19055 15845
rect 19095 15805 19105 15845
rect 19145 15805 19155 15845
rect 19195 15805 19205 15845
rect 19245 15805 19255 15845
rect 19295 15805 19305 15845
rect 19345 15805 19355 15845
rect 19395 15805 19405 15845
rect 19445 15805 19455 15845
rect 19495 15805 19505 15845
rect 19545 15805 19555 15845
rect 19595 15805 19605 15845
rect 19645 15805 19655 15845
rect 19695 15805 19705 15845
rect 19745 15805 19755 15845
rect 19795 15805 19805 15845
rect 19845 15805 19855 15845
rect 19895 15805 19905 15845
rect 19945 15805 19955 15845
rect 19995 15805 20005 15845
rect 20045 15805 20055 15845
rect 20095 15805 20105 15845
rect 20145 15805 20155 15845
rect 20195 15805 20205 15845
rect 20245 15805 20255 15845
rect 20295 15805 20305 15845
rect 20345 15805 20355 15845
rect 20395 15805 20405 15845
rect 20445 15805 20455 15845
rect 20495 15805 20505 15845
rect 20545 15805 20555 15845
rect 20595 15805 20605 15845
rect 20645 15805 20655 15845
rect 20695 15805 20705 15845
rect 20745 15805 20755 15845
rect 20795 15805 20805 15845
rect 20845 15805 20855 15845
rect 20895 15805 20905 15845
rect 20945 15805 20955 15845
rect 20995 15805 21005 15845
rect 21045 15805 21055 15845
rect 21095 15805 21105 15845
rect 21145 15805 21155 15845
rect 21195 15805 21205 15845
rect 21245 15805 21255 15845
rect 21295 15805 21305 15845
rect 21345 15805 21355 15845
rect 21395 15805 21405 15845
rect 21445 15805 21455 15845
rect 21495 15805 21505 15845
rect 21545 15805 21555 15845
rect 21595 15805 21605 15845
rect 21645 15805 21655 15845
rect 21695 15805 21705 15845
rect 21745 15805 21755 15845
rect 21795 15805 21805 15845
rect 21845 15805 21855 15845
rect 21895 15805 21905 15845
rect 21945 15805 21955 15845
rect 21995 15805 22005 15845
rect 22045 15805 22055 15845
rect 22095 15805 22105 15845
rect 22145 15805 22155 15845
rect 22195 15805 22205 15845
rect 22245 15805 22255 15845
rect 22295 15805 22305 15845
rect 22345 15805 22355 15845
rect 22395 15805 22405 15845
rect 22445 15805 22455 15845
rect 22495 15805 22505 15845
rect 22545 15805 22555 15845
rect 22595 15805 22605 15845
rect 22645 15805 22655 15845
rect 22695 15805 22705 15845
rect 22745 15805 22755 15845
rect 22795 15805 22805 15845
rect 22845 15805 22855 15845
rect 22895 15805 22905 15845
rect 22945 15805 22955 15845
rect 22995 15805 23005 15845
rect 23045 15805 23055 15845
rect 23095 15805 23105 15845
rect 23145 15805 23155 15845
rect 23195 15805 23205 15845
rect 23245 15805 23255 15845
rect 23295 15805 23305 15845
rect 23345 15805 23355 15845
rect 23395 15805 23405 15845
rect 23445 15805 23455 15845
rect 23495 15805 23505 15845
rect 23545 15805 23555 15845
rect 23595 15805 23605 15845
rect 23645 15805 23655 15845
rect 23695 15805 23705 15845
rect 23745 15805 23755 15845
rect 23795 15805 23805 15845
rect 23845 15805 23855 15845
rect 23895 15805 23905 15845
rect 23945 15805 23955 15845
rect 23995 15805 24005 15845
rect 24045 15805 24055 15845
rect 24095 15805 24105 15845
rect 24145 15805 24155 15845
rect 24195 15805 24205 15845
rect 24245 15805 24255 15845
rect 24295 15805 24305 15845
rect 24345 15805 24355 15845
rect 24395 15805 24405 15845
rect 24445 15805 24455 15845
rect 24495 15805 24505 15845
rect 24545 15805 24555 15845
rect 24595 15805 24605 15845
rect 24645 15805 24655 15845
rect 24695 15805 24705 15845
rect 24745 15805 24755 15845
rect 24795 15805 24805 15845
rect 24845 15805 24855 15845
rect 24895 15805 24905 15845
rect 24945 15805 24955 15845
rect 24995 15805 25005 15845
rect 25045 15805 25055 15845
rect 25095 15805 25105 15845
rect 25145 15805 25155 15845
rect 25195 15805 25205 15845
rect 25245 15805 25255 15845
rect 25295 15805 25305 15845
rect 25345 15805 25355 15845
rect 25395 15805 25405 15845
rect 25445 15805 25455 15845
rect 25495 15805 25505 15845
rect 25545 15805 25555 15845
rect 25595 15805 25605 15845
rect 25645 15805 25655 15845
rect 25695 15805 25705 15845
rect 25745 15805 25755 15845
rect 25795 15805 25805 15845
rect 25845 15805 25855 15845
rect 25895 15805 25905 15845
rect 25945 15805 25955 15845
rect 25995 15805 26005 15845
rect 26045 15805 26055 15845
rect 26095 15805 26105 15845
rect 26145 15805 26155 15845
rect 26195 15805 26205 15845
rect 26245 15805 26255 15845
rect 26295 15805 26305 15845
rect 26345 15805 26355 15845
rect 26395 15805 26405 15845
rect 26445 15805 26455 15845
rect 26495 15805 26505 15845
rect 26545 15805 26555 15845
rect 26595 15805 26605 15845
rect 26645 15805 26655 15845
rect 26695 15805 26705 15845
rect 26745 15805 26755 15845
rect 26795 15805 26805 15845
rect 26845 15805 26855 15845
rect 26895 15805 26905 15845
rect 26945 15805 26955 15845
rect 26995 15805 27005 15845
rect 27045 15805 27055 15845
rect 27095 15805 27105 15845
rect 27145 15805 27155 15845
rect 27195 15805 27205 15845
rect 27245 15805 27255 15845
rect 27295 15805 27305 15845
rect 27345 15805 27355 15845
rect 27395 15805 27405 15845
rect 27445 15805 27455 15845
rect 27495 15805 27505 15845
rect 27545 15805 27555 15845
rect 27595 15805 27605 15845
rect 27645 15805 27655 15845
rect 27695 15805 27705 15845
rect 27745 15805 27755 15845
rect 27795 15805 27805 15845
rect 27845 15805 27855 15845
rect 27895 15805 27905 15845
rect 27945 15805 27955 15845
rect 27995 15805 28005 15845
rect 28045 15805 28055 15845
rect 28095 15805 28105 15845
rect 28145 15805 28155 15845
rect 28195 15805 28205 15845
rect 28245 15805 28255 15845
rect 28295 15805 28305 15845
rect 28345 15805 28355 15845
rect 28395 15805 28405 15845
rect 28445 15805 28455 15845
rect 28495 15805 28505 15845
rect 28545 15805 28555 15845
rect 28595 15805 28605 15845
rect 28645 15805 28655 15845
rect 28695 15805 28705 15845
rect 28745 15805 28755 15845
rect 28795 15805 28805 15845
rect 28845 15805 28855 15845
rect 28895 15805 28905 15845
rect 28945 15805 28955 15845
rect 28995 15805 29005 15845
rect 29045 15805 29055 15845
rect 29095 15805 29105 15845
rect 29145 15805 29155 15845
rect 29195 15805 29205 15845
rect 29245 15805 29255 15845
rect 29295 15805 29305 15845
rect 29345 15805 29355 15845
rect 29395 15805 29405 15845
rect 29445 15805 29455 15845
rect 29495 15805 29505 15845
rect 29545 15805 29555 15845
rect 29595 15805 29605 15845
rect 29645 15805 29655 15845
rect 29695 15805 29705 15845
rect 29745 15805 29755 15845
rect 29795 15805 29805 15845
rect 29845 15805 29855 15845
rect 29895 15805 29905 15845
rect 29945 15805 29955 15845
rect 29995 15805 30005 15845
rect 30045 15805 30055 15845
rect 30095 15805 30105 15845
rect 30145 15805 30155 15845
rect 30195 15805 30205 15845
rect 30245 15805 30255 15845
rect 30295 15805 30305 15845
rect 30345 15805 30355 15845
rect 30395 15805 30405 15845
rect 30445 15805 30455 15845
rect 30495 15805 30505 15845
rect 30545 15805 30555 15845
rect 30595 15805 30605 15845
rect 30645 15805 30655 15845
rect 30695 15805 30705 15845
rect 30745 15805 30755 15845
rect 30795 15805 30805 15845
rect 30845 15805 30855 15845
rect 30895 15805 30905 15845
rect 30945 15805 30955 15845
rect 30995 15805 31005 15845
rect 31045 15805 31055 15845
rect 31095 15805 31105 15845
rect 31145 15805 31155 15845
rect 31195 15805 31205 15845
rect 31245 15805 31255 15845
rect 31295 15805 31305 15845
rect 31345 15805 31355 15845
rect 31395 15805 31405 15845
rect 31445 15805 31455 15845
rect 31495 15805 31505 15845
rect 31545 15805 31555 15845
rect 31595 15805 31605 15845
rect 31645 15805 31655 15845
rect 31695 15805 31705 15845
rect 31745 15805 31755 15845
rect 31795 15805 31805 15845
rect 31845 15805 31855 15845
rect 31895 15805 31905 15845
rect 31945 15805 31955 15845
rect 31995 15805 32005 15845
rect 32045 15805 32055 15845
rect 32095 15805 32105 15845
rect 32145 15805 32155 15845
rect 32195 15805 32205 15845
rect 32245 15805 32255 15845
rect 32295 15805 32305 15845
rect 32345 15805 32355 15845
rect 32395 15805 32405 15845
rect 32445 15805 32455 15845
rect 32495 15805 32505 15845
rect 32545 15805 32555 15845
rect 32595 15805 32605 15845
rect 32645 15805 32655 15845
rect 32695 15805 32705 15845
rect 32745 15805 32755 15845
rect 32795 15805 32805 15845
rect 32845 15805 32855 15845
rect 32895 15805 32905 15845
rect 32945 15805 32955 15845
rect 32995 15805 33005 15845
rect 33045 15805 33055 15845
rect 33095 15805 33105 15845
rect 33145 15805 33155 15845
rect 33195 15805 33205 15845
rect 33245 15805 33255 15845
rect 33295 15805 33305 15845
rect 33345 15805 33355 15845
rect 33395 15805 33405 15845
rect 33445 15805 33455 15845
rect 33495 15805 33505 15845
rect 33545 15805 33555 15845
rect 33595 15805 33605 15845
rect 33645 15805 33655 15845
rect 33695 15805 33705 15845
rect 33745 15805 33755 15845
rect 33795 15805 33805 15845
rect 33845 15805 33855 15845
rect 33895 15805 33905 15845
rect 33945 15805 33955 15845
rect 33995 15805 34005 15845
rect 34045 15805 34055 15845
rect 34095 15805 34105 15845
rect 34145 15805 34155 15845
rect 34195 15805 34205 15845
rect 34245 15805 34255 15845
rect 34295 15805 34305 15845
rect 34345 15805 34355 15845
rect 34395 15805 34405 15845
rect 34445 15805 34455 15845
rect 34495 15805 34505 15845
rect 34545 15805 34555 15845
rect 34595 15805 34605 15845
rect 34645 15805 34655 15845
rect 34695 15805 34705 15845
rect 34745 15805 34755 15845
rect 34795 15805 34805 15845
rect 34845 15805 34855 15845
rect 34895 15805 34905 15845
rect 34945 15805 34955 15845
rect 34995 15805 35005 15845
rect 35045 15805 35055 15845
rect 35095 15805 35105 15845
rect 35145 15805 35155 15845
rect 35195 15805 35205 15845
rect 35245 15805 35255 15845
rect 35295 15805 35305 15845
rect 35345 15805 35355 15845
rect 35395 15805 35405 15845
rect 35445 15805 35455 15845
rect 35495 15805 35505 15845
rect 35545 15805 35555 15845
rect 35595 15805 35605 15845
rect 35645 15805 35655 15845
rect 35695 15805 35705 15845
rect 35745 15805 35755 15845
rect 35795 15805 35805 15845
rect 35845 15805 35855 15845
rect 35895 15805 35905 15845
rect 35945 15805 35955 15845
rect 35995 15805 36005 15845
rect 36045 15805 36055 15845
rect 36095 15805 36105 15845
rect 36145 15805 36155 15845
rect 36195 15805 36205 15845
rect 36245 15805 36255 15845
rect 36295 15805 36305 15845
rect 36345 15805 36355 15845
rect 36395 15805 36405 15845
rect 36445 15805 36455 15845
rect 36495 15805 36505 15845
rect 36545 15805 36555 15845
rect 36595 15805 36605 15845
rect 36645 15805 36655 15845
rect 36695 15805 36705 15845
rect 36745 15805 36755 15845
rect 36795 15805 36805 15845
rect 36845 15805 36855 15845
rect 36895 15805 36905 15845
rect 36945 15805 36955 15845
rect 36995 15805 37005 15845
rect 37045 15805 37055 15845
rect 37095 15805 37105 15845
rect 37145 15805 37155 15845
rect 37195 15805 37205 15845
rect 37245 15805 37255 15845
rect 37295 15805 37305 15845
rect 37345 15805 37355 15845
rect 37395 15805 37405 15845
rect 37445 15805 37455 15845
rect 37495 15805 37505 15845
rect 37545 15805 37555 15845
rect 37595 15805 37605 15845
rect 37645 15805 37655 15845
rect 37695 15805 37705 15845
rect 37745 15805 37755 15845
rect 37795 15805 37805 15845
rect 37845 15805 37855 15845
rect 37895 15805 37905 15845
rect 37945 15805 37955 15845
rect 37995 15805 38005 15845
rect 38045 15805 38055 15845
rect 38095 15805 38105 15845
rect 38145 15805 38155 15845
rect 38195 15805 38205 15845
rect 38245 15805 38255 15845
rect 38295 15805 38305 15845
rect 38345 15805 38355 15845
rect 38395 15805 38405 15845
rect 38445 15805 38455 15845
rect 38495 15805 38505 15845
rect 38545 15805 38555 15845
rect 38595 15805 38605 15845
rect 38645 15805 38655 15845
rect 38695 15805 38705 15845
rect 38745 15805 38755 15845
rect 38795 15805 38805 15845
rect 38845 15805 38855 15845
rect 38895 15805 38905 15845
rect 38945 15805 38955 15845
rect 38995 15805 39005 15845
rect 39045 15805 39055 15845
rect 39095 15805 39105 15845
rect 39145 15805 39155 15845
rect 39195 15805 39205 15845
rect 39245 15805 39255 15845
rect 39295 15805 39305 15845
rect 39345 15805 39355 15845
rect 39395 15805 39405 15845
rect 39445 15805 39455 15845
rect 39495 15805 39505 15845
rect 39545 15805 39555 15845
rect 39595 15805 39605 15845
rect 39645 15805 39655 15845
rect 39695 15805 39705 15845
rect 39745 15805 39750 15845
rect 0 15800 39750 15805
rect -3500 15745 -50 15750
rect -3500 15705 -3495 15745
rect -3455 15705 -3295 15745
rect -3255 15705 -3095 15745
rect -3055 15705 -1595 15745
rect -1555 15705 -1195 15745
rect -1155 15705 -1095 15745
rect -1055 15705 -995 15745
rect -955 15705 -895 15745
rect -855 15705 -695 15745
rect -655 15705 -595 15745
rect -555 15705 -495 15745
rect -455 15705 -295 15745
rect -255 15705 -195 15745
rect -155 15705 -95 15745
rect -55 15705 -50 15745
rect -3500 15700 -50 15705
rect 0 15745 40900 15750
rect 0 15705 5 15745
rect 45 15705 55 15745
rect 95 15705 105 15745
rect 145 15705 155 15745
rect 195 15705 205 15745
rect 245 15705 255 15745
rect 295 15705 305 15745
rect 345 15705 355 15745
rect 395 15705 405 15745
rect 445 15705 455 15745
rect 495 15705 505 15745
rect 545 15705 555 15745
rect 595 15705 605 15745
rect 645 15705 655 15745
rect 695 15705 705 15745
rect 745 15705 755 15745
rect 795 15705 805 15745
rect 845 15705 855 15745
rect 895 15705 905 15745
rect 945 15705 955 15745
rect 995 15705 1005 15745
rect 1045 15705 1055 15745
rect 1095 15705 1105 15745
rect 1145 15705 1155 15745
rect 1195 15705 1205 15745
rect 1245 15705 1255 15745
rect 1295 15705 1305 15745
rect 1345 15705 1355 15745
rect 1395 15705 1405 15745
rect 1445 15705 1455 15745
rect 1495 15705 1505 15745
rect 1545 15705 1555 15745
rect 1595 15705 1605 15745
rect 1645 15705 1655 15745
rect 1695 15705 1705 15745
rect 1745 15705 1755 15745
rect 1795 15705 1805 15745
rect 1845 15705 1855 15745
rect 1895 15705 1905 15745
rect 1945 15705 1955 15745
rect 1995 15705 2005 15745
rect 2045 15705 2055 15745
rect 2095 15705 2105 15745
rect 2145 15705 2155 15745
rect 2195 15705 2205 15745
rect 2245 15705 2255 15745
rect 2295 15705 2305 15745
rect 2345 15705 2355 15745
rect 2395 15705 2405 15745
rect 2445 15705 2455 15745
rect 2495 15705 2505 15745
rect 2545 15705 2555 15745
rect 2595 15705 2605 15745
rect 2645 15705 2655 15745
rect 2695 15705 2705 15745
rect 2745 15705 2755 15745
rect 2795 15705 2805 15745
rect 2845 15705 2855 15745
rect 2895 15705 2905 15745
rect 2945 15705 2955 15745
rect 2995 15705 3005 15745
rect 3045 15705 3055 15745
rect 3095 15705 3105 15745
rect 3145 15705 3155 15745
rect 3195 15705 3205 15745
rect 3245 15705 3255 15745
rect 3295 15705 3305 15745
rect 3345 15705 3355 15745
rect 3395 15705 3405 15745
rect 3445 15705 3455 15745
rect 3495 15705 3505 15745
rect 3545 15705 3555 15745
rect 3595 15705 3605 15745
rect 3645 15705 3655 15745
rect 3695 15705 3705 15745
rect 3745 15705 3755 15745
rect 3795 15705 3805 15745
rect 3845 15705 3855 15745
rect 3895 15705 3905 15745
rect 3945 15705 3955 15745
rect 3995 15705 4005 15745
rect 4045 15705 4055 15745
rect 4095 15705 4105 15745
rect 4145 15705 4155 15745
rect 4195 15705 4205 15745
rect 4245 15705 4255 15745
rect 4295 15705 4305 15745
rect 4345 15705 4355 15745
rect 4395 15705 4405 15745
rect 4445 15705 4455 15745
rect 4495 15705 4505 15745
rect 4545 15705 4555 15745
rect 4595 15705 4605 15745
rect 4645 15705 4655 15745
rect 4695 15705 4705 15745
rect 4745 15705 4755 15745
rect 4795 15705 4805 15745
rect 4845 15705 4855 15745
rect 4895 15705 4905 15745
rect 4945 15705 4955 15745
rect 4995 15705 5005 15745
rect 5045 15705 5055 15745
rect 5095 15705 5105 15745
rect 5145 15705 5155 15745
rect 5195 15705 5205 15745
rect 5245 15705 5255 15745
rect 5295 15705 5305 15745
rect 5345 15705 5355 15745
rect 5395 15705 5405 15745
rect 5445 15705 5455 15745
rect 5495 15705 5505 15745
rect 5545 15705 5555 15745
rect 5595 15705 5605 15745
rect 5645 15705 5655 15745
rect 5695 15705 5705 15745
rect 5745 15705 5755 15745
rect 5795 15705 5805 15745
rect 5845 15705 5855 15745
rect 5895 15705 5905 15745
rect 5945 15705 5955 15745
rect 5995 15705 6005 15745
rect 6045 15705 6055 15745
rect 6095 15705 6105 15745
rect 6145 15705 6155 15745
rect 6195 15705 6205 15745
rect 6245 15705 6255 15745
rect 6295 15705 6305 15745
rect 6345 15705 6355 15745
rect 6395 15705 6405 15745
rect 6445 15705 6455 15745
rect 6495 15705 6505 15745
rect 6545 15705 6555 15745
rect 6595 15705 6605 15745
rect 6645 15705 6655 15745
rect 6695 15705 6705 15745
rect 6745 15705 6755 15745
rect 6795 15705 6805 15745
rect 6845 15705 6855 15745
rect 6895 15705 6905 15745
rect 6945 15705 6955 15745
rect 6995 15705 7005 15745
rect 7045 15705 7055 15745
rect 7095 15705 7105 15745
rect 7145 15705 7155 15745
rect 7195 15705 7205 15745
rect 7245 15705 7255 15745
rect 7295 15705 7305 15745
rect 7345 15705 7355 15745
rect 7395 15705 7405 15745
rect 7445 15705 7455 15745
rect 7495 15705 7505 15745
rect 7545 15705 7555 15745
rect 7595 15705 7605 15745
rect 7645 15705 7655 15745
rect 7695 15705 7705 15745
rect 7745 15705 7755 15745
rect 7795 15705 7805 15745
rect 7845 15705 7855 15745
rect 7895 15705 7905 15745
rect 7945 15705 7955 15745
rect 7995 15705 8005 15745
rect 8045 15705 8055 15745
rect 8095 15705 8105 15745
rect 8145 15705 8155 15745
rect 8195 15705 8205 15745
rect 8245 15705 8255 15745
rect 8295 15705 8305 15745
rect 8345 15705 8355 15745
rect 8395 15705 8405 15745
rect 8445 15705 8455 15745
rect 8495 15705 8505 15745
rect 8545 15705 8555 15745
rect 8595 15705 8605 15745
rect 8645 15705 8655 15745
rect 8695 15705 8705 15745
rect 8745 15705 8755 15745
rect 8795 15705 8805 15745
rect 8845 15705 8855 15745
rect 8895 15705 8905 15745
rect 8945 15705 8955 15745
rect 8995 15705 9005 15745
rect 9045 15705 9055 15745
rect 9095 15705 9105 15745
rect 9145 15705 9155 15745
rect 9195 15705 9205 15745
rect 9245 15705 9255 15745
rect 9295 15705 9305 15745
rect 9345 15705 9355 15745
rect 9395 15705 9405 15745
rect 9445 15705 9455 15745
rect 9495 15705 9505 15745
rect 9545 15705 9555 15745
rect 9595 15705 9605 15745
rect 9645 15705 9655 15745
rect 9695 15705 9705 15745
rect 9745 15705 9755 15745
rect 9795 15705 9805 15745
rect 9845 15705 9855 15745
rect 9895 15705 9905 15745
rect 9945 15705 9955 15745
rect 9995 15705 10005 15745
rect 10045 15705 10055 15745
rect 10095 15705 10105 15745
rect 10145 15705 10155 15745
rect 10195 15705 10205 15745
rect 10245 15705 10255 15745
rect 10295 15705 10305 15745
rect 10345 15705 10355 15745
rect 10395 15705 10405 15745
rect 10445 15705 10455 15745
rect 10495 15705 10505 15745
rect 10545 15705 10555 15745
rect 10595 15705 10605 15745
rect 10645 15705 10655 15745
rect 10695 15705 10705 15745
rect 10745 15705 10755 15745
rect 10795 15705 10805 15745
rect 10845 15705 10855 15745
rect 10895 15705 10905 15745
rect 10945 15705 10955 15745
rect 10995 15705 11005 15745
rect 11045 15705 11055 15745
rect 11095 15705 11105 15745
rect 11145 15705 11155 15745
rect 11195 15705 11205 15745
rect 11245 15705 11255 15745
rect 11295 15705 11305 15745
rect 11345 15705 11355 15745
rect 11395 15705 11405 15745
rect 11445 15705 11455 15745
rect 11495 15705 11505 15745
rect 11545 15705 11555 15745
rect 11595 15705 11605 15745
rect 11645 15705 11655 15745
rect 11695 15705 11705 15745
rect 11745 15705 11755 15745
rect 11795 15705 11805 15745
rect 11845 15705 11855 15745
rect 11895 15705 11905 15745
rect 11945 15705 11955 15745
rect 11995 15705 12005 15745
rect 12045 15705 12055 15745
rect 12095 15705 12105 15745
rect 12145 15705 12155 15745
rect 12195 15705 12205 15745
rect 12245 15705 12255 15745
rect 12295 15705 12305 15745
rect 12345 15705 12355 15745
rect 12395 15705 12405 15745
rect 12445 15705 12455 15745
rect 12495 15705 12505 15745
rect 12545 15705 12555 15745
rect 12595 15705 12605 15745
rect 12645 15705 12655 15745
rect 12695 15705 12705 15745
rect 12745 15705 12755 15745
rect 12795 15705 12805 15745
rect 12845 15705 12855 15745
rect 12895 15705 12905 15745
rect 12945 15705 12955 15745
rect 12995 15705 13005 15745
rect 13045 15705 13055 15745
rect 13095 15705 13105 15745
rect 13145 15705 13155 15745
rect 13195 15705 13205 15745
rect 13245 15705 13255 15745
rect 13295 15705 13305 15745
rect 13345 15705 13355 15745
rect 13395 15705 13405 15745
rect 13445 15705 13455 15745
rect 13495 15705 13505 15745
rect 13545 15705 13555 15745
rect 13595 15705 13605 15745
rect 13645 15705 13655 15745
rect 13695 15705 13705 15745
rect 13745 15705 13755 15745
rect 13795 15705 13805 15745
rect 13845 15705 13855 15745
rect 13895 15705 13905 15745
rect 13945 15705 13955 15745
rect 13995 15705 14005 15745
rect 14045 15705 14055 15745
rect 14095 15705 14105 15745
rect 14145 15705 14155 15745
rect 14195 15705 14205 15745
rect 14245 15705 14255 15745
rect 14295 15705 14305 15745
rect 14345 15705 14355 15745
rect 14395 15705 14405 15745
rect 14445 15705 14455 15745
rect 14495 15705 14505 15745
rect 14545 15705 14555 15745
rect 14595 15705 14605 15745
rect 14645 15705 14655 15745
rect 14695 15705 14705 15745
rect 14745 15705 14755 15745
rect 14795 15705 14805 15745
rect 14845 15705 14855 15745
rect 14895 15705 14905 15745
rect 14945 15705 14955 15745
rect 14995 15705 15005 15745
rect 15045 15705 15055 15745
rect 15095 15705 15105 15745
rect 15145 15705 15155 15745
rect 15195 15705 15205 15745
rect 15245 15705 15255 15745
rect 15295 15705 15305 15745
rect 15345 15705 15355 15745
rect 15395 15705 15405 15745
rect 15445 15705 15455 15745
rect 15495 15705 15505 15745
rect 15545 15705 15555 15745
rect 15595 15705 15605 15745
rect 15645 15705 15655 15745
rect 15695 15705 15705 15745
rect 15745 15705 15755 15745
rect 15795 15705 15805 15745
rect 15845 15705 15855 15745
rect 15895 15705 15905 15745
rect 15945 15705 15955 15745
rect 15995 15705 16005 15745
rect 16045 15705 16055 15745
rect 16095 15705 16105 15745
rect 16145 15705 16155 15745
rect 16195 15705 16205 15745
rect 16245 15705 16255 15745
rect 16295 15705 16305 15745
rect 16345 15705 16355 15745
rect 16395 15705 16405 15745
rect 16445 15705 16455 15745
rect 16495 15705 16505 15745
rect 16545 15705 16555 15745
rect 16595 15705 16605 15745
rect 16645 15705 16655 15745
rect 16695 15705 16705 15745
rect 16745 15705 16755 15745
rect 16795 15705 16805 15745
rect 16845 15705 16855 15745
rect 16895 15705 16905 15745
rect 16945 15705 16955 15745
rect 16995 15705 17005 15745
rect 17045 15705 17055 15745
rect 17095 15705 17105 15745
rect 17145 15705 17155 15745
rect 17195 15705 17205 15745
rect 17245 15705 17255 15745
rect 17295 15705 17305 15745
rect 17345 15705 17355 15745
rect 17395 15705 17405 15745
rect 17445 15705 17455 15745
rect 17495 15705 17505 15745
rect 17545 15705 17555 15745
rect 17595 15705 17605 15745
rect 17645 15705 17655 15745
rect 17695 15705 17705 15745
rect 17745 15705 17755 15745
rect 17795 15705 17805 15745
rect 17845 15705 17855 15745
rect 17895 15705 17905 15745
rect 17945 15705 17955 15745
rect 17995 15705 18005 15745
rect 18045 15705 18055 15745
rect 18095 15705 18105 15745
rect 18145 15705 18155 15745
rect 18195 15705 18205 15745
rect 18245 15705 18255 15745
rect 18295 15705 18305 15745
rect 18345 15705 18355 15745
rect 18395 15705 18405 15745
rect 18445 15705 18455 15745
rect 18495 15705 18505 15745
rect 18545 15705 18555 15745
rect 18595 15705 18605 15745
rect 18645 15705 18655 15745
rect 18695 15705 18705 15745
rect 18745 15705 18755 15745
rect 18795 15705 18805 15745
rect 18845 15705 18855 15745
rect 18895 15705 18905 15745
rect 18945 15705 18955 15745
rect 18995 15705 19005 15745
rect 19045 15705 19055 15745
rect 19095 15705 19105 15745
rect 19145 15705 19155 15745
rect 19195 15705 19205 15745
rect 19245 15705 19255 15745
rect 19295 15705 19305 15745
rect 19345 15705 19355 15745
rect 19395 15705 19405 15745
rect 19445 15705 19455 15745
rect 19495 15705 19505 15745
rect 19545 15705 19555 15745
rect 19595 15705 19605 15745
rect 19645 15705 19655 15745
rect 19695 15705 19705 15745
rect 19745 15705 19755 15745
rect 19795 15705 19805 15745
rect 19845 15705 19855 15745
rect 19895 15705 19905 15745
rect 19945 15705 19955 15745
rect 19995 15705 20005 15745
rect 20045 15705 20055 15745
rect 20095 15705 20105 15745
rect 20145 15705 20155 15745
rect 20195 15705 20205 15745
rect 20245 15705 20255 15745
rect 20295 15705 20305 15745
rect 20345 15705 20355 15745
rect 20395 15705 20405 15745
rect 20445 15705 20455 15745
rect 20495 15705 20505 15745
rect 20545 15705 20555 15745
rect 20595 15705 20605 15745
rect 20645 15705 20655 15745
rect 20695 15705 20705 15745
rect 20745 15705 20755 15745
rect 20795 15705 20805 15745
rect 20845 15705 20855 15745
rect 20895 15705 20905 15745
rect 20945 15705 20955 15745
rect 20995 15705 21005 15745
rect 21045 15705 21055 15745
rect 21095 15705 21105 15745
rect 21145 15705 21155 15745
rect 21195 15705 21205 15745
rect 21245 15705 21255 15745
rect 21295 15705 21305 15745
rect 21345 15705 21355 15745
rect 21395 15705 21405 15745
rect 21445 15705 21455 15745
rect 21495 15705 21505 15745
rect 21545 15705 21555 15745
rect 21595 15705 21605 15745
rect 21645 15705 21655 15745
rect 21695 15705 21705 15745
rect 21745 15705 21755 15745
rect 21795 15705 21805 15745
rect 21845 15705 21855 15745
rect 21895 15705 21905 15745
rect 21945 15705 21955 15745
rect 21995 15705 22005 15745
rect 22045 15705 22055 15745
rect 22095 15705 22105 15745
rect 22145 15705 22155 15745
rect 22195 15705 22205 15745
rect 22245 15705 22255 15745
rect 22295 15705 22305 15745
rect 22345 15705 22355 15745
rect 22395 15705 22405 15745
rect 22445 15705 22455 15745
rect 22495 15705 22505 15745
rect 22545 15705 22555 15745
rect 22595 15705 22605 15745
rect 22645 15705 22655 15745
rect 22695 15705 22705 15745
rect 22745 15705 22755 15745
rect 22795 15705 22805 15745
rect 22845 15705 22855 15745
rect 22895 15705 22905 15745
rect 22945 15705 22955 15745
rect 22995 15705 23005 15745
rect 23045 15705 23055 15745
rect 23095 15705 23105 15745
rect 23145 15705 23155 15745
rect 23195 15705 23205 15745
rect 23245 15705 23255 15745
rect 23295 15705 23305 15745
rect 23345 15705 23355 15745
rect 23395 15705 23405 15745
rect 23445 15705 23455 15745
rect 23495 15705 23505 15745
rect 23545 15705 23555 15745
rect 23595 15705 23605 15745
rect 23645 15705 23655 15745
rect 23695 15705 23705 15745
rect 23745 15705 23755 15745
rect 23795 15705 23805 15745
rect 23845 15705 23855 15745
rect 23895 15705 23905 15745
rect 23945 15705 23955 15745
rect 23995 15705 24005 15745
rect 24045 15705 24055 15745
rect 24095 15705 24105 15745
rect 24145 15705 24155 15745
rect 24195 15705 24205 15745
rect 24245 15705 24255 15745
rect 24295 15705 24305 15745
rect 24345 15705 24355 15745
rect 24395 15705 24405 15745
rect 24445 15705 24455 15745
rect 24495 15705 24505 15745
rect 24545 15705 24555 15745
rect 24595 15705 24605 15745
rect 24645 15705 24655 15745
rect 24695 15705 24705 15745
rect 24745 15705 24755 15745
rect 24795 15705 24805 15745
rect 24845 15705 24855 15745
rect 24895 15705 24905 15745
rect 24945 15705 24955 15745
rect 24995 15705 25005 15745
rect 25045 15705 25055 15745
rect 25095 15705 25105 15745
rect 25145 15705 25155 15745
rect 25195 15705 25205 15745
rect 25245 15705 25255 15745
rect 25295 15705 25305 15745
rect 25345 15705 25355 15745
rect 25395 15705 25405 15745
rect 25445 15705 25455 15745
rect 25495 15705 25505 15745
rect 25545 15705 25555 15745
rect 25595 15705 25605 15745
rect 25645 15705 25655 15745
rect 25695 15705 25705 15745
rect 25745 15705 25755 15745
rect 25795 15705 25805 15745
rect 25845 15705 25855 15745
rect 25895 15705 25905 15745
rect 25945 15705 25955 15745
rect 25995 15705 26005 15745
rect 26045 15705 26055 15745
rect 26095 15705 26105 15745
rect 26145 15705 26155 15745
rect 26195 15705 26205 15745
rect 26245 15705 26255 15745
rect 26295 15705 26305 15745
rect 26345 15705 26355 15745
rect 26395 15705 26405 15745
rect 26445 15705 26455 15745
rect 26495 15705 26505 15745
rect 26545 15705 26555 15745
rect 26595 15705 26605 15745
rect 26645 15705 26655 15745
rect 26695 15705 26705 15745
rect 26745 15705 26755 15745
rect 26795 15705 26805 15745
rect 26845 15705 26855 15745
rect 26895 15705 26905 15745
rect 26945 15705 26955 15745
rect 26995 15705 27005 15745
rect 27045 15705 27055 15745
rect 27095 15705 27105 15745
rect 27145 15705 27155 15745
rect 27195 15705 27205 15745
rect 27245 15705 27255 15745
rect 27295 15705 27305 15745
rect 27345 15705 27355 15745
rect 27395 15705 27405 15745
rect 27445 15705 27455 15745
rect 27495 15705 27505 15745
rect 27545 15705 27555 15745
rect 27595 15705 27605 15745
rect 27645 15705 27655 15745
rect 27695 15705 27705 15745
rect 27745 15705 27755 15745
rect 27795 15705 27805 15745
rect 27845 15705 27855 15745
rect 27895 15705 27905 15745
rect 27945 15705 27955 15745
rect 27995 15705 28005 15745
rect 28045 15705 28055 15745
rect 28095 15705 28105 15745
rect 28145 15705 28155 15745
rect 28195 15705 28205 15745
rect 28245 15705 28255 15745
rect 28295 15705 28305 15745
rect 28345 15705 28355 15745
rect 28395 15705 28405 15745
rect 28445 15705 28455 15745
rect 28495 15705 28505 15745
rect 28545 15705 28555 15745
rect 28595 15705 28605 15745
rect 28645 15705 28655 15745
rect 28695 15705 28705 15745
rect 28745 15705 28755 15745
rect 28795 15705 28805 15745
rect 28845 15705 28855 15745
rect 28895 15705 28905 15745
rect 28945 15705 28955 15745
rect 28995 15705 29005 15745
rect 29045 15705 29055 15745
rect 29095 15705 29105 15745
rect 29145 15705 29155 15745
rect 29195 15705 29205 15745
rect 29245 15705 29255 15745
rect 29295 15705 29305 15745
rect 29345 15705 29355 15745
rect 29395 15705 29405 15745
rect 29445 15705 29455 15745
rect 29495 15705 29505 15745
rect 29545 15705 29555 15745
rect 29595 15705 29605 15745
rect 29645 15705 29655 15745
rect 29695 15705 29705 15745
rect 29745 15705 29755 15745
rect 29795 15705 29805 15745
rect 29845 15705 29855 15745
rect 29895 15705 29905 15745
rect 29945 15705 29955 15745
rect 29995 15705 30005 15745
rect 30045 15705 30055 15745
rect 30095 15705 30105 15745
rect 30145 15705 30155 15745
rect 30195 15705 30205 15745
rect 30245 15705 30255 15745
rect 30295 15705 30305 15745
rect 30345 15705 30355 15745
rect 30395 15705 30405 15745
rect 30445 15705 30455 15745
rect 30495 15705 30505 15745
rect 30545 15705 30555 15745
rect 30595 15705 30605 15745
rect 30645 15705 30655 15745
rect 30695 15705 30705 15745
rect 30745 15705 30755 15745
rect 30795 15705 30805 15745
rect 30845 15705 30855 15745
rect 30895 15705 30905 15745
rect 30945 15705 30955 15745
rect 30995 15705 31005 15745
rect 31045 15705 31055 15745
rect 31095 15705 31105 15745
rect 31145 15705 31155 15745
rect 31195 15705 31205 15745
rect 31245 15705 31255 15745
rect 31295 15705 31305 15745
rect 31345 15705 31355 15745
rect 31395 15705 31405 15745
rect 31445 15705 31455 15745
rect 31495 15705 31505 15745
rect 31545 15705 31555 15745
rect 31595 15705 31605 15745
rect 31645 15705 31655 15745
rect 31695 15705 31705 15745
rect 31745 15705 31755 15745
rect 31795 15705 31805 15745
rect 31845 15705 31855 15745
rect 31895 15705 31905 15745
rect 31945 15705 31955 15745
rect 31995 15705 32005 15745
rect 32045 15705 32055 15745
rect 32095 15705 32105 15745
rect 32145 15705 32155 15745
rect 32195 15705 32205 15745
rect 32245 15705 32255 15745
rect 32295 15705 32305 15745
rect 32345 15705 32355 15745
rect 32395 15705 32405 15745
rect 32445 15705 32455 15745
rect 32495 15705 32505 15745
rect 32545 15705 32555 15745
rect 32595 15705 32605 15745
rect 32645 15705 32655 15745
rect 32695 15705 32705 15745
rect 32745 15705 32755 15745
rect 32795 15705 32805 15745
rect 32845 15705 32855 15745
rect 32895 15705 32905 15745
rect 32945 15705 32955 15745
rect 32995 15705 33005 15745
rect 33045 15705 33055 15745
rect 33095 15705 33105 15745
rect 33145 15705 33155 15745
rect 33195 15705 33205 15745
rect 33245 15705 33255 15745
rect 33295 15705 33305 15745
rect 33345 15705 33355 15745
rect 33395 15705 33405 15745
rect 33445 15705 33455 15745
rect 33495 15705 33505 15745
rect 33545 15705 33555 15745
rect 33595 15705 33605 15745
rect 33645 15705 33655 15745
rect 33695 15705 33705 15745
rect 33745 15705 33755 15745
rect 33795 15705 33805 15745
rect 33845 15705 33855 15745
rect 33895 15705 33905 15745
rect 33945 15705 33955 15745
rect 33995 15705 34005 15745
rect 34045 15705 34055 15745
rect 34095 15705 34105 15745
rect 34145 15705 34155 15745
rect 34195 15705 34205 15745
rect 34245 15705 34255 15745
rect 34295 15705 34305 15745
rect 34345 15705 34355 15745
rect 34395 15705 34405 15745
rect 34445 15705 34455 15745
rect 34495 15705 34505 15745
rect 34545 15705 34555 15745
rect 34595 15705 34605 15745
rect 34645 15705 34655 15745
rect 34695 15705 34705 15745
rect 34745 15705 34755 15745
rect 34795 15705 34805 15745
rect 34845 15705 34855 15745
rect 34895 15705 34905 15745
rect 34945 15705 34955 15745
rect 34995 15705 35005 15745
rect 35045 15705 35055 15745
rect 35095 15705 35105 15745
rect 35145 15705 35155 15745
rect 35195 15705 35205 15745
rect 35245 15705 35255 15745
rect 35295 15705 35305 15745
rect 35345 15705 35355 15745
rect 35395 15705 35405 15745
rect 35445 15705 35455 15745
rect 35495 15705 35505 15745
rect 35545 15705 35555 15745
rect 35595 15705 35605 15745
rect 35645 15705 35655 15745
rect 35695 15705 35705 15745
rect 35745 15705 35755 15745
rect 35795 15705 35805 15745
rect 35845 15705 35855 15745
rect 35895 15705 35905 15745
rect 35945 15705 35955 15745
rect 35995 15705 36005 15745
rect 36045 15705 36055 15745
rect 36095 15705 36105 15745
rect 36145 15705 36155 15745
rect 36195 15705 36205 15745
rect 36245 15705 36255 15745
rect 36295 15705 36305 15745
rect 36345 15705 36355 15745
rect 36395 15705 36405 15745
rect 36445 15705 36455 15745
rect 36495 15705 36505 15745
rect 36545 15705 36555 15745
rect 36595 15705 36605 15745
rect 36645 15705 36655 15745
rect 36695 15705 36705 15745
rect 36745 15705 36755 15745
rect 36795 15705 36805 15745
rect 36845 15705 36855 15745
rect 36895 15705 36905 15745
rect 36945 15705 36955 15745
rect 36995 15705 37005 15745
rect 37045 15705 37055 15745
rect 37095 15705 37105 15745
rect 37145 15705 37155 15745
rect 37195 15705 37205 15745
rect 37245 15705 37255 15745
rect 37295 15705 37305 15745
rect 37345 15705 37355 15745
rect 37395 15705 37405 15745
rect 37445 15705 37455 15745
rect 37495 15705 37505 15745
rect 37545 15705 37555 15745
rect 37595 15705 37605 15745
rect 37645 15705 37655 15745
rect 37695 15705 37705 15745
rect 37745 15705 37755 15745
rect 37795 15705 37805 15745
rect 37845 15705 37855 15745
rect 37895 15705 37905 15745
rect 37945 15705 37955 15745
rect 37995 15705 38005 15745
rect 38045 15705 38055 15745
rect 38095 15705 38105 15745
rect 38145 15705 38155 15745
rect 38195 15705 38205 15745
rect 38245 15705 38255 15745
rect 38295 15705 38305 15745
rect 38345 15705 38355 15745
rect 38395 15705 38405 15745
rect 38445 15705 38455 15745
rect 38495 15705 38505 15745
rect 38545 15705 38555 15745
rect 38595 15705 38605 15745
rect 38645 15705 38655 15745
rect 38695 15705 38705 15745
rect 38745 15705 38755 15745
rect 38795 15705 38805 15745
rect 38845 15705 38855 15745
rect 38895 15705 38905 15745
rect 38945 15705 38955 15745
rect 38995 15705 39005 15745
rect 39045 15705 39055 15745
rect 39095 15705 39105 15745
rect 39145 15705 39155 15745
rect 39195 15705 39205 15745
rect 39245 15705 39255 15745
rect 39295 15705 39305 15745
rect 39345 15705 39355 15745
rect 39395 15705 39405 15745
rect 39445 15705 39455 15745
rect 39495 15705 39505 15745
rect 39545 15705 39555 15745
rect 39595 15705 39605 15745
rect 39645 15705 39655 15745
rect 39695 15705 39705 15745
rect 39745 15705 39905 15745
rect 39945 15705 39955 15745
rect 39995 15705 40005 15745
rect 40045 15705 40055 15745
rect 40095 15705 40105 15745
rect 40145 15705 40155 15745
rect 40195 15705 40205 15745
rect 40245 15705 40255 15745
rect 40295 15705 40305 15745
rect 40345 15705 40355 15745
rect 40395 15705 40405 15745
rect 40445 15705 40455 15745
rect 40495 15705 40505 15745
rect 40545 15705 40555 15745
rect 40595 15705 40605 15745
rect 40645 15705 40655 15745
rect 40695 15705 40705 15745
rect 40745 15705 40755 15745
rect 40795 15705 40805 15745
rect 40845 15705 40855 15745
rect 40895 15705 40900 15745
rect 0 15700 40900 15705
rect -3500 15345 0 15350
rect -3500 15305 -3495 15345
rect -3455 15305 -3295 15345
rect -3255 15305 -3095 15345
rect -3055 15305 -1595 15345
rect -1555 15305 -1095 15345
rect -1055 15305 -895 15345
rect -855 15305 -695 15345
rect -655 15305 -495 15345
rect -455 15305 -295 15345
rect -255 15305 -95 15345
rect -55 15305 0 15345
rect -3500 15295 0 15305
rect -3500 15255 -3495 15295
rect -3455 15255 -3295 15295
rect -3255 15255 -3095 15295
rect -3055 15255 -1595 15295
rect -1555 15255 -1095 15295
rect -1055 15255 -895 15295
rect -855 15255 -695 15295
rect -655 15255 -495 15295
rect -455 15255 -295 15295
rect -255 15255 -95 15295
rect -55 15255 0 15295
rect -3500 15245 0 15255
rect -3500 15205 -3495 15245
rect -3455 15205 -3295 15245
rect -3255 15205 -3095 15245
rect -3055 15205 -1595 15245
rect -1555 15205 -1095 15245
rect -1055 15205 -895 15245
rect -855 15205 -695 15245
rect -655 15205 -495 15245
rect -455 15205 -295 15245
rect -255 15205 -95 15245
rect -55 15205 0 15245
rect -3500 15200 0 15205
rect -200 14645 0 14650
rect -200 14605 -195 14645
rect -155 14605 0 14645
rect -200 14600 0 14605
rect -400 14245 0 14250
rect -400 14205 -395 14245
rect -355 14205 0 14245
rect -400 14200 0 14205
rect -600 14045 0 14050
rect -600 14005 -595 14045
rect -555 14005 0 14045
rect -600 14000 0 14005
rect -3500 13645 0 13650
rect -3500 13605 -3495 13645
rect -3455 13605 -3295 13645
rect -3255 13605 -3095 13645
rect -3055 13605 -1595 13645
rect -1555 13605 -1095 13645
rect -1055 13605 -895 13645
rect -855 13605 -695 13645
rect -655 13605 -495 13645
rect -455 13605 -295 13645
rect -255 13605 -95 13645
rect -55 13605 0 13645
rect -3500 13595 0 13605
rect -3500 13555 -3495 13595
rect -3455 13555 -3295 13595
rect -3255 13555 -3095 13595
rect -3055 13555 -1595 13595
rect -1555 13555 -1095 13595
rect -1055 13555 -895 13595
rect -855 13555 -695 13595
rect -655 13555 -495 13595
rect -455 13555 -295 13595
rect -255 13555 -95 13595
rect -55 13555 0 13595
rect -3500 13545 0 13555
rect -3500 13505 -3495 13545
rect -3455 13505 -3295 13545
rect -3255 13505 -3095 13545
rect -3055 13505 -1595 13545
rect -1555 13505 -1095 13545
rect -1055 13505 -895 13545
rect -855 13505 -695 13545
rect -655 13505 -495 13545
rect -455 13505 -295 13545
rect -255 13505 -95 13545
rect -55 13505 0 13545
rect -3500 13500 0 13505
rect -800 13145 0 13150
rect -800 13105 -795 13145
rect -755 13105 0 13145
rect -800 13100 0 13105
rect -1000 12945 0 12950
rect -1000 12905 -995 12945
rect -955 12905 0 12945
rect -1000 12900 0 12905
rect -1200 12545 0 12550
rect -1200 12505 -1195 12545
rect -1155 12505 0 12545
rect -1200 12500 0 12505
rect -1300 12445 0 12450
rect -1300 12405 -1295 12445
rect -1255 12405 0 12445
rect -1300 12400 0 12405
rect -1400 12345 0 12350
rect -1400 12305 -1395 12345
rect -1355 12305 0 12345
rect -1400 12300 0 12305
rect -1500 12245 0 12250
rect -1500 12205 -1495 12245
rect -1455 12205 0 12245
rect -1500 12200 0 12205
rect -3500 11945 0 11950
rect -3500 11905 -3495 11945
rect -3455 11905 -3295 11945
rect -3255 11905 -3095 11945
rect -3055 11905 -1595 11945
rect -1555 11905 -1095 11945
rect -1055 11905 -895 11945
rect -855 11905 -695 11945
rect -655 11905 -495 11945
rect -455 11905 -295 11945
rect -255 11905 -95 11945
rect -55 11905 0 11945
rect -3500 11895 0 11905
rect -3500 11855 -3495 11895
rect -3455 11855 -3295 11895
rect -3255 11855 -3095 11895
rect -3055 11855 -1595 11895
rect -1555 11855 -1095 11895
rect -1055 11855 -895 11895
rect -855 11855 -695 11895
rect -655 11855 -495 11895
rect -455 11855 -295 11895
rect -255 11855 -95 11895
rect -55 11855 0 11895
rect -3500 11845 0 11855
rect -3500 11805 -3495 11845
rect -3455 11805 -3295 11845
rect -3255 11805 -3095 11845
rect -3055 11805 -1595 11845
rect -1555 11805 -1095 11845
rect -1055 11805 -895 11845
rect -855 11805 -695 11845
rect -655 11805 -495 11845
rect -455 11805 -295 11845
rect -255 11805 -95 11845
rect -55 11805 0 11845
rect -3500 11800 0 11805
rect -3200 11445 0 11450
rect -3200 11405 -3195 11445
rect -3155 11405 0 11445
rect -3200 11400 0 11405
rect 39750 11345 39900 11350
rect 39750 11305 39805 11345
rect 39845 11305 39900 11345
rect 39750 11300 39900 11305
rect 39750 11245 40900 11250
rect 39750 11205 39905 11245
rect 39945 11205 39955 11245
rect 39995 11205 40005 11245
rect 40045 11205 40055 11245
rect 40095 11205 40105 11245
rect 40145 11205 40155 11245
rect 40195 11205 40205 11245
rect 40245 11205 40255 11245
rect 40295 11205 40305 11245
rect 40345 11205 40355 11245
rect 40395 11205 40405 11245
rect 40445 11205 40455 11245
rect 40495 11205 40505 11245
rect 40545 11205 40555 11245
rect 40595 11205 40605 11245
rect 40645 11205 40655 11245
rect 40695 11205 40705 11245
rect 40745 11205 40755 11245
rect 40795 11205 40805 11245
rect 40845 11205 40855 11245
rect 40895 11205 40900 11245
rect 39750 11195 40900 11205
rect 39750 11155 39905 11195
rect 39945 11155 39955 11195
rect 39995 11155 40005 11195
rect 40045 11155 40055 11195
rect 40095 11155 40105 11195
rect 40145 11155 40155 11195
rect 40195 11155 40205 11195
rect 40245 11155 40255 11195
rect 40295 11155 40305 11195
rect 40345 11155 40355 11195
rect 40395 11155 40405 11195
rect 40445 11155 40455 11195
rect 40495 11155 40505 11195
rect 40545 11155 40555 11195
rect 40595 11155 40605 11195
rect 40645 11155 40655 11195
rect 40695 11155 40705 11195
rect 40745 11155 40755 11195
rect 40795 11155 40805 11195
rect 40845 11155 40855 11195
rect 40895 11155 40900 11195
rect 39750 11145 40900 11155
rect 39750 11105 39905 11145
rect 39945 11105 39955 11145
rect 39995 11105 40005 11145
rect 40045 11105 40055 11145
rect 40095 11105 40105 11145
rect 40145 11105 40155 11145
rect 40195 11105 40205 11145
rect 40245 11105 40255 11145
rect 40295 11105 40305 11145
rect 40345 11105 40355 11145
rect 40395 11105 40405 11145
rect 40445 11105 40455 11145
rect 40495 11105 40505 11145
rect 40545 11105 40555 11145
rect 40595 11105 40605 11145
rect 40645 11105 40655 11145
rect 40695 11105 40705 11145
rect 40745 11105 40755 11145
rect 40795 11105 40805 11145
rect 40845 11105 40855 11145
rect 40895 11105 40900 11145
rect 39750 11095 40900 11105
rect 39750 11055 39905 11095
rect 39945 11055 39955 11095
rect 39995 11055 40005 11095
rect 40045 11055 40055 11095
rect 40095 11055 40105 11095
rect 40145 11055 40155 11095
rect 40195 11055 40205 11095
rect 40245 11055 40255 11095
rect 40295 11055 40305 11095
rect 40345 11055 40355 11095
rect 40395 11055 40405 11095
rect 40445 11055 40455 11095
rect 40495 11055 40505 11095
rect 40545 11055 40555 11095
rect 40595 11055 40605 11095
rect 40645 11055 40655 11095
rect 40695 11055 40705 11095
rect 40745 11055 40755 11095
rect 40795 11055 40805 11095
rect 40845 11055 40855 11095
rect 40895 11055 40900 11095
rect 39750 11045 40900 11055
rect 39750 11005 39905 11045
rect 39945 11005 39955 11045
rect 39995 11005 40005 11045
rect 40045 11005 40055 11045
rect 40095 11005 40105 11045
rect 40145 11005 40155 11045
rect 40195 11005 40205 11045
rect 40245 11005 40255 11045
rect 40295 11005 40305 11045
rect 40345 11005 40355 11045
rect 40395 11005 40405 11045
rect 40445 11005 40455 11045
rect 40495 11005 40505 11045
rect 40545 11005 40555 11045
rect 40595 11005 40605 11045
rect 40645 11005 40655 11045
rect 40695 11005 40705 11045
rect 40745 11005 40755 11045
rect 40795 11005 40805 11045
rect 40845 11005 40855 11045
rect 40895 11005 40900 11045
rect 39750 11000 40900 11005
rect 39750 10945 39900 10950
rect 39750 10905 39805 10945
rect 39845 10905 39900 10945
rect 39750 10900 39900 10905
rect -3400 10845 0 10850
rect -3400 10805 -3395 10845
rect -3355 10805 0 10845
rect -3400 10800 0 10805
rect -3100 10645 0 10650
rect -3100 10605 -2995 10645
rect -2955 10605 -2795 10645
rect -2755 10605 -2595 10645
rect -2555 10605 -2395 10645
rect -2355 10605 -2195 10645
rect -2155 10605 -1995 10645
rect -1955 10605 -1695 10645
rect -1655 10605 0 10645
rect -3100 10595 0 10605
rect -3100 10555 -2995 10595
rect -2955 10555 -2795 10595
rect -2755 10555 -2595 10595
rect -2555 10555 -2395 10595
rect -2355 10555 -2195 10595
rect -2155 10555 -1995 10595
rect -1955 10555 -1695 10595
rect -1655 10555 0 10595
rect -3100 10545 0 10555
rect -3100 10505 -2995 10545
rect -2955 10505 -2795 10545
rect -2755 10505 -2595 10545
rect -2555 10505 -2395 10545
rect -2355 10505 -2195 10545
rect -2155 10505 -1995 10545
rect -1955 10505 -1695 10545
rect -1655 10505 0 10545
rect -3100 10500 0 10505
rect -1800 10245 0 10250
rect -1800 10205 -1795 10245
rect -1755 10205 0 10245
rect -1800 10200 0 10205
rect -1900 10145 0 10150
rect -1900 10105 -1895 10145
rect -1855 10105 0 10145
rect -1900 10100 0 10105
rect -2100 9745 0 9750
rect -2100 9705 -2095 9745
rect -2055 9705 0 9745
rect -2100 9700 0 9705
rect -2300 9545 0 9550
rect -2300 9505 -2295 9545
rect -2255 9505 0 9545
rect -2300 9500 0 9505
rect -3100 9345 0 9350
rect -3100 9305 -2995 9345
rect -2955 9305 -2795 9345
rect -2755 9305 -2595 9345
rect -2555 9305 -2395 9345
rect -2355 9305 -2195 9345
rect -2155 9305 -1995 9345
rect -1955 9305 -1695 9345
rect -1655 9305 0 9345
rect -3100 9295 0 9305
rect -3100 9255 -2995 9295
rect -2955 9255 -2795 9295
rect -2755 9255 -2595 9295
rect -2555 9255 -2395 9295
rect -2355 9255 -2195 9295
rect -2155 9255 -1995 9295
rect -1955 9255 -1695 9295
rect -1655 9255 0 9295
rect -3100 9245 0 9255
rect -3100 9205 -2995 9245
rect -2955 9205 -2795 9245
rect -2755 9205 -2595 9245
rect -2555 9205 -2395 9245
rect -2355 9205 -2195 9245
rect -2155 9205 -1995 9245
rect -1955 9205 -1695 9245
rect -1655 9205 0 9245
rect -3100 9200 0 9205
rect -2500 9045 0 9050
rect -2500 9005 -2495 9045
rect -2455 9005 0 9045
rect -2500 9000 0 9005
rect -2700 8845 0 8850
rect -2700 8805 -2695 8845
rect -2655 8805 0 8845
rect -2700 8800 0 8805
rect -2900 8445 0 8450
rect -2900 8405 -2895 8445
rect -2855 8405 0 8445
rect -2900 8400 0 8405
rect -3100 8045 0 8050
rect -3100 8005 -2995 8045
rect -2955 8005 -2795 8045
rect -2755 8005 -2595 8045
rect -2555 8005 -2395 8045
rect -2355 8005 -2195 8045
rect -2155 8005 -1995 8045
rect -1955 8005 -1695 8045
rect -1655 8005 0 8045
rect -3100 7995 0 8005
rect -3100 7955 -2995 7995
rect -2955 7955 -2795 7995
rect -2755 7955 -2595 7995
rect -2555 7955 -2395 7995
rect -2355 7955 -2195 7995
rect -2155 7955 -1995 7995
rect -1955 7955 -1695 7995
rect -1655 7955 0 7995
rect -3100 7945 0 7955
rect -3100 7905 -2995 7945
rect -2955 7905 -2795 7945
rect -2755 7905 -2595 7945
rect -2555 7905 -2395 7945
rect -2355 7905 -2195 7945
rect -2155 7905 -1995 7945
rect -1955 7905 -1695 7945
rect -1655 7905 0 7945
rect -3100 7900 0 7905
rect -3100 7745 0 7750
rect -3100 7705 -2995 7745
rect -2955 7705 -2795 7745
rect -2755 7705 -2595 7745
rect -2555 7705 -2395 7745
rect -2355 7705 -2195 7745
rect -2155 7705 -1995 7745
rect -1955 7705 -1695 7745
rect -1655 7705 0 7745
rect -3100 7695 0 7705
rect -3100 7655 -2995 7695
rect -2955 7655 -2795 7695
rect -2755 7655 -2595 7695
rect -2555 7655 -2395 7695
rect -2355 7655 -2195 7695
rect -2155 7655 -1995 7695
rect -1955 7655 -1695 7695
rect -1655 7655 0 7695
rect -3100 7645 0 7655
rect -3100 7605 -2995 7645
rect -2955 7605 -2795 7645
rect -2755 7605 -2595 7645
rect -2555 7605 -2395 7645
rect -2355 7605 -2195 7645
rect -2155 7605 -1995 7645
rect -1955 7605 -1695 7645
rect -1655 7605 0 7645
rect -3100 7600 0 7605
rect -2900 7245 0 7250
rect -2900 7205 -2895 7245
rect -2855 7205 0 7245
rect -2900 7200 0 7205
rect -2700 6845 0 6850
rect -2700 6805 -2695 6845
rect -2655 6805 0 6845
rect -2700 6800 0 6805
rect -2500 6645 0 6650
rect -2500 6605 -2495 6645
rect -2455 6605 0 6645
rect -2500 6600 0 6605
rect -3100 6445 0 6450
rect -3100 6405 -2995 6445
rect -2955 6405 -2795 6445
rect -2755 6405 -2595 6445
rect -2555 6405 -2395 6445
rect -2355 6405 -2195 6445
rect -2155 6405 -1995 6445
rect -1955 6405 -1695 6445
rect -1655 6405 0 6445
rect -3100 6395 0 6405
rect -3100 6355 -2995 6395
rect -2955 6355 -2795 6395
rect -2755 6355 -2595 6395
rect -2555 6355 -2395 6395
rect -2355 6355 -2195 6395
rect -2155 6355 -1995 6395
rect -1955 6355 -1695 6395
rect -1655 6355 0 6395
rect -3100 6345 0 6355
rect -3100 6305 -2995 6345
rect -2955 6305 -2795 6345
rect -2755 6305 -2595 6345
rect -2555 6305 -2395 6345
rect -2355 6305 -2195 6345
rect -2155 6305 -1995 6345
rect -1955 6305 -1695 6345
rect -1655 6305 0 6345
rect -3100 6300 0 6305
rect -2300 6145 0 6150
rect -2300 6105 -2295 6145
rect -2255 6105 0 6145
rect -2300 6100 0 6105
rect -2100 5945 0 5950
rect -2100 5905 -2095 5945
rect -2055 5905 0 5945
rect -2100 5900 0 5905
rect -1900 5545 0 5550
rect -1900 5505 -1895 5545
rect -1855 5505 0 5545
rect -1900 5500 0 5505
rect -1800 5445 0 5450
rect -1800 5405 -1795 5445
rect -1755 5405 0 5445
rect -1800 5400 0 5405
rect -3100 5145 0 5150
rect -3100 5105 -2995 5145
rect -2955 5105 -2795 5145
rect -2755 5105 -2595 5145
rect -2555 5105 -2395 5145
rect -2355 5105 -2195 5145
rect -2155 5105 -1995 5145
rect -1955 5105 -1695 5145
rect -1655 5105 0 5145
rect -3100 5095 0 5105
rect -3100 5055 -2995 5095
rect -2955 5055 -2795 5095
rect -2755 5055 -2595 5095
rect -2555 5055 -2395 5095
rect -2355 5055 -2195 5095
rect -2155 5055 -1995 5095
rect -1955 5055 -1695 5095
rect -1655 5055 0 5095
rect -3100 5045 0 5055
rect -3100 5005 -2995 5045
rect -2955 5005 -2795 5045
rect -2755 5005 -2595 5045
rect -2555 5005 -2395 5045
rect -2355 5005 -2195 5045
rect -2155 5005 -1995 5045
rect -1955 5005 -1695 5045
rect -1655 5005 0 5045
rect -3100 5000 0 5005
rect -3400 4845 0 4850
rect -3400 4805 -3395 4845
rect -3355 4805 0 4845
rect -3400 4800 0 4805
rect 39750 4745 39900 4750
rect 39750 4705 39805 4745
rect 39845 4705 39900 4745
rect 39750 4700 39900 4705
rect 39750 4645 40900 4650
rect 39750 4605 39905 4645
rect 39945 4605 39955 4645
rect 39995 4605 40005 4645
rect 40045 4605 40055 4645
rect 40095 4605 40105 4645
rect 40145 4605 40155 4645
rect 40195 4605 40205 4645
rect 40245 4605 40255 4645
rect 40295 4605 40305 4645
rect 40345 4605 40355 4645
rect 40395 4605 40405 4645
rect 40445 4605 40455 4645
rect 40495 4605 40505 4645
rect 40545 4605 40555 4645
rect 40595 4605 40605 4645
rect 40645 4605 40655 4645
rect 40695 4605 40705 4645
rect 40745 4605 40755 4645
rect 40795 4605 40805 4645
rect 40845 4605 40855 4645
rect 40895 4605 40900 4645
rect 39750 4595 40900 4605
rect 39750 4555 39905 4595
rect 39945 4555 39955 4595
rect 39995 4555 40005 4595
rect 40045 4555 40055 4595
rect 40095 4555 40105 4595
rect 40145 4555 40155 4595
rect 40195 4555 40205 4595
rect 40245 4555 40255 4595
rect 40295 4555 40305 4595
rect 40345 4555 40355 4595
rect 40395 4555 40405 4595
rect 40445 4555 40455 4595
rect 40495 4555 40505 4595
rect 40545 4555 40555 4595
rect 40595 4555 40605 4595
rect 40645 4555 40655 4595
rect 40695 4555 40705 4595
rect 40745 4555 40755 4595
rect 40795 4555 40805 4595
rect 40845 4555 40855 4595
rect 40895 4555 40900 4595
rect 39750 4545 40900 4555
rect 39750 4505 39905 4545
rect 39945 4505 39955 4545
rect 39995 4505 40005 4545
rect 40045 4505 40055 4545
rect 40095 4505 40105 4545
rect 40145 4505 40155 4545
rect 40195 4505 40205 4545
rect 40245 4505 40255 4545
rect 40295 4505 40305 4545
rect 40345 4505 40355 4545
rect 40395 4505 40405 4545
rect 40445 4505 40455 4545
rect 40495 4505 40505 4545
rect 40545 4505 40555 4545
rect 40595 4505 40605 4545
rect 40645 4505 40655 4545
rect 40695 4505 40705 4545
rect 40745 4505 40755 4545
rect 40795 4505 40805 4545
rect 40845 4505 40855 4545
rect 40895 4505 40900 4545
rect 39750 4495 40900 4505
rect 39750 4455 39905 4495
rect 39945 4455 39955 4495
rect 39995 4455 40005 4495
rect 40045 4455 40055 4495
rect 40095 4455 40105 4495
rect 40145 4455 40155 4495
rect 40195 4455 40205 4495
rect 40245 4455 40255 4495
rect 40295 4455 40305 4495
rect 40345 4455 40355 4495
rect 40395 4455 40405 4495
rect 40445 4455 40455 4495
rect 40495 4455 40505 4495
rect 40545 4455 40555 4495
rect 40595 4455 40605 4495
rect 40645 4455 40655 4495
rect 40695 4455 40705 4495
rect 40745 4455 40755 4495
rect 40795 4455 40805 4495
rect 40845 4455 40855 4495
rect 40895 4455 40900 4495
rect 39750 4445 40900 4455
rect 39750 4405 39905 4445
rect 39945 4405 39955 4445
rect 39995 4405 40005 4445
rect 40045 4405 40055 4445
rect 40095 4405 40105 4445
rect 40145 4405 40155 4445
rect 40195 4405 40205 4445
rect 40245 4405 40255 4445
rect 40295 4405 40305 4445
rect 40345 4405 40355 4445
rect 40395 4405 40405 4445
rect 40445 4405 40455 4445
rect 40495 4405 40505 4445
rect 40545 4405 40555 4445
rect 40595 4405 40605 4445
rect 40645 4405 40655 4445
rect 40695 4405 40705 4445
rect 40745 4405 40755 4445
rect 40795 4405 40805 4445
rect 40845 4405 40855 4445
rect 40895 4405 40900 4445
rect 39750 4400 40900 4405
rect 39750 4345 39900 4350
rect 39750 4305 39805 4345
rect 39845 4305 39900 4345
rect 39750 4300 39900 4305
rect -3200 4245 0 4250
rect -3200 4205 -3195 4245
rect -3155 4205 0 4245
rect -3200 4200 0 4205
rect -3500 3845 0 3850
rect -3500 3805 -3495 3845
rect -3455 3805 -3295 3845
rect -3255 3805 -3095 3845
rect -3055 3805 -1595 3845
rect -1555 3805 -1095 3845
rect -1055 3805 -895 3845
rect -855 3805 -695 3845
rect -655 3805 -495 3845
rect -455 3805 -295 3845
rect -255 3805 -95 3845
rect -55 3805 0 3845
rect -3500 3795 0 3805
rect -3500 3755 -3495 3795
rect -3455 3755 -3295 3795
rect -3255 3755 -3095 3795
rect -3055 3755 -1595 3795
rect -1555 3755 -1095 3795
rect -1055 3755 -895 3795
rect -855 3755 -695 3795
rect -655 3755 -495 3795
rect -455 3755 -295 3795
rect -255 3755 -95 3795
rect -55 3755 0 3795
rect -3500 3745 0 3755
rect -3500 3705 -3495 3745
rect -3455 3705 -3295 3745
rect -3255 3705 -3095 3745
rect -3055 3705 -1595 3745
rect -1555 3705 -1095 3745
rect -1055 3705 -895 3745
rect -855 3705 -695 3745
rect -655 3705 -495 3745
rect -455 3705 -295 3745
rect -255 3705 -95 3745
rect -55 3705 0 3745
rect -3500 3700 0 3705
rect -1500 3445 0 3450
rect -1500 3405 -1495 3445
rect -1455 3405 0 3445
rect -1500 3400 0 3405
rect -1400 3345 0 3350
rect -1400 3305 -1395 3345
rect -1355 3305 0 3345
rect -1400 3300 0 3305
rect -1300 3245 0 3250
rect -1300 3205 -1295 3245
rect -1255 3205 0 3245
rect -1300 3200 0 3205
rect -1200 3145 0 3150
rect -1200 3105 -1195 3145
rect -1155 3105 0 3145
rect -1200 3100 0 3105
rect -1000 2745 0 2750
rect -1000 2705 -995 2745
rect -955 2705 0 2745
rect -1000 2700 0 2705
rect -800 2545 0 2550
rect -800 2505 -795 2545
rect -755 2505 0 2545
rect -800 2500 0 2505
rect -3500 2145 0 2150
rect -3500 2105 -3495 2145
rect -3455 2105 -3295 2145
rect -3255 2105 -3095 2145
rect -3055 2105 -1595 2145
rect -1555 2105 -1095 2145
rect -1055 2105 -895 2145
rect -855 2105 -695 2145
rect -655 2105 -495 2145
rect -455 2105 -295 2145
rect -255 2105 -95 2145
rect -55 2105 0 2145
rect -3500 2095 0 2105
rect -3500 2055 -3495 2095
rect -3455 2055 -3295 2095
rect -3255 2055 -3095 2095
rect -3055 2055 -1595 2095
rect -1555 2055 -1095 2095
rect -1055 2055 -895 2095
rect -855 2055 -695 2095
rect -655 2055 -495 2095
rect -455 2055 -295 2095
rect -255 2055 -95 2095
rect -55 2055 0 2095
rect -3500 2045 0 2055
rect -3500 2005 -3495 2045
rect -3455 2005 -3295 2045
rect -3255 2005 -3095 2045
rect -3055 2005 -1595 2045
rect -1555 2005 -1095 2045
rect -1055 2005 -895 2045
rect -855 2005 -695 2045
rect -655 2005 -495 2045
rect -455 2005 -295 2045
rect -255 2005 -95 2045
rect -55 2005 0 2045
rect -3500 2000 0 2005
rect -600 1645 0 1650
rect -600 1605 -595 1645
rect -555 1605 0 1645
rect -600 1600 0 1605
rect -400 1445 0 1450
rect -400 1405 -395 1445
rect -355 1405 0 1445
rect -400 1400 0 1405
rect -200 1045 0 1050
rect -200 1005 -195 1045
rect -155 1005 0 1045
rect -200 1000 0 1005
rect -3500 445 0 450
rect -3500 405 -3495 445
rect -3455 405 -3295 445
rect -3255 405 -3095 445
rect -3055 405 -1595 445
rect -1555 405 -1095 445
rect -1055 405 -895 445
rect -855 405 -695 445
rect -655 405 -495 445
rect -455 405 -295 445
rect -255 405 -95 445
rect -55 405 0 445
rect -3500 395 0 405
rect -3500 355 -3495 395
rect -3455 355 -3295 395
rect -3255 355 -3095 395
rect -3055 355 -1595 395
rect -1555 355 -1095 395
rect -1055 355 -895 395
rect -855 355 -695 395
rect -655 355 -495 395
rect -455 355 -295 395
rect -255 355 -95 395
rect -55 355 0 395
rect -3500 345 0 355
rect -3500 305 -3495 345
rect -3455 305 -3295 345
rect -3255 305 -3095 345
rect -3055 305 -1595 345
rect -1555 305 -1095 345
rect -1055 305 -895 345
rect -855 305 -695 345
rect -655 305 -495 345
rect -455 305 -295 345
rect -255 305 -95 345
rect -55 305 0 345
rect -3500 300 0 305
<< via3 >>
rect 5 18105 45 18145
rect 55 18105 95 18145
rect 105 18105 145 18145
rect 155 18105 195 18145
rect 205 18105 245 18145
rect 255 18105 295 18145
rect 305 18105 345 18145
rect 355 18105 395 18145
rect 405 18105 445 18145
rect 455 18105 495 18145
rect 505 18105 545 18145
rect 555 18105 595 18145
rect 605 18105 645 18145
rect 655 18105 695 18145
rect 705 18105 745 18145
rect 755 18105 795 18145
rect 805 18105 845 18145
rect 855 18105 895 18145
rect 905 18105 945 18145
rect 955 18105 995 18145
rect 1005 18105 1045 18145
rect 1055 18105 1095 18145
rect 1105 18105 1145 18145
rect 1155 18105 1195 18145
rect 1205 18105 1245 18145
rect 1255 18105 1295 18145
rect 1305 18105 1345 18145
rect 1355 18105 1395 18145
rect 1405 18105 1445 18145
rect 1455 18105 1495 18145
rect 1505 18105 1545 18145
rect 1555 18105 1595 18145
rect 1605 18105 1645 18145
rect 1655 18105 1695 18145
rect 1705 18105 1745 18145
rect 1755 18105 1795 18145
rect 1805 18105 1845 18145
rect 1855 18105 1895 18145
rect 1905 18105 1945 18145
rect 1955 18105 1995 18145
rect 2005 18105 2045 18145
rect 2055 18105 2095 18145
rect 2105 18105 2145 18145
rect 2155 18105 2195 18145
rect 2205 18105 2245 18145
rect 2255 18105 2295 18145
rect 2305 18105 2345 18145
rect 2355 18105 2395 18145
rect 2405 18105 2445 18145
rect 2455 18105 2495 18145
rect 2505 18105 2545 18145
rect 2555 18105 2595 18145
rect 2605 18105 2645 18145
rect 2655 18105 2695 18145
rect 2705 18105 2745 18145
rect 2755 18105 2795 18145
rect 2805 18105 2845 18145
rect 2855 18105 2895 18145
rect 2905 18105 2945 18145
rect 2955 18105 2995 18145
rect 3005 18105 3045 18145
rect 3055 18105 3095 18145
rect 3105 18105 3145 18145
rect 3155 18105 3195 18145
rect 3205 18105 3245 18145
rect 3255 18105 3295 18145
rect 3305 18105 3345 18145
rect 3355 18105 3395 18145
rect 3405 18105 3445 18145
rect 3455 18105 3495 18145
rect 3505 18105 3545 18145
rect 3555 18105 3595 18145
rect 3605 18105 3645 18145
rect 3655 18105 3695 18145
rect 3705 18105 3745 18145
rect 3755 18105 3795 18145
rect 3805 18105 3845 18145
rect 3855 18105 3895 18145
rect 3905 18105 3945 18145
rect 3955 18105 3995 18145
rect 4005 18105 4045 18145
rect 4055 18105 4095 18145
rect 4105 18105 4145 18145
rect 4155 18105 4195 18145
rect 4205 18105 4245 18145
rect 4255 18105 4295 18145
rect 4305 18105 4345 18145
rect 4355 18105 4395 18145
rect 4405 18105 4445 18145
rect 4455 18105 4495 18145
rect 4505 18105 4545 18145
rect 4555 18105 4595 18145
rect 4605 18105 4645 18145
rect 4655 18105 4695 18145
rect 4705 18105 4745 18145
rect 4755 18105 4795 18145
rect 4805 18105 4845 18145
rect 4855 18105 4895 18145
rect 4905 18105 4945 18145
rect 4955 18105 4995 18145
rect 5005 18105 5045 18145
rect 5055 18105 5095 18145
rect 5105 18105 5145 18145
rect 5155 18105 5195 18145
rect 5205 18105 5245 18145
rect 5255 18105 5295 18145
rect 5305 18105 5345 18145
rect 5355 18105 5395 18145
rect 5405 18105 5445 18145
rect 5455 18105 5495 18145
rect 5505 18105 5545 18145
rect 5555 18105 5595 18145
rect 5605 18105 5645 18145
rect 5655 18105 5695 18145
rect 5705 18105 5745 18145
rect 5755 18105 5795 18145
rect 5805 18105 5845 18145
rect 5855 18105 5895 18145
rect 5905 18105 5945 18145
rect 5955 18105 5995 18145
rect 6005 18105 6045 18145
rect 6055 18105 6095 18145
rect 6105 18105 6145 18145
rect 6155 18105 6195 18145
rect 6205 18105 6245 18145
rect 6255 18105 6295 18145
rect 6305 18105 6345 18145
rect 6355 18105 6395 18145
rect 6405 18105 6445 18145
rect 6455 18105 6495 18145
rect 6505 18105 6545 18145
rect 6555 18105 6595 18145
rect 6605 18105 6645 18145
rect 6655 18105 6695 18145
rect 6705 18105 6745 18145
rect 6755 18105 6795 18145
rect 6805 18105 6845 18145
rect 6855 18105 6895 18145
rect 6905 18105 6945 18145
rect 6955 18105 6995 18145
rect 7005 18105 7045 18145
rect 7055 18105 7095 18145
rect 7105 18105 7145 18145
rect 7155 18105 7195 18145
rect 7205 18105 7245 18145
rect 7255 18105 7295 18145
rect 7305 18105 7345 18145
rect 7355 18105 7395 18145
rect 7405 18105 7445 18145
rect 7455 18105 7495 18145
rect 7505 18105 7545 18145
rect 7555 18105 7595 18145
rect 7605 18105 7645 18145
rect 7655 18105 7695 18145
rect 7705 18105 7745 18145
rect 7755 18105 7795 18145
rect 7805 18105 7845 18145
rect 7855 18105 7895 18145
rect 7905 18105 7945 18145
rect 7955 18105 7995 18145
rect 8005 18105 8045 18145
rect 8055 18105 8095 18145
rect 8105 18105 8145 18145
rect 8155 18105 8195 18145
rect 8205 18105 8245 18145
rect 8255 18105 8295 18145
rect 8305 18105 8345 18145
rect 8355 18105 8395 18145
rect 8405 18105 8445 18145
rect 8455 18105 8495 18145
rect 8505 18105 8545 18145
rect 8555 18105 8595 18145
rect 8605 18105 8645 18145
rect 8655 18105 8695 18145
rect 8705 18105 8745 18145
rect 8755 18105 8795 18145
rect 8805 18105 8845 18145
rect 8855 18105 8895 18145
rect 8905 18105 8945 18145
rect 8955 18105 8995 18145
rect 9005 18105 9045 18145
rect 9055 18105 9095 18145
rect 9105 18105 9145 18145
rect 9155 18105 9195 18145
rect 9205 18105 9245 18145
rect 9255 18105 9295 18145
rect 9305 18105 9345 18145
rect 9355 18105 9395 18145
rect 9405 18105 9445 18145
rect 9455 18105 9495 18145
rect 9505 18105 9545 18145
rect 9555 18105 9595 18145
rect 9605 18105 9645 18145
rect 9655 18105 9695 18145
rect 9705 18105 9745 18145
rect 9755 18105 9795 18145
rect 9805 18105 9845 18145
rect 9855 18105 9895 18145
rect 9905 18105 9945 18145
rect 9955 18105 9995 18145
rect 10005 18105 10045 18145
rect 10055 18105 10095 18145
rect 10105 18105 10145 18145
rect 10155 18105 10195 18145
rect 10205 18105 10245 18145
rect 10255 18105 10295 18145
rect 10305 18105 10345 18145
rect 10355 18105 10395 18145
rect 10405 18105 10445 18145
rect 10455 18105 10495 18145
rect 10505 18105 10545 18145
rect 10555 18105 10595 18145
rect 10605 18105 10645 18145
rect 10655 18105 10695 18145
rect 10705 18105 10745 18145
rect 10755 18105 10795 18145
rect 10805 18105 10845 18145
rect 10855 18105 10895 18145
rect 10905 18105 10945 18145
rect 10955 18105 10995 18145
rect 11005 18105 11045 18145
rect 11055 18105 11095 18145
rect 11105 18105 11145 18145
rect 11155 18105 11195 18145
rect 11205 18105 11245 18145
rect 11255 18105 11295 18145
rect 11305 18105 11345 18145
rect 11355 18105 11395 18145
rect 11405 18105 11445 18145
rect 11455 18105 11495 18145
rect 11505 18105 11545 18145
rect 11555 18105 11595 18145
rect 11605 18105 11645 18145
rect 11655 18105 11695 18145
rect 11705 18105 11745 18145
rect 11755 18105 11795 18145
rect 11805 18105 11845 18145
rect 11855 18105 11895 18145
rect 11905 18105 11945 18145
rect 11955 18105 11995 18145
rect 12005 18105 12045 18145
rect 12055 18105 12095 18145
rect 12105 18105 12145 18145
rect 12155 18105 12195 18145
rect 12205 18105 12245 18145
rect 12255 18105 12295 18145
rect 12305 18105 12345 18145
rect 12355 18105 12395 18145
rect 12405 18105 12445 18145
rect 12455 18105 12495 18145
rect 12505 18105 12545 18145
rect 12555 18105 12595 18145
rect 12605 18105 12645 18145
rect 12655 18105 12695 18145
rect 12705 18105 12745 18145
rect 12755 18105 12795 18145
rect 12805 18105 12845 18145
rect 12855 18105 12895 18145
rect 12905 18105 12945 18145
rect 12955 18105 12995 18145
rect 13005 18105 13045 18145
rect 13055 18105 13095 18145
rect 13105 18105 13145 18145
rect 13155 18105 13195 18145
rect 13205 18105 13245 18145
rect 13255 18105 13295 18145
rect 13305 18105 13345 18145
rect 13355 18105 13395 18145
rect 13405 18105 13445 18145
rect 13455 18105 13495 18145
rect 13505 18105 13545 18145
rect 13555 18105 13595 18145
rect 13605 18105 13645 18145
rect 13655 18105 13695 18145
rect 13705 18105 13745 18145
rect 13755 18105 13795 18145
rect 13805 18105 13845 18145
rect 13855 18105 13895 18145
rect 13905 18105 13945 18145
rect 13955 18105 13995 18145
rect 14005 18105 14045 18145
rect 14055 18105 14095 18145
rect 14105 18105 14145 18145
rect 14155 18105 14195 18145
rect 14205 18105 14245 18145
rect 14255 18105 14295 18145
rect 14305 18105 14345 18145
rect 14355 18105 14395 18145
rect 14405 18105 14445 18145
rect 14455 18105 14495 18145
rect 14505 18105 14545 18145
rect 14555 18105 14595 18145
rect 14605 18105 14645 18145
rect 14655 18105 14695 18145
rect 14705 18105 14745 18145
rect 14755 18105 14795 18145
rect 14805 18105 14845 18145
rect 14855 18105 14895 18145
rect 14905 18105 14945 18145
rect 14955 18105 14995 18145
rect 15005 18105 15045 18145
rect 15055 18105 15095 18145
rect 15105 18105 15145 18145
rect 15155 18105 15195 18145
rect 15205 18105 15245 18145
rect 15255 18105 15295 18145
rect 15305 18105 15345 18145
rect 15355 18105 15395 18145
rect 15405 18105 15445 18145
rect 15455 18105 15495 18145
rect 15505 18105 15545 18145
rect 15555 18105 15595 18145
rect 15605 18105 15645 18145
rect 15655 18105 15695 18145
rect 15705 18105 15745 18145
rect 15755 18105 15795 18145
rect 15805 18105 15845 18145
rect 15855 18105 15895 18145
rect 15905 18105 15945 18145
rect 15955 18105 15995 18145
rect 16005 18105 16045 18145
rect 16055 18105 16095 18145
rect 16105 18105 16145 18145
rect 16155 18105 16195 18145
rect 16205 18105 16245 18145
rect 16255 18105 16295 18145
rect 16305 18105 16345 18145
rect 16355 18105 16395 18145
rect 16405 18105 16445 18145
rect 16455 18105 16495 18145
rect 16505 18105 16545 18145
rect 16555 18105 16595 18145
rect 16605 18105 16645 18145
rect 16655 18105 16695 18145
rect 16705 18105 16745 18145
rect 16755 18105 16795 18145
rect 16805 18105 16845 18145
rect 16855 18105 16895 18145
rect 16905 18105 16945 18145
rect 16955 18105 16995 18145
rect 17005 18105 17045 18145
rect 17055 18105 17095 18145
rect 17105 18105 17145 18145
rect 17155 18105 17195 18145
rect 17205 18105 17245 18145
rect 17255 18105 17295 18145
rect 17305 18105 17345 18145
rect 17355 18105 17395 18145
rect 17405 18105 17445 18145
rect 17455 18105 17495 18145
rect 17505 18105 17545 18145
rect 17555 18105 17595 18145
rect 17605 18105 17645 18145
rect 17655 18105 17695 18145
rect 17705 18105 17745 18145
rect 17755 18105 17795 18145
rect 17805 18105 17845 18145
rect 17855 18105 17895 18145
rect 17905 18105 17945 18145
rect 17955 18105 17995 18145
rect 18005 18105 18045 18145
rect 18055 18105 18095 18145
rect 18105 18105 18145 18145
rect 18155 18105 18195 18145
rect 18205 18105 18245 18145
rect 18255 18105 18295 18145
rect 18305 18105 18345 18145
rect 18355 18105 18395 18145
rect 18405 18105 18445 18145
rect 18455 18105 18495 18145
rect 18505 18105 18545 18145
rect 18555 18105 18595 18145
rect 18605 18105 18645 18145
rect 18655 18105 18695 18145
rect 18705 18105 18745 18145
rect 18755 18105 18795 18145
rect 18805 18105 18845 18145
rect 18855 18105 18895 18145
rect 18905 18105 18945 18145
rect 18955 18105 18995 18145
rect 19005 18105 19045 18145
rect 19055 18105 19095 18145
rect 19105 18105 19145 18145
rect 19155 18105 19195 18145
rect 19205 18105 19245 18145
rect 19255 18105 19295 18145
rect 19305 18105 19345 18145
rect 19355 18105 19395 18145
rect 19405 18105 19445 18145
rect 19455 18105 19495 18145
rect 19505 18105 19545 18145
rect 19555 18105 19595 18145
rect 19605 18105 19645 18145
rect 19655 18105 19695 18145
rect 19705 18105 19745 18145
rect 19755 18105 19795 18145
rect 19805 18105 19845 18145
rect 19855 18105 19895 18145
rect 19905 18105 19945 18145
rect 19955 18105 19995 18145
rect 20005 18105 20045 18145
rect 20055 18105 20095 18145
rect 20105 18105 20145 18145
rect 20155 18105 20195 18145
rect 20205 18105 20245 18145
rect 20255 18105 20295 18145
rect 20305 18105 20345 18145
rect 20355 18105 20395 18145
rect 20405 18105 20445 18145
rect 20455 18105 20495 18145
rect 20505 18105 20545 18145
rect 20555 18105 20595 18145
rect 20605 18105 20645 18145
rect 20655 18105 20695 18145
rect 20705 18105 20745 18145
rect 20755 18105 20795 18145
rect 20805 18105 20845 18145
rect 20855 18105 20895 18145
rect 20905 18105 20945 18145
rect 20955 18105 20995 18145
rect 21005 18105 21045 18145
rect 21055 18105 21095 18145
rect 21105 18105 21145 18145
rect 21155 18105 21195 18145
rect 21205 18105 21245 18145
rect 21255 18105 21295 18145
rect 21305 18105 21345 18145
rect 21355 18105 21395 18145
rect 21405 18105 21445 18145
rect 21455 18105 21495 18145
rect 21505 18105 21545 18145
rect 21555 18105 21595 18145
rect 21605 18105 21645 18145
rect 21655 18105 21695 18145
rect 21705 18105 21745 18145
rect 21755 18105 21795 18145
rect 21805 18105 21845 18145
rect 21855 18105 21895 18145
rect 21905 18105 21945 18145
rect 21955 18105 21995 18145
rect 22005 18105 22045 18145
rect 22055 18105 22095 18145
rect 22105 18105 22145 18145
rect 22155 18105 22195 18145
rect 22205 18105 22245 18145
rect 22255 18105 22295 18145
rect 22305 18105 22345 18145
rect 22355 18105 22395 18145
rect 22405 18105 22445 18145
rect 22455 18105 22495 18145
rect 22505 18105 22545 18145
rect 22555 18105 22595 18145
rect 22605 18105 22645 18145
rect 22655 18105 22695 18145
rect 22705 18105 22745 18145
rect 22755 18105 22795 18145
rect 22805 18105 22845 18145
rect 22855 18105 22895 18145
rect 22905 18105 22945 18145
rect 22955 18105 22995 18145
rect 23005 18105 23045 18145
rect 23055 18105 23095 18145
rect 23105 18105 23145 18145
rect 23155 18105 23195 18145
rect 23205 18105 23245 18145
rect 23255 18105 23295 18145
rect 23305 18105 23345 18145
rect 23355 18105 23395 18145
rect 23405 18105 23445 18145
rect 23455 18105 23495 18145
rect 23505 18105 23545 18145
rect 23555 18105 23595 18145
rect 23605 18105 23645 18145
rect 23655 18105 23695 18145
rect 23705 18105 23745 18145
rect 23755 18105 23795 18145
rect 23805 18105 23845 18145
rect 23855 18105 23895 18145
rect 23905 18105 23945 18145
rect 23955 18105 23995 18145
rect 24005 18105 24045 18145
rect 24055 18105 24095 18145
rect 24105 18105 24145 18145
rect 24155 18105 24195 18145
rect 24205 18105 24245 18145
rect 24255 18105 24295 18145
rect 24305 18105 24345 18145
rect 24355 18105 24395 18145
rect 24405 18105 24445 18145
rect 24455 18105 24495 18145
rect 24505 18105 24545 18145
rect 24555 18105 24595 18145
rect 24605 18105 24645 18145
rect 24655 18105 24695 18145
rect 24705 18105 24745 18145
rect 24755 18105 24795 18145
rect 24805 18105 24845 18145
rect 24855 18105 24895 18145
rect 24905 18105 24945 18145
rect 24955 18105 24995 18145
rect 25005 18105 25045 18145
rect 25055 18105 25095 18145
rect 25105 18105 25145 18145
rect 25155 18105 25195 18145
rect 25205 18105 25245 18145
rect 25255 18105 25295 18145
rect 25305 18105 25345 18145
rect 25355 18105 25395 18145
rect 25405 18105 25445 18145
rect 25455 18105 25495 18145
rect 25505 18105 25545 18145
rect 25555 18105 25595 18145
rect 25605 18105 25645 18145
rect 25655 18105 25695 18145
rect 25705 18105 25745 18145
rect 25755 18105 25795 18145
rect 25805 18105 25845 18145
rect 25855 18105 25895 18145
rect 25905 18105 25945 18145
rect 25955 18105 25995 18145
rect 26005 18105 26045 18145
rect 26055 18105 26095 18145
rect 26105 18105 26145 18145
rect 26155 18105 26195 18145
rect 26205 18105 26245 18145
rect 26255 18105 26295 18145
rect 26305 18105 26345 18145
rect 26355 18105 26395 18145
rect 26405 18105 26445 18145
rect 26455 18105 26495 18145
rect 26505 18105 26545 18145
rect 26555 18105 26595 18145
rect 26605 18105 26645 18145
rect 26655 18105 26695 18145
rect 26705 18105 26745 18145
rect 26755 18105 26795 18145
rect 26805 18105 26845 18145
rect 26855 18105 26895 18145
rect 26905 18105 26945 18145
rect 26955 18105 26995 18145
rect 27005 18105 27045 18145
rect 27055 18105 27095 18145
rect 27105 18105 27145 18145
rect 27155 18105 27195 18145
rect 27205 18105 27245 18145
rect 27255 18105 27295 18145
rect 27305 18105 27345 18145
rect 27355 18105 27395 18145
rect 27405 18105 27445 18145
rect 27455 18105 27495 18145
rect 27505 18105 27545 18145
rect 27555 18105 27595 18145
rect 27605 18105 27645 18145
rect 27655 18105 27695 18145
rect 27705 18105 27745 18145
rect 27755 18105 27795 18145
rect 27805 18105 27845 18145
rect 27855 18105 27895 18145
rect 27905 18105 27945 18145
rect 27955 18105 27995 18145
rect 28005 18105 28045 18145
rect 28055 18105 28095 18145
rect 28105 18105 28145 18145
rect 28155 18105 28195 18145
rect 28205 18105 28245 18145
rect 28255 18105 28295 18145
rect 28305 18105 28345 18145
rect 28355 18105 28395 18145
rect 28405 18105 28445 18145
rect 28455 18105 28495 18145
rect 28505 18105 28545 18145
rect 28555 18105 28595 18145
rect 28605 18105 28645 18145
rect 28655 18105 28695 18145
rect 28705 18105 28745 18145
rect 28755 18105 28795 18145
rect 28805 18105 28845 18145
rect 28855 18105 28895 18145
rect 28905 18105 28945 18145
rect 28955 18105 28995 18145
rect 29005 18105 29045 18145
rect 29055 18105 29095 18145
rect 29105 18105 29145 18145
rect 29155 18105 29195 18145
rect 29205 18105 29245 18145
rect 29255 18105 29295 18145
rect 29305 18105 29345 18145
rect 29355 18105 29395 18145
rect 29405 18105 29445 18145
rect 29455 18105 29495 18145
rect 29505 18105 29545 18145
rect 29555 18105 29595 18145
rect 29605 18105 29645 18145
rect 29655 18105 29695 18145
rect 29705 18105 29745 18145
rect 29755 18105 29795 18145
rect 29805 18105 29845 18145
rect 29855 18105 29895 18145
rect 29905 18105 29945 18145
rect 29955 18105 29995 18145
rect 30005 18105 30045 18145
rect 30055 18105 30095 18145
rect 30105 18105 30145 18145
rect 30155 18105 30195 18145
rect 30205 18105 30245 18145
rect 30255 18105 30295 18145
rect 30305 18105 30345 18145
rect 30355 18105 30395 18145
rect 30405 18105 30445 18145
rect 30455 18105 30495 18145
rect 30505 18105 30545 18145
rect 30555 18105 30595 18145
rect 30605 18105 30645 18145
rect 30655 18105 30695 18145
rect 30705 18105 30745 18145
rect 30755 18105 30795 18145
rect 30805 18105 30845 18145
rect 30855 18105 30895 18145
rect 30905 18105 30945 18145
rect 30955 18105 30995 18145
rect 31005 18105 31045 18145
rect 31055 18105 31095 18145
rect 31105 18105 31145 18145
rect 31155 18105 31195 18145
rect 31205 18105 31245 18145
rect 31255 18105 31295 18145
rect 31305 18105 31345 18145
rect 31355 18105 31395 18145
rect 31405 18105 31445 18145
rect 31455 18105 31495 18145
rect 31505 18105 31545 18145
rect 31555 18105 31595 18145
rect 31605 18105 31645 18145
rect 31655 18105 31695 18145
rect 31705 18105 31745 18145
rect 31755 18105 31795 18145
rect 31805 18105 31845 18145
rect 31855 18105 31895 18145
rect 31905 18105 31945 18145
rect 31955 18105 31995 18145
rect 32005 18105 32045 18145
rect 32055 18105 32095 18145
rect 32105 18105 32145 18145
rect 32155 18105 32195 18145
rect 32205 18105 32245 18145
rect 32255 18105 32295 18145
rect 32305 18105 32345 18145
rect 32355 18105 32395 18145
rect 32405 18105 32445 18145
rect 32455 18105 32495 18145
rect 32505 18105 32545 18145
rect 32555 18105 32595 18145
rect 32605 18105 32645 18145
rect 32655 18105 32695 18145
rect 32705 18105 32745 18145
rect 32755 18105 32795 18145
rect 32805 18105 32845 18145
rect 32855 18105 32895 18145
rect 32905 18105 32945 18145
rect 32955 18105 32995 18145
rect 33005 18105 33045 18145
rect 33055 18105 33095 18145
rect 33105 18105 33145 18145
rect 33155 18105 33195 18145
rect 33205 18105 33245 18145
rect 33255 18105 33295 18145
rect 33305 18105 33345 18145
rect 33355 18105 33395 18145
rect 33405 18105 33445 18145
rect 33455 18105 33495 18145
rect 33505 18105 33545 18145
rect 33555 18105 33595 18145
rect 33605 18105 33645 18145
rect 33655 18105 33695 18145
rect 33705 18105 33745 18145
rect 33755 18105 33795 18145
rect 33805 18105 33845 18145
rect 33855 18105 33895 18145
rect 33905 18105 33945 18145
rect 33955 18105 33995 18145
rect 34005 18105 34045 18145
rect 34055 18105 34095 18145
rect 34105 18105 34145 18145
rect 34155 18105 34195 18145
rect 34205 18105 34245 18145
rect 34255 18105 34295 18145
rect 34305 18105 34345 18145
rect 34355 18105 34395 18145
rect 34405 18105 34445 18145
rect 34455 18105 34495 18145
rect 34505 18105 34545 18145
rect 34555 18105 34595 18145
rect 34605 18105 34645 18145
rect 34655 18105 34695 18145
rect 34705 18105 34745 18145
rect 34755 18105 34795 18145
rect 34805 18105 34845 18145
rect 34855 18105 34895 18145
rect 34905 18105 34945 18145
rect 34955 18105 34995 18145
rect 35005 18105 35045 18145
rect 35055 18105 35095 18145
rect 35105 18105 35145 18145
rect 35155 18105 35195 18145
rect 35205 18105 35245 18145
rect 35255 18105 35295 18145
rect 35305 18105 35345 18145
rect 35355 18105 35395 18145
rect 35405 18105 35445 18145
rect 35455 18105 35495 18145
rect 35505 18105 35545 18145
rect 35555 18105 35595 18145
rect 35605 18105 35645 18145
rect 35655 18105 35695 18145
rect 35705 18105 35745 18145
rect 35755 18105 35795 18145
rect 35805 18105 35845 18145
rect 35855 18105 35895 18145
rect 35905 18105 35945 18145
rect 35955 18105 35995 18145
rect 36005 18105 36045 18145
rect 36055 18105 36095 18145
rect 36105 18105 36145 18145
rect 36155 18105 36195 18145
rect 36205 18105 36245 18145
rect 36255 18105 36295 18145
rect 36305 18105 36345 18145
rect 36355 18105 36395 18145
rect 36405 18105 36445 18145
rect 36455 18105 36495 18145
rect 36505 18105 36545 18145
rect 36555 18105 36595 18145
rect 36605 18105 36645 18145
rect 36655 18105 36695 18145
rect 36705 18105 36745 18145
rect 36755 18105 36795 18145
rect 36805 18105 36845 18145
rect 36855 18105 36895 18145
rect 36905 18105 36945 18145
rect 36955 18105 36995 18145
rect 37005 18105 37045 18145
rect 37055 18105 37095 18145
rect 37105 18105 37145 18145
rect 37155 18105 37195 18145
rect 37205 18105 37245 18145
rect 37255 18105 37295 18145
rect 37305 18105 37345 18145
rect 37355 18105 37395 18145
rect 37405 18105 37445 18145
rect 37455 18105 37495 18145
rect 37505 18105 37545 18145
rect 37555 18105 37595 18145
rect 37605 18105 37645 18145
rect 37655 18105 37695 18145
rect 37705 18105 37745 18145
rect 37755 18105 37795 18145
rect 37805 18105 37845 18145
rect 37855 18105 37895 18145
rect 37905 18105 37945 18145
rect 37955 18105 37995 18145
rect 38005 18105 38045 18145
rect 38055 18105 38095 18145
rect 38105 18105 38145 18145
rect 38155 18105 38195 18145
rect 38205 18105 38245 18145
rect 38255 18105 38295 18145
rect 38305 18105 38345 18145
rect 38355 18105 38395 18145
rect 38405 18105 38445 18145
rect 38455 18105 38495 18145
rect 38505 18105 38545 18145
rect 38555 18105 38595 18145
rect 38605 18105 38645 18145
rect 38655 18105 38695 18145
rect 38705 18105 38745 18145
rect 38755 18105 38795 18145
rect 38805 18105 38845 18145
rect 38855 18105 38895 18145
rect 38905 18105 38945 18145
rect 38955 18105 38995 18145
rect 39005 18105 39045 18145
rect 39055 18105 39095 18145
rect 39105 18105 39145 18145
rect 39155 18105 39195 18145
rect 39205 18105 39245 18145
rect 39255 18105 39295 18145
rect 39305 18105 39345 18145
rect 39355 18105 39395 18145
rect 39405 18105 39445 18145
rect 39455 18105 39495 18145
rect 39505 18105 39545 18145
rect 39555 18105 39595 18145
rect 39605 18105 39645 18145
rect 39655 18105 39695 18145
rect 39705 18105 39745 18145
rect 39905 18105 39945 18145
rect 39955 18105 39995 18145
rect 40005 18105 40045 18145
rect 40055 18105 40095 18145
rect 40105 18105 40145 18145
rect 40155 18105 40195 18145
rect 40205 18105 40245 18145
rect 40255 18105 40295 18145
rect 40305 18105 40345 18145
rect 40355 18105 40395 18145
rect 40405 18105 40445 18145
rect 40455 18105 40495 18145
rect 40505 18105 40545 18145
rect 40555 18105 40595 18145
rect 40605 18105 40645 18145
rect 40655 18105 40695 18145
rect 40705 18105 40745 18145
rect 40755 18105 40795 18145
rect 40805 18105 40845 18145
rect 40855 18105 40895 18145
rect 5 18005 45 18045
rect 55 18005 95 18045
rect 105 18005 145 18045
rect 155 18005 195 18045
rect 205 18005 245 18045
rect 255 18005 295 18045
rect 305 18005 345 18045
rect 355 18005 395 18045
rect 405 18005 445 18045
rect 455 18005 495 18045
rect 505 18005 545 18045
rect 555 18005 595 18045
rect 605 18005 645 18045
rect 655 18005 695 18045
rect 705 18005 745 18045
rect 755 18005 795 18045
rect 805 18005 845 18045
rect 855 18005 895 18045
rect 905 18005 945 18045
rect 955 18005 995 18045
rect 1005 18005 1045 18045
rect 1055 18005 1095 18045
rect 1105 18005 1145 18045
rect 1155 18005 1195 18045
rect 1205 18005 1245 18045
rect 1255 18005 1295 18045
rect 1305 18005 1345 18045
rect 1355 18005 1395 18045
rect 1405 18005 1445 18045
rect 1455 18005 1495 18045
rect 1505 18005 1545 18045
rect 1555 18005 1595 18045
rect 1605 18005 1645 18045
rect 1655 18005 1695 18045
rect 1705 18005 1745 18045
rect 1755 18005 1795 18045
rect 1805 18005 1845 18045
rect 1855 18005 1895 18045
rect 1905 18005 1945 18045
rect 1955 18005 1995 18045
rect 2005 18005 2045 18045
rect 2055 18005 2095 18045
rect 2105 18005 2145 18045
rect 2155 18005 2195 18045
rect 2205 18005 2245 18045
rect 2255 18005 2295 18045
rect 2305 18005 2345 18045
rect 2355 18005 2395 18045
rect 2405 18005 2445 18045
rect 2455 18005 2495 18045
rect 2505 18005 2545 18045
rect 2555 18005 2595 18045
rect 2605 18005 2645 18045
rect 2655 18005 2695 18045
rect 2705 18005 2745 18045
rect 2755 18005 2795 18045
rect 2805 18005 2845 18045
rect 2855 18005 2895 18045
rect 2905 18005 2945 18045
rect 2955 18005 2995 18045
rect 3005 18005 3045 18045
rect 3055 18005 3095 18045
rect 3105 18005 3145 18045
rect 3155 18005 3195 18045
rect 3205 18005 3245 18045
rect 3255 18005 3295 18045
rect 3305 18005 3345 18045
rect 3355 18005 3395 18045
rect 3405 18005 3445 18045
rect 3455 18005 3495 18045
rect 3505 18005 3545 18045
rect 3555 18005 3595 18045
rect 3605 18005 3645 18045
rect 3655 18005 3695 18045
rect 3705 18005 3745 18045
rect 3755 18005 3795 18045
rect 3805 18005 3845 18045
rect 3855 18005 3895 18045
rect 3905 18005 3945 18045
rect 3955 18005 3995 18045
rect 4005 18005 4045 18045
rect 4055 18005 4095 18045
rect 4105 18005 4145 18045
rect 4155 18005 4195 18045
rect 4205 18005 4245 18045
rect 4255 18005 4295 18045
rect 4305 18005 4345 18045
rect 4355 18005 4395 18045
rect 4405 18005 4445 18045
rect 4455 18005 4495 18045
rect 4505 18005 4545 18045
rect 4555 18005 4595 18045
rect 4605 18005 4645 18045
rect 4655 18005 4695 18045
rect 4705 18005 4745 18045
rect 4755 18005 4795 18045
rect 4805 18005 4845 18045
rect 4855 18005 4895 18045
rect 4905 18005 4945 18045
rect 4955 18005 4995 18045
rect 5005 18005 5045 18045
rect 5055 18005 5095 18045
rect 5105 18005 5145 18045
rect 5155 18005 5195 18045
rect 5205 18005 5245 18045
rect 5255 18005 5295 18045
rect 5305 18005 5345 18045
rect 5355 18005 5395 18045
rect 5405 18005 5445 18045
rect 5455 18005 5495 18045
rect 5505 18005 5545 18045
rect 5555 18005 5595 18045
rect 5605 18005 5645 18045
rect 5655 18005 5695 18045
rect 5705 18005 5745 18045
rect 5755 18005 5795 18045
rect 5805 18005 5845 18045
rect 5855 18005 5895 18045
rect 5905 18005 5945 18045
rect 5955 18005 5995 18045
rect 6005 18005 6045 18045
rect 6055 18005 6095 18045
rect 6105 18005 6145 18045
rect 6155 18005 6195 18045
rect 6205 18005 6245 18045
rect 6255 18005 6295 18045
rect 6305 18005 6345 18045
rect 6355 18005 6395 18045
rect 6405 18005 6445 18045
rect 6455 18005 6495 18045
rect 6505 18005 6545 18045
rect 6555 18005 6595 18045
rect 6605 18005 6645 18045
rect 6655 18005 6695 18045
rect 6705 18005 6745 18045
rect 6755 18005 6795 18045
rect 6805 18005 6845 18045
rect 6855 18005 6895 18045
rect 6905 18005 6945 18045
rect 6955 18005 6995 18045
rect 7005 18005 7045 18045
rect 7055 18005 7095 18045
rect 7105 18005 7145 18045
rect 7155 18005 7195 18045
rect 7205 18005 7245 18045
rect 7255 18005 7295 18045
rect 7305 18005 7345 18045
rect 7355 18005 7395 18045
rect 7405 18005 7445 18045
rect 7455 18005 7495 18045
rect 7505 18005 7545 18045
rect 7555 18005 7595 18045
rect 7605 18005 7645 18045
rect 7655 18005 7695 18045
rect 7705 18005 7745 18045
rect 7755 18005 7795 18045
rect 7805 18005 7845 18045
rect 7855 18005 7895 18045
rect 7905 18005 7945 18045
rect 7955 18005 7995 18045
rect 8005 18005 8045 18045
rect 8055 18005 8095 18045
rect 8105 18005 8145 18045
rect 8155 18005 8195 18045
rect 8205 18005 8245 18045
rect 8255 18005 8295 18045
rect 8305 18005 8345 18045
rect 8355 18005 8395 18045
rect 8405 18005 8445 18045
rect 8455 18005 8495 18045
rect 8505 18005 8545 18045
rect 8555 18005 8595 18045
rect 8605 18005 8645 18045
rect 8655 18005 8695 18045
rect 8705 18005 8745 18045
rect 8755 18005 8795 18045
rect 8805 18005 8845 18045
rect 8855 18005 8895 18045
rect 8905 18005 8945 18045
rect 8955 18005 8995 18045
rect 9005 18005 9045 18045
rect 9055 18005 9095 18045
rect 9105 18005 9145 18045
rect 9155 18005 9195 18045
rect 9205 18005 9245 18045
rect 9255 18005 9295 18045
rect 9305 18005 9345 18045
rect 9355 18005 9395 18045
rect 9405 18005 9445 18045
rect 9455 18005 9495 18045
rect 9505 18005 9545 18045
rect 9555 18005 9595 18045
rect 9605 18005 9645 18045
rect 9655 18005 9695 18045
rect 9705 18005 9745 18045
rect 9755 18005 9795 18045
rect 9805 18005 9845 18045
rect 9855 18005 9895 18045
rect 9905 18005 9945 18045
rect 9955 18005 9995 18045
rect 10005 18005 10045 18045
rect 10055 18005 10095 18045
rect 10105 18005 10145 18045
rect 10155 18005 10195 18045
rect 10205 18005 10245 18045
rect 10255 18005 10295 18045
rect 10305 18005 10345 18045
rect 10355 18005 10395 18045
rect 10405 18005 10445 18045
rect 10455 18005 10495 18045
rect 10505 18005 10545 18045
rect 10555 18005 10595 18045
rect 10605 18005 10645 18045
rect 10655 18005 10695 18045
rect 10705 18005 10745 18045
rect 10755 18005 10795 18045
rect 10805 18005 10845 18045
rect 10855 18005 10895 18045
rect 10905 18005 10945 18045
rect 10955 18005 10995 18045
rect 11005 18005 11045 18045
rect 11055 18005 11095 18045
rect 11105 18005 11145 18045
rect 11155 18005 11195 18045
rect 11205 18005 11245 18045
rect 11255 18005 11295 18045
rect 11305 18005 11345 18045
rect 11355 18005 11395 18045
rect 11405 18005 11445 18045
rect 11455 18005 11495 18045
rect 11505 18005 11545 18045
rect 11555 18005 11595 18045
rect 11605 18005 11645 18045
rect 11655 18005 11695 18045
rect 11705 18005 11745 18045
rect 11755 18005 11795 18045
rect 11805 18005 11845 18045
rect 11855 18005 11895 18045
rect 11905 18005 11945 18045
rect 11955 18005 11995 18045
rect 12005 18005 12045 18045
rect 12055 18005 12095 18045
rect 12105 18005 12145 18045
rect 12155 18005 12195 18045
rect 12205 18005 12245 18045
rect 12255 18005 12295 18045
rect 12305 18005 12345 18045
rect 12355 18005 12395 18045
rect 12405 18005 12445 18045
rect 12455 18005 12495 18045
rect 12505 18005 12545 18045
rect 12555 18005 12595 18045
rect 12605 18005 12645 18045
rect 12655 18005 12695 18045
rect 12705 18005 12745 18045
rect 12755 18005 12795 18045
rect 12805 18005 12845 18045
rect 12855 18005 12895 18045
rect 12905 18005 12945 18045
rect 12955 18005 12995 18045
rect 13005 18005 13045 18045
rect 13055 18005 13095 18045
rect 13105 18005 13145 18045
rect 13155 18005 13195 18045
rect 13205 18005 13245 18045
rect 13255 18005 13295 18045
rect 13305 18005 13345 18045
rect 13355 18005 13395 18045
rect 13405 18005 13445 18045
rect 13455 18005 13495 18045
rect 13505 18005 13545 18045
rect 13555 18005 13595 18045
rect 13605 18005 13645 18045
rect 13655 18005 13695 18045
rect 13705 18005 13745 18045
rect 13755 18005 13795 18045
rect 13805 18005 13845 18045
rect 13855 18005 13895 18045
rect 13905 18005 13945 18045
rect 13955 18005 13995 18045
rect 14005 18005 14045 18045
rect 14055 18005 14095 18045
rect 14105 18005 14145 18045
rect 14155 18005 14195 18045
rect 14205 18005 14245 18045
rect 14255 18005 14295 18045
rect 14305 18005 14345 18045
rect 14355 18005 14395 18045
rect 14405 18005 14445 18045
rect 14455 18005 14495 18045
rect 14505 18005 14545 18045
rect 14555 18005 14595 18045
rect 14605 18005 14645 18045
rect 14655 18005 14695 18045
rect 14705 18005 14745 18045
rect 14755 18005 14795 18045
rect 14805 18005 14845 18045
rect 14855 18005 14895 18045
rect 14905 18005 14945 18045
rect 14955 18005 14995 18045
rect 15005 18005 15045 18045
rect 15055 18005 15095 18045
rect 15105 18005 15145 18045
rect 15155 18005 15195 18045
rect 15205 18005 15245 18045
rect 15255 18005 15295 18045
rect 15305 18005 15345 18045
rect 15355 18005 15395 18045
rect 15405 18005 15445 18045
rect 15455 18005 15495 18045
rect 15505 18005 15545 18045
rect 15555 18005 15595 18045
rect 15605 18005 15645 18045
rect 15655 18005 15695 18045
rect 15705 18005 15745 18045
rect 15755 18005 15795 18045
rect 15805 18005 15845 18045
rect 15855 18005 15895 18045
rect 15905 18005 15945 18045
rect 15955 18005 15995 18045
rect 16005 18005 16045 18045
rect 16055 18005 16095 18045
rect 16105 18005 16145 18045
rect 16155 18005 16195 18045
rect 16205 18005 16245 18045
rect 16255 18005 16295 18045
rect 16305 18005 16345 18045
rect 16355 18005 16395 18045
rect 16405 18005 16445 18045
rect 16455 18005 16495 18045
rect 16505 18005 16545 18045
rect 16555 18005 16595 18045
rect 16605 18005 16645 18045
rect 16655 18005 16695 18045
rect 16705 18005 16745 18045
rect 16755 18005 16795 18045
rect 16805 18005 16845 18045
rect 16855 18005 16895 18045
rect 16905 18005 16945 18045
rect 16955 18005 16995 18045
rect 17005 18005 17045 18045
rect 17055 18005 17095 18045
rect 17105 18005 17145 18045
rect 17155 18005 17195 18045
rect 17205 18005 17245 18045
rect 17255 18005 17295 18045
rect 17305 18005 17345 18045
rect 17355 18005 17395 18045
rect 17405 18005 17445 18045
rect 17455 18005 17495 18045
rect 17505 18005 17545 18045
rect 17555 18005 17595 18045
rect 17605 18005 17645 18045
rect 17655 18005 17695 18045
rect 17705 18005 17745 18045
rect 17755 18005 17795 18045
rect 17805 18005 17845 18045
rect 17855 18005 17895 18045
rect 17905 18005 17945 18045
rect 17955 18005 17995 18045
rect 18005 18005 18045 18045
rect 18055 18005 18095 18045
rect 18105 18005 18145 18045
rect 18155 18005 18195 18045
rect 18205 18005 18245 18045
rect 18255 18005 18295 18045
rect 18305 18005 18345 18045
rect 18355 18005 18395 18045
rect 18405 18005 18445 18045
rect 18455 18005 18495 18045
rect 18505 18005 18545 18045
rect 18555 18005 18595 18045
rect 18605 18005 18645 18045
rect 18655 18005 18695 18045
rect 18705 18005 18745 18045
rect 18755 18005 18795 18045
rect 18805 18005 18845 18045
rect 18855 18005 18895 18045
rect 18905 18005 18945 18045
rect 18955 18005 18995 18045
rect 19005 18005 19045 18045
rect 19055 18005 19095 18045
rect 19105 18005 19145 18045
rect 19155 18005 19195 18045
rect 19205 18005 19245 18045
rect 19255 18005 19295 18045
rect 19305 18005 19345 18045
rect 19355 18005 19395 18045
rect 19405 18005 19445 18045
rect 19455 18005 19495 18045
rect 19505 18005 19545 18045
rect 19555 18005 19595 18045
rect 19605 18005 19645 18045
rect 19655 18005 19695 18045
rect 19705 18005 19745 18045
rect 19755 18005 19795 18045
rect 19805 18005 19845 18045
rect 19855 18005 19895 18045
rect 19905 18005 19945 18045
rect 19955 18005 19995 18045
rect 20005 18005 20045 18045
rect 20055 18005 20095 18045
rect 20105 18005 20145 18045
rect 20155 18005 20195 18045
rect 20205 18005 20245 18045
rect 20255 18005 20295 18045
rect 20305 18005 20345 18045
rect 20355 18005 20395 18045
rect 20405 18005 20445 18045
rect 20455 18005 20495 18045
rect 20505 18005 20545 18045
rect 20555 18005 20595 18045
rect 20605 18005 20645 18045
rect 20655 18005 20695 18045
rect 20705 18005 20745 18045
rect 20755 18005 20795 18045
rect 20805 18005 20845 18045
rect 20855 18005 20895 18045
rect 20905 18005 20945 18045
rect 20955 18005 20995 18045
rect 21005 18005 21045 18045
rect 21055 18005 21095 18045
rect 21105 18005 21145 18045
rect 21155 18005 21195 18045
rect 21205 18005 21245 18045
rect 21255 18005 21295 18045
rect 21305 18005 21345 18045
rect 21355 18005 21395 18045
rect 21405 18005 21445 18045
rect 21455 18005 21495 18045
rect 21505 18005 21545 18045
rect 21555 18005 21595 18045
rect 21605 18005 21645 18045
rect 21655 18005 21695 18045
rect 21705 18005 21745 18045
rect 21755 18005 21795 18045
rect 21805 18005 21845 18045
rect 21855 18005 21895 18045
rect 21905 18005 21945 18045
rect 21955 18005 21995 18045
rect 22005 18005 22045 18045
rect 22055 18005 22095 18045
rect 22105 18005 22145 18045
rect 22155 18005 22195 18045
rect 22205 18005 22245 18045
rect 22255 18005 22295 18045
rect 22305 18005 22345 18045
rect 22355 18005 22395 18045
rect 22405 18005 22445 18045
rect 22455 18005 22495 18045
rect 22505 18005 22545 18045
rect 22555 18005 22595 18045
rect 22605 18005 22645 18045
rect 22655 18005 22695 18045
rect 22705 18005 22745 18045
rect 22755 18005 22795 18045
rect 22805 18005 22845 18045
rect 22855 18005 22895 18045
rect 22905 18005 22945 18045
rect 22955 18005 22995 18045
rect 23005 18005 23045 18045
rect 23055 18005 23095 18045
rect 23105 18005 23145 18045
rect 23155 18005 23195 18045
rect 23205 18005 23245 18045
rect 23255 18005 23295 18045
rect 23305 18005 23345 18045
rect 23355 18005 23395 18045
rect 23405 18005 23445 18045
rect 23455 18005 23495 18045
rect 23505 18005 23545 18045
rect 23555 18005 23595 18045
rect 23605 18005 23645 18045
rect 23655 18005 23695 18045
rect 23705 18005 23745 18045
rect 23755 18005 23795 18045
rect 23805 18005 23845 18045
rect 23855 18005 23895 18045
rect 23905 18005 23945 18045
rect 23955 18005 23995 18045
rect 24005 18005 24045 18045
rect 24055 18005 24095 18045
rect 24105 18005 24145 18045
rect 24155 18005 24195 18045
rect 24205 18005 24245 18045
rect 24255 18005 24295 18045
rect 24305 18005 24345 18045
rect 24355 18005 24395 18045
rect 24405 18005 24445 18045
rect 24455 18005 24495 18045
rect 24505 18005 24545 18045
rect 24555 18005 24595 18045
rect 24605 18005 24645 18045
rect 24655 18005 24695 18045
rect 24705 18005 24745 18045
rect 24755 18005 24795 18045
rect 24805 18005 24845 18045
rect 24855 18005 24895 18045
rect 24905 18005 24945 18045
rect 24955 18005 24995 18045
rect 25005 18005 25045 18045
rect 25055 18005 25095 18045
rect 25105 18005 25145 18045
rect 25155 18005 25195 18045
rect 25205 18005 25245 18045
rect 25255 18005 25295 18045
rect 25305 18005 25345 18045
rect 25355 18005 25395 18045
rect 25405 18005 25445 18045
rect 25455 18005 25495 18045
rect 25505 18005 25545 18045
rect 25555 18005 25595 18045
rect 25605 18005 25645 18045
rect 25655 18005 25695 18045
rect 25705 18005 25745 18045
rect 25755 18005 25795 18045
rect 25805 18005 25845 18045
rect 25855 18005 25895 18045
rect 25905 18005 25945 18045
rect 25955 18005 25995 18045
rect 26005 18005 26045 18045
rect 26055 18005 26095 18045
rect 26105 18005 26145 18045
rect 26155 18005 26195 18045
rect 26205 18005 26245 18045
rect 26255 18005 26295 18045
rect 26305 18005 26345 18045
rect 26355 18005 26395 18045
rect 26405 18005 26445 18045
rect 26455 18005 26495 18045
rect 26505 18005 26545 18045
rect 26555 18005 26595 18045
rect 26605 18005 26645 18045
rect 26655 18005 26695 18045
rect 26705 18005 26745 18045
rect 26755 18005 26795 18045
rect 26805 18005 26845 18045
rect 26855 18005 26895 18045
rect 26905 18005 26945 18045
rect 26955 18005 26995 18045
rect 27005 18005 27045 18045
rect 27055 18005 27095 18045
rect 27105 18005 27145 18045
rect 27155 18005 27195 18045
rect 27205 18005 27245 18045
rect 27255 18005 27295 18045
rect 27305 18005 27345 18045
rect 27355 18005 27395 18045
rect 27405 18005 27445 18045
rect 27455 18005 27495 18045
rect 27505 18005 27545 18045
rect 27555 18005 27595 18045
rect 27605 18005 27645 18045
rect 27655 18005 27695 18045
rect 27705 18005 27745 18045
rect 27755 18005 27795 18045
rect 27805 18005 27845 18045
rect 27855 18005 27895 18045
rect 27905 18005 27945 18045
rect 27955 18005 27995 18045
rect 28005 18005 28045 18045
rect 28055 18005 28095 18045
rect 28105 18005 28145 18045
rect 28155 18005 28195 18045
rect 28205 18005 28245 18045
rect 28255 18005 28295 18045
rect 28305 18005 28345 18045
rect 28355 18005 28395 18045
rect 28405 18005 28445 18045
rect 28455 18005 28495 18045
rect 28505 18005 28545 18045
rect 28555 18005 28595 18045
rect 28605 18005 28645 18045
rect 28655 18005 28695 18045
rect 28705 18005 28745 18045
rect 28755 18005 28795 18045
rect 28805 18005 28845 18045
rect 28855 18005 28895 18045
rect 28905 18005 28945 18045
rect 28955 18005 28995 18045
rect 29005 18005 29045 18045
rect 29055 18005 29095 18045
rect 29105 18005 29145 18045
rect 29155 18005 29195 18045
rect 29205 18005 29245 18045
rect 29255 18005 29295 18045
rect 29305 18005 29345 18045
rect 29355 18005 29395 18045
rect 29405 18005 29445 18045
rect 29455 18005 29495 18045
rect 29505 18005 29545 18045
rect 29555 18005 29595 18045
rect 29605 18005 29645 18045
rect 29655 18005 29695 18045
rect 29705 18005 29745 18045
rect 29755 18005 29795 18045
rect 29805 18005 29845 18045
rect 29855 18005 29895 18045
rect 29905 18005 29945 18045
rect 29955 18005 29995 18045
rect 30005 18005 30045 18045
rect 30055 18005 30095 18045
rect 30105 18005 30145 18045
rect 30155 18005 30195 18045
rect 30205 18005 30245 18045
rect 30255 18005 30295 18045
rect 30305 18005 30345 18045
rect 30355 18005 30395 18045
rect 30405 18005 30445 18045
rect 30455 18005 30495 18045
rect 30505 18005 30545 18045
rect 30555 18005 30595 18045
rect 30605 18005 30645 18045
rect 30655 18005 30695 18045
rect 30705 18005 30745 18045
rect 30755 18005 30795 18045
rect 30805 18005 30845 18045
rect 30855 18005 30895 18045
rect 30905 18005 30945 18045
rect 30955 18005 30995 18045
rect 31005 18005 31045 18045
rect 31055 18005 31095 18045
rect 31105 18005 31145 18045
rect 31155 18005 31195 18045
rect 31205 18005 31245 18045
rect 31255 18005 31295 18045
rect 31305 18005 31345 18045
rect 31355 18005 31395 18045
rect 31405 18005 31445 18045
rect 31455 18005 31495 18045
rect 31505 18005 31545 18045
rect 31555 18005 31595 18045
rect 31605 18005 31645 18045
rect 31655 18005 31695 18045
rect 31705 18005 31745 18045
rect 31755 18005 31795 18045
rect 31805 18005 31845 18045
rect 31855 18005 31895 18045
rect 31905 18005 31945 18045
rect 31955 18005 31995 18045
rect 32005 18005 32045 18045
rect 32055 18005 32095 18045
rect 32105 18005 32145 18045
rect 32155 18005 32195 18045
rect 32205 18005 32245 18045
rect 32255 18005 32295 18045
rect 32305 18005 32345 18045
rect 32355 18005 32395 18045
rect 32405 18005 32445 18045
rect 32455 18005 32495 18045
rect 32505 18005 32545 18045
rect 32555 18005 32595 18045
rect 32605 18005 32645 18045
rect 32655 18005 32695 18045
rect 32705 18005 32745 18045
rect 32755 18005 32795 18045
rect 32805 18005 32845 18045
rect 32855 18005 32895 18045
rect 32905 18005 32945 18045
rect 32955 18005 32995 18045
rect 33005 18005 33045 18045
rect 33055 18005 33095 18045
rect 33105 18005 33145 18045
rect 33155 18005 33195 18045
rect 33205 18005 33245 18045
rect 33255 18005 33295 18045
rect 33305 18005 33345 18045
rect 33355 18005 33395 18045
rect 33405 18005 33445 18045
rect 33455 18005 33495 18045
rect 33505 18005 33545 18045
rect 33555 18005 33595 18045
rect 33605 18005 33645 18045
rect 33655 18005 33695 18045
rect 33705 18005 33745 18045
rect 33755 18005 33795 18045
rect 33805 18005 33845 18045
rect 33855 18005 33895 18045
rect 33905 18005 33945 18045
rect 33955 18005 33995 18045
rect 34005 18005 34045 18045
rect 34055 18005 34095 18045
rect 34105 18005 34145 18045
rect 34155 18005 34195 18045
rect 34205 18005 34245 18045
rect 34255 18005 34295 18045
rect 34305 18005 34345 18045
rect 34355 18005 34395 18045
rect 34405 18005 34445 18045
rect 34455 18005 34495 18045
rect 34505 18005 34545 18045
rect 34555 18005 34595 18045
rect 34605 18005 34645 18045
rect 34655 18005 34695 18045
rect 34705 18005 34745 18045
rect 34755 18005 34795 18045
rect 34805 18005 34845 18045
rect 34855 18005 34895 18045
rect 34905 18005 34945 18045
rect 34955 18005 34995 18045
rect 35005 18005 35045 18045
rect 35055 18005 35095 18045
rect 35105 18005 35145 18045
rect 35155 18005 35195 18045
rect 35205 18005 35245 18045
rect 35255 18005 35295 18045
rect 35305 18005 35345 18045
rect 35355 18005 35395 18045
rect 35405 18005 35445 18045
rect 35455 18005 35495 18045
rect 35505 18005 35545 18045
rect 35555 18005 35595 18045
rect 35605 18005 35645 18045
rect 35655 18005 35695 18045
rect 35705 18005 35745 18045
rect 35755 18005 35795 18045
rect 35805 18005 35845 18045
rect 35855 18005 35895 18045
rect 35905 18005 35945 18045
rect 35955 18005 35995 18045
rect 36005 18005 36045 18045
rect 36055 18005 36095 18045
rect 36105 18005 36145 18045
rect 36155 18005 36195 18045
rect 36205 18005 36245 18045
rect 36255 18005 36295 18045
rect 36305 18005 36345 18045
rect 36355 18005 36395 18045
rect 36405 18005 36445 18045
rect 36455 18005 36495 18045
rect 36505 18005 36545 18045
rect 36555 18005 36595 18045
rect 36605 18005 36645 18045
rect 36655 18005 36695 18045
rect 36705 18005 36745 18045
rect 36755 18005 36795 18045
rect 36805 18005 36845 18045
rect 36855 18005 36895 18045
rect 36905 18005 36945 18045
rect 36955 18005 36995 18045
rect 37005 18005 37045 18045
rect 37055 18005 37095 18045
rect 37105 18005 37145 18045
rect 37155 18005 37195 18045
rect 37205 18005 37245 18045
rect 37255 18005 37295 18045
rect 37305 18005 37345 18045
rect 37355 18005 37395 18045
rect 37405 18005 37445 18045
rect 37455 18005 37495 18045
rect 37505 18005 37545 18045
rect 37555 18005 37595 18045
rect 37605 18005 37645 18045
rect 37655 18005 37695 18045
rect 37705 18005 37745 18045
rect 37755 18005 37795 18045
rect 37805 18005 37845 18045
rect 37855 18005 37895 18045
rect 37905 18005 37945 18045
rect 37955 18005 37995 18045
rect 38005 18005 38045 18045
rect 38055 18005 38095 18045
rect 38105 18005 38145 18045
rect 38155 18005 38195 18045
rect 38205 18005 38245 18045
rect 38255 18005 38295 18045
rect 38305 18005 38345 18045
rect 38355 18005 38395 18045
rect 38405 18005 38445 18045
rect 38455 18005 38495 18045
rect 38505 18005 38545 18045
rect 38555 18005 38595 18045
rect 38605 18005 38645 18045
rect 38655 18005 38695 18045
rect 38705 18005 38745 18045
rect 38755 18005 38795 18045
rect 38805 18005 38845 18045
rect 38855 18005 38895 18045
rect 38905 18005 38945 18045
rect 38955 18005 38995 18045
rect 39005 18005 39045 18045
rect 39055 18005 39095 18045
rect 39105 18005 39145 18045
rect 39155 18005 39195 18045
rect 39205 18005 39245 18045
rect 39255 18005 39295 18045
rect 39305 18005 39345 18045
rect 39355 18005 39395 18045
rect 39405 18005 39445 18045
rect 39455 18005 39495 18045
rect 39505 18005 39545 18045
rect 39555 18005 39595 18045
rect 39605 18005 39645 18045
rect 39655 18005 39695 18045
rect 39705 18005 39745 18045
rect -2695 17005 -2655 17045
rect 105 17005 145 17045
rect 155 17005 195 17045
rect 205 17005 245 17045
rect 255 17005 295 17045
rect 305 17005 345 17045
rect 355 17005 395 17045
rect 405 17005 445 17045
rect 455 17005 495 17045
rect 505 17005 545 17045
rect 555 17005 595 17045
rect 605 17005 645 17045
rect 655 17005 695 17045
rect 705 17005 745 17045
rect 755 17005 795 17045
rect 805 17005 845 17045
rect 855 17005 895 17045
rect 905 17005 945 17045
rect 955 17005 995 17045
rect 1005 17005 1045 17045
rect 1055 17005 1095 17045
rect 1105 17005 1145 17045
rect 1155 17005 1195 17045
rect 1205 17005 1245 17045
rect 1255 17005 1295 17045
rect 1305 17005 1345 17045
rect 1355 17005 1395 17045
rect 1405 17005 1445 17045
rect 1455 17005 1495 17045
rect 1505 17005 1545 17045
rect 1555 17005 1595 17045
rect 1605 17005 1645 17045
rect 1655 17005 1695 17045
rect 1705 17005 1745 17045
rect 1755 17005 1795 17045
rect 1805 17005 1845 17045
rect 1855 17005 1895 17045
rect 1905 17005 1945 17045
rect 1955 17005 1995 17045
rect 2005 17005 2045 17045
rect 2055 17005 2095 17045
rect 2105 17005 2145 17045
rect 2155 17005 2195 17045
rect 2205 17005 2245 17045
rect 2255 17005 2295 17045
rect 2305 17005 2345 17045
rect 2355 17005 2395 17045
rect 2405 17005 2445 17045
rect 2455 17005 2495 17045
rect 2505 17005 2545 17045
rect 2555 17005 2595 17045
rect 2605 17005 2645 17045
rect 2655 17005 2695 17045
rect 2705 17005 2745 17045
rect 2755 17005 2795 17045
rect 2805 17005 2845 17045
rect 2855 17005 2895 17045
rect 2905 17005 2945 17045
rect 2955 17005 2995 17045
rect 3005 17005 3045 17045
rect 3055 17005 3095 17045
rect 3105 17005 3145 17045
rect 3155 17005 3195 17045
rect 3205 17005 3245 17045
rect 3255 17005 3295 17045
rect 3305 17005 3345 17045
rect 3355 17005 3395 17045
rect 3405 17005 3445 17045
rect 3455 17005 3495 17045
rect 3505 17005 3545 17045
rect 3555 17005 3595 17045
rect 3605 17005 3645 17045
rect 3655 17005 3695 17045
rect 3705 17005 3745 17045
rect 3755 17005 3795 17045
rect 3805 17005 3845 17045
rect 3855 17005 3895 17045
rect 3905 17005 3945 17045
rect 3955 17005 3995 17045
rect 4005 17005 4045 17045
rect 4055 17005 4095 17045
rect 4105 17005 4145 17045
rect 4155 17005 4195 17045
rect 4205 17005 4245 17045
rect 4255 17005 4295 17045
rect 4305 17005 4345 17045
rect 4355 17005 4395 17045
rect 4405 17005 4445 17045
rect 4455 17005 4495 17045
rect 4505 17005 4545 17045
rect 4555 17005 4595 17045
rect 4605 17005 4645 17045
rect 4655 17005 4695 17045
rect 4705 17005 4745 17045
rect 4755 17005 4795 17045
rect 4805 17005 4845 17045
rect 4855 17005 4895 17045
rect 4905 17005 4945 17045
rect 4955 17005 4995 17045
rect 5005 17005 5045 17045
rect 5055 17005 5095 17045
rect 5105 17005 5145 17045
rect 5155 17005 5195 17045
rect 5205 17005 5245 17045
rect 5255 17005 5295 17045
rect 5305 17005 5345 17045
rect 5355 17005 5395 17045
rect 5405 17005 5445 17045
rect 5455 17005 5495 17045
rect 5505 17005 5545 17045
rect 5555 17005 5595 17045
rect 5605 17005 5645 17045
rect 5655 17005 5695 17045
rect 5705 17005 5745 17045
rect 5755 17005 5795 17045
rect 5805 17005 5845 17045
rect 5855 17005 5895 17045
rect 5905 17005 5945 17045
rect 5955 17005 5995 17045
rect 6005 17005 6045 17045
rect 6055 17005 6095 17045
rect 6105 17005 6145 17045
rect 6155 17005 6195 17045
rect 6205 17005 6245 17045
rect 6255 17005 6295 17045
rect 6305 17005 6345 17045
rect 6355 17005 6395 17045
rect 6405 17005 6445 17045
rect 6455 17005 6495 17045
rect 6505 17005 6545 17045
rect 6555 17005 6595 17045
rect 6605 17005 6645 17045
rect 6655 17005 6695 17045
rect 6705 17005 6745 17045
rect 6755 17005 6795 17045
rect 6805 17005 6845 17045
rect 6855 17005 6895 17045
rect 6905 17005 6945 17045
rect 6955 17005 6995 17045
rect 7005 17005 7045 17045
rect 7055 17005 7095 17045
rect 7105 17005 7145 17045
rect 7155 17005 7195 17045
rect 7205 17005 7245 17045
rect 7255 17005 7295 17045
rect 7305 17005 7345 17045
rect 7355 17005 7395 17045
rect 7405 17005 7445 17045
rect 7455 17005 7495 17045
rect 7505 17005 7545 17045
rect 7555 17005 7595 17045
rect 7605 17005 7645 17045
rect 7655 17005 7695 17045
rect 7705 17005 7745 17045
rect 7755 17005 7795 17045
rect 7805 17005 7845 17045
rect 7855 17005 7895 17045
rect 7905 17005 7945 17045
rect 7955 17005 7995 17045
rect 8005 17005 8045 17045
rect 8055 17005 8095 17045
rect 8105 17005 8145 17045
rect 8155 17005 8195 17045
rect 8205 17005 8245 17045
rect 8255 17005 8295 17045
rect 8305 17005 8345 17045
rect 8355 17005 8395 17045
rect 8405 17005 8445 17045
rect 8455 17005 8495 17045
rect 8505 17005 8545 17045
rect 8555 17005 8595 17045
rect 8605 17005 8645 17045
rect 8655 17005 8695 17045
rect 8705 17005 8745 17045
rect 8755 17005 8795 17045
rect 8805 17005 8845 17045
rect 8855 17005 8895 17045
rect 8905 17005 8945 17045
rect 8955 17005 8995 17045
rect 9005 17005 9045 17045
rect 9055 17005 9095 17045
rect 9105 17005 9145 17045
rect 9155 17005 9195 17045
rect 9205 17005 9245 17045
rect 9255 17005 9295 17045
rect 9305 17005 9345 17045
rect 9355 17005 9395 17045
rect 9405 17005 9445 17045
rect 9455 17005 9495 17045
rect 9505 17005 9545 17045
rect 9555 17005 9595 17045
rect 9605 17005 9645 17045
rect 9655 17005 9695 17045
rect 9705 17005 9745 17045
rect 9755 17005 9795 17045
rect 9805 17005 9845 17045
rect 9855 17005 9895 17045
rect 9905 17005 9945 17045
rect 9955 17005 9995 17045
rect 10005 17005 10045 17045
rect 10055 17005 10095 17045
rect 10105 17005 10145 17045
rect 10155 17005 10195 17045
rect 10205 17005 10245 17045
rect 10255 17005 10295 17045
rect 10305 17005 10345 17045
rect 10355 17005 10395 17045
rect 10405 17005 10445 17045
rect 10455 17005 10495 17045
rect 10505 17005 10545 17045
rect 10555 17005 10595 17045
rect 10605 17005 10645 17045
rect 10655 17005 10695 17045
rect 10705 17005 10745 17045
rect 10755 17005 10795 17045
rect 10805 17005 10845 17045
rect 10855 17005 10895 17045
rect 10905 17005 10945 17045
rect 10955 17005 10995 17045
rect 11005 17005 11045 17045
rect 11055 17005 11095 17045
rect 11105 17005 11145 17045
rect 11155 17005 11195 17045
rect 11205 17005 11245 17045
rect 11255 17005 11295 17045
rect 11305 17005 11345 17045
rect 11355 17005 11395 17045
rect 11405 17005 11445 17045
rect 11455 17005 11495 17045
rect 11505 17005 11545 17045
rect 11555 17005 11595 17045
rect 11605 17005 11645 17045
rect 11655 17005 11695 17045
rect 11705 17005 11745 17045
rect 11755 17005 11795 17045
rect 11805 17005 11845 17045
rect 11855 17005 11895 17045
rect 11905 17005 11945 17045
rect 11955 17005 11995 17045
rect 12005 17005 12045 17045
rect 12055 17005 12095 17045
rect 12105 17005 12145 17045
rect 12155 17005 12195 17045
rect 12205 17005 12245 17045
rect 12255 17005 12295 17045
rect 12305 17005 12345 17045
rect 12355 17005 12395 17045
rect 12405 17005 12445 17045
rect 12455 17005 12495 17045
rect 12505 17005 12545 17045
rect 12555 17005 12595 17045
rect 12605 17005 12645 17045
rect 12655 17005 12695 17045
rect 12705 17005 12745 17045
rect 12755 17005 12795 17045
rect 12805 17005 12845 17045
rect 12855 17005 12895 17045
rect 12905 17005 12945 17045
rect 12955 17005 12995 17045
rect 13005 17005 13045 17045
rect 13055 17005 13095 17045
rect 13105 17005 13145 17045
rect 13155 17005 13195 17045
rect 13205 17005 13245 17045
rect 13255 17005 13295 17045
rect 13305 17005 13345 17045
rect 13355 17005 13395 17045
rect 13405 17005 13445 17045
rect 13455 17005 13495 17045
rect 13505 17005 13545 17045
rect 13555 17005 13595 17045
rect 13605 17005 13645 17045
rect 13655 17005 13695 17045
rect 13705 17005 13745 17045
rect 13755 17005 13795 17045
rect 13805 17005 13845 17045
rect 13855 17005 13895 17045
rect 13905 17005 13945 17045
rect 13955 17005 13995 17045
rect 14005 17005 14045 17045
rect 14055 17005 14095 17045
rect 14105 17005 14145 17045
rect 14155 17005 14195 17045
rect 14205 17005 14245 17045
rect 14255 17005 14295 17045
rect 14305 17005 14345 17045
rect 14355 17005 14395 17045
rect 14405 17005 14445 17045
rect 14455 17005 14495 17045
rect 14505 17005 14545 17045
rect 14555 17005 14595 17045
rect 14605 17005 14645 17045
rect 14655 17005 14695 17045
rect 14705 17005 14745 17045
rect 14755 17005 14795 17045
rect 14805 17005 14845 17045
rect 14855 17005 14895 17045
rect 14905 17005 14945 17045
rect 14955 17005 14995 17045
rect 15005 17005 15045 17045
rect 15055 17005 15095 17045
rect 15105 17005 15145 17045
rect 15155 17005 15195 17045
rect 15205 17005 15245 17045
rect 15255 17005 15295 17045
rect 15305 17005 15345 17045
rect 15355 17005 15395 17045
rect 15405 17005 15445 17045
rect 15455 17005 15495 17045
rect 15505 17005 15545 17045
rect 15555 17005 15595 17045
rect 15605 17005 15645 17045
rect 15655 17005 15695 17045
rect 15705 17005 15745 17045
rect 15755 17005 15795 17045
rect 15805 17005 15845 17045
rect 15855 17005 15895 17045
rect 15905 17005 15945 17045
rect 15955 17005 15995 17045
rect 16005 17005 16045 17045
rect 16055 17005 16095 17045
rect 16105 17005 16145 17045
rect 16155 17005 16195 17045
rect 16205 17005 16245 17045
rect 16255 17005 16295 17045
rect 16305 17005 16345 17045
rect 16355 17005 16395 17045
rect 16405 17005 16445 17045
rect 16455 17005 16495 17045
rect 16505 17005 16545 17045
rect 16555 17005 16595 17045
rect 16605 17005 16645 17045
rect 16655 17005 16695 17045
rect 16705 17005 16745 17045
rect 16755 17005 16795 17045
rect 16805 17005 16845 17045
rect 16855 17005 16895 17045
rect 16905 17005 16945 17045
rect 16955 17005 16995 17045
rect 17005 17005 17045 17045
rect 17055 17005 17095 17045
rect 17105 17005 17145 17045
rect 17155 17005 17195 17045
rect 17205 17005 17245 17045
rect 17255 17005 17295 17045
rect 17305 17005 17345 17045
rect 17355 17005 17395 17045
rect 17405 17005 17445 17045
rect 17455 17005 17495 17045
rect 17505 17005 17545 17045
rect 17555 17005 17595 17045
rect 17605 17005 17645 17045
rect 17655 17005 17695 17045
rect 17705 17005 17745 17045
rect 17755 17005 17795 17045
rect 17805 17005 17845 17045
rect 17855 17005 17895 17045
rect 17905 17005 17945 17045
rect 17955 17005 17995 17045
rect 18005 17005 18045 17045
rect 18055 17005 18095 17045
rect 18105 17005 18145 17045
rect 18155 17005 18195 17045
rect 18205 17005 18245 17045
rect 18255 17005 18295 17045
rect 18305 17005 18345 17045
rect 18355 17005 18395 17045
rect 18405 17005 18445 17045
rect 18455 17005 18495 17045
rect 18505 17005 18545 17045
rect 18555 17005 18595 17045
rect 18605 17005 18645 17045
rect 18655 17005 18695 17045
rect 18705 17005 18745 17045
rect 18755 17005 18795 17045
rect 18805 17005 18845 17045
rect 18855 17005 18895 17045
rect 18905 17005 18945 17045
rect 18955 17005 18995 17045
rect 19005 17005 19045 17045
rect 19055 17005 19095 17045
rect 19105 17005 19145 17045
rect 19155 17005 19195 17045
rect 19205 17005 19245 17045
rect 19255 17005 19295 17045
rect 19305 17005 19345 17045
rect 19355 17005 19395 17045
rect 19405 17005 19445 17045
rect 19455 17005 19495 17045
rect 19505 17005 19545 17045
rect 19555 17005 19595 17045
rect 19605 17005 19645 17045
rect 19655 17005 19695 17045
rect 19705 17005 19745 17045
rect 19755 17005 19795 17045
rect 19805 17005 19845 17045
rect 19855 17005 19895 17045
rect 19905 17005 19945 17045
rect 19955 17005 19995 17045
rect 20005 17005 20045 17045
rect 20055 17005 20095 17045
rect 20105 17005 20145 17045
rect 20155 17005 20195 17045
rect 20205 17005 20245 17045
rect 20255 17005 20295 17045
rect 20305 17005 20345 17045
rect 20355 17005 20395 17045
rect 20405 17005 20445 17045
rect 20455 17005 20495 17045
rect 20505 17005 20545 17045
rect 20555 17005 20595 17045
rect 20605 17005 20645 17045
rect 20655 17005 20695 17045
rect 20705 17005 20745 17045
rect 20755 17005 20795 17045
rect 20805 17005 20845 17045
rect 20855 17005 20895 17045
rect 20905 17005 20945 17045
rect 20955 17005 20995 17045
rect 21005 17005 21045 17045
rect 21055 17005 21095 17045
rect 21105 17005 21145 17045
rect 21155 17005 21195 17045
rect 21205 17005 21245 17045
rect 21255 17005 21295 17045
rect 21305 17005 21345 17045
rect 21355 17005 21395 17045
rect 21405 17005 21445 17045
rect 21455 17005 21495 17045
rect 21505 17005 21545 17045
rect 21555 17005 21595 17045
rect 21605 17005 21645 17045
rect 21655 17005 21695 17045
rect 21705 17005 21745 17045
rect 21755 17005 21795 17045
rect 21805 17005 21845 17045
rect 21855 17005 21895 17045
rect 21905 17005 21945 17045
rect 21955 17005 21995 17045
rect 22005 17005 22045 17045
rect 22055 17005 22095 17045
rect 22105 17005 22145 17045
rect 22155 17005 22195 17045
rect 22205 17005 22245 17045
rect 22255 17005 22295 17045
rect 22305 17005 22345 17045
rect 22355 17005 22395 17045
rect 22405 17005 22445 17045
rect 22455 17005 22495 17045
rect 22505 17005 22545 17045
rect 22555 17005 22595 17045
rect 22605 17005 22645 17045
rect 22655 17005 22695 17045
rect 22705 17005 22745 17045
rect 22755 17005 22795 17045
rect 22805 17005 22845 17045
rect 22855 17005 22895 17045
rect 22905 17005 22945 17045
rect 22955 17005 22995 17045
rect 23005 17005 23045 17045
rect 23055 17005 23095 17045
rect 23105 17005 23145 17045
rect 23155 17005 23195 17045
rect 23205 17005 23245 17045
rect 23255 17005 23295 17045
rect 23305 17005 23345 17045
rect 23355 17005 23395 17045
rect 23405 17005 23445 17045
rect 23455 17005 23495 17045
rect 23505 17005 23545 17045
rect 23555 17005 23595 17045
rect 23605 17005 23645 17045
rect 23655 17005 23695 17045
rect 23705 17005 23745 17045
rect 23755 17005 23795 17045
rect 23805 17005 23845 17045
rect 23855 17005 23895 17045
rect 23905 17005 23945 17045
rect 23955 17005 23995 17045
rect 24005 17005 24045 17045
rect 24055 17005 24095 17045
rect 24105 17005 24145 17045
rect 24155 17005 24195 17045
rect 24205 17005 24245 17045
rect 24255 17005 24295 17045
rect 24305 17005 24345 17045
rect 24355 17005 24395 17045
rect 24405 17005 24445 17045
rect 24455 17005 24495 17045
rect 24505 17005 24545 17045
rect 24555 17005 24595 17045
rect 24605 17005 24645 17045
rect 24655 17005 24695 17045
rect 24705 17005 24745 17045
rect 24755 17005 24795 17045
rect 24805 17005 24845 17045
rect 24855 17005 24895 17045
rect 24905 17005 24945 17045
rect 24955 17005 24995 17045
rect 25005 17005 25045 17045
rect 25055 17005 25095 17045
rect 25105 17005 25145 17045
rect 25155 17005 25195 17045
rect 25205 17005 25245 17045
rect 25255 17005 25295 17045
rect 25305 17005 25345 17045
rect 25355 17005 25395 17045
rect 25405 17005 25445 17045
rect 25455 17005 25495 17045
rect 25505 17005 25545 17045
rect 25555 17005 25595 17045
rect 25605 17005 25645 17045
rect 25655 17005 25695 17045
rect 25705 17005 25745 17045
rect 25755 17005 25795 17045
rect 25805 17005 25845 17045
rect 25855 17005 25895 17045
rect 25905 17005 25945 17045
rect 25955 17005 25995 17045
rect 26005 17005 26045 17045
rect 26055 17005 26095 17045
rect 26105 17005 26145 17045
rect 26155 17005 26195 17045
rect 26205 17005 26245 17045
rect 26255 17005 26295 17045
rect 26305 17005 26345 17045
rect 26355 17005 26395 17045
rect 26405 17005 26445 17045
rect 26455 17005 26495 17045
rect 26505 17005 26545 17045
rect 26555 17005 26595 17045
rect 26605 17005 26645 17045
rect 26655 17005 26695 17045
rect 26705 17005 26745 17045
rect 26755 17005 26795 17045
rect 26805 17005 26845 17045
rect 26855 17005 26895 17045
rect 26905 17005 26945 17045
rect 26955 17005 26995 17045
rect 27005 17005 27045 17045
rect 27055 17005 27095 17045
rect 27105 17005 27145 17045
rect 27155 17005 27195 17045
rect 27205 17005 27245 17045
rect 27255 17005 27295 17045
rect 27305 17005 27345 17045
rect 27355 17005 27395 17045
rect 27405 17005 27445 17045
rect 27455 17005 27495 17045
rect 27505 17005 27545 17045
rect 27555 17005 27595 17045
rect 27605 17005 27645 17045
rect 27655 17005 27695 17045
rect 27705 17005 27745 17045
rect 27755 17005 27795 17045
rect 27805 17005 27845 17045
rect 27855 17005 27895 17045
rect 27905 17005 27945 17045
rect 27955 17005 27995 17045
rect 28005 17005 28045 17045
rect 28055 17005 28095 17045
rect 28105 17005 28145 17045
rect 28155 17005 28195 17045
rect 28205 17005 28245 17045
rect 28255 17005 28295 17045
rect 28305 17005 28345 17045
rect 28355 17005 28395 17045
rect 28405 17005 28445 17045
rect 28455 17005 28495 17045
rect 28505 17005 28545 17045
rect 28555 17005 28595 17045
rect 28605 17005 28645 17045
rect 28655 17005 28695 17045
rect 28705 17005 28745 17045
rect 28755 17005 28795 17045
rect 28805 17005 28845 17045
rect 28855 17005 28895 17045
rect 28905 17005 28945 17045
rect 28955 17005 28995 17045
rect 29005 17005 29045 17045
rect 29055 17005 29095 17045
rect 29105 17005 29145 17045
rect 29155 17005 29195 17045
rect 29205 17005 29245 17045
rect 29255 17005 29295 17045
rect 29305 17005 29345 17045
rect 29355 17005 29395 17045
rect 29405 17005 29445 17045
rect 29455 17005 29495 17045
rect 29505 17005 29545 17045
rect 29555 17005 29595 17045
rect 29605 17005 29645 17045
rect 29655 17005 29695 17045
rect 29705 17005 29745 17045
rect 29755 17005 29795 17045
rect 29805 17005 29845 17045
rect 29855 17005 29895 17045
rect 29905 17005 29945 17045
rect 29955 17005 29995 17045
rect 30005 17005 30045 17045
rect 30055 17005 30095 17045
rect 30105 17005 30145 17045
rect 30155 17005 30195 17045
rect 30205 17005 30245 17045
rect 30255 17005 30295 17045
rect 30305 17005 30345 17045
rect 30355 17005 30395 17045
rect 30405 17005 30445 17045
rect 30455 17005 30495 17045
rect 30505 17005 30545 17045
rect 30555 17005 30595 17045
rect 30605 17005 30645 17045
rect 30655 17005 30695 17045
rect 30705 17005 30745 17045
rect 30755 17005 30795 17045
rect 30805 17005 30845 17045
rect 30855 17005 30895 17045
rect 30905 17005 30945 17045
rect 30955 17005 30995 17045
rect 31005 17005 31045 17045
rect 31055 17005 31095 17045
rect 31105 17005 31145 17045
rect 31155 17005 31195 17045
rect 31205 17005 31245 17045
rect 31255 17005 31295 17045
rect 31305 17005 31345 17045
rect 31355 17005 31395 17045
rect 31405 17005 31445 17045
rect 31455 17005 31495 17045
rect 31505 17005 31545 17045
rect 31555 17005 31595 17045
rect 31605 17005 31645 17045
rect 31655 17005 31695 17045
rect 31705 17005 31745 17045
rect 31755 17005 31795 17045
rect 31805 17005 31845 17045
rect 31855 17005 31895 17045
rect 31905 17005 31945 17045
rect 31955 17005 31995 17045
rect 32005 17005 32045 17045
rect 32055 17005 32095 17045
rect 32105 17005 32145 17045
rect 32155 17005 32195 17045
rect 32205 17005 32245 17045
rect 32255 17005 32295 17045
rect 32305 17005 32345 17045
rect 32355 17005 32395 17045
rect 32405 17005 32445 17045
rect 32455 17005 32495 17045
rect 32505 17005 32545 17045
rect 32555 17005 32595 17045
rect 32605 17005 32645 17045
rect 32655 17005 32695 17045
rect 32705 17005 32745 17045
rect 32755 17005 32795 17045
rect 32805 17005 32845 17045
rect 32855 17005 32895 17045
rect 32905 17005 32945 17045
rect 32955 17005 32995 17045
rect 33005 17005 33045 17045
rect 33055 17005 33095 17045
rect 33105 17005 33145 17045
rect 33155 17005 33195 17045
rect 33205 17005 33245 17045
rect 33255 17005 33295 17045
rect 33305 17005 33345 17045
rect 33355 17005 33395 17045
rect 33405 17005 33445 17045
rect 33455 17005 33495 17045
rect 33505 17005 33545 17045
rect 33555 17005 33595 17045
rect 33605 17005 33645 17045
rect 33655 17005 33695 17045
rect 33705 17005 33745 17045
rect 33755 17005 33795 17045
rect 33805 17005 33845 17045
rect 33855 17005 33895 17045
rect 33905 17005 33945 17045
rect 33955 17005 33995 17045
rect 34005 17005 34045 17045
rect 34055 17005 34095 17045
rect 34105 17005 34145 17045
rect 34155 17005 34195 17045
rect 34205 17005 34245 17045
rect 34255 17005 34295 17045
rect 34305 17005 34345 17045
rect 34355 17005 34395 17045
rect 34405 17005 34445 17045
rect 34455 17005 34495 17045
rect 34505 17005 34545 17045
rect 34555 17005 34595 17045
rect 34605 17005 34645 17045
rect 34655 17005 34695 17045
rect 34705 17005 34745 17045
rect 34755 17005 34795 17045
rect 34805 17005 34845 17045
rect 34855 17005 34895 17045
rect 34905 17005 34945 17045
rect 34955 17005 34995 17045
rect 35005 17005 35045 17045
rect 35055 17005 35095 17045
rect 35105 17005 35145 17045
rect 35155 17005 35195 17045
rect 35205 17005 35245 17045
rect 35255 17005 35295 17045
rect 35305 17005 35345 17045
rect 35355 17005 35395 17045
rect 35405 17005 35445 17045
rect 35455 17005 35495 17045
rect 35505 17005 35545 17045
rect 35555 17005 35595 17045
rect 35605 17005 35645 17045
rect 35655 17005 35695 17045
rect 35705 17005 35745 17045
rect 35755 17005 35795 17045
rect 35805 17005 35845 17045
rect 35855 17005 35895 17045
rect 35905 17005 35945 17045
rect 35955 17005 35995 17045
rect 36005 17005 36045 17045
rect 36055 17005 36095 17045
rect 36105 17005 36145 17045
rect 36155 17005 36195 17045
rect 36205 17005 36245 17045
rect 36255 17005 36295 17045
rect 36305 17005 36345 17045
rect 36355 17005 36395 17045
rect 36405 17005 36445 17045
rect 36455 17005 36495 17045
rect 36505 17005 36545 17045
rect 36555 17005 36595 17045
rect 36605 17005 36645 17045
rect 36655 17005 36695 17045
rect 36705 17005 36745 17045
rect 36755 17005 36795 17045
rect 36805 17005 36845 17045
rect 36855 17005 36895 17045
rect 36905 17005 36945 17045
rect 36955 17005 36995 17045
rect 37005 17005 37045 17045
rect 37055 17005 37095 17045
rect 37105 17005 37145 17045
rect 37155 17005 37195 17045
rect 37205 17005 37245 17045
rect 37255 17005 37295 17045
rect 37305 17005 37345 17045
rect 37355 17005 37395 17045
rect 37405 17005 37445 17045
rect 37455 17005 37495 17045
rect 37505 17005 37545 17045
rect 37555 17005 37595 17045
rect 37605 17005 37645 17045
rect 37655 17005 37695 17045
rect 37705 17005 37745 17045
rect 37755 17005 37795 17045
rect 37805 17005 37845 17045
rect 37855 17005 37895 17045
rect 37905 17005 37945 17045
rect 37955 17005 37995 17045
rect 38005 17005 38045 17045
rect 38055 17005 38095 17045
rect 38105 17005 38145 17045
rect 38155 17005 38195 17045
rect 38205 17005 38245 17045
rect 38255 17005 38295 17045
rect 38305 17005 38345 17045
rect 38355 17005 38395 17045
rect 38405 17005 38445 17045
rect 38455 17005 38495 17045
rect 38505 17005 38545 17045
rect 38555 17005 38595 17045
rect 38605 17005 38645 17045
rect 38655 17005 38695 17045
rect 38705 17005 38745 17045
rect 38755 17005 38795 17045
rect 38805 17005 38845 17045
rect 38855 17005 38895 17045
rect 38905 17005 38945 17045
rect 38955 17005 38995 17045
rect 39005 17005 39045 17045
rect 39055 17005 39095 17045
rect 39105 17005 39145 17045
rect 39155 17005 39195 17045
rect 39205 17005 39245 17045
rect 39255 17005 39295 17045
rect 39305 17005 39345 17045
rect 39355 17005 39395 17045
rect 39405 17005 39445 17045
rect 39455 17005 39495 17045
rect 39505 17005 39545 17045
rect 39555 17005 39595 17045
rect 39605 17005 39645 17045
rect 39655 17005 39695 17045
rect 39705 17005 39745 17045
rect -3495 16940 -3455 16945
rect -3495 16910 -3490 16940
rect -3490 16910 -3460 16940
rect -3460 16910 -3455 16940
rect -3495 16905 -3455 16910
rect -3295 16940 -3255 16945
rect -3295 16910 -3290 16940
rect -3290 16910 -3260 16940
rect -3260 16910 -3255 16940
rect -3295 16905 -3255 16910
rect -3095 16940 -3055 16945
rect -3095 16910 -3090 16940
rect -3090 16910 -3060 16940
rect -3060 16910 -3055 16940
rect -3095 16905 -3055 16910
rect -1595 16940 -1555 16945
rect -1595 16910 -1590 16940
rect -1590 16910 -1560 16940
rect -1560 16910 -1555 16940
rect -1595 16905 -1555 16910
rect -1195 16940 -1155 16945
rect -1195 16910 -1190 16940
rect -1190 16910 -1160 16940
rect -1160 16910 -1155 16940
rect -1195 16905 -1155 16910
rect -1095 16940 -1055 16945
rect -1095 16910 -1090 16940
rect -1090 16910 -1060 16940
rect -1060 16910 -1055 16940
rect -1095 16905 -1055 16910
rect -995 16940 -955 16945
rect -995 16910 -990 16940
rect -990 16910 -960 16940
rect -960 16910 -955 16940
rect -995 16905 -955 16910
rect -895 16940 -855 16945
rect -895 16910 -890 16940
rect -890 16910 -860 16940
rect -860 16910 -855 16940
rect -895 16905 -855 16910
rect -795 16940 -755 16945
rect -795 16910 -790 16940
rect -790 16910 -760 16940
rect -760 16910 -755 16940
rect -795 16905 -755 16910
rect -695 16940 -655 16945
rect -695 16910 -690 16940
rect -690 16910 -660 16940
rect -660 16910 -655 16940
rect -695 16905 -655 16910
rect -595 16940 -555 16945
rect -595 16910 -590 16940
rect -590 16910 -560 16940
rect -560 16910 -555 16940
rect -595 16905 -555 16910
rect -495 16940 -455 16945
rect -495 16910 -490 16940
rect -490 16910 -460 16940
rect -460 16910 -455 16940
rect -495 16905 -455 16910
rect -395 16940 -355 16945
rect -395 16910 -390 16940
rect -390 16910 -360 16940
rect -360 16910 -355 16940
rect -395 16905 -355 16910
rect -295 16940 -255 16945
rect -295 16910 -290 16940
rect -290 16910 -260 16940
rect -260 16910 -255 16940
rect -295 16905 -255 16910
rect -195 16940 -155 16945
rect -195 16910 -190 16940
rect -190 16910 -160 16940
rect -160 16910 -155 16940
rect -195 16905 -155 16910
rect -95 16940 -55 16945
rect -95 16910 -90 16940
rect -90 16910 -60 16940
rect -60 16910 -55 16940
rect -95 16905 -55 16910
rect 5 16905 45 16945
rect 55 16905 95 16945
rect 105 16905 145 16945
rect 155 16905 195 16945
rect 205 16905 245 16945
rect 255 16905 295 16945
rect 305 16905 345 16945
rect 355 16905 395 16945
rect 405 16905 445 16945
rect 455 16905 495 16945
rect 505 16905 545 16945
rect 555 16905 595 16945
rect 605 16905 645 16945
rect 655 16905 695 16945
rect 705 16905 745 16945
rect 755 16905 795 16945
rect 805 16905 845 16945
rect 855 16905 895 16945
rect 905 16905 945 16945
rect 955 16905 995 16945
rect 1005 16905 1045 16945
rect 1055 16905 1095 16945
rect 1105 16905 1145 16945
rect 1155 16905 1195 16945
rect 1205 16905 1245 16945
rect 1255 16905 1295 16945
rect 1305 16905 1345 16945
rect 1355 16905 1395 16945
rect 1405 16905 1445 16945
rect 1455 16905 1495 16945
rect 1505 16905 1545 16945
rect 1555 16905 1595 16945
rect 1605 16905 1645 16945
rect 1655 16905 1695 16945
rect 1705 16905 1745 16945
rect 1755 16905 1795 16945
rect 1805 16905 1845 16945
rect 1855 16905 1895 16945
rect 1905 16905 1945 16945
rect 1955 16905 1995 16945
rect 2005 16905 2045 16945
rect 2055 16905 2095 16945
rect 2105 16905 2145 16945
rect 2155 16905 2195 16945
rect 2205 16905 2245 16945
rect 2255 16905 2295 16945
rect 2305 16905 2345 16945
rect 2355 16905 2395 16945
rect 2405 16905 2445 16945
rect 2455 16905 2495 16945
rect 2505 16905 2545 16945
rect 2555 16905 2595 16945
rect 2605 16905 2645 16945
rect 2655 16905 2695 16945
rect 2705 16905 2745 16945
rect 2755 16905 2795 16945
rect 2805 16905 2845 16945
rect 2855 16905 2895 16945
rect 2905 16905 2945 16945
rect 2955 16905 2995 16945
rect 3005 16905 3045 16945
rect 3055 16905 3095 16945
rect 3105 16905 3145 16945
rect 3155 16905 3195 16945
rect 3205 16905 3245 16945
rect 3255 16905 3295 16945
rect 3305 16905 3345 16945
rect 3355 16905 3395 16945
rect 3405 16905 3445 16945
rect 3455 16905 3495 16945
rect 3505 16905 3545 16945
rect 3555 16905 3595 16945
rect 3605 16905 3645 16945
rect 3655 16905 3695 16945
rect 3705 16905 3745 16945
rect 3755 16905 3795 16945
rect 3805 16905 3845 16945
rect 3855 16905 3895 16945
rect 3905 16905 3945 16945
rect 3955 16905 3995 16945
rect 4005 16905 4045 16945
rect 4055 16905 4095 16945
rect 4105 16905 4145 16945
rect 4155 16905 4195 16945
rect 4205 16905 4245 16945
rect 4255 16905 4295 16945
rect 4305 16905 4345 16945
rect 4355 16905 4395 16945
rect 4405 16905 4445 16945
rect 4455 16905 4495 16945
rect 4505 16905 4545 16945
rect 4555 16905 4595 16945
rect 4605 16905 4645 16945
rect 4655 16905 4695 16945
rect 4705 16905 4745 16945
rect 4755 16905 4795 16945
rect 4805 16905 4845 16945
rect 4855 16905 4895 16945
rect 4905 16905 4945 16945
rect 4955 16905 4995 16945
rect 5005 16905 5045 16945
rect 5055 16905 5095 16945
rect 5105 16905 5145 16945
rect 5155 16905 5195 16945
rect 5205 16905 5245 16945
rect 5255 16905 5295 16945
rect 5305 16905 5345 16945
rect 5355 16905 5395 16945
rect 5405 16905 5445 16945
rect 5455 16905 5495 16945
rect 5505 16905 5545 16945
rect 5555 16905 5595 16945
rect 5605 16905 5645 16945
rect 5655 16905 5695 16945
rect 5705 16905 5745 16945
rect 5755 16905 5795 16945
rect 5805 16905 5845 16945
rect 5855 16905 5895 16945
rect 5905 16905 5945 16945
rect 5955 16905 5995 16945
rect 6005 16905 6045 16945
rect 6055 16905 6095 16945
rect 6105 16905 6145 16945
rect 6155 16905 6195 16945
rect 6205 16905 6245 16945
rect 6255 16905 6295 16945
rect 6305 16905 6345 16945
rect 6355 16905 6395 16945
rect 6405 16905 6445 16945
rect 6455 16905 6495 16945
rect 6505 16905 6545 16945
rect 6555 16905 6595 16945
rect 6605 16905 6645 16945
rect 6655 16905 6695 16945
rect 6705 16905 6745 16945
rect 6755 16905 6795 16945
rect 6805 16905 6845 16945
rect 6855 16905 6895 16945
rect 6905 16905 6945 16945
rect 6955 16905 6995 16945
rect 7005 16905 7045 16945
rect 7055 16905 7095 16945
rect 7105 16905 7145 16945
rect 7155 16905 7195 16945
rect 7205 16905 7245 16945
rect 7255 16905 7295 16945
rect 7305 16905 7345 16945
rect 7355 16905 7395 16945
rect 7405 16905 7445 16945
rect 7455 16905 7495 16945
rect 7505 16905 7545 16945
rect 7555 16905 7595 16945
rect 7605 16905 7645 16945
rect 7655 16905 7695 16945
rect 7705 16905 7745 16945
rect 7755 16905 7795 16945
rect 7805 16905 7845 16945
rect 7855 16905 7895 16945
rect 7905 16905 7945 16945
rect 7955 16905 7995 16945
rect 8005 16905 8045 16945
rect 8055 16905 8095 16945
rect 8105 16905 8145 16945
rect 8155 16905 8195 16945
rect 8205 16905 8245 16945
rect 8255 16905 8295 16945
rect 8305 16905 8345 16945
rect 8355 16905 8395 16945
rect 8405 16905 8445 16945
rect 8455 16905 8495 16945
rect 8505 16905 8545 16945
rect 8555 16905 8595 16945
rect 8605 16905 8645 16945
rect 8655 16905 8695 16945
rect 8705 16905 8745 16945
rect 8755 16905 8795 16945
rect 8805 16905 8845 16945
rect 8855 16905 8895 16945
rect 8905 16905 8945 16945
rect 8955 16905 8995 16945
rect 9005 16905 9045 16945
rect 9055 16905 9095 16945
rect 9105 16905 9145 16945
rect 9155 16905 9195 16945
rect 9205 16905 9245 16945
rect 9255 16905 9295 16945
rect 9305 16905 9345 16945
rect 9355 16905 9395 16945
rect 9405 16905 9445 16945
rect 9455 16905 9495 16945
rect 9505 16905 9545 16945
rect 9555 16905 9595 16945
rect 9605 16905 9645 16945
rect 9655 16905 9695 16945
rect 9705 16905 9745 16945
rect 9755 16905 9795 16945
rect 9805 16905 9845 16945
rect 9855 16905 9895 16945
rect 9905 16905 9945 16945
rect 9955 16905 9995 16945
rect 10005 16905 10045 16945
rect 10055 16905 10095 16945
rect 10105 16905 10145 16945
rect 10155 16905 10195 16945
rect 10205 16905 10245 16945
rect 10255 16905 10295 16945
rect 10305 16905 10345 16945
rect 10355 16905 10395 16945
rect 10405 16905 10445 16945
rect 10455 16905 10495 16945
rect 10505 16905 10545 16945
rect 10555 16905 10595 16945
rect 10605 16905 10645 16945
rect 10655 16905 10695 16945
rect 10705 16905 10745 16945
rect 10755 16905 10795 16945
rect 10805 16905 10845 16945
rect 10855 16905 10895 16945
rect 10905 16905 10945 16945
rect 10955 16905 10995 16945
rect 11005 16905 11045 16945
rect 11055 16905 11095 16945
rect 11105 16905 11145 16945
rect 11155 16905 11195 16945
rect 11205 16905 11245 16945
rect 11255 16905 11295 16945
rect 11305 16905 11345 16945
rect 11355 16905 11395 16945
rect 11405 16905 11445 16945
rect 11455 16905 11495 16945
rect 11505 16905 11545 16945
rect 11555 16905 11595 16945
rect 11605 16905 11645 16945
rect 11655 16905 11695 16945
rect 11705 16905 11745 16945
rect 11755 16905 11795 16945
rect 11805 16905 11845 16945
rect 11855 16905 11895 16945
rect 11905 16905 11945 16945
rect 11955 16905 11995 16945
rect 12005 16905 12045 16945
rect 12055 16905 12095 16945
rect 12105 16905 12145 16945
rect 12155 16905 12195 16945
rect 12205 16905 12245 16945
rect 12255 16905 12295 16945
rect 12305 16905 12345 16945
rect 12355 16905 12395 16945
rect 12405 16905 12445 16945
rect 12455 16905 12495 16945
rect 12505 16905 12545 16945
rect 12555 16905 12595 16945
rect 12605 16905 12645 16945
rect 12655 16905 12695 16945
rect 12705 16905 12745 16945
rect 12755 16905 12795 16945
rect 12805 16905 12845 16945
rect 12855 16905 12895 16945
rect 12905 16905 12945 16945
rect 12955 16905 12995 16945
rect 13005 16905 13045 16945
rect 13055 16905 13095 16945
rect 13105 16905 13145 16945
rect 13155 16905 13195 16945
rect 13205 16905 13245 16945
rect 13255 16905 13295 16945
rect 13305 16905 13345 16945
rect 13355 16905 13395 16945
rect 13405 16905 13445 16945
rect 13455 16905 13495 16945
rect 13505 16905 13545 16945
rect 13555 16905 13595 16945
rect 13605 16905 13645 16945
rect 13655 16905 13695 16945
rect 13705 16905 13745 16945
rect 13755 16905 13795 16945
rect 13805 16905 13845 16945
rect 13855 16905 13895 16945
rect 13905 16905 13945 16945
rect 13955 16905 13995 16945
rect 14005 16905 14045 16945
rect 14055 16905 14095 16945
rect 14105 16905 14145 16945
rect 14155 16905 14195 16945
rect 14205 16905 14245 16945
rect 14255 16905 14295 16945
rect 14305 16905 14345 16945
rect 14355 16905 14395 16945
rect 14405 16905 14445 16945
rect 14455 16905 14495 16945
rect 14505 16905 14545 16945
rect 14555 16905 14595 16945
rect 14605 16905 14645 16945
rect 14655 16905 14695 16945
rect 14705 16905 14745 16945
rect 14755 16905 14795 16945
rect 14805 16905 14845 16945
rect 14855 16905 14895 16945
rect 14905 16905 14945 16945
rect 14955 16905 14995 16945
rect 15005 16905 15045 16945
rect 15055 16905 15095 16945
rect 15105 16905 15145 16945
rect 15155 16905 15195 16945
rect 15205 16905 15245 16945
rect 15255 16905 15295 16945
rect 15305 16905 15345 16945
rect 15355 16905 15395 16945
rect 15405 16905 15445 16945
rect 15455 16905 15495 16945
rect 15505 16905 15545 16945
rect 15555 16905 15595 16945
rect 15605 16905 15645 16945
rect 15655 16905 15695 16945
rect 15705 16905 15745 16945
rect 15755 16905 15795 16945
rect 15805 16905 15845 16945
rect 15855 16905 15895 16945
rect 15905 16905 15945 16945
rect 15955 16905 15995 16945
rect 16005 16905 16045 16945
rect 16055 16905 16095 16945
rect 16105 16905 16145 16945
rect 16155 16905 16195 16945
rect 16205 16905 16245 16945
rect 16255 16905 16295 16945
rect 16305 16905 16345 16945
rect 16355 16905 16395 16945
rect 16405 16905 16445 16945
rect 16455 16905 16495 16945
rect 16505 16905 16545 16945
rect 16555 16905 16595 16945
rect 16605 16905 16645 16945
rect 16655 16905 16695 16945
rect 16705 16905 16745 16945
rect 16755 16905 16795 16945
rect 16805 16905 16845 16945
rect 16855 16905 16895 16945
rect 16905 16905 16945 16945
rect 16955 16905 16995 16945
rect 17005 16905 17045 16945
rect 17055 16905 17095 16945
rect 17105 16905 17145 16945
rect 17155 16905 17195 16945
rect 17205 16905 17245 16945
rect 17255 16905 17295 16945
rect 17305 16905 17345 16945
rect 17355 16905 17395 16945
rect 17405 16905 17445 16945
rect 17455 16905 17495 16945
rect 17505 16905 17545 16945
rect 17555 16905 17595 16945
rect 17605 16905 17645 16945
rect 17655 16905 17695 16945
rect 17705 16905 17745 16945
rect 17755 16905 17795 16945
rect 17805 16905 17845 16945
rect 17855 16905 17895 16945
rect 17905 16905 17945 16945
rect 17955 16905 17995 16945
rect 18005 16905 18045 16945
rect 18055 16905 18095 16945
rect 18105 16905 18145 16945
rect 18155 16905 18195 16945
rect 18205 16905 18245 16945
rect 18255 16905 18295 16945
rect 18305 16905 18345 16945
rect 18355 16905 18395 16945
rect 18405 16905 18445 16945
rect 18455 16905 18495 16945
rect 18505 16905 18545 16945
rect 18555 16905 18595 16945
rect 18605 16905 18645 16945
rect 18655 16905 18695 16945
rect 18705 16905 18745 16945
rect 18755 16905 18795 16945
rect 18805 16905 18845 16945
rect 18855 16905 18895 16945
rect 18905 16905 18945 16945
rect 18955 16905 18995 16945
rect 19005 16905 19045 16945
rect 19055 16905 19095 16945
rect 19105 16905 19145 16945
rect 19155 16905 19195 16945
rect 19205 16905 19245 16945
rect 19255 16905 19295 16945
rect 19305 16905 19345 16945
rect 19355 16905 19395 16945
rect 19405 16905 19445 16945
rect 19455 16905 19495 16945
rect 19505 16905 19545 16945
rect 19555 16905 19595 16945
rect 19605 16905 19645 16945
rect 19655 16905 19695 16945
rect 19705 16905 19745 16945
rect 19755 16905 19795 16945
rect 19805 16905 19845 16945
rect 19855 16905 19895 16945
rect 19905 16905 19945 16945
rect 19955 16905 19995 16945
rect 20005 16905 20045 16945
rect 20055 16905 20095 16945
rect 20105 16905 20145 16945
rect 20155 16905 20195 16945
rect 20205 16905 20245 16945
rect 20255 16905 20295 16945
rect 20305 16905 20345 16945
rect 20355 16905 20395 16945
rect 20405 16905 20445 16945
rect 20455 16905 20495 16945
rect 20505 16905 20545 16945
rect 20555 16905 20595 16945
rect 20605 16905 20645 16945
rect 20655 16905 20695 16945
rect 20705 16905 20745 16945
rect 20755 16905 20795 16945
rect 20805 16905 20845 16945
rect 20855 16905 20895 16945
rect 20905 16905 20945 16945
rect 20955 16905 20995 16945
rect 21005 16905 21045 16945
rect 21055 16905 21095 16945
rect 21105 16905 21145 16945
rect 21155 16905 21195 16945
rect 21205 16905 21245 16945
rect 21255 16905 21295 16945
rect 21305 16905 21345 16945
rect 21355 16905 21395 16945
rect 21405 16905 21445 16945
rect 21455 16905 21495 16945
rect 21505 16905 21545 16945
rect 21555 16905 21595 16945
rect 21605 16905 21645 16945
rect 21655 16905 21695 16945
rect 21705 16905 21745 16945
rect 21755 16905 21795 16945
rect 21805 16905 21845 16945
rect 21855 16905 21895 16945
rect 21905 16905 21945 16945
rect 21955 16905 21995 16945
rect 22005 16905 22045 16945
rect 22055 16905 22095 16945
rect 22105 16905 22145 16945
rect 22155 16905 22195 16945
rect 22205 16905 22245 16945
rect 22255 16905 22295 16945
rect 22305 16905 22345 16945
rect 22355 16905 22395 16945
rect 22405 16905 22445 16945
rect 22455 16905 22495 16945
rect 22505 16905 22545 16945
rect 22555 16905 22595 16945
rect 22605 16905 22645 16945
rect 22655 16905 22695 16945
rect 22705 16905 22745 16945
rect 22755 16905 22795 16945
rect 22805 16905 22845 16945
rect 22855 16905 22895 16945
rect 22905 16905 22945 16945
rect 22955 16905 22995 16945
rect 23005 16905 23045 16945
rect 23055 16905 23095 16945
rect 23105 16905 23145 16945
rect 23155 16905 23195 16945
rect 23205 16905 23245 16945
rect 23255 16905 23295 16945
rect 23305 16905 23345 16945
rect 23355 16905 23395 16945
rect 23405 16905 23445 16945
rect 23455 16905 23495 16945
rect 23505 16905 23545 16945
rect 23555 16905 23595 16945
rect 23605 16905 23645 16945
rect 23655 16905 23695 16945
rect 23705 16905 23745 16945
rect 23755 16905 23795 16945
rect 23805 16905 23845 16945
rect 23855 16905 23895 16945
rect 23905 16905 23945 16945
rect 23955 16905 23995 16945
rect 24005 16905 24045 16945
rect 24055 16905 24095 16945
rect 24105 16905 24145 16945
rect 24155 16905 24195 16945
rect 24205 16905 24245 16945
rect 24255 16905 24295 16945
rect 24305 16905 24345 16945
rect 24355 16905 24395 16945
rect 24405 16905 24445 16945
rect 24455 16905 24495 16945
rect 24505 16905 24545 16945
rect 24555 16905 24595 16945
rect 24605 16905 24645 16945
rect 24655 16905 24695 16945
rect 24705 16905 24745 16945
rect 24755 16905 24795 16945
rect 24805 16905 24845 16945
rect 24855 16905 24895 16945
rect 24905 16905 24945 16945
rect 24955 16905 24995 16945
rect 25005 16905 25045 16945
rect 25055 16905 25095 16945
rect 25105 16905 25145 16945
rect 25155 16905 25195 16945
rect 25205 16905 25245 16945
rect 25255 16905 25295 16945
rect 25305 16905 25345 16945
rect 25355 16905 25395 16945
rect 25405 16905 25445 16945
rect 25455 16905 25495 16945
rect 25505 16905 25545 16945
rect 25555 16905 25595 16945
rect 25605 16905 25645 16945
rect 25655 16905 25695 16945
rect 25705 16905 25745 16945
rect 25755 16905 25795 16945
rect 25805 16905 25845 16945
rect 25855 16905 25895 16945
rect 25905 16905 25945 16945
rect 25955 16905 25995 16945
rect 26005 16905 26045 16945
rect 26055 16905 26095 16945
rect 26105 16905 26145 16945
rect 26155 16905 26195 16945
rect 26205 16905 26245 16945
rect 26255 16905 26295 16945
rect 26305 16905 26345 16945
rect 26355 16905 26395 16945
rect 26405 16905 26445 16945
rect 26455 16905 26495 16945
rect 26505 16905 26545 16945
rect 26555 16905 26595 16945
rect 26605 16905 26645 16945
rect 26655 16905 26695 16945
rect 26705 16905 26745 16945
rect 26755 16905 26795 16945
rect 26805 16905 26845 16945
rect 26855 16905 26895 16945
rect 26905 16905 26945 16945
rect 26955 16905 26995 16945
rect 27005 16905 27045 16945
rect 27055 16905 27095 16945
rect 27105 16905 27145 16945
rect 27155 16905 27195 16945
rect 27205 16905 27245 16945
rect 27255 16905 27295 16945
rect 27305 16905 27345 16945
rect 27355 16905 27395 16945
rect 27405 16905 27445 16945
rect 27455 16905 27495 16945
rect 27505 16905 27545 16945
rect 27555 16905 27595 16945
rect 27605 16905 27645 16945
rect 27655 16905 27695 16945
rect 27705 16905 27745 16945
rect 27755 16905 27795 16945
rect 27805 16905 27845 16945
rect 27855 16905 27895 16945
rect 27905 16905 27945 16945
rect 27955 16905 27995 16945
rect 28005 16905 28045 16945
rect 28055 16905 28095 16945
rect 28105 16905 28145 16945
rect 28155 16905 28195 16945
rect 28205 16905 28245 16945
rect 28255 16905 28295 16945
rect 28305 16905 28345 16945
rect 28355 16905 28395 16945
rect 28405 16905 28445 16945
rect 28455 16905 28495 16945
rect 28505 16905 28545 16945
rect 28555 16905 28595 16945
rect 28605 16905 28645 16945
rect 28655 16905 28695 16945
rect 28705 16905 28745 16945
rect 28755 16905 28795 16945
rect 28805 16905 28845 16945
rect 28855 16905 28895 16945
rect 28905 16905 28945 16945
rect 28955 16905 28995 16945
rect 29005 16905 29045 16945
rect 29055 16905 29095 16945
rect 29105 16905 29145 16945
rect 29155 16905 29195 16945
rect 29205 16905 29245 16945
rect 29255 16905 29295 16945
rect 29305 16905 29345 16945
rect 29355 16905 29395 16945
rect 29405 16905 29445 16945
rect 29455 16905 29495 16945
rect 29505 16905 29545 16945
rect 29555 16905 29595 16945
rect 29605 16905 29645 16945
rect 29655 16905 29695 16945
rect 29705 16905 29745 16945
rect 29755 16905 29795 16945
rect 29805 16905 29845 16945
rect 29855 16905 29895 16945
rect 29905 16905 29945 16945
rect 29955 16905 29995 16945
rect 30005 16905 30045 16945
rect 30055 16905 30095 16945
rect 30105 16905 30145 16945
rect 30155 16905 30195 16945
rect 30205 16905 30245 16945
rect 30255 16905 30295 16945
rect 30305 16905 30345 16945
rect 30355 16905 30395 16945
rect 30405 16905 30445 16945
rect 30455 16905 30495 16945
rect 30505 16905 30545 16945
rect 30555 16905 30595 16945
rect 30605 16905 30645 16945
rect 30655 16905 30695 16945
rect 30705 16905 30745 16945
rect 30755 16905 30795 16945
rect 30805 16905 30845 16945
rect 30855 16905 30895 16945
rect 30905 16905 30945 16945
rect 30955 16905 30995 16945
rect 31005 16905 31045 16945
rect 31055 16905 31095 16945
rect 31105 16905 31145 16945
rect 31155 16905 31195 16945
rect 31205 16905 31245 16945
rect 31255 16905 31295 16945
rect 31305 16905 31345 16945
rect 31355 16905 31395 16945
rect 31405 16905 31445 16945
rect 31455 16905 31495 16945
rect 31505 16905 31545 16945
rect 31555 16905 31595 16945
rect 31605 16905 31645 16945
rect 31655 16905 31695 16945
rect 31705 16905 31745 16945
rect 31755 16905 31795 16945
rect 31805 16905 31845 16945
rect 31855 16905 31895 16945
rect 31905 16905 31945 16945
rect 31955 16905 31995 16945
rect 32005 16905 32045 16945
rect 32055 16905 32095 16945
rect 32105 16905 32145 16945
rect 32155 16905 32195 16945
rect 32205 16905 32245 16945
rect 32255 16905 32295 16945
rect 32305 16905 32345 16945
rect 32355 16905 32395 16945
rect 32405 16905 32445 16945
rect 32455 16905 32495 16945
rect 32505 16905 32545 16945
rect 32555 16905 32595 16945
rect 32605 16905 32645 16945
rect 32655 16905 32695 16945
rect 32705 16905 32745 16945
rect 32755 16905 32795 16945
rect 32805 16905 32845 16945
rect 32855 16905 32895 16945
rect 32905 16905 32945 16945
rect 32955 16905 32995 16945
rect 33005 16905 33045 16945
rect 33055 16905 33095 16945
rect 33105 16905 33145 16945
rect 33155 16905 33195 16945
rect 33205 16905 33245 16945
rect 33255 16905 33295 16945
rect 33305 16905 33345 16945
rect 33355 16905 33395 16945
rect 33405 16905 33445 16945
rect 33455 16905 33495 16945
rect 33505 16905 33545 16945
rect 33555 16905 33595 16945
rect 33605 16905 33645 16945
rect 33655 16905 33695 16945
rect 33705 16905 33745 16945
rect 33755 16905 33795 16945
rect 33805 16905 33845 16945
rect 33855 16905 33895 16945
rect 33905 16905 33945 16945
rect 33955 16905 33995 16945
rect 34005 16905 34045 16945
rect 34055 16905 34095 16945
rect 34105 16905 34145 16945
rect 34155 16905 34195 16945
rect 34205 16905 34245 16945
rect 34255 16905 34295 16945
rect 34305 16905 34345 16945
rect 34355 16905 34395 16945
rect 34405 16905 34445 16945
rect 34455 16905 34495 16945
rect 34505 16905 34545 16945
rect 34555 16905 34595 16945
rect 34605 16905 34645 16945
rect 34655 16905 34695 16945
rect 34705 16905 34745 16945
rect 34755 16905 34795 16945
rect 34805 16905 34845 16945
rect 34855 16905 34895 16945
rect 34905 16905 34945 16945
rect 34955 16905 34995 16945
rect 35005 16905 35045 16945
rect 35055 16905 35095 16945
rect 35105 16905 35145 16945
rect 35155 16905 35195 16945
rect 35205 16905 35245 16945
rect 35255 16905 35295 16945
rect 35305 16905 35345 16945
rect 35355 16905 35395 16945
rect 35405 16905 35445 16945
rect 35455 16905 35495 16945
rect 35505 16905 35545 16945
rect 35555 16905 35595 16945
rect 35605 16905 35645 16945
rect 35655 16905 35695 16945
rect 35705 16905 35745 16945
rect 35755 16905 35795 16945
rect 35805 16905 35845 16945
rect 35855 16905 35895 16945
rect 35905 16905 35945 16945
rect 35955 16905 35995 16945
rect 36005 16905 36045 16945
rect 36055 16905 36095 16945
rect 36105 16905 36145 16945
rect 36155 16905 36195 16945
rect 36205 16905 36245 16945
rect 36255 16905 36295 16945
rect 36305 16905 36345 16945
rect 36355 16905 36395 16945
rect 36405 16905 36445 16945
rect 36455 16905 36495 16945
rect 36505 16905 36545 16945
rect 36555 16905 36595 16945
rect 36605 16905 36645 16945
rect 36655 16905 36695 16945
rect 36705 16905 36745 16945
rect 36755 16905 36795 16945
rect 36805 16905 36845 16945
rect 36855 16905 36895 16945
rect 36905 16905 36945 16945
rect 36955 16905 36995 16945
rect 37005 16905 37045 16945
rect 37055 16905 37095 16945
rect 37105 16905 37145 16945
rect 37155 16905 37195 16945
rect 37205 16905 37245 16945
rect 37255 16905 37295 16945
rect 37305 16905 37345 16945
rect 37355 16905 37395 16945
rect 37405 16905 37445 16945
rect 37455 16905 37495 16945
rect 37505 16905 37545 16945
rect 37555 16905 37595 16945
rect 37605 16905 37645 16945
rect 37655 16905 37695 16945
rect 37705 16905 37745 16945
rect 37755 16905 37795 16945
rect 37805 16905 37845 16945
rect 37855 16905 37895 16945
rect 37905 16905 37945 16945
rect 37955 16905 37995 16945
rect 38005 16905 38045 16945
rect 38055 16905 38095 16945
rect 38105 16905 38145 16945
rect 38155 16905 38195 16945
rect 38205 16905 38245 16945
rect 38255 16905 38295 16945
rect 38305 16905 38345 16945
rect 38355 16905 38395 16945
rect 38405 16905 38445 16945
rect 38455 16905 38495 16945
rect 38505 16905 38545 16945
rect 38555 16905 38595 16945
rect 38605 16905 38645 16945
rect 38655 16905 38695 16945
rect 38705 16905 38745 16945
rect 38755 16905 38795 16945
rect 38805 16905 38845 16945
rect 38855 16905 38895 16945
rect 38905 16905 38945 16945
rect 38955 16905 38995 16945
rect 39005 16905 39045 16945
rect 39055 16905 39095 16945
rect 39105 16905 39145 16945
rect 39155 16905 39195 16945
rect 39205 16905 39245 16945
rect 39255 16905 39295 16945
rect 39305 16905 39345 16945
rect 39355 16905 39395 16945
rect 39405 16905 39445 16945
rect 39455 16905 39495 16945
rect 39505 16905 39545 16945
rect 39555 16905 39595 16945
rect 39605 16905 39645 16945
rect 39655 16905 39695 16945
rect 39705 16905 39745 16945
rect 39905 16905 39945 16945
rect 39955 16905 39995 16945
rect 40005 16905 40045 16945
rect 40055 16905 40095 16945
rect 40105 16905 40145 16945
rect 40155 16905 40195 16945
rect 40205 16905 40245 16945
rect 40255 16905 40295 16945
rect 40305 16905 40345 16945
rect 40355 16905 40395 16945
rect 40405 16905 40445 16945
rect 40455 16905 40495 16945
rect 40505 16905 40545 16945
rect 40555 16905 40595 16945
rect 40605 16905 40645 16945
rect 40655 16905 40695 16945
rect 40705 16905 40745 16945
rect 40755 16905 40795 16945
rect 40805 16905 40845 16945
rect 40855 16905 40895 16945
rect -395 16805 -355 16845
rect 105 16805 145 16845
rect 155 16805 195 16845
rect 205 16805 245 16845
rect 255 16805 295 16845
rect 305 16805 345 16845
rect 355 16805 395 16845
rect 405 16805 445 16845
rect 455 16805 495 16845
rect 505 16805 545 16845
rect 555 16805 595 16845
rect 605 16805 645 16845
rect 655 16805 695 16845
rect 705 16805 745 16845
rect 755 16805 795 16845
rect 805 16805 845 16845
rect 855 16805 895 16845
rect 905 16805 945 16845
rect 955 16805 995 16845
rect 1005 16805 1045 16845
rect 1055 16805 1095 16845
rect 1105 16805 1145 16845
rect 1155 16805 1195 16845
rect 1205 16805 1245 16845
rect 1255 16805 1295 16845
rect 1305 16805 1345 16845
rect 1355 16805 1395 16845
rect 1405 16805 1445 16845
rect 1455 16805 1495 16845
rect 1505 16805 1545 16845
rect 1555 16805 1595 16845
rect 1605 16805 1645 16845
rect 1655 16805 1695 16845
rect 1705 16805 1745 16845
rect 1755 16805 1795 16845
rect 1805 16805 1845 16845
rect 1855 16805 1895 16845
rect 1905 16805 1945 16845
rect 1955 16805 1995 16845
rect 2005 16805 2045 16845
rect 2055 16805 2095 16845
rect 2105 16805 2145 16845
rect 2155 16805 2195 16845
rect 2205 16805 2245 16845
rect 2255 16805 2295 16845
rect 2305 16805 2345 16845
rect 2355 16805 2395 16845
rect 2405 16805 2445 16845
rect 2455 16805 2495 16845
rect 2505 16805 2545 16845
rect 2555 16805 2595 16845
rect 2605 16805 2645 16845
rect 2655 16805 2695 16845
rect 2705 16805 2745 16845
rect 2755 16805 2795 16845
rect 2805 16805 2845 16845
rect 2855 16805 2895 16845
rect 2905 16805 2945 16845
rect 2955 16805 2995 16845
rect 3005 16805 3045 16845
rect 3055 16805 3095 16845
rect 3105 16805 3145 16845
rect 3155 16805 3195 16845
rect 3205 16805 3245 16845
rect 3255 16805 3295 16845
rect 3305 16805 3345 16845
rect 3355 16805 3395 16845
rect 3405 16805 3445 16845
rect 3455 16805 3495 16845
rect 3505 16805 3545 16845
rect 3555 16805 3595 16845
rect 3605 16805 3645 16845
rect 3655 16805 3695 16845
rect 3705 16805 3745 16845
rect 3755 16805 3795 16845
rect 3805 16805 3845 16845
rect 3855 16805 3895 16845
rect 3905 16805 3945 16845
rect 3955 16805 3995 16845
rect 4005 16805 4045 16845
rect 4055 16805 4095 16845
rect 4105 16805 4145 16845
rect 4155 16805 4195 16845
rect 4205 16805 4245 16845
rect 4255 16805 4295 16845
rect 4305 16805 4345 16845
rect 4355 16805 4395 16845
rect 4405 16805 4445 16845
rect 4455 16805 4495 16845
rect 4505 16805 4545 16845
rect 4555 16805 4595 16845
rect 4605 16805 4645 16845
rect 4655 16805 4695 16845
rect 4705 16805 4745 16845
rect 4755 16805 4795 16845
rect 4805 16805 4845 16845
rect 4855 16805 4895 16845
rect 4905 16805 4945 16845
rect 4955 16805 4995 16845
rect 5005 16805 5045 16845
rect 5055 16805 5095 16845
rect 5105 16805 5145 16845
rect 5155 16805 5195 16845
rect 5205 16805 5245 16845
rect 5255 16805 5295 16845
rect 5305 16805 5345 16845
rect 5355 16805 5395 16845
rect 5405 16805 5445 16845
rect 5455 16805 5495 16845
rect 5505 16805 5545 16845
rect 5555 16805 5595 16845
rect 5605 16805 5645 16845
rect 5655 16805 5695 16845
rect 5705 16805 5745 16845
rect 5755 16805 5795 16845
rect 5805 16805 5845 16845
rect 5855 16805 5895 16845
rect 5905 16805 5945 16845
rect 5955 16805 5995 16845
rect 6005 16805 6045 16845
rect 6055 16805 6095 16845
rect 6105 16805 6145 16845
rect 6155 16805 6195 16845
rect 6205 16805 6245 16845
rect 6255 16805 6295 16845
rect 6305 16805 6345 16845
rect 6355 16805 6395 16845
rect 6405 16805 6445 16845
rect 6455 16805 6495 16845
rect 6505 16805 6545 16845
rect 6555 16805 6595 16845
rect 6605 16805 6645 16845
rect 6655 16805 6695 16845
rect 6705 16805 6745 16845
rect 6755 16805 6795 16845
rect 6805 16805 6845 16845
rect 6855 16805 6895 16845
rect 6905 16805 6945 16845
rect 6955 16805 6995 16845
rect 7005 16805 7045 16845
rect 7055 16805 7095 16845
rect 7105 16805 7145 16845
rect 7155 16805 7195 16845
rect 7205 16805 7245 16845
rect 7255 16805 7295 16845
rect 7305 16805 7345 16845
rect 7355 16805 7395 16845
rect 7405 16805 7445 16845
rect 7455 16805 7495 16845
rect 7505 16805 7545 16845
rect 7555 16805 7595 16845
rect 7605 16805 7645 16845
rect 7655 16805 7695 16845
rect 7705 16805 7745 16845
rect 7755 16805 7795 16845
rect 7805 16805 7845 16845
rect 7855 16805 7895 16845
rect 7905 16805 7945 16845
rect 7955 16805 7995 16845
rect 8005 16805 8045 16845
rect 8055 16805 8095 16845
rect 8105 16805 8145 16845
rect 8155 16805 8195 16845
rect 8205 16805 8245 16845
rect 8255 16805 8295 16845
rect 8305 16805 8345 16845
rect 8355 16805 8395 16845
rect 8405 16805 8445 16845
rect 8455 16805 8495 16845
rect 8505 16805 8545 16845
rect 8555 16805 8595 16845
rect 8605 16805 8645 16845
rect 8655 16805 8695 16845
rect 8705 16805 8745 16845
rect 8755 16805 8795 16845
rect 8805 16805 8845 16845
rect 8855 16805 8895 16845
rect 8905 16805 8945 16845
rect 8955 16805 8995 16845
rect 9005 16805 9045 16845
rect 9055 16805 9095 16845
rect 9105 16805 9145 16845
rect 9155 16805 9195 16845
rect 9205 16805 9245 16845
rect 9255 16805 9295 16845
rect 9305 16805 9345 16845
rect 9355 16805 9395 16845
rect 9405 16805 9445 16845
rect 9455 16805 9495 16845
rect 9505 16805 9545 16845
rect 9555 16805 9595 16845
rect 9605 16805 9645 16845
rect 9655 16805 9695 16845
rect 9705 16805 9745 16845
rect 9755 16805 9795 16845
rect 9805 16805 9845 16845
rect 9855 16805 9895 16845
rect 9905 16805 9945 16845
rect 9955 16805 9995 16845
rect 10005 16805 10045 16845
rect 10055 16805 10095 16845
rect 10105 16805 10145 16845
rect 10155 16805 10195 16845
rect 10205 16805 10245 16845
rect 10255 16805 10295 16845
rect 10305 16805 10345 16845
rect 10355 16805 10395 16845
rect 10405 16805 10445 16845
rect 10455 16805 10495 16845
rect 10505 16805 10545 16845
rect 10555 16805 10595 16845
rect 10605 16805 10645 16845
rect 10655 16805 10695 16845
rect 10705 16805 10745 16845
rect 10755 16805 10795 16845
rect 10805 16805 10845 16845
rect 10855 16805 10895 16845
rect 10905 16805 10945 16845
rect 10955 16805 10995 16845
rect 11005 16805 11045 16845
rect 11055 16805 11095 16845
rect 11105 16805 11145 16845
rect 11155 16805 11195 16845
rect 11205 16805 11245 16845
rect 11255 16805 11295 16845
rect 11305 16805 11345 16845
rect 11355 16805 11395 16845
rect 11405 16805 11445 16845
rect 11455 16805 11495 16845
rect 11505 16805 11545 16845
rect 11555 16805 11595 16845
rect 11605 16805 11645 16845
rect 11655 16805 11695 16845
rect 11705 16805 11745 16845
rect 11755 16805 11795 16845
rect 11805 16805 11845 16845
rect 11855 16805 11895 16845
rect 11905 16805 11945 16845
rect 11955 16805 11995 16845
rect 12005 16805 12045 16845
rect 12055 16805 12095 16845
rect 12105 16805 12145 16845
rect 12155 16805 12195 16845
rect 12205 16805 12245 16845
rect 12255 16805 12295 16845
rect 12305 16805 12345 16845
rect 12355 16805 12395 16845
rect 12405 16805 12445 16845
rect 12455 16805 12495 16845
rect 12505 16805 12545 16845
rect 12555 16805 12595 16845
rect 12605 16805 12645 16845
rect 12655 16805 12695 16845
rect 12705 16805 12745 16845
rect 12755 16805 12795 16845
rect 12805 16805 12845 16845
rect 12855 16805 12895 16845
rect 12905 16805 12945 16845
rect 12955 16805 12995 16845
rect 13005 16805 13045 16845
rect 13055 16805 13095 16845
rect 13105 16805 13145 16845
rect 13155 16805 13195 16845
rect 13205 16805 13245 16845
rect 13255 16805 13295 16845
rect 13305 16805 13345 16845
rect 13355 16805 13395 16845
rect 13405 16805 13445 16845
rect 13455 16805 13495 16845
rect 13505 16805 13545 16845
rect 13555 16805 13595 16845
rect 13605 16805 13645 16845
rect 13655 16805 13695 16845
rect 13705 16805 13745 16845
rect 13755 16805 13795 16845
rect 13805 16805 13845 16845
rect 13855 16805 13895 16845
rect 13905 16805 13945 16845
rect 13955 16805 13995 16845
rect 14005 16805 14045 16845
rect 14055 16805 14095 16845
rect 14105 16805 14145 16845
rect 14155 16805 14195 16845
rect 14205 16805 14245 16845
rect 14255 16805 14295 16845
rect 14305 16805 14345 16845
rect 14355 16805 14395 16845
rect 14405 16805 14445 16845
rect 14455 16805 14495 16845
rect 14505 16805 14545 16845
rect 14555 16805 14595 16845
rect 14605 16805 14645 16845
rect 14655 16805 14695 16845
rect 14705 16805 14745 16845
rect 14755 16805 14795 16845
rect 14805 16805 14845 16845
rect 14855 16805 14895 16845
rect 14905 16805 14945 16845
rect 14955 16805 14995 16845
rect 15005 16805 15045 16845
rect 15055 16805 15095 16845
rect 15105 16805 15145 16845
rect 15155 16805 15195 16845
rect 15205 16805 15245 16845
rect 15255 16805 15295 16845
rect 15305 16805 15345 16845
rect 15355 16805 15395 16845
rect 15405 16805 15445 16845
rect 15455 16805 15495 16845
rect 15505 16805 15545 16845
rect 15555 16805 15595 16845
rect 15605 16805 15645 16845
rect 15655 16805 15695 16845
rect 15705 16805 15745 16845
rect 15755 16805 15795 16845
rect 15805 16805 15845 16845
rect 15855 16805 15895 16845
rect 15905 16805 15945 16845
rect 15955 16805 15995 16845
rect 16005 16805 16045 16845
rect 16055 16805 16095 16845
rect 16105 16805 16145 16845
rect 16155 16805 16195 16845
rect 16205 16805 16245 16845
rect 16255 16805 16295 16845
rect 16305 16805 16345 16845
rect 16355 16805 16395 16845
rect 16405 16805 16445 16845
rect 16455 16805 16495 16845
rect 16505 16805 16545 16845
rect 16555 16805 16595 16845
rect 16605 16805 16645 16845
rect 16655 16805 16695 16845
rect 16705 16805 16745 16845
rect 16755 16805 16795 16845
rect 16805 16805 16845 16845
rect 16855 16805 16895 16845
rect 16905 16805 16945 16845
rect 16955 16805 16995 16845
rect 17005 16805 17045 16845
rect 17055 16805 17095 16845
rect 17105 16805 17145 16845
rect 17155 16805 17195 16845
rect 17205 16805 17245 16845
rect 17255 16805 17295 16845
rect 17305 16805 17345 16845
rect 17355 16805 17395 16845
rect 17405 16805 17445 16845
rect 17455 16805 17495 16845
rect 17505 16805 17545 16845
rect 17555 16805 17595 16845
rect 17605 16805 17645 16845
rect 17655 16805 17695 16845
rect 17705 16805 17745 16845
rect 17755 16805 17795 16845
rect 17805 16805 17845 16845
rect 17855 16805 17895 16845
rect 17905 16805 17945 16845
rect 17955 16805 17995 16845
rect 18005 16805 18045 16845
rect 18055 16805 18095 16845
rect 18105 16805 18145 16845
rect 18155 16805 18195 16845
rect 18205 16805 18245 16845
rect 18255 16805 18295 16845
rect 18305 16805 18345 16845
rect 18355 16805 18395 16845
rect 18405 16805 18445 16845
rect 18455 16805 18495 16845
rect 18505 16805 18545 16845
rect 18555 16805 18595 16845
rect 18605 16805 18645 16845
rect 18655 16805 18695 16845
rect 18705 16805 18745 16845
rect 18755 16805 18795 16845
rect 18805 16805 18845 16845
rect 18855 16805 18895 16845
rect 18905 16805 18945 16845
rect 18955 16805 18995 16845
rect 19005 16805 19045 16845
rect 19055 16805 19095 16845
rect 19105 16805 19145 16845
rect 19155 16805 19195 16845
rect 19205 16805 19245 16845
rect 19255 16805 19295 16845
rect 19305 16805 19345 16845
rect 19355 16805 19395 16845
rect 19405 16805 19445 16845
rect 19455 16805 19495 16845
rect 19505 16805 19545 16845
rect 19555 16805 19595 16845
rect 19605 16805 19645 16845
rect 19655 16805 19695 16845
rect 19705 16805 19745 16845
rect 19755 16805 19795 16845
rect 19805 16805 19845 16845
rect 19855 16805 19895 16845
rect 19905 16805 19945 16845
rect 19955 16805 19995 16845
rect 20005 16805 20045 16845
rect 20055 16805 20095 16845
rect 20105 16805 20145 16845
rect 20155 16805 20195 16845
rect 20205 16805 20245 16845
rect 20255 16805 20295 16845
rect 20305 16805 20345 16845
rect 20355 16805 20395 16845
rect 20405 16805 20445 16845
rect 20455 16805 20495 16845
rect 20505 16805 20545 16845
rect 20555 16805 20595 16845
rect 20605 16805 20645 16845
rect 20655 16805 20695 16845
rect 20705 16805 20745 16845
rect 20755 16805 20795 16845
rect 20805 16805 20845 16845
rect 20855 16805 20895 16845
rect 20905 16805 20945 16845
rect 20955 16805 20995 16845
rect 21005 16805 21045 16845
rect 21055 16805 21095 16845
rect 21105 16805 21145 16845
rect 21155 16805 21195 16845
rect 21205 16805 21245 16845
rect 21255 16805 21295 16845
rect 21305 16805 21345 16845
rect 21355 16805 21395 16845
rect 21405 16805 21445 16845
rect 21455 16805 21495 16845
rect 21505 16805 21545 16845
rect 21555 16805 21595 16845
rect 21605 16805 21645 16845
rect 21655 16805 21695 16845
rect 21705 16805 21745 16845
rect 21755 16805 21795 16845
rect 21805 16805 21845 16845
rect 21855 16805 21895 16845
rect 21905 16805 21945 16845
rect 21955 16805 21995 16845
rect 22005 16805 22045 16845
rect 22055 16805 22095 16845
rect 22105 16805 22145 16845
rect 22155 16805 22195 16845
rect 22205 16805 22245 16845
rect 22255 16805 22295 16845
rect 22305 16805 22345 16845
rect 22355 16805 22395 16845
rect 22405 16805 22445 16845
rect 22455 16805 22495 16845
rect 22505 16805 22545 16845
rect 22555 16805 22595 16845
rect 22605 16805 22645 16845
rect 22655 16805 22695 16845
rect 22705 16805 22745 16845
rect 22755 16805 22795 16845
rect 22805 16805 22845 16845
rect 22855 16805 22895 16845
rect 22905 16805 22945 16845
rect 22955 16805 22995 16845
rect 23005 16805 23045 16845
rect 23055 16805 23095 16845
rect 23105 16805 23145 16845
rect 23155 16805 23195 16845
rect 23205 16805 23245 16845
rect 23255 16805 23295 16845
rect 23305 16805 23345 16845
rect 23355 16805 23395 16845
rect 23405 16805 23445 16845
rect 23455 16805 23495 16845
rect 23505 16805 23545 16845
rect 23555 16805 23595 16845
rect 23605 16805 23645 16845
rect 23655 16805 23695 16845
rect 23705 16805 23745 16845
rect 23755 16805 23795 16845
rect 23805 16805 23845 16845
rect 23855 16805 23895 16845
rect 23905 16805 23945 16845
rect 23955 16805 23995 16845
rect 24005 16805 24045 16845
rect 24055 16805 24095 16845
rect 24105 16805 24145 16845
rect 24155 16805 24195 16845
rect 24205 16805 24245 16845
rect 24255 16805 24295 16845
rect 24305 16805 24345 16845
rect 24355 16805 24395 16845
rect 24405 16805 24445 16845
rect 24455 16805 24495 16845
rect 24505 16805 24545 16845
rect 24555 16805 24595 16845
rect 24605 16805 24645 16845
rect 24655 16805 24695 16845
rect 24705 16805 24745 16845
rect 24755 16805 24795 16845
rect 24805 16805 24845 16845
rect 24855 16805 24895 16845
rect 24905 16805 24945 16845
rect 24955 16805 24995 16845
rect 25005 16805 25045 16845
rect 25055 16805 25095 16845
rect 25105 16805 25145 16845
rect 25155 16805 25195 16845
rect 25205 16805 25245 16845
rect 25255 16805 25295 16845
rect 25305 16805 25345 16845
rect 25355 16805 25395 16845
rect 25405 16805 25445 16845
rect 25455 16805 25495 16845
rect 25505 16805 25545 16845
rect 25555 16805 25595 16845
rect 25605 16805 25645 16845
rect 25655 16805 25695 16845
rect 25705 16805 25745 16845
rect 25755 16805 25795 16845
rect 25805 16805 25845 16845
rect 25855 16805 25895 16845
rect 25905 16805 25945 16845
rect 25955 16805 25995 16845
rect 26005 16805 26045 16845
rect 26055 16805 26095 16845
rect 26105 16805 26145 16845
rect 26155 16805 26195 16845
rect 26205 16805 26245 16845
rect 26255 16805 26295 16845
rect 26305 16805 26345 16845
rect 26355 16805 26395 16845
rect 26405 16805 26445 16845
rect 26455 16805 26495 16845
rect 26505 16805 26545 16845
rect 26555 16805 26595 16845
rect 26605 16805 26645 16845
rect 26655 16805 26695 16845
rect 26705 16805 26745 16845
rect 26755 16805 26795 16845
rect 26805 16805 26845 16845
rect 26855 16805 26895 16845
rect 26905 16805 26945 16845
rect 26955 16805 26995 16845
rect 27005 16805 27045 16845
rect 27055 16805 27095 16845
rect 27105 16805 27145 16845
rect 27155 16805 27195 16845
rect 27205 16805 27245 16845
rect 27255 16805 27295 16845
rect 27305 16805 27345 16845
rect 27355 16805 27395 16845
rect 27405 16805 27445 16845
rect 27455 16805 27495 16845
rect 27505 16805 27545 16845
rect 27555 16805 27595 16845
rect 27605 16805 27645 16845
rect 27655 16805 27695 16845
rect 27705 16805 27745 16845
rect 27755 16805 27795 16845
rect 27805 16805 27845 16845
rect 27855 16805 27895 16845
rect 27905 16805 27945 16845
rect 27955 16805 27995 16845
rect 28005 16805 28045 16845
rect 28055 16805 28095 16845
rect 28105 16805 28145 16845
rect 28155 16805 28195 16845
rect 28205 16805 28245 16845
rect 28255 16805 28295 16845
rect 28305 16805 28345 16845
rect 28355 16805 28395 16845
rect 28405 16805 28445 16845
rect 28455 16805 28495 16845
rect 28505 16805 28545 16845
rect 28555 16805 28595 16845
rect 28605 16805 28645 16845
rect 28655 16805 28695 16845
rect 28705 16805 28745 16845
rect 28755 16805 28795 16845
rect 28805 16805 28845 16845
rect 28855 16805 28895 16845
rect 28905 16805 28945 16845
rect 28955 16805 28995 16845
rect 29005 16805 29045 16845
rect 29055 16805 29095 16845
rect 29105 16805 29145 16845
rect 29155 16805 29195 16845
rect 29205 16805 29245 16845
rect 29255 16805 29295 16845
rect 29305 16805 29345 16845
rect 29355 16805 29395 16845
rect 29405 16805 29445 16845
rect 29455 16805 29495 16845
rect 29505 16805 29545 16845
rect 29555 16805 29595 16845
rect 29605 16805 29645 16845
rect 29655 16805 29695 16845
rect 29705 16805 29745 16845
rect 29755 16805 29795 16845
rect 29805 16805 29845 16845
rect 29855 16805 29895 16845
rect 29905 16805 29945 16845
rect 29955 16805 29995 16845
rect 30005 16805 30045 16845
rect 30055 16805 30095 16845
rect 30105 16805 30145 16845
rect 30155 16805 30195 16845
rect 30205 16805 30245 16845
rect 30255 16805 30295 16845
rect 30305 16805 30345 16845
rect 30355 16805 30395 16845
rect 30405 16805 30445 16845
rect 30455 16805 30495 16845
rect 30505 16805 30545 16845
rect 30555 16805 30595 16845
rect 30605 16805 30645 16845
rect 30655 16805 30695 16845
rect 30705 16805 30745 16845
rect 30755 16805 30795 16845
rect 30805 16805 30845 16845
rect 30855 16805 30895 16845
rect 30905 16805 30945 16845
rect 30955 16805 30995 16845
rect 31005 16805 31045 16845
rect 31055 16805 31095 16845
rect 31105 16805 31145 16845
rect 31155 16805 31195 16845
rect 31205 16805 31245 16845
rect 31255 16805 31295 16845
rect 31305 16805 31345 16845
rect 31355 16805 31395 16845
rect 31405 16805 31445 16845
rect 31455 16805 31495 16845
rect 31505 16805 31545 16845
rect 31555 16805 31595 16845
rect 31605 16805 31645 16845
rect 31655 16805 31695 16845
rect 31705 16805 31745 16845
rect 31755 16805 31795 16845
rect 31805 16805 31845 16845
rect 31855 16805 31895 16845
rect 31905 16805 31945 16845
rect 31955 16805 31995 16845
rect 32005 16805 32045 16845
rect 32055 16805 32095 16845
rect 32105 16805 32145 16845
rect 32155 16805 32195 16845
rect 32205 16805 32245 16845
rect 32255 16805 32295 16845
rect 32305 16805 32345 16845
rect 32355 16805 32395 16845
rect 32405 16805 32445 16845
rect 32455 16805 32495 16845
rect 32505 16805 32545 16845
rect 32555 16805 32595 16845
rect 32605 16805 32645 16845
rect 32655 16805 32695 16845
rect 32705 16805 32745 16845
rect 32755 16805 32795 16845
rect 32805 16805 32845 16845
rect 32855 16805 32895 16845
rect 32905 16805 32945 16845
rect 32955 16805 32995 16845
rect 33005 16805 33045 16845
rect 33055 16805 33095 16845
rect 33105 16805 33145 16845
rect 33155 16805 33195 16845
rect 33205 16805 33245 16845
rect 33255 16805 33295 16845
rect 33305 16805 33345 16845
rect 33355 16805 33395 16845
rect 33405 16805 33445 16845
rect 33455 16805 33495 16845
rect 33505 16805 33545 16845
rect 33555 16805 33595 16845
rect 33605 16805 33645 16845
rect 33655 16805 33695 16845
rect 33705 16805 33745 16845
rect 33755 16805 33795 16845
rect 33805 16805 33845 16845
rect 33855 16805 33895 16845
rect 33905 16805 33945 16845
rect 33955 16805 33995 16845
rect 34005 16805 34045 16845
rect 34055 16805 34095 16845
rect 34105 16805 34145 16845
rect 34155 16805 34195 16845
rect 34205 16805 34245 16845
rect 34255 16805 34295 16845
rect 34305 16805 34345 16845
rect 34355 16805 34395 16845
rect 34405 16805 34445 16845
rect 34455 16805 34495 16845
rect 34505 16805 34545 16845
rect 34555 16805 34595 16845
rect 34605 16805 34645 16845
rect 34655 16805 34695 16845
rect 34705 16805 34745 16845
rect 34755 16805 34795 16845
rect 34805 16805 34845 16845
rect 34855 16805 34895 16845
rect 34905 16805 34945 16845
rect 34955 16805 34995 16845
rect 35005 16805 35045 16845
rect 35055 16805 35095 16845
rect 35105 16805 35145 16845
rect 35155 16805 35195 16845
rect 35205 16805 35245 16845
rect 35255 16805 35295 16845
rect 35305 16805 35345 16845
rect 35355 16805 35395 16845
rect 35405 16805 35445 16845
rect 35455 16805 35495 16845
rect 35505 16805 35545 16845
rect 35555 16805 35595 16845
rect 35605 16805 35645 16845
rect 35655 16805 35695 16845
rect 35705 16805 35745 16845
rect 35755 16805 35795 16845
rect 35805 16805 35845 16845
rect 35855 16805 35895 16845
rect 35905 16805 35945 16845
rect 35955 16805 35995 16845
rect 36005 16805 36045 16845
rect 36055 16805 36095 16845
rect 36105 16805 36145 16845
rect 36155 16805 36195 16845
rect 36205 16805 36245 16845
rect 36255 16805 36295 16845
rect 36305 16805 36345 16845
rect 36355 16805 36395 16845
rect 36405 16805 36445 16845
rect 36455 16805 36495 16845
rect 36505 16805 36545 16845
rect 36555 16805 36595 16845
rect 36605 16805 36645 16845
rect 36655 16805 36695 16845
rect 36705 16805 36745 16845
rect 36755 16805 36795 16845
rect 36805 16805 36845 16845
rect 36855 16805 36895 16845
rect 36905 16805 36945 16845
rect 36955 16805 36995 16845
rect 37005 16805 37045 16845
rect 37055 16805 37095 16845
rect 37105 16805 37145 16845
rect 37155 16805 37195 16845
rect 37205 16805 37245 16845
rect 37255 16805 37295 16845
rect 37305 16805 37345 16845
rect 37355 16805 37395 16845
rect 37405 16805 37445 16845
rect 37455 16805 37495 16845
rect 37505 16805 37545 16845
rect 37555 16805 37595 16845
rect 37605 16805 37645 16845
rect 37655 16805 37695 16845
rect 37705 16805 37745 16845
rect 37755 16805 37795 16845
rect 37805 16805 37845 16845
rect 37855 16805 37895 16845
rect 37905 16805 37945 16845
rect 37955 16805 37995 16845
rect 38005 16805 38045 16845
rect 38055 16805 38095 16845
rect 38105 16805 38145 16845
rect 38155 16805 38195 16845
rect 38205 16805 38245 16845
rect 38255 16805 38295 16845
rect 38305 16805 38345 16845
rect 38355 16805 38395 16845
rect 38405 16805 38445 16845
rect 38455 16805 38495 16845
rect 38505 16805 38545 16845
rect 38555 16805 38595 16845
rect 38605 16805 38645 16845
rect 38655 16805 38695 16845
rect 38705 16805 38745 16845
rect 38755 16805 38795 16845
rect 38805 16805 38845 16845
rect 38855 16805 38895 16845
rect 38905 16805 38945 16845
rect 38955 16805 38995 16845
rect 39005 16805 39045 16845
rect 39055 16805 39095 16845
rect 39105 16805 39145 16845
rect 39155 16805 39195 16845
rect 39205 16805 39245 16845
rect 39255 16805 39295 16845
rect 39305 16805 39345 16845
rect 39355 16805 39395 16845
rect 39405 16805 39445 16845
rect 39455 16805 39495 16845
rect 39505 16805 39545 16845
rect 39555 16805 39595 16845
rect 39605 16805 39645 16845
rect 39655 16805 39695 16845
rect 39705 16805 39745 16845
rect 5 15805 45 15845
rect 55 15805 95 15845
rect 105 15805 145 15845
rect 155 15805 195 15845
rect 205 15805 245 15845
rect 255 15805 295 15845
rect 305 15805 345 15845
rect 355 15805 395 15845
rect 405 15805 445 15845
rect 455 15805 495 15845
rect 505 15805 545 15845
rect 555 15805 595 15845
rect 605 15805 645 15845
rect 655 15805 695 15845
rect 705 15805 745 15845
rect 755 15805 795 15845
rect 805 15805 845 15845
rect 855 15805 895 15845
rect 905 15805 945 15845
rect 955 15805 995 15845
rect 1005 15805 1045 15845
rect 1055 15805 1095 15845
rect 1105 15805 1145 15845
rect 1155 15805 1195 15845
rect 1205 15805 1245 15845
rect 1255 15805 1295 15845
rect 1305 15805 1345 15845
rect 1355 15805 1395 15845
rect 1405 15805 1445 15845
rect 1455 15805 1495 15845
rect 1505 15805 1545 15845
rect 1555 15805 1595 15845
rect 1605 15805 1645 15845
rect 1655 15805 1695 15845
rect 1705 15805 1745 15845
rect 1755 15805 1795 15845
rect 1805 15805 1845 15845
rect 1855 15805 1895 15845
rect 1905 15805 1945 15845
rect 1955 15805 1995 15845
rect 2005 15805 2045 15845
rect 2055 15805 2095 15845
rect 2105 15805 2145 15845
rect 2155 15805 2195 15845
rect 2205 15805 2245 15845
rect 2255 15805 2295 15845
rect 2305 15805 2345 15845
rect 2355 15805 2395 15845
rect 2405 15805 2445 15845
rect 2455 15805 2495 15845
rect 2505 15805 2545 15845
rect 2555 15805 2595 15845
rect 2605 15805 2645 15845
rect 2655 15805 2695 15845
rect 2705 15805 2745 15845
rect 2755 15805 2795 15845
rect 2805 15805 2845 15845
rect 2855 15805 2895 15845
rect 2905 15805 2945 15845
rect 2955 15805 2995 15845
rect 3005 15805 3045 15845
rect 3055 15805 3095 15845
rect 3105 15805 3145 15845
rect 3155 15805 3195 15845
rect 3205 15805 3245 15845
rect 3255 15805 3295 15845
rect 3305 15805 3345 15845
rect 3355 15805 3395 15845
rect 3405 15805 3445 15845
rect 3455 15805 3495 15845
rect 3505 15805 3545 15845
rect 3555 15805 3595 15845
rect 3605 15805 3645 15845
rect 3655 15805 3695 15845
rect 3705 15805 3745 15845
rect 3755 15805 3795 15845
rect 3805 15805 3845 15845
rect 3855 15805 3895 15845
rect 3905 15805 3945 15845
rect 3955 15805 3995 15845
rect 4005 15805 4045 15845
rect 4055 15805 4095 15845
rect 4105 15805 4145 15845
rect 4155 15805 4195 15845
rect 4205 15805 4245 15845
rect 4255 15805 4295 15845
rect 4305 15805 4345 15845
rect 4355 15805 4395 15845
rect 4405 15805 4445 15845
rect 4455 15805 4495 15845
rect 4505 15805 4545 15845
rect 4555 15805 4595 15845
rect 4605 15805 4645 15845
rect 4655 15805 4695 15845
rect 4705 15805 4745 15845
rect 4755 15805 4795 15845
rect 4805 15805 4845 15845
rect 4855 15805 4895 15845
rect 4905 15805 4945 15845
rect 4955 15805 4995 15845
rect 5005 15805 5045 15845
rect 5055 15805 5095 15845
rect 5105 15805 5145 15845
rect 5155 15805 5195 15845
rect 5205 15805 5245 15845
rect 5255 15805 5295 15845
rect 5305 15805 5345 15845
rect 5355 15805 5395 15845
rect 5405 15805 5445 15845
rect 5455 15805 5495 15845
rect 5505 15805 5545 15845
rect 5555 15805 5595 15845
rect 5605 15805 5645 15845
rect 5655 15805 5695 15845
rect 5705 15805 5745 15845
rect 5755 15805 5795 15845
rect 5805 15805 5845 15845
rect 5855 15805 5895 15845
rect 5905 15805 5945 15845
rect 5955 15805 5995 15845
rect 6005 15805 6045 15845
rect 6055 15805 6095 15845
rect 6105 15805 6145 15845
rect 6155 15805 6195 15845
rect 6205 15805 6245 15845
rect 6255 15805 6295 15845
rect 6305 15805 6345 15845
rect 6355 15805 6395 15845
rect 6405 15805 6445 15845
rect 6455 15805 6495 15845
rect 6505 15805 6545 15845
rect 6555 15805 6595 15845
rect 6605 15805 6645 15845
rect 6655 15805 6695 15845
rect 6705 15805 6745 15845
rect 6755 15805 6795 15845
rect 6805 15805 6845 15845
rect 6855 15805 6895 15845
rect 6905 15805 6945 15845
rect 6955 15805 6995 15845
rect 7005 15805 7045 15845
rect 7055 15805 7095 15845
rect 7105 15805 7145 15845
rect 7155 15805 7195 15845
rect 7205 15805 7245 15845
rect 7255 15805 7295 15845
rect 7305 15805 7345 15845
rect 7355 15805 7395 15845
rect 7405 15805 7445 15845
rect 7455 15805 7495 15845
rect 7505 15805 7545 15845
rect 7555 15805 7595 15845
rect 7605 15805 7645 15845
rect 7655 15805 7695 15845
rect 7705 15805 7745 15845
rect 7755 15805 7795 15845
rect 7805 15805 7845 15845
rect 7855 15805 7895 15845
rect 7905 15805 7945 15845
rect 7955 15805 7995 15845
rect 8005 15805 8045 15845
rect 8055 15805 8095 15845
rect 8105 15805 8145 15845
rect 8155 15805 8195 15845
rect 8205 15805 8245 15845
rect 8255 15805 8295 15845
rect 8305 15805 8345 15845
rect 8355 15805 8395 15845
rect 8405 15805 8445 15845
rect 8455 15805 8495 15845
rect 8505 15805 8545 15845
rect 8555 15805 8595 15845
rect 8605 15805 8645 15845
rect 8655 15805 8695 15845
rect 8705 15805 8745 15845
rect 8755 15805 8795 15845
rect 8805 15805 8845 15845
rect 8855 15805 8895 15845
rect 8905 15805 8945 15845
rect 8955 15805 8995 15845
rect 9005 15805 9045 15845
rect 9055 15805 9095 15845
rect 9105 15805 9145 15845
rect 9155 15805 9195 15845
rect 9205 15805 9245 15845
rect 9255 15805 9295 15845
rect 9305 15805 9345 15845
rect 9355 15805 9395 15845
rect 9405 15805 9445 15845
rect 9455 15805 9495 15845
rect 9505 15805 9545 15845
rect 9555 15805 9595 15845
rect 9605 15805 9645 15845
rect 9655 15805 9695 15845
rect 9705 15805 9745 15845
rect 9755 15805 9795 15845
rect 9805 15805 9845 15845
rect 9855 15805 9895 15845
rect 9905 15805 9945 15845
rect 9955 15805 9995 15845
rect 10005 15805 10045 15845
rect 10055 15805 10095 15845
rect 10105 15805 10145 15845
rect 10155 15805 10195 15845
rect 10205 15805 10245 15845
rect 10255 15805 10295 15845
rect 10305 15805 10345 15845
rect 10355 15805 10395 15845
rect 10405 15805 10445 15845
rect 10455 15805 10495 15845
rect 10505 15805 10545 15845
rect 10555 15805 10595 15845
rect 10605 15805 10645 15845
rect 10655 15805 10695 15845
rect 10705 15805 10745 15845
rect 10755 15805 10795 15845
rect 10805 15805 10845 15845
rect 10855 15805 10895 15845
rect 10905 15805 10945 15845
rect 10955 15805 10995 15845
rect 11005 15805 11045 15845
rect 11055 15805 11095 15845
rect 11105 15805 11145 15845
rect 11155 15805 11195 15845
rect 11205 15805 11245 15845
rect 11255 15805 11295 15845
rect 11305 15805 11345 15845
rect 11355 15805 11395 15845
rect 11405 15805 11445 15845
rect 11455 15805 11495 15845
rect 11505 15805 11545 15845
rect 11555 15805 11595 15845
rect 11605 15805 11645 15845
rect 11655 15805 11695 15845
rect 11705 15805 11745 15845
rect 11755 15805 11795 15845
rect 11805 15805 11845 15845
rect 11855 15805 11895 15845
rect 11905 15805 11945 15845
rect 11955 15805 11995 15845
rect 12005 15805 12045 15845
rect 12055 15805 12095 15845
rect 12105 15805 12145 15845
rect 12155 15805 12195 15845
rect 12205 15805 12245 15845
rect 12255 15805 12295 15845
rect 12305 15805 12345 15845
rect 12355 15805 12395 15845
rect 12405 15805 12445 15845
rect 12455 15805 12495 15845
rect 12505 15805 12545 15845
rect 12555 15805 12595 15845
rect 12605 15805 12645 15845
rect 12655 15805 12695 15845
rect 12705 15805 12745 15845
rect 12755 15805 12795 15845
rect 12805 15805 12845 15845
rect 12855 15805 12895 15845
rect 12905 15805 12945 15845
rect 12955 15805 12995 15845
rect 13005 15805 13045 15845
rect 13055 15805 13095 15845
rect 13105 15805 13145 15845
rect 13155 15805 13195 15845
rect 13205 15805 13245 15845
rect 13255 15805 13295 15845
rect 13305 15805 13345 15845
rect 13355 15805 13395 15845
rect 13405 15805 13445 15845
rect 13455 15805 13495 15845
rect 13505 15805 13545 15845
rect 13555 15805 13595 15845
rect 13605 15805 13645 15845
rect 13655 15805 13695 15845
rect 13705 15805 13745 15845
rect 13755 15805 13795 15845
rect 13805 15805 13845 15845
rect 13855 15805 13895 15845
rect 13905 15805 13945 15845
rect 13955 15805 13995 15845
rect 14005 15805 14045 15845
rect 14055 15805 14095 15845
rect 14105 15805 14145 15845
rect 14155 15805 14195 15845
rect 14205 15805 14245 15845
rect 14255 15805 14295 15845
rect 14305 15805 14345 15845
rect 14355 15805 14395 15845
rect 14405 15805 14445 15845
rect 14455 15805 14495 15845
rect 14505 15805 14545 15845
rect 14555 15805 14595 15845
rect 14605 15805 14645 15845
rect 14655 15805 14695 15845
rect 14705 15805 14745 15845
rect 14755 15805 14795 15845
rect 14805 15805 14845 15845
rect 14855 15805 14895 15845
rect 14905 15805 14945 15845
rect 14955 15805 14995 15845
rect 15005 15805 15045 15845
rect 15055 15805 15095 15845
rect 15105 15805 15145 15845
rect 15155 15805 15195 15845
rect 15205 15805 15245 15845
rect 15255 15805 15295 15845
rect 15305 15805 15345 15845
rect 15355 15805 15395 15845
rect 15405 15805 15445 15845
rect 15455 15805 15495 15845
rect 15505 15805 15545 15845
rect 15555 15805 15595 15845
rect 15605 15805 15645 15845
rect 15655 15805 15695 15845
rect 15705 15805 15745 15845
rect 15755 15805 15795 15845
rect 15805 15805 15845 15845
rect 15855 15805 15895 15845
rect 15905 15805 15945 15845
rect 15955 15805 15995 15845
rect 16005 15805 16045 15845
rect 16055 15805 16095 15845
rect 16105 15805 16145 15845
rect 16155 15805 16195 15845
rect 16205 15805 16245 15845
rect 16255 15805 16295 15845
rect 16305 15805 16345 15845
rect 16355 15805 16395 15845
rect 16405 15805 16445 15845
rect 16455 15805 16495 15845
rect 16505 15805 16545 15845
rect 16555 15805 16595 15845
rect 16605 15805 16645 15845
rect 16655 15805 16695 15845
rect 16705 15805 16745 15845
rect 16755 15805 16795 15845
rect 16805 15805 16845 15845
rect 16855 15805 16895 15845
rect 16905 15805 16945 15845
rect 16955 15805 16995 15845
rect 17005 15805 17045 15845
rect 17055 15805 17095 15845
rect 17105 15805 17145 15845
rect 17155 15805 17195 15845
rect 17205 15805 17245 15845
rect 17255 15805 17295 15845
rect 17305 15805 17345 15845
rect 17355 15805 17395 15845
rect 17405 15805 17445 15845
rect 17455 15805 17495 15845
rect 17505 15805 17545 15845
rect 17555 15805 17595 15845
rect 17605 15805 17645 15845
rect 17655 15805 17695 15845
rect 17705 15805 17745 15845
rect 17755 15805 17795 15845
rect 17805 15805 17845 15845
rect 17855 15805 17895 15845
rect 17905 15805 17945 15845
rect 17955 15805 17995 15845
rect 18005 15805 18045 15845
rect 18055 15805 18095 15845
rect 18105 15805 18145 15845
rect 18155 15805 18195 15845
rect 18205 15805 18245 15845
rect 18255 15805 18295 15845
rect 18305 15805 18345 15845
rect 18355 15805 18395 15845
rect 18405 15805 18445 15845
rect 18455 15805 18495 15845
rect 18505 15805 18545 15845
rect 18555 15805 18595 15845
rect 18605 15805 18645 15845
rect 18655 15805 18695 15845
rect 18705 15805 18745 15845
rect 18755 15805 18795 15845
rect 18805 15805 18845 15845
rect 18855 15805 18895 15845
rect 18905 15805 18945 15845
rect 18955 15805 18995 15845
rect 19005 15805 19045 15845
rect 19055 15805 19095 15845
rect 19105 15805 19145 15845
rect 19155 15805 19195 15845
rect 19205 15805 19245 15845
rect 19255 15805 19295 15845
rect 19305 15805 19345 15845
rect 19355 15805 19395 15845
rect 19405 15805 19445 15845
rect 19455 15805 19495 15845
rect 19505 15805 19545 15845
rect 19555 15805 19595 15845
rect 19605 15805 19645 15845
rect 19655 15805 19695 15845
rect 19705 15805 19745 15845
rect 19755 15805 19795 15845
rect 19805 15805 19845 15845
rect 19855 15805 19895 15845
rect 19905 15805 19945 15845
rect 19955 15805 19995 15845
rect 20005 15805 20045 15845
rect 20055 15805 20095 15845
rect 20105 15805 20145 15845
rect 20155 15805 20195 15845
rect 20205 15805 20245 15845
rect 20255 15805 20295 15845
rect 20305 15805 20345 15845
rect 20355 15805 20395 15845
rect 20405 15805 20445 15845
rect 20455 15805 20495 15845
rect 20505 15805 20545 15845
rect 20555 15805 20595 15845
rect 20605 15805 20645 15845
rect 20655 15805 20695 15845
rect 20705 15805 20745 15845
rect 20755 15805 20795 15845
rect 20805 15805 20845 15845
rect 20855 15805 20895 15845
rect 20905 15805 20945 15845
rect 20955 15805 20995 15845
rect 21005 15805 21045 15845
rect 21055 15805 21095 15845
rect 21105 15805 21145 15845
rect 21155 15805 21195 15845
rect 21205 15805 21245 15845
rect 21255 15805 21295 15845
rect 21305 15805 21345 15845
rect 21355 15805 21395 15845
rect 21405 15805 21445 15845
rect 21455 15805 21495 15845
rect 21505 15805 21545 15845
rect 21555 15805 21595 15845
rect 21605 15805 21645 15845
rect 21655 15805 21695 15845
rect 21705 15805 21745 15845
rect 21755 15805 21795 15845
rect 21805 15805 21845 15845
rect 21855 15805 21895 15845
rect 21905 15805 21945 15845
rect 21955 15805 21995 15845
rect 22005 15805 22045 15845
rect 22055 15805 22095 15845
rect 22105 15805 22145 15845
rect 22155 15805 22195 15845
rect 22205 15805 22245 15845
rect 22255 15805 22295 15845
rect 22305 15805 22345 15845
rect 22355 15805 22395 15845
rect 22405 15805 22445 15845
rect 22455 15805 22495 15845
rect 22505 15805 22545 15845
rect 22555 15805 22595 15845
rect 22605 15805 22645 15845
rect 22655 15805 22695 15845
rect 22705 15805 22745 15845
rect 22755 15805 22795 15845
rect 22805 15805 22845 15845
rect 22855 15805 22895 15845
rect 22905 15805 22945 15845
rect 22955 15805 22995 15845
rect 23005 15805 23045 15845
rect 23055 15805 23095 15845
rect 23105 15805 23145 15845
rect 23155 15805 23195 15845
rect 23205 15805 23245 15845
rect 23255 15805 23295 15845
rect 23305 15805 23345 15845
rect 23355 15805 23395 15845
rect 23405 15805 23445 15845
rect 23455 15805 23495 15845
rect 23505 15805 23545 15845
rect 23555 15805 23595 15845
rect 23605 15805 23645 15845
rect 23655 15805 23695 15845
rect 23705 15805 23745 15845
rect 23755 15805 23795 15845
rect 23805 15805 23845 15845
rect 23855 15805 23895 15845
rect 23905 15805 23945 15845
rect 23955 15805 23995 15845
rect 24005 15805 24045 15845
rect 24055 15805 24095 15845
rect 24105 15805 24145 15845
rect 24155 15805 24195 15845
rect 24205 15805 24245 15845
rect 24255 15805 24295 15845
rect 24305 15805 24345 15845
rect 24355 15805 24395 15845
rect 24405 15805 24445 15845
rect 24455 15805 24495 15845
rect 24505 15805 24545 15845
rect 24555 15805 24595 15845
rect 24605 15805 24645 15845
rect 24655 15805 24695 15845
rect 24705 15805 24745 15845
rect 24755 15805 24795 15845
rect 24805 15805 24845 15845
rect 24855 15805 24895 15845
rect 24905 15805 24945 15845
rect 24955 15805 24995 15845
rect 25005 15805 25045 15845
rect 25055 15805 25095 15845
rect 25105 15805 25145 15845
rect 25155 15805 25195 15845
rect 25205 15805 25245 15845
rect 25255 15805 25295 15845
rect 25305 15805 25345 15845
rect 25355 15805 25395 15845
rect 25405 15805 25445 15845
rect 25455 15805 25495 15845
rect 25505 15805 25545 15845
rect 25555 15805 25595 15845
rect 25605 15805 25645 15845
rect 25655 15805 25695 15845
rect 25705 15805 25745 15845
rect 25755 15805 25795 15845
rect 25805 15805 25845 15845
rect 25855 15805 25895 15845
rect 25905 15805 25945 15845
rect 25955 15805 25995 15845
rect 26005 15805 26045 15845
rect 26055 15805 26095 15845
rect 26105 15805 26145 15845
rect 26155 15805 26195 15845
rect 26205 15805 26245 15845
rect 26255 15805 26295 15845
rect 26305 15805 26345 15845
rect 26355 15805 26395 15845
rect 26405 15805 26445 15845
rect 26455 15805 26495 15845
rect 26505 15805 26545 15845
rect 26555 15805 26595 15845
rect 26605 15805 26645 15845
rect 26655 15805 26695 15845
rect 26705 15805 26745 15845
rect 26755 15805 26795 15845
rect 26805 15805 26845 15845
rect 26855 15805 26895 15845
rect 26905 15805 26945 15845
rect 26955 15805 26995 15845
rect 27005 15805 27045 15845
rect 27055 15805 27095 15845
rect 27105 15805 27145 15845
rect 27155 15805 27195 15845
rect 27205 15805 27245 15845
rect 27255 15805 27295 15845
rect 27305 15805 27345 15845
rect 27355 15805 27395 15845
rect 27405 15805 27445 15845
rect 27455 15805 27495 15845
rect 27505 15805 27545 15845
rect 27555 15805 27595 15845
rect 27605 15805 27645 15845
rect 27655 15805 27695 15845
rect 27705 15805 27745 15845
rect 27755 15805 27795 15845
rect 27805 15805 27845 15845
rect 27855 15805 27895 15845
rect 27905 15805 27945 15845
rect 27955 15805 27995 15845
rect 28005 15805 28045 15845
rect 28055 15805 28095 15845
rect 28105 15805 28145 15845
rect 28155 15805 28195 15845
rect 28205 15805 28245 15845
rect 28255 15805 28295 15845
rect 28305 15805 28345 15845
rect 28355 15805 28395 15845
rect 28405 15805 28445 15845
rect 28455 15805 28495 15845
rect 28505 15805 28545 15845
rect 28555 15805 28595 15845
rect 28605 15805 28645 15845
rect 28655 15805 28695 15845
rect 28705 15805 28745 15845
rect 28755 15805 28795 15845
rect 28805 15805 28845 15845
rect 28855 15805 28895 15845
rect 28905 15805 28945 15845
rect 28955 15805 28995 15845
rect 29005 15805 29045 15845
rect 29055 15805 29095 15845
rect 29105 15805 29145 15845
rect 29155 15805 29195 15845
rect 29205 15805 29245 15845
rect 29255 15805 29295 15845
rect 29305 15805 29345 15845
rect 29355 15805 29395 15845
rect 29405 15805 29445 15845
rect 29455 15805 29495 15845
rect 29505 15805 29545 15845
rect 29555 15805 29595 15845
rect 29605 15805 29645 15845
rect 29655 15805 29695 15845
rect 29705 15805 29745 15845
rect 29755 15805 29795 15845
rect 29805 15805 29845 15845
rect 29855 15805 29895 15845
rect 29905 15805 29945 15845
rect 29955 15805 29995 15845
rect 30005 15805 30045 15845
rect 30055 15805 30095 15845
rect 30105 15805 30145 15845
rect 30155 15805 30195 15845
rect 30205 15805 30245 15845
rect 30255 15805 30295 15845
rect 30305 15805 30345 15845
rect 30355 15805 30395 15845
rect 30405 15805 30445 15845
rect 30455 15805 30495 15845
rect 30505 15805 30545 15845
rect 30555 15805 30595 15845
rect 30605 15805 30645 15845
rect 30655 15805 30695 15845
rect 30705 15805 30745 15845
rect 30755 15805 30795 15845
rect 30805 15805 30845 15845
rect 30855 15805 30895 15845
rect 30905 15805 30945 15845
rect 30955 15805 30995 15845
rect 31005 15805 31045 15845
rect 31055 15805 31095 15845
rect 31105 15805 31145 15845
rect 31155 15805 31195 15845
rect 31205 15805 31245 15845
rect 31255 15805 31295 15845
rect 31305 15805 31345 15845
rect 31355 15805 31395 15845
rect 31405 15805 31445 15845
rect 31455 15805 31495 15845
rect 31505 15805 31545 15845
rect 31555 15805 31595 15845
rect 31605 15805 31645 15845
rect 31655 15805 31695 15845
rect 31705 15805 31745 15845
rect 31755 15805 31795 15845
rect 31805 15805 31845 15845
rect 31855 15805 31895 15845
rect 31905 15805 31945 15845
rect 31955 15805 31995 15845
rect 32005 15805 32045 15845
rect 32055 15805 32095 15845
rect 32105 15805 32145 15845
rect 32155 15805 32195 15845
rect 32205 15805 32245 15845
rect 32255 15805 32295 15845
rect 32305 15805 32345 15845
rect 32355 15805 32395 15845
rect 32405 15805 32445 15845
rect 32455 15805 32495 15845
rect 32505 15805 32545 15845
rect 32555 15805 32595 15845
rect 32605 15805 32645 15845
rect 32655 15805 32695 15845
rect 32705 15805 32745 15845
rect 32755 15805 32795 15845
rect 32805 15805 32845 15845
rect 32855 15805 32895 15845
rect 32905 15805 32945 15845
rect 32955 15805 32995 15845
rect 33005 15805 33045 15845
rect 33055 15805 33095 15845
rect 33105 15805 33145 15845
rect 33155 15805 33195 15845
rect 33205 15805 33245 15845
rect 33255 15805 33295 15845
rect 33305 15805 33345 15845
rect 33355 15805 33395 15845
rect 33405 15805 33445 15845
rect 33455 15805 33495 15845
rect 33505 15805 33545 15845
rect 33555 15805 33595 15845
rect 33605 15805 33645 15845
rect 33655 15805 33695 15845
rect 33705 15805 33745 15845
rect 33755 15805 33795 15845
rect 33805 15805 33845 15845
rect 33855 15805 33895 15845
rect 33905 15805 33945 15845
rect 33955 15805 33995 15845
rect 34005 15805 34045 15845
rect 34055 15805 34095 15845
rect 34105 15805 34145 15845
rect 34155 15805 34195 15845
rect 34205 15805 34245 15845
rect 34255 15805 34295 15845
rect 34305 15805 34345 15845
rect 34355 15805 34395 15845
rect 34405 15805 34445 15845
rect 34455 15805 34495 15845
rect 34505 15805 34545 15845
rect 34555 15805 34595 15845
rect 34605 15805 34645 15845
rect 34655 15805 34695 15845
rect 34705 15805 34745 15845
rect 34755 15805 34795 15845
rect 34805 15805 34845 15845
rect 34855 15805 34895 15845
rect 34905 15805 34945 15845
rect 34955 15805 34995 15845
rect 35005 15805 35045 15845
rect 35055 15805 35095 15845
rect 35105 15805 35145 15845
rect 35155 15805 35195 15845
rect 35205 15805 35245 15845
rect 35255 15805 35295 15845
rect 35305 15805 35345 15845
rect 35355 15805 35395 15845
rect 35405 15805 35445 15845
rect 35455 15805 35495 15845
rect 35505 15805 35545 15845
rect 35555 15805 35595 15845
rect 35605 15805 35645 15845
rect 35655 15805 35695 15845
rect 35705 15805 35745 15845
rect 35755 15805 35795 15845
rect 35805 15805 35845 15845
rect 35855 15805 35895 15845
rect 35905 15805 35945 15845
rect 35955 15805 35995 15845
rect 36005 15805 36045 15845
rect 36055 15805 36095 15845
rect 36105 15805 36145 15845
rect 36155 15805 36195 15845
rect 36205 15805 36245 15845
rect 36255 15805 36295 15845
rect 36305 15805 36345 15845
rect 36355 15805 36395 15845
rect 36405 15805 36445 15845
rect 36455 15805 36495 15845
rect 36505 15805 36545 15845
rect 36555 15805 36595 15845
rect 36605 15805 36645 15845
rect 36655 15805 36695 15845
rect 36705 15805 36745 15845
rect 36755 15805 36795 15845
rect 36805 15805 36845 15845
rect 36855 15805 36895 15845
rect 36905 15805 36945 15845
rect 36955 15805 36995 15845
rect 37005 15805 37045 15845
rect 37055 15805 37095 15845
rect 37105 15805 37145 15845
rect 37155 15805 37195 15845
rect 37205 15805 37245 15845
rect 37255 15805 37295 15845
rect 37305 15805 37345 15845
rect 37355 15805 37395 15845
rect 37405 15805 37445 15845
rect 37455 15805 37495 15845
rect 37505 15805 37545 15845
rect 37555 15805 37595 15845
rect 37605 15805 37645 15845
rect 37655 15805 37695 15845
rect 37705 15805 37745 15845
rect 37755 15805 37795 15845
rect 37805 15805 37845 15845
rect 37855 15805 37895 15845
rect 37905 15805 37945 15845
rect 37955 15805 37995 15845
rect 38005 15805 38045 15845
rect 38055 15805 38095 15845
rect 38105 15805 38145 15845
rect 38155 15805 38195 15845
rect 38205 15805 38245 15845
rect 38255 15805 38295 15845
rect 38305 15805 38345 15845
rect 38355 15805 38395 15845
rect 38405 15805 38445 15845
rect 38455 15805 38495 15845
rect 38505 15805 38545 15845
rect 38555 15805 38595 15845
rect 38605 15805 38645 15845
rect 38655 15805 38695 15845
rect 38705 15805 38745 15845
rect 38755 15805 38795 15845
rect 38805 15805 38845 15845
rect 38855 15805 38895 15845
rect 38905 15805 38945 15845
rect 38955 15805 38995 15845
rect 39005 15805 39045 15845
rect 39055 15805 39095 15845
rect 39105 15805 39145 15845
rect 39155 15805 39195 15845
rect 39205 15805 39245 15845
rect 39255 15805 39295 15845
rect 39305 15805 39345 15845
rect 39355 15805 39395 15845
rect 39405 15805 39445 15845
rect 39455 15805 39495 15845
rect 39505 15805 39545 15845
rect 39555 15805 39595 15845
rect 39605 15805 39645 15845
rect 39655 15805 39695 15845
rect 39705 15805 39745 15845
rect -3495 15740 -3455 15745
rect -3495 15710 -3490 15740
rect -3490 15710 -3460 15740
rect -3460 15710 -3455 15740
rect -3495 15705 -3455 15710
rect -3295 15740 -3255 15745
rect -3295 15710 -3290 15740
rect -3290 15710 -3260 15740
rect -3260 15710 -3255 15740
rect -3295 15705 -3255 15710
rect -3095 15740 -3055 15745
rect -3095 15710 -3090 15740
rect -3090 15710 -3060 15740
rect -3060 15710 -3055 15740
rect -3095 15705 -3055 15710
rect -1595 15740 -1555 15745
rect -1595 15710 -1590 15740
rect -1590 15710 -1560 15740
rect -1560 15710 -1555 15740
rect -1595 15705 -1555 15710
rect -1195 15740 -1155 15745
rect -1195 15710 -1190 15740
rect -1190 15710 -1160 15740
rect -1160 15710 -1155 15740
rect -1195 15705 -1155 15710
rect -1095 15740 -1055 15745
rect -1095 15710 -1090 15740
rect -1090 15710 -1060 15740
rect -1060 15710 -1055 15740
rect -1095 15705 -1055 15710
rect -995 15740 -955 15745
rect -995 15710 -990 15740
rect -990 15710 -960 15740
rect -960 15710 -955 15740
rect -995 15705 -955 15710
rect -895 15740 -855 15745
rect -895 15710 -890 15740
rect -890 15710 -860 15740
rect -860 15710 -855 15740
rect -895 15705 -855 15710
rect -695 15740 -655 15745
rect -695 15710 -690 15740
rect -690 15710 -660 15740
rect -660 15710 -655 15740
rect -695 15705 -655 15710
rect -595 15740 -555 15745
rect -595 15710 -590 15740
rect -590 15710 -560 15740
rect -560 15710 -555 15740
rect -595 15705 -555 15710
rect -495 15740 -455 15745
rect -495 15710 -490 15740
rect -490 15710 -460 15740
rect -460 15710 -455 15740
rect -495 15705 -455 15710
rect -295 15740 -255 15745
rect -295 15710 -290 15740
rect -290 15710 -260 15740
rect -260 15710 -255 15740
rect -295 15705 -255 15710
rect -195 15740 -155 15745
rect -195 15710 -190 15740
rect -190 15710 -160 15740
rect -160 15710 -155 15740
rect -195 15705 -155 15710
rect -95 15740 -55 15745
rect -95 15710 -90 15740
rect -90 15710 -60 15740
rect -60 15710 -55 15740
rect -95 15705 -55 15710
rect 5 15705 45 15745
rect 55 15705 95 15745
rect 105 15705 145 15745
rect 155 15705 195 15745
rect 205 15705 245 15745
rect 255 15705 295 15745
rect 305 15705 345 15745
rect 355 15705 395 15745
rect 405 15705 445 15745
rect 455 15705 495 15745
rect 505 15705 545 15745
rect 555 15705 595 15745
rect 605 15705 645 15745
rect 655 15705 695 15745
rect 705 15705 745 15745
rect 755 15705 795 15745
rect 805 15705 845 15745
rect 855 15705 895 15745
rect 905 15705 945 15745
rect 955 15705 995 15745
rect 1005 15705 1045 15745
rect 1055 15705 1095 15745
rect 1105 15705 1145 15745
rect 1155 15705 1195 15745
rect 1205 15705 1245 15745
rect 1255 15705 1295 15745
rect 1305 15705 1345 15745
rect 1355 15705 1395 15745
rect 1405 15705 1445 15745
rect 1455 15705 1495 15745
rect 1505 15705 1545 15745
rect 1555 15705 1595 15745
rect 1605 15705 1645 15745
rect 1655 15705 1695 15745
rect 1705 15705 1745 15745
rect 1755 15705 1795 15745
rect 1805 15705 1845 15745
rect 1855 15705 1895 15745
rect 1905 15705 1945 15745
rect 1955 15705 1995 15745
rect 2005 15705 2045 15745
rect 2055 15705 2095 15745
rect 2105 15705 2145 15745
rect 2155 15705 2195 15745
rect 2205 15705 2245 15745
rect 2255 15705 2295 15745
rect 2305 15705 2345 15745
rect 2355 15705 2395 15745
rect 2405 15705 2445 15745
rect 2455 15705 2495 15745
rect 2505 15705 2545 15745
rect 2555 15705 2595 15745
rect 2605 15705 2645 15745
rect 2655 15705 2695 15745
rect 2705 15705 2745 15745
rect 2755 15705 2795 15745
rect 2805 15705 2845 15745
rect 2855 15705 2895 15745
rect 2905 15705 2945 15745
rect 2955 15705 2995 15745
rect 3005 15705 3045 15745
rect 3055 15705 3095 15745
rect 3105 15705 3145 15745
rect 3155 15705 3195 15745
rect 3205 15705 3245 15745
rect 3255 15705 3295 15745
rect 3305 15705 3345 15745
rect 3355 15705 3395 15745
rect 3405 15705 3445 15745
rect 3455 15705 3495 15745
rect 3505 15705 3545 15745
rect 3555 15705 3595 15745
rect 3605 15705 3645 15745
rect 3655 15705 3695 15745
rect 3705 15705 3745 15745
rect 3755 15705 3795 15745
rect 3805 15705 3845 15745
rect 3855 15705 3895 15745
rect 3905 15705 3945 15745
rect 3955 15705 3995 15745
rect 4005 15705 4045 15745
rect 4055 15705 4095 15745
rect 4105 15705 4145 15745
rect 4155 15705 4195 15745
rect 4205 15705 4245 15745
rect 4255 15705 4295 15745
rect 4305 15705 4345 15745
rect 4355 15705 4395 15745
rect 4405 15705 4445 15745
rect 4455 15705 4495 15745
rect 4505 15705 4545 15745
rect 4555 15705 4595 15745
rect 4605 15705 4645 15745
rect 4655 15705 4695 15745
rect 4705 15705 4745 15745
rect 4755 15705 4795 15745
rect 4805 15705 4845 15745
rect 4855 15705 4895 15745
rect 4905 15705 4945 15745
rect 4955 15705 4995 15745
rect 5005 15705 5045 15745
rect 5055 15705 5095 15745
rect 5105 15705 5145 15745
rect 5155 15705 5195 15745
rect 5205 15705 5245 15745
rect 5255 15705 5295 15745
rect 5305 15705 5345 15745
rect 5355 15705 5395 15745
rect 5405 15705 5445 15745
rect 5455 15705 5495 15745
rect 5505 15705 5545 15745
rect 5555 15705 5595 15745
rect 5605 15705 5645 15745
rect 5655 15705 5695 15745
rect 5705 15705 5745 15745
rect 5755 15705 5795 15745
rect 5805 15705 5845 15745
rect 5855 15705 5895 15745
rect 5905 15705 5945 15745
rect 5955 15705 5995 15745
rect 6005 15705 6045 15745
rect 6055 15705 6095 15745
rect 6105 15705 6145 15745
rect 6155 15705 6195 15745
rect 6205 15705 6245 15745
rect 6255 15705 6295 15745
rect 6305 15705 6345 15745
rect 6355 15705 6395 15745
rect 6405 15705 6445 15745
rect 6455 15705 6495 15745
rect 6505 15705 6545 15745
rect 6555 15705 6595 15745
rect 6605 15705 6645 15745
rect 6655 15705 6695 15745
rect 6705 15705 6745 15745
rect 6755 15705 6795 15745
rect 6805 15705 6845 15745
rect 6855 15705 6895 15745
rect 6905 15705 6945 15745
rect 6955 15705 6995 15745
rect 7005 15705 7045 15745
rect 7055 15705 7095 15745
rect 7105 15705 7145 15745
rect 7155 15705 7195 15745
rect 7205 15705 7245 15745
rect 7255 15705 7295 15745
rect 7305 15705 7345 15745
rect 7355 15705 7395 15745
rect 7405 15705 7445 15745
rect 7455 15705 7495 15745
rect 7505 15705 7545 15745
rect 7555 15705 7595 15745
rect 7605 15705 7645 15745
rect 7655 15705 7695 15745
rect 7705 15705 7745 15745
rect 7755 15705 7795 15745
rect 7805 15705 7845 15745
rect 7855 15705 7895 15745
rect 7905 15705 7945 15745
rect 7955 15705 7995 15745
rect 8005 15705 8045 15745
rect 8055 15705 8095 15745
rect 8105 15705 8145 15745
rect 8155 15705 8195 15745
rect 8205 15705 8245 15745
rect 8255 15705 8295 15745
rect 8305 15705 8345 15745
rect 8355 15705 8395 15745
rect 8405 15705 8445 15745
rect 8455 15705 8495 15745
rect 8505 15705 8545 15745
rect 8555 15705 8595 15745
rect 8605 15705 8645 15745
rect 8655 15705 8695 15745
rect 8705 15705 8745 15745
rect 8755 15705 8795 15745
rect 8805 15705 8845 15745
rect 8855 15705 8895 15745
rect 8905 15705 8945 15745
rect 8955 15705 8995 15745
rect 9005 15705 9045 15745
rect 9055 15705 9095 15745
rect 9105 15705 9145 15745
rect 9155 15705 9195 15745
rect 9205 15705 9245 15745
rect 9255 15705 9295 15745
rect 9305 15705 9345 15745
rect 9355 15705 9395 15745
rect 9405 15705 9445 15745
rect 9455 15705 9495 15745
rect 9505 15705 9545 15745
rect 9555 15705 9595 15745
rect 9605 15705 9645 15745
rect 9655 15705 9695 15745
rect 9705 15705 9745 15745
rect 9755 15705 9795 15745
rect 9805 15705 9845 15745
rect 9855 15705 9895 15745
rect 9905 15705 9945 15745
rect 9955 15705 9995 15745
rect 10005 15705 10045 15745
rect 10055 15705 10095 15745
rect 10105 15705 10145 15745
rect 10155 15705 10195 15745
rect 10205 15705 10245 15745
rect 10255 15705 10295 15745
rect 10305 15705 10345 15745
rect 10355 15705 10395 15745
rect 10405 15705 10445 15745
rect 10455 15705 10495 15745
rect 10505 15705 10545 15745
rect 10555 15705 10595 15745
rect 10605 15705 10645 15745
rect 10655 15705 10695 15745
rect 10705 15705 10745 15745
rect 10755 15705 10795 15745
rect 10805 15705 10845 15745
rect 10855 15705 10895 15745
rect 10905 15705 10945 15745
rect 10955 15705 10995 15745
rect 11005 15705 11045 15745
rect 11055 15705 11095 15745
rect 11105 15705 11145 15745
rect 11155 15705 11195 15745
rect 11205 15705 11245 15745
rect 11255 15705 11295 15745
rect 11305 15705 11345 15745
rect 11355 15705 11395 15745
rect 11405 15705 11445 15745
rect 11455 15705 11495 15745
rect 11505 15705 11545 15745
rect 11555 15705 11595 15745
rect 11605 15705 11645 15745
rect 11655 15705 11695 15745
rect 11705 15705 11745 15745
rect 11755 15705 11795 15745
rect 11805 15705 11845 15745
rect 11855 15705 11895 15745
rect 11905 15705 11945 15745
rect 11955 15705 11995 15745
rect 12005 15705 12045 15745
rect 12055 15705 12095 15745
rect 12105 15705 12145 15745
rect 12155 15705 12195 15745
rect 12205 15705 12245 15745
rect 12255 15705 12295 15745
rect 12305 15705 12345 15745
rect 12355 15705 12395 15745
rect 12405 15705 12445 15745
rect 12455 15705 12495 15745
rect 12505 15705 12545 15745
rect 12555 15705 12595 15745
rect 12605 15705 12645 15745
rect 12655 15705 12695 15745
rect 12705 15705 12745 15745
rect 12755 15705 12795 15745
rect 12805 15705 12845 15745
rect 12855 15705 12895 15745
rect 12905 15705 12945 15745
rect 12955 15705 12995 15745
rect 13005 15705 13045 15745
rect 13055 15705 13095 15745
rect 13105 15705 13145 15745
rect 13155 15705 13195 15745
rect 13205 15705 13245 15745
rect 13255 15705 13295 15745
rect 13305 15705 13345 15745
rect 13355 15705 13395 15745
rect 13405 15705 13445 15745
rect 13455 15705 13495 15745
rect 13505 15705 13545 15745
rect 13555 15705 13595 15745
rect 13605 15705 13645 15745
rect 13655 15705 13695 15745
rect 13705 15705 13745 15745
rect 13755 15705 13795 15745
rect 13805 15705 13845 15745
rect 13855 15705 13895 15745
rect 13905 15705 13945 15745
rect 13955 15705 13995 15745
rect 14005 15705 14045 15745
rect 14055 15705 14095 15745
rect 14105 15705 14145 15745
rect 14155 15705 14195 15745
rect 14205 15705 14245 15745
rect 14255 15705 14295 15745
rect 14305 15705 14345 15745
rect 14355 15705 14395 15745
rect 14405 15705 14445 15745
rect 14455 15705 14495 15745
rect 14505 15705 14545 15745
rect 14555 15705 14595 15745
rect 14605 15705 14645 15745
rect 14655 15705 14695 15745
rect 14705 15705 14745 15745
rect 14755 15705 14795 15745
rect 14805 15705 14845 15745
rect 14855 15705 14895 15745
rect 14905 15705 14945 15745
rect 14955 15705 14995 15745
rect 15005 15705 15045 15745
rect 15055 15705 15095 15745
rect 15105 15705 15145 15745
rect 15155 15705 15195 15745
rect 15205 15705 15245 15745
rect 15255 15705 15295 15745
rect 15305 15705 15345 15745
rect 15355 15705 15395 15745
rect 15405 15705 15445 15745
rect 15455 15705 15495 15745
rect 15505 15705 15545 15745
rect 15555 15705 15595 15745
rect 15605 15705 15645 15745
rect 15655 15705 15695 15745
rect 15705 15705 15745 15745
rect 15755 15705 15795 15745
rect 15805 15705 15845 15745
rect 15855 15705 15895 15745
rect 15905 15705 15945 15745
rect 15955 15705 15995 15745
rect 16005 15705 16045 15745
rect 16055 15705 16095 15745
rect 16105 15705 16145 15745
rect 16155 15705 16195 15745
rect 16205 15705 16245 15745
rect 16255 15705 16295 15745
rect 16305 15705 16345 15745
rect 16355 15705 16395 15745
rect 16405 15705 16445 15745
rect 16455 15705 16495 15745
rect 16505 15705 16545 15745
rect 16555 15705 16595 15745
rect 16605 15705 16645 15745
rect 16655 15705 16695 15745
rect 16705 15705 16745 15745
rect 16755 15705 16795 15745
rect 16805 15705 16845 15745
rect 16855 15705 16895 15745
rect 16905 15705 16945 15745
rect 16955 15705 16995 15745
rect 17005 15705 17045 15745
rect 17055 15705 17095 15745
rect 17105 15705 17145 15745
rect 17155 15705 17195 15745
rect 17205 15705 17245 15745
rect 17255 15705 17295 15745
rect 17305 15705 17345 15745
rect 17355 15705 17395 15745
rect 17405 15705 17445 15745
rect 17455 15705 17495 15745
rect 17505 15705 17545 15745
rect 17555 15705 17595 15745
rect 17605 15705 17645 15745
rect 17655 15705 17695 15745
rect 17705 15705 17745 15745
rect 17755 15705 17795 15745
rect 17805 15705 17845 15745
rect 17855 15705 17895 15745
rect 17905 15705 17945 15745
rect 17955 15705 17995 15745
rect 18005 15705 18045 15745
rect 18055 15705 18095 15745
rect 18105 15705 18145 15745
rect 18155 15705 18195 15745
rect 18205 15705 18245 15745
rect 18255 15705 18295 15745
rect 18305 15705 18345 15745
rect 18355 15705 18395 15745
rect 18405 15705 18445 15745
rect 18455 15705 18495 15745
rect 18505 15705 18545 15745
rect 18555 15705 18595 15745
rect 18605 15705 18645 15745
rect 18655 15705 18695 15745
rect 18705 15705 18745 15745
rect 18755 15705 18795 15745
rect 18805 15705 18845 15745
rect 18855 15705 18895 15745
rect 18905 15705 18945 15745
rect 18955 15705 18995 15745
rect 19005 15705 19045 15745
rect 19055 15705 19095 15745
rect 19105 15705 19145 15745
rect 19155 15705 19195 15745
rect 19205 15705 19245 15745
rect 19255 15705 19295 15745
rect 19305 15705 19345 15745
rect 19355 15705 19395 15745
rect 19405 15705 19445 15745
rect 19455 15705 19495 15745
rect 19505 15705 19545 15745
rect 19555 15705 19595 15745
rect 19605 15705 19645 15745
rect 19655 15705 19695 15745
rect 19705 15705 19745 15745
rect 19755 15705 19795 15745
rect 19805 15705 19845 15745
rect 19855 15705 19895 15745
rect 19905 15705 19945 15745
rect 19955 15705 19995 15745
rect 20005 15705 20045 15745
rect 20055 15705 20095 15745
rect 20105 15705 20145 15745
rect 20155 15705 20195 15745
rect 20205 15705 20245 15745
rect 20255 15705 20295 15745
rect 20305 15705 20345 15745
rect 20355 15705 20395 15745
rect 20405 15705 20445 15745
rect 20455 15705 20495 15745
rect 20505 15705 20545 15745
rect 20555 15705 20595 15745
rect 20605 15705 20645 15745
rect 20655 15705 20695 15745
rect 20705 15705 20745 15745
rect 20755 15705 20795 15745
rect 20805 15705 20845 15745
rect 20855 15705 20895 15745
rect 20905 15705 20945 15745
rect 20955 15705 20995 15745
rect 21005 15705 21045 15745
rect 21055 15705 21095 15745
rect 21105 15705 21145 15745
rect 21155 15705 21195 15745
rect 21205 15705 21245 15745
rect 21255 15705 21295 15745
rect 21305 15705 21345 15745
rect 21355 15705 21395 15745
rect 21405 15705 21445 15745
rect 21455 15705 21495 15745
rect 21505 15705 21545 15745
rect 21555 15705 21595 15745
rect 21605 15705 21645 15745
rect 21655 15705 21695 15745
rect 21705 15705 21745 15745
rect 21755 15705 21795 15745
rect 21805 15705 21845 15745
rect 21855 15705 21895 15745
rect 21905 15705 21945 15745
rect 21955 15705 21995 15745
rect 22005 15705 22045 15745
rect 22055 15705 22095 15745
rect 22105 15705 22145 15745
rect 22155 15705 22195 15745
rect 22205 15705 22245 15745
rect 22255 15705 22295 15745
rect 22305 15705 22345 15745
rect 22355 15705 22395 15745
rect 22405 15705 22445 15745
rect 22455 15705 22495 15745
rect 22505 15705 22545 15745
rect 22555 15705 22595 15745
rect 22605 15705 22645 15745
rect 22655 15705 22695 15745
rect 22705 15705 22745 15745
rect 22755 15705 22795 15745
rect 22805 15705 22845 15745
rect 22855 15705 22895 15745
rect 22905 15705 22945 15745
rect 22955 15705 22995 15745
rect 23005 15705 23045 15745
rect 23055 15705 23095 15745
rect 23105 15705 23145 15745
rect 23155 15705 23195 15745
rect 23205 15705 23245 15745
rect 23255 15705 23295 15745
rect 23305 15705 23345 15745
rect 23355 15705 23395 15745
rect 23405 15705 23445 15745
rect 23455 15705 23495 15745
rect 23505 15705 23545 15745
rect 23555 15705 23595 15745
rect 23605 15705 23645 15745
rect 23655 15705 23695 15745
rect 23705 15705 23745 15745
rect 23755 15705 23795 15745
rect 23805 15705 23845 15745
rect 23855 15705 23895 15745
rect 23905 15705 23945 15745
rect 23955 15705 23995 15745
rect 24005 15705 24045 15745
rect 24055 15705 24095 15745
rect 24105 15705 24145 15745
rect 24155 15705 24195 15745
rect 24205 15705 24245 15745
rect 24255 15705 24295 15745
rect 24305 15705 24345 15745
rect 24355 15705 24395 15745
rect 24405 15705 24445 15745
rect 24455 15705 24495 15745
rect 24505 15705 24545 15745
rect 24555 15705 24595 15745
rect 24605 15705 24645 15745
rect 24655 15705 24695 15745
rect 24705 15705 24745 15745
rect 24755 15705 24795 15745
rect 24805 15705 24845 15745
rect 24855 15705 24895 15745
rect 24905 15705 24945 15745
rect 24955 15705 24995 15745
rect 25005 15705 25045 15745
rect 25055 15705 25095 15745
rect 25105 15705 25145 15745
rect 25155 15705 25195 15745
rect 25205 15705 25245 15745
rect 25255 15705 25295 15745
rect 25305 15705 25345 15745
rect 25355 15705 25395 15745
rect 25405 15705 25445 15745
rect 25455 15705 25495 15745
rect 25505 15705 25545 15745
rect 25555 15705 25595 15745
rect 25605 15705 25645 15745
rect 25655 15705 25695 15745
rect 25705 15705 25745 15745
rect 25755 15705 25795 15745
rect 25805 15705 25845 15745
rect 25855 15705 25895 15745
rect 25905 15705 25945 15745
rect 25955 15705 25995 15745
rect 26005 15705 26045 15745
rect 26055 15705 26095 15745
rect 26105 15705 26145 15745
rect 26155 15705 26195 15745
rect 26205 15705 26245 15745
rect 26255 15705 26295 15745
rect 26305 15705 26345 15745
rect 26355 15705 26395 15745
rect 26405 15705 26445 15745
rect 26455 15705 26495 15745
rect 26505 15705 26545 15745
rect 26555 15705 26595 15745
rect 26605 15705 26645 15745
rect 26655 15705 26695 15745
rect 26705 15705 26745 15745
rect 26755 15705 26795 15745
rect 26805 15705 26845 15745
rect 26855 15705 26895 15745
rect 26905 15705 26945 15745
rect 26955 15705 26995 15745
rect 27005 15705 27045 15745
rect 27055 15705 27095 15745
rect 27105 15705 27145 15745
rect 27155 15705 27195 15745
rect 27205 15705 27245 15745
rect 27255 15705 27295 15745
rect 27305 15705 27345 15745
rect 27355 15705 27395 15745
rect 27405 15705 27445 15745
rect 27455 15705 27495 15745
rect 27505 15705 27545 15745
rect 27555 15705 27595 15745
rect 27605 15705 27645 15745
rect 27655 15705 27695 15745
rect 27705 15705 27745 15745
rect 27755 15705 27795 15745
rect 27805 15705 27845 15745
rect 27855 15705 27895 15745
rect 27905 15705 27945 15745
rect 27955 15705 27995 15745
rect 28005 15705 28045 15745
rect 28055 15705 28095 15745
rect 28105 15705 28145 15745
rect 28155 15705 28195 15745
rect 28205 15705 28245 15745
rect 28255 15705 28295 15745
rect 28305 15705 28345 15745
rect 28355 15705 28395 15745
rect 28405 15705 28445 15745
rect 28455 15705 28495 15745
rect 28505 15705 28545 15745
rect 28555 15705 28595 15745
rect 28605 15705 28645 15745
rect 28655 15705 28695 15745
rect 28705 15705 28745 15745
rect 28755 15705 28795 15745
rect 28805 15705 28845 15745
rect 28855 15705 28895 15745
rect 28905 15705 28945 15745
rect 28955 15705 28995 15745
rect 29005 15705 29045 15745
rect 29055 15705 29095 15745
rect 29105 15705 29145 15745
rect 29155 15705 29195 15745
rect 29205 15705 29245 15745
rect 29255 15705 29295 15745
rect 29305 15705 29345 15745
rect 29355 15705 29395 15745
rect 29405 15705 29445 15745
rect 29455 15705 29495 15745
rect 29505 15705 29545 15745
rect 29555 15705 29595 15745
rect 29605 15705 29645 15745
rect 29655 15705 29695 15745
rect 29705 15705 29745 15745
rect 29755 15705 29795 15745
rect 29805 15705 29845 15745
rect 29855 15705 29895 15745
rect 29905 15705 29945 15745
rect 29955 15705 29995 15745
rect 30005 15705 30045 15745
rect 30055 15705 30095 15745
rect 30105 15705 30145 15745
rect 30155 15705 30195 15745
rect 30205 15705 30245 15745
rect 30255 15705 30295 15745
rect 30305 15705 30345 15745
rect 30355 15705 30395 15745
rect 30405 15705 30445 15745
rect 30455 15705 30495 15745
rect 30505 15705 30545 15745
rect 30555 15705 30595 15745
rect 30605 15705 30645 15745
rect 30655 15705 30695 15745
rect 30705 15705 30745 15745
rect 30755 15705 30795 15745
rect 30805 15705 30845 15745
rect 30855 15705 30895 15745
rect 30905 15705 30945 15745
rect 30955 15705 30995 15745
rect 31005 15705 31045 15745
rect 31055 15705 31095 15745
rect 31105 15705 31145 15745
rect 31155 15705 31195 15745
rect 31205 15705 31245 15745
rect 31255 15705 31295 15745
rect 31305 15705 31345 15745
rect 31355 15705 31395 15745
rect 31405 15705 31445 15745
rect 31455 15705 31495 15745
rect 31505 15705 31545 15745
rect 31555 15705 31595 15745
rect 31605 15705 31645 15745
rect 31655 15705 31695 15745
rect 31705 15705 31745 15745
rect 31755 15705 31795 15745
rect 31805 15705 31845 15745
rect 31855 15705 31895 15745
rect 31905 15705 31945 15745
rect 31955 15705 31995 15745
rect 32005 15705 32045 15745
rect 32055 15705 32095 15745
rect 32105 15705 32145 15745
rect 32155 15705 32195 15745
rect 32205 15705 32245 15745
rect 32255 15705 32295 15745
rect 32305 15705 32345 15745
rect 32355 15705 32395 15745
rect 32405 15705 32445 15745
rect 32455 15705 32495 15745
rect 32505 15705 32545 15745
rect 32555 15705 32595 15745
rect 32605 15705 32645 15745
rect 32655 15705 32695 15745
rect 32705 15705 32745 15745
rect 32755 15705 32795 15745
rect 32805 15705 32845 15745
rect 32855 15705 32895 15745
rect 32905 15705 32945 15745
rect 32955 15705 32995 15745
rect 33005 15705 33045 15745
rect 33055 15705 33095 15745
rect 33105 15705 33145 15745
rect 33155 15705 33195 15745
rect 33205 15705 33245 15745
rect 33255 15705 33295 15745
rect 33305 15705 33345 15745
rect 33355 15705 33395 15745
rect 33405 15705 33445 15745
rect 33455 15705 33495 15745
rect 33505 15705 33545 15745
rect 33555 15705 33595 15745
rect 33605 15705 33645 15745
rect 33655 15705 33695 15745
rect 33705 15705 33745 15745
rect 33755 15705 33795 15745
rect 33805 15705 33845 15745
rect 33855 15705 33895 15745
rect 33905 15705 33945 15745
rect 33955 15705 33995 15745
rect 34005 15705 34045 15745
rect 34055 15705 34095 15745
rect 34105 15705 34145 15745
rect 34155 15705 34195 15745
rect 34205 15705 34245 15745
rect 34255 15705 34295 15745
rect 34305 15705 34345 15745
rect 34355 15705 34395 15745
rect 34405 15705 34445 15745
rect 34455 15705 34495 15745
rect 34505 15705 34545 15745
rect 34555 15705 34595 15745
rect 34605 15705 34645 15745
rect 34655 15705 34695 15745
rect 34705 15705 34745 15745
rect 34755 15705 34795 15745
rect 34805 15705 34845 15745
rect 34855 15705 34895 15745
rect 34905 15705 34945 15745
rect 34955 15705 34995 15745
rect 35005 15705 35045 15745
rect 35055 15705 35095 15745
rect 35105 15705 35145 15745
rect 35155 15705 35195 15745
rect 35205 15705 35245 15745
rect 35255 15705 35295 15745
rect 35305 15705 35345 15745
rect 35355 15705 35395 15745
rect 35405 15705 35445 15745
rect 35455 15705 35495 15745
rect 35505 15705 35545 15745
rect 35555 15705 35595 15745
rect 35605 15705 35645 15745
rect 35655 15705 35695 15745
rect 35705 15705 35745 15745
rect 35755 15705 35795 15745
rect 35805 15705 35845 15745
rect 35855 15705 35895 15745
rect 35905 15705 35945 15745
rect 35955 15705 35995 15745
rect 36005 15705 36045 15745
rect 36055 15705 36095 15745
rect 36105 15705 36145 15745
rect 36155 15705 36195 15745
rect 36205 15705 36245 15745
rect 36255 15705 36295 15745
rect 36305 15705 36345 15745
rect 36355 15705 36395 15745
rect 36405 15705 36445 15745
rect 36455 15705 36495 15745
rect 36505 15705 36545 15745
rect 36555 15705 36595 15745
rect 36605 15705 36645 15745
rect 36655 15705 36695 15745
rect 36705 15705 36745 15745
rect 36755 15705 36795 15745
rect 36805 15705 36845 15745
rect 36855 15705 36895 15745
rect 36905 15705 36945 15745
rect 36955 15705 36995 15745
rect 37005 15705 37045 15745
rect 37055 15705 37095 15745
rect 37105 15705 37145 15745
rect 37155 15705 37195 15745
rect 37205 15705 37245 15745
rect 37255 15705 37295 15745
rect 37305 15705 37345 15745
rect 37355 15705 37395 15745
rect 37405 15705 37445 15745
rect 37455 15705 37495 15745
rect 37505 15705 37545 15745
rect 37555 15705 37595 15745
rect 37605 15705 37645 15745
rect 37655 15705 37695 15745
rect 37705 15705 37745 15745
rect 37755 15705 37795 15745
rect 37805 15705 37845 15745
rect 37855 15705 37895 15745
rect 37905 15705 37945 15745
rect 37955 15705 37995 15745
rect 38005 15705 38045 15745
rect 38055 15705 38095 15745
rect 38105 15705 38145 15745
rect 38155 15705 38195 15745
rect 38205 15705 38245 15745
rect 38255 15705 38295 15745
rect 38305 15705 38345 15745
rect 38355 15705 38395 15745
rect 38405 15705 38445 15745
rect 38455 15705 38495 15745
rect 38505 15705 38545 15745
rect 38555 15705 38595 15745
rect 38605 15705 38645 15745
rect 38655 15705 38695 15745
rect 38705 15705 38745 15745
rect 38755 15705 38795 15745
rect 38805 15705 38845 15745
rect 38855 15705 38895 15745
rect 38905 15705 38945 15745
rect 38955 15705 38995 15745
rect 39005 15705 39045 15745
rect 39055 15705 39095 15745
rect 39105 15705 39145 15745
rect 39155 15705 39195 15745
rect 39205 15705 39245 15745
rect 39255 15705 39295 15745
rect 39305 15705 39345 15745
rect 39355 15705 39395 15745
rect 39405 15705 39445 15745
rect 39455 15705 39495 15745
rect 39505 15705 39545 15745
rect 39555 15705 39595 15745
rect 39605 15705 39645 15745
rect 39655 15705 39695 15745
rect 39705 15705 39745 15745
rect 39905 15705 39945 15745
rect 39955 15705 39995 15745
rect 40005 15705 40045 15745
rect 40055 15705 40095 15745
rect 40105 15705 40145 15745
rect 40155 15705 40195 15745
rect 40205 15705 40245 15745
rect 40255 15705 40295 15745
rect 40305 15705 40345 15745
rect 40355 15705 40395 15745
rect 40405 15705 40445 15745
rect 40455 15705 40495 15745
rect 40505 15705 40545 15745
rect 40555 15705 40595 15745
rect 40605 15705 40645 15745
rect 40655 15705 40695 15745
rect 40705 15705 40745 15745
rect 40755 15705 40795 15745
rect 40805 15705 40845 15745
rect 40855 15705 40895 15745
rect -3495 15340 -3455 15345
rect -3495 15310 -3490 15340
rect -3490 15310 -3460 15340
rect -3460 15310 -3455 15340
rect -3495 15305 -3455 15310
rect -3295 15340 -3255 15345
rect -3295 15310 -3290 15340
rect -3290 15310 -3260 15340
rect -3260 15310 -3255 15340
rect -3295 15305 -3255 15310
rect -3095 15340 -3055 15345
rect -3095 15310 -3090 15340
rect -3090 15310 -3060 15340
rect -3060 15310 -3055 15340
rect -3095 15305 -3055 15310
rect -1595 15340 -1555 15345
rect -1595 15310 -1590 15340
rect -1590 15310 -1560 15340
rect -1560 15310 -1555 15340
rect -1595 15305 -1555 15310
rect -1095 15340 -1055 15345
rect -1095 15310 -1090 15340
rect -1090 15310 -1060 15340
rect -1060 15310 -1055 15340
rect -1095 15305 -1055 15310
rect -895 15340 -855 15345
rect -895 15310 -890 15340
rect -890 15310 -860 15340
rect -860 15310 -855 15340
rect -895 15305 -855 15310
rect -695 15340 -655 15345
rect -695 15310 -690 15340
rect -690 15310 -660 15340
rect -660 15310 -655 15340
rect -695 15305 -655 15310
rect -495 15340 -455 15345
rect -495 15310 -490 15340
rect -490 15310 -460 15340
rect -460 15310 -455 15340
rect -495 15305 -455 15310
rect -295 15340 -255 15345
rect -295 15310 -290 15340
rect -290 15310 -260 15340
rect -260 15310 -255 15340
rect -295 15305 -255 15310
rect -95 15340 -55 15345
rect -95 15310 -90 15340
rect -90 15310 -60 15340
rect -60 15310 -55 15340
rect -95 15305 -55 15310
rect -3495 15290 -3455 15295
rect -3495 15260 -3490 15290
rect -3490 15260 -3460 15290
rect -3460 15260 -3455 15290
rect -3495 15255 -3455 15260
rect -3295 15290 -3255 15295
rect -3295 15260 -3290 15290
rect -3290 15260 -3260 15290
rect -3260 15260 -3255 15290
rect -3295 15255 -3255 15260
rect -3095 15290 -3055 15295
rect -3095 15260 -3090 15290
rect -3090 15260 -3060 15290
rect -3060 15260 -3055 15290
rect -3095 15255 -3055 15260
rect -1595 15290 -1555 15295
rect -1595 15260 -1590 15290
rect -1590 15260 -1560 15290
rect -1560 15260 -1555 15290
rect -1595 15255 -1555 15260
rect -1095 15290 -1055 15295
rect -1095 15260 -1090 15290
rect -1090 15260 -1060 15290
rect -1060 15260 -1055 15290
rect -1095 15255 -1055 15260
rect -895 15290 -855 15295
rect -895 15260 -890 15290
rect -890 15260 -860 15290
rect -860 15260 -855 15290
rect -895 15255 -855 15260
rect -695 15290 -655 15295
rect -695 15260 -690 15290
rect -690 15260 -660 15290
rect -660 15260 -655 15290
rect -695 15255 -655 15260
rect -495 15290 -455 15295
rect -495 15260 -490 15290
rect -490 15260 -460 15290
rect -460 15260 -455 15290
rect -495 15255 -455 15260
rect -295 15290 -255 15295
rect -295 15260 -290 15290
rect -290 15260 -260 15290
rect -260 15260 -255 15290
rect -295 15255 -255 15260
rect -95 15290 -55 15295
rect -95 15260 -90 15290
rect -90 15260 -60 15290
rect -60 15260 -55 15290
rect -95 15255 -55 15260
rect -3495 15240 -3455 15245
rect -3495 15210 -3490 15240
rect -3490 15210 -3460 15240
rect -3460 15210 -3455 15240
rect -3495 15205 -3455 15210
rect -3295 15240 -3255 15245
rect -3295 15210 -3290 15240
rect -3290 15210 -3260 15240
rect -3260 15210 -3255 15240
rect -3295 15205 -3255 15210
rect -3095 15240 -3055 15245
rect -3095 15210 -3090 15240
rect -3090 15210 -3060 15240
rect -3060 15210 -3055 15240
rect -3095 15205 -3055 15210
rect -1595 15240 -1555 15245
rect -1595 15210 -1590 15240
rect -1590 15210 -1560 15240
rect -1560 15210 -1555 15240
rect -1595 15205 -1555 15210
rect -1095 15240 -1055 15245
rect -1095 15210 -1090 15240
rect -1090 15210 -1060 15240
rect -1060 15210 -1055 15240
rect -1095 15205 -1055 15210
rect -895 15240 -855 15245
rect -895 15210 -890 15240
rect -890 15210 -860 15240
rect -860 15210 -855 15240
rect -895 15205 -855 15210
rect -695 15240 -655 15245
rect -695 15210 -690 15240
rect -690 15210 -660 15240
rect -660 15210 -655 15240
rect -695 15205 -655 15210
rect -495 15240 -455 15245
rect -495 15210 -490 15240
rect -490 15210 -460 15240
rect -460 15210 -455 15240
rect -495 15205 -455 15210
rect -295 15240 -255 15245
rect -295 15210 -290 15240
rect -290 15210 -260 15240
rect -260 15210 -255 15240
rect -295 15205 -255 15210
rect -95 15240 -55 15245
rect -95 15210 -90 15240
rect -90 15210 -60 15240
rect -60 15210 -55 15240
rect -95 15205 -55 15210
rect -195 14605 -155 14645
rect -395 14205 -355 14245
rect -595 14005 -555 14045
rect -3495 13640 -3455 13645
rect -3495 13610 -3490 13640
rect -3490 13610 -3460 13640
rect -3460 13610 -3455 13640
rect -3495 13605 -3455 13610
rect -3295 13640 -3255 13645
rect -3295 13610 -3290 13640
rect -3290 13610 -3260 13640
rect -3260 13610 -3255 13640
rect -3295 13605 -3255 13610
rect -3095 13640 -3055 13645
rect -3095 13610 -3090 13640
rect -3090 13610 -3060 13640
rect -3060 13610 -3055 13640
rect -3095 13605 -3055 13610
rect -1595 13640 -1555 13645
rect -1595 13610 -1590 13640
rect -1590 13610 -1560 13640
rect -1560 13610 -1555 13640
rect -1595 13605 -1555 13610
rect -1095 13640 -1055 13645
rect -1095 13610 -1090 13640
rect -1090 13610 -1060 13640
rect -1060 13610 -1055 13640
rect -1095 13605 -1055 13610
rect -895 13640 -855 13645
rect -895 13610 -890 13640
rect -890 13610 -860 13640
rect -860 13610 -855 13640
rect -895 13605 -855 13610
rect -695 13640 -655 13645
rect -695 13610 -690 13640
rect -690 13610 -660 13640
rect -660 13610 -655 13640
rect -695 13605 -655 13610
rect -495 13640 -455 13645
rect -495 13610 -490 13640
rect -490 13610 -460 13640
rect -460 13610 -455 13640
rect -495 13605 -455 13610
rect -295 13640 -255 13645
rect -295 13610 -290 13640
rect -290 13610 -260 13640
rect -260 13610 -255 13640
rect -295 13605 -255 13610
rect -95 13640 -55 13645
rect -95 13610 -90 13640
rect -90 13610 -60 13640
rect -60 13610 -55 13640
rect -95 13605 -55 13610
rect -3495 13590 -3455 13595
rect -3495 13560 -3490 13590
rect -3490 13560 -3460 13590
rect -3460 13560 -3455 13590
rect -3495 13555 -3455 13560
rect -3295 13590 -3255 13595
rect -3295 13560 -3290 13590
rect -3290 13560 -3260 13590
rect -3260 13560 -3255 13590
rect -3295 13555 -3255 13560
rect -3095 13590 -3055 13595
rect -3095 13560 -3090 13590
rect -3090 13560 -3060 13590
rect -3060 13560 -3055 13590
rect -3095 13555 -3055 13560
rect -1595 13590 -1555 13595
rect -1595 13560 -1590 13590
rect -1590 13560 -1560 13590
rect -1560 13560 -1555 13590
rect -1595 13555 -1555 13560
rect -1095 13590 -1055 13595
rect -1095 13560 -1090 13590
rect -1090 13560 -1060 13590
rect -1060 13560 -1055 13590
rect -1095 13555 -1055 13560
rect -895 13590 -855 13595
rect -895 13560 -890 13590
rect -890 13560 -860 13590
rect -860 13560 -855 13590
rect -895 13555 -855 13560
rect -695 13590 -655 13595
rect -695 13560 -690 13590
rect -690 13560 -660 13590
rect -660 13560 -655 13590
rect -695 13555 -655 13560
rect -495 13590 -455 13595
rect -495 13560 -490 13590
rect -490 13560 -460 13590
rect -460 13560 -455 13590
rect -495 13555 -455 13560
rect -295 13590 -255 13595
rect -295 13560 -290 13590
rect -290 13560 -260 13590
rect -260 13560 -255 13590
rect -295 13555 -255 13560
rect -95 13590 -55 13595
rect -95 13560 -90 13590
rect -90 13560 -60 13590
rect -60 13560 -55 13590
rect -95 13555 -55 13560
rect -3495 13540 -3455 13545
rect -3495 13510 -3490 13540
rect -3490 13510 -3460 13540
rect -3460 13510 -3455 13540
rect -3495 13505 -3455 13510
rect -3295 13540 -3255 13545
rect -3295 13510 -3290 13540
rect -3290 13510 -3260 13540
rect -3260 13510 -3255 13540
rect -3295 13505 -3255 13510
rect -3095 13540 -3055 13545
rect -3095 13510 -3090 13540
rect -3090 13510 -3060 13540
rect -3060 13510 -3055 13540
rect -3095 13505 -3055 13510
rect -1595 13540 -1555 13545
rect -1595 13510 -1590 13540
rect -1590 13510 -1560 13540
rect -1560 13510 -1555 13540
rect -1595 13505 -1555 13510
rect -1095 13540 -1055 13545
rect -1095 13510 -1090 13540
rect -1090 13510 -1060 13540
rect -1060 13510 -1055 13540
rect -1095 13505 -1055 13510
rect -895 13540 -855 13545
rect -895 13510 -890 13540
rect -890 13510 -860 13540
rect -860 13510 -855 13540
rect -895 13505 -855 13510
rect -695 13540 -655 13545
rect -695 13510 -690 13540
rect -690 13510 -660 13540
rect -660 13510 -655 13540
rect -695 13505 -655 13510
rect -495 13540 -455 13545
rect -495 13510 -490 13540
rect -490 13510 -460 13540
rect -460 13510 -455 13540
rect -495 13505 -455 13510
rect -295 13540 -255 13545
rect -295 13510 -290 13540
rect -290 13510 -260 13540
rect -260 13510 -255 13540
rect -295 13505 -255 13510
rect -95 13540 -55 13545
rect -95 13510 -90 13540
rect -90 13510 -60 13540
rect -60 13510 -55 13540
rect -95 13505 -55 13510
rect -795 13105 -755 13145
rect -995 12905 -955 12945
rect -1195 12505 -1155 12545
rect -1295 12405 -1255 12445
rect -1395 12305 -1355 12345
rect -1495 12205 -1455 12245
rect -3495 11940 -3455 11945
rect -3495 11910 -3490 11940
rect -3490 11910 -3460 11940
rect -3460 11910 -3455 11940
rect -3495 11905 -3455 11910
rect -3295 11940 -3255 11945
rect -3295 11910 -3290 11940
rect -3290 11910 -3260 11940
rect -3260 11910 -3255 11940
rect -3295 11905 -3255 11910
rect -3095 11940 -3055 11945
rect -3095 11910 -3090 11940
rect -3090 11910 -3060 11940
rect -3060 11910 -3055 11940
rect -3095 11905 -3055 11910
rect -1595 11940 -1555 11945
rect -1595 11910 -1590 11940
rect -1590 11910 -1560 11940
rect -1560 11910 -1555 11940
rect -1595 11905 -1555 11910
rect -1095 11940 -1055 11945
rect -1095 11910 -1090 11940
rect -1090 11910 -1060 11940
rect -1060 11910 -1055 11940
rect -1095 11905 -1055 11910
rect -895 11940 -855 11945
rect -895 11910 -890 11940
rect -890 11910 -860 11940
rect -860 11910 -855 11940
rect -895 11905 -855 11910
rect -695 11940 -655 11945
rect -695 11910 -690 11940
rect -690 11910 -660 11940
rect -660 11910 -655 11940
rect -695 11905 -655 11910
rect -495 11940 -455 11945
rect -495 11910 -490 11940
rect -490 11910 -460 11940
rect -460 11910 -455 11940
rect -495 11905 -455 11910
rect -295 11940 -255 11945
rect -295 11910 -290 11940
rect -290 11910 -260 11940
rect -260 11910 -255 11940
rect -295 11905 -255 11910
rect -95 11940 -55 11945
rect -95 11910 -90 11940
rect -90 11910 -60 11940
rect -60 11910 -55 11940
rect -95 11905 -55 11910
rect -3495 11890 -3455 11895
rect -3495 11860 -3490 11890
rect -3490 11860 -3460 11890
rect -3460 11860 -3455 11890
rect -3495 11855 -3455 11860
rect -3295 11890 -3255 11895
rect -3295 11860 -3290 11890
rect -3290 11860 -3260 11890
rect -3260 11860 -3255 11890
rect -3295 11855 -3255 11860
rect -3095 11890 -3055 11895
rect -3095 11860 -3090 11890
rect -3090 11860 -3060 11890
rect -3060 11860 -3055 11890
rect -3095 11855 -3055 11860
rect -1595 11890 -1555 11895
rect -1595 11860 -1590 11890
rect -1590 11860 -1560 11890
rect -1560 11860 -1555 11890
rect -1595 11855 -1555 11860
rect -1095 11890 -1055 11895
rect -1095 11860 -1090 11890
rect -1090 11860 -1060 11890
rect -1060 11860 -1055 11890
rect -1095 11855 -1055 11860
rect -895 11890 -855 11895
rect -895 11860 -890 11890
rect -890 11860 -860 11890
rect -860 11860 -855 11890
rect -895 11855 -855 11860
rect -695 11890 -655 11895
rect -695 11860 -690 11890
rect -690 11860 -660 11890
rect -660 11860 -655 11890
rect -695 11855 -655 11860
rect -495 11890 -455 11895
rect -495 11860 -490 11890
rect -490 11860 -460 11890
rect -460 11860 -455 11890
rect -495 11855 -455 11860
rect -295 11890 -255 11895
rect -295 11860 -290 11890
rect -290 11860 -260 11890
rect -260 11860 -255 11890
rect -295 11855 -255 11860
rect -95 11890 -55 11895
rect -95 11860 -90 11890
rect -90 11860 -60 11890
rect -60 11860 -55 11890
rect -95 11855 -55 11860
rect -3495 11840 -3455 11845
rect -3495 11810 -3490 11840
rect -3490 11810 -3460 11840
rect -3460 11810 -3455 11840
rect -3495 11805 -3455 11810
rect -3295 11840 -3255 11845
rect -3295 11810 -3290 11840
rect -3290 11810 -3260 11840
rect -3260 11810 -3255 11840
rect -3295 11805 -3255 11810
rect -3095 11840 -3055 11845
rect -3095 11810 -3090 11840
rect -3090 11810 -3060 11840
rect -3060 11810 -3055 11840
rect -3095 11805 -3055 11810
rect -1595 11840 -1555 11845
rect -1595 11810 -1590 11840
rect -1590 11810 -1560 11840
rect -1560 11810 -1555 11840
rect -1595 11805 -1555 11810
rect -1095 11840 -1055 11845
rect -1095 11810 -1090 11840
rect -1090 11810 -1060 11840
rect -1060 11810 -1055 11840
rect -1095 11805 -1055 11810
rect -895 11840 -855 11845
rect -895 11810 -890 11840
rect -890 11810 -860 11840
rect -860 11810 -855 11840
rect -895 11805 -855 11810
rect -695 11840 -655 11845
rect -695 11810 -690 11840
rect -690 11810 -660 11840
rect -660 11810 -655 11840
rect -695 11805 -655 11810
rect -495 11840 -455 11845
rect -495 11810 -490 11840
rect -490 11810 -460 11840
rect -460 11810 -455 11840
rect -495 11805 -455 11810
rect -295 11840 -255 11845
rect -295 11810 -290 11840
rect -290 11810 -260 11840
rect -260 11810 -255 11840
rect -295 11805 -255 11810
rect -95 11840 -55 11845
rect -95 11810 -90 11840
rect -90 11810 -60 11840
rect -60 11810 -55 11840
rect -95 11805 -55 11810
rect -3195 11405 -3155 11445
rect 39805 11340 39845 11345
rect 39805 11310 39810 11340
rect 39810 11310 39840 11340
rect 39840 11310 39845 11340
rect 39805 11305 39845 11310
rect 39905 11240 39945 11245
rect 39905 11210 39910 11240
rect 39910 11210 39940 11240
rect 39940 11210 39945 11240
rect 39905 11205 39945 11210
rect 39955 11240 39995 11245
rect 39955 11210 39960 11240
rect 39960 11210 39990 11240
rect 39990 11210 39995 11240
rect 39955 11205 39995 11210
rect 40005 11240 40045 11245
rect 40005 11210 40010 11240
rect 40010 11210 40040 11240
rect 40040 11210 40045 11240
rect 40005 11205 40045 11210
rect 40055 11240 40095 11245
rect 40055 11210 40060 11240
rect 40060 11210 40090 11240
rect 40090 11210 40095 11240
rect 40055 11205 40095 11210
rect 40105 11240 40145 11245
rect 40105 11210 40110 11240
rect 40110 11210 40140 11240
rect 40140 11210 40145 11240
rect 40105 11205 40145 11210
rect 40155 11240 40195 11245
rect 40155 11210 40160 11240
rect 40160 11210 40190 11240
rect 40190 11210 40195 11240
rect 40155 11205 40195 11210
rect 40205 11240 40245 11245
rect 40205 11210 40210 11240
rect 40210 11210 40240 11240
rect 40240 11210 40245 11240
rect 40205 11205 40245 11210
rect 40255 11240 40295 11245
rect 40255 11210 40260 11240
rect 40260 11210 40290 11240
rect 40290 11210 40295 11240
rect 40255 11205 40295 11210
rect 40305 11240 40345 11245
rect 40305 11210 40310 11240
rect 40310 11210 40340 11240
rect 40340 11210 40345 11240
rect 40305 11205 40345 11210
rect 40355 11240 40395 11245
rect 40355 11210 40360 11240
rect 40360 11210 40390 11240
rect 40390 11210 40395 11240
rect 40355 11205 40395 11210
rect 40405 11240 40445 11245
rect 40405 11210 40410 11240
rect 40410 11210 40440 11240
rect 40440 11210 40445 11240
rect 40405 11205 40445 11210
rect 40455 11240 40495 11245
rect 40455 11210 40460 11240
rect 40460 11210 40490 11240
rect 40490 11210 40495 11240
rect 40455 11205 40495 11210
rect 40505 11240 40545 11245
rect 40505 11210 40510 11240
rect 40510 11210 40540 11240
rect 40540 11210 40545 11240
rect 40505 11205 40545 11210
rect 40555 11240 40595 11245
rect 40555 11210 40560 11240
rect 40560 11210 40590 11240
rect 40590 11210 40595 11240
rect 40555 11205 40595 11210
rect 40605 11240 40645 11245
rect 40605 11210 40610 11240
rect 40610 11210 40640 11240
rect 40640 11210 40645 11240
rect 40605 11205 40645 11210
rect 40655 11240 40695 11245
rect 40655 11210 40660 11240
rect 40660 11210 40690 11240
rect 40690 11210 40695 11240
rect 40655 11205 40695 11210
rect 40705 11240 40745 11245
rect 40705 11210 40710 11240
rect 40710 11210 40740 11240
rect 40740 11210 40745 11240
rect 40705 11205 40745 11210
rect 40755 11240 40795 11245
rect 40755 11210 40760 11240
rect 40760 11210 40790 11240
rect 40790 11210 40795 11240
rect 40755 11205 40795 11210
rect 40805 11240 40845 11245
rect 40805 11210 40810 11240
rect 40810 11210 40840 11240
rect 40840 11210 40845 11240
rect 40805 11205 40845 11210
rect 40855 11240 40895 11245
rect 40855 11210 40860 11240
rect 40860 11210 40890 11240
rect 40890 11210 40895 11240
rect 40855 11205 40895 11210
rect 39905 11190 39945 11195
rect 39905 11160 39910 11190
rect 39910 11160 39940 11190
rect 39940 11160 39945 11190
rect 39905 11155 39945 11160
rect 39955 11190 39995 11195
rect 39955 11160 39960 11190
rect 39960 11160 39990 11190
rect 39990 11160 39995 11190
rect 39955 11155 39995 11160
rect 40005 11190 40045 11195
rect 40005 11160 40010 11190
rect 40010 11160 40040 11190
rect 40040 11160 40045 11190
rect 40005 11155 40045 11160
rect 40055 11190 40095 11195
rect 40055 11160 40060 11190
rect 40060 11160 40090 11190
rect 40090 11160 40095 11190
rect 40055 11155 40095 11160
rect 40105 11190 40145 11195
rect 40105 11160 40110 11190
rect 40110 11160 40140 11190
rect 40140 11160 40145 11190
rect 40105 11155 40145 11160
rect 40155 11190 40195 11195
rect 40155 11160 40160 11190
rect 40160 11160 40190 11190
rect 40190 11160 40195 11190
rect 40155 11155 40195 11160
rect 40205 11190 40245 11195
rect 40205 11160 40210 11190
rect 40210 11160 40240 11190
rect 40240 11160 40245 11190
rect 40205 11155 40245 11160
rect 40255 11190 40295 11195
rect 40255 11160 40260 11190
rect 40260 11160 40290 11190
rect 40290 11160 40295 11190
rect 40255 11155 40295 11160
rect 40305 11190 40345 11195
rect 40305 11160 40310 11190
rect 40310 11160 40340 11190
rect 40340 11160 40345 11190
rect 40305 11155 40345 11160
rect 40355 11190 40395 11195
rect 40355 11160 40360 11190
rect 40360 11160 40390 11190
rect 40390 11160 40395 11190
rect 40355 11155 40395 11160
rect 40405 11190 40445 11195
rect 40405 11160 40410 11190
rect 40410 11160 40440 11190
rect 40440 11160 40445 11190
rect 40405 11155 40445 11160
rect 40455 11190 40495 11195
rect 40455 11160 40460 11190
rect 40460 11160 40490 11190
rect 40490 11160 40495 11190
rect 40455 11155 40495 11160
rect 40505 11190 40545 11195
rect 40505 11160 40510 11190
rect 40510 11160 40540 11190
rect 40540 11160 40545 11190
rect 40505 11155 40545 11160
rect 40555 11190 40595 11195
rect 40555 11160 40560 11190
rect 40560 11160 40590 11190
rect 40590 11160 40595 11190
rect 40555 11155 40595 11160
rect 40605 11190 40645 11195
rect 40605 11160 40610 11190
rect 40610 11160 40640 11190
rect 40640 11160 40645 11190
rect 40605 11155 40645 11160
rect 40655 11190 40695 11195
rect 40655 11160 40660 11190
rect 40660 11160 40690 11190
rect 40690 11160 40695 11190
rect 40655 11155 40695 11160
rect 40705 11190 40745 11195
rect 40705 11160 40710 11190
rect 40710 11160 40740 11190
rect 40740 11160 40745 11190
rect 40705 11155 40745 11160
rect 40755 11190 40795 11195
rect 40755 11160 40760 11190
rect 40760 11160 40790 11190
rect 40790 11160 40795 11190
rect 40755 11155 40795 11160
rect 40805 11190 40845 11195
rect 40805 11160 40810 11190
rect 40810 11160 40840 11190
rect 40840 11160 40845 11190
rect 40805 11155 40845 11160
rect 40855 11190 40895 11195
rect 40855 11160 40860 11190
rect 40860 11160 40890 11190
rect 40890 11160 40895 11190
rect 40855 11155 40895 11160
rect 39905 11140 39945 11145
rect 39905 11110 39910 11140
rect 39910 11110 39940 11140
rect 39940 11110 39945 11140
rect 39905 11105 39945 11110
rect 39955 11140 39995 11145
rect 39955 11110 39960 11140
rect 39960 11110 39990 11140
rect 39990 11110 39995 11140
rect 39955 11105 39995 11110
rect 40005 11140 40045 11145
rect 40005 11110 40010 11140
rect 40010 11110 40040 11140
rect 40040 11110 40045 11140
rect 40005 11105 40045 11110
rect 40055 11140 40095 11145
rect 40055 11110 40060 11140
rect 40060 11110 40090 11140
rect 40090 11110 40095 11140
rect 40055 11105 40095 11110
rect 40105 11140 40145 11145
rect 40105 11110 40110 11140
rect 40110 11110 40140 11140
rect 40140 11110 40145 11140
rect 40105 11105 40145 11110
rect 40155 11140 40195 11145
rect 40155 11110 40160 11140
rect 40160 11110 40190 11140
rect 40190 11110 40195 11140
rect 40155 11105 40195 11110
rect 40205 11140 40245 11145
rect 40205 11110 40210 11140
rect 40210 11110 40240 11140
rect 40240 11110 40245 11140
rect 40205 11105 40245 11110
rect 40255 11140 40295 11145
rect 40255 11110 40260 11140
rect 40260 11110 40290 11140
rect 40290 11110 40295 11140
rect 40255 11105 40295 11110
rect 40305 11140 40345 11145
rect 40305 11110 40310 11140
rect 40310 11110 40340 11140
rect 40340 11110 40345 11140
rect 40305 11105 40345 11110
rect 40355 11140 40395 11145
rect 40355 11110 40360 11140
rect 40360 11110 40390 11140
rect 40390 11110 40395 11140
rect 40355 11105 40395 11110
rect 40405 11140 40445 11145
rect 40405 11110 40410 11140
rect 40410 11110 40440 11140
rect 40440 11110 40445 11140
rect 40405 11105 40445 11110
rect 40455 11140 40495 11145
rect 40455 11110 40460 11140
rect 40460 11110 40490 11140
rect 40490 11110 40495 11140
rect 40455 11105 40495 11110
rect 40505 11140 40545 11145
rect 40505 11110 40510 11140
rect 40510 11110 40540 11140
rect 40540 11110 40545 11140
rect 40505 11105 40545 11110
rect 40555 11140 40595 11145
rect 40555 11110 40560 11140
rect 40560 11110 40590 11140
rect 40590 11110 40595 11140
rect 40555 11105 40595 11110
rect 40605 11140 40645 11145
rect 40605 11110 40610 11140
rect 40610 11110 40640 11140
rect 40640 11110 40645 11140
rect 40605 11105 40645 11110
rect 40655 11140 40695 11145
rect 40655 11110 40660 11140
rect 40660 11110 40690 11140
rect 40690 11110 40695 11140
rect 40655 11105 40695 11110
rect 40705 11140 40745 11145
rect 40705 11110 40710 11140
rect 40710 11110 40740 11140
rect 40740 11110 40745 11140
rect 40705 11105 40745 11110
rect 40755 11140 40795 11145
rect 40755 11110 40760 11140
rect 40760 11110 40790 11140
rect 40790 11110 40795 11140
rect 40755 11105 40795 11110
rect 40805 11140 40845 11145
rect 40805 11110 40810 11140
rect 40810 11110 40840 11140
rect 40840 11110 40845 11140
rect 40805 11105 40845 11110
rect 40855 11140 40895 11145
rect 40855 11110 40860 11140
rect 40860 11110 40890 11140
rect 40890 11110 40895 11140
rect 40855 11105 40895 11110
rect 39905 11090 39945 11095
rect 39905 11060 39910 11090
rect 39910 11060 39940 11090
rect 39940 11060 39945 11090
rect 39905 11055 39945 11060
rect 39955 11090 39995 11095
rect 39955 11060 39960 11090
rect 39960 11060 39990 11090
rect 39990 11060 39995 11090
rect 39955 11055 39995 11060
rect 40005 11090 40045 11095
rect 40005 11060 40010 11090
rect 40010 11060 40040 11090
rect 40040 11060 40045 11090
rect 40005 11055 40045 11060
rect 40055 11090 40095 11095
rect 40055 11060 40060 11090
rect 40060 11060 40090 11090
rect 40090 11060 40095 11090
rect 40055 11055 40095 11060
rect 40105 11090 40145 11095
rect 40105 11060 40110 11090
rect 40110 11060 40140 11090
rect 40140 11060 40145 11090
rect 40105 11055 40145 11060
rect 40155 11090 40195 11095
rect 40155 11060 40160 11090
rect 40160 11060 40190 11090
rect 40190 11060 40195 11090
rect 40155 11055 40195 11060
rect 40205 11090 40245 11095
rect 40205 11060 40210 11090
rect 40210 11060 40240 11090
rect 40240 11060 40245 11090
rect 40205 11055 40245 11060
rect 40255 11090 40295 11095
rect 40255 11060 40260 11090
rect 40260 11060 40290 11090
rect 40290 11060 40295 11090
rect 40255 11055 40295 11060
rect 40305 11090 40345 11095
rect 40305 11060 40310 11090
rect 40310 11060 40340 11090
rect 40340 11060 40345 11090
rect 40305 11055 40345 11060
rect 40355 11090 40395 11095
rect 40355 11060 40360 11090
rect 40360 11060 40390 11090
rect 40390 11060 40395 11090
rect 40355 11055 40395 11060
rect 40405 11090 40445 11095
rect 40405 11060 40410 11090
rect 40410 11060 40440 11090
rect 40440 11060 40445 11090
rect 40405 11055 40445 11060
rect 40455 11090 40495 11095
rect 40455 11060 40460 11090
rect 40460 11060 40490 11090
rect 40490 11060 40495 11090
rect 40455 11055 40495 11060
rect 40505 11090 40545 11095
rect 40505 11060 40510 11090
rect 40510 11060 40540 11090
rect 40540 11060 40545 11090
rect 40505 11055 40545 11060
rect 40555 11090 40595 11095
rect 40555 11060 40560 11090
rect 40560 11060 40590 11090
rect 40590 11060 40595 11090
rect 40555 11055 40595 11060
rect 40605 11090 40645 11095
rect 40605 11060 40610 11090
rect 40610 11060 40640 11090
rect 40640 11060 40645 11090
rect 40605 11055 40645 11060
rect 40655 11090 40695 11095
rect 40655 11060 40660 11090
rect 40660 11060 40690 11090
rect 40690 11060 40695 11090
rect 40655 11055 40695 11060
rect 40705 11090 40745 11095
rect 40705 11060 40710 11090
rect 40710 11060 40740 11090
rect 40740 11060 40745 11090
rect 40705 11055 40745 11060
rect 40755 11090 40795 11095
rect 40755 11060 40760 11090
rect 40760 11060 40790 11090
rect 40790 11060 40795 11090
rect 40755 11055 40795 11060
rect 40805 11090 40845 11095
rect 40805 11060 40810 11090
rect 40810 11060 40840 11090
rect 40840 11060 40845 11090
rect 40805 11055 40845 11060
rect 40855 11090 40895 11095
rect 40855 11060 40860 11090
rect 40860 11060 40890 11090
rect 40890 11060 40895 11090
rect 40855 11055 40895 11060
rect 39905 11040 39945 11045
rect 39905 11010 39910 11040
rect 39910 11010 39940 11040
rect 39940 11010 39945 11040
rect 39905 11005 39945 11010
rect 39955 11040 39995 11045
rect 39955 11010 39960 11040
rect 39960 11010 39990 11040
rect 39990 11010 39995 11040
rect 39955 11005 39995 11010
rect 40005 11040 40045 11045
rect 40005 11010 40010 11040
rect 40010 11010 40040 11040
rect 40040 11010 40045 11040
rect 40005 11005 40045 11010
rect 40055 11040 40095 11045
rect 40055 11010 40060 11040
rect 40060 11010 40090 11040
rect 40090 11010 40095 11040
rect 40055 11005 40095 11010
rect 40105 11040 40145 11045
rect 40105 11010 40110 11040
rect 40110 11010 40140 11040
rect 40140 11010 40145 11040
rect 40105 11005 40145 11010
rect 40155 11040 40195 11045
rect 40155 11010 40160 11040
rect 40160 11010 40190 11040
rect 40190 11010 40195 11040
rect 40155 11005 40195 11010
rect 40205 11040 40245 11045
rect 40205 11010 40210 11040
rect 40210 11010 40240 11040
rect 40240 11010 40245 11040
rect 40205 11005 40245 11010
rect 40255 11040 40295 11045
rect 40255 11010 40260 11040
rect 40260 11010 40290 11040
rect 40290 11010 40295 11040
rect 40255 11005 40295 11010
rect 40305 11040 40345 11045
rect 40305 11010 40310 11040
rect 40310 11010 40340 11040
rect 40340 11010 40345 11040
rect 40305 11005 40345 11010
rect 40355 11040 40395 11045
rect 40355 11010 40360 11040
rect 40360 11010 40390 11040
rect 40390 11010 40395 11040
rect 40355 11005 40395 11010
rect 40405 11040 40445 11045
rect 40405 11010 40410 11040
rect 40410 11010 40440 11040
rect 40440 11010 40445 11040
rect 40405 11005 40445 11010
rect 40455 11040 40495 11045
rect 40455 11010 40460 11040
rect 40460 11010 40490 11040
rect 40490 11010 40495 11040
rect 40455 11005 40495 11010
rect 40505 11040 40545 11045
rect 40505 11010 40510 11040
rect 40510 11010 40540 11040
rect 40540 11010 40545 11040
rect 40505 11005 40545 11010
rect 40555 11040 40595 11045
rect 40555 11010 40560 11040
rect 40560 11010 40590 11040
rect 40590 11010 40595 11040
rect 40555 11005 40595 11010
rect 40605 11040 40645 11045
rect 40605 11010 40610 11040
rect 40610 11010 40640 11040
rect 40640 11010 40645 11040
rect 40605 11005 40645 11010
rect 40655 11040 40695 11045
rect 40655 11010 40660 11040
rect 40660 11010 40690 11040
rect 40690 11010 40695 11040
rect 40655 11005 40695 11010
rect 40705 11040 40745 11045
rect 40705 11010 40710 11040
rect 40710 11010 40740 11040
rect 40740 11010 40745 11040
rect 40705 11005 40745 11010
rect 40755 11040 40795 11045
rect 40755 11010 40760 11040
rect 40760 11010 40790 11040
rect 40790 11010 40795 11040
rect 40755 11005 40795 11010
rect 40805 11040 40845 11045
rect 40805 11010 40810 11040
rect 40810 11010 40840 11040
rect 40840 11010 40845 11040
rect 40805 11005 40845 11010
rect 40855 11040 40895 11045
rect 40855 11010 40860 11040
rect 40860 11010 40890 11040
rect 40890 11010 40895 11040
rect 40855 11005 40895 11010
rect 39805 10940 39845 10945
rect 39805 10910 39810 10940
rect 39810 10910 39840 10940
rect 39840 10910 39845 10940
rect 39805 10905 39845 10910
rect -3395 10805 -3355 10845
rect -2995 10640 -2955 10645
rect -2995 10610 -2990 10640
rect -2990 10610 -2960 10640
rect -2960 10610 -2955 10640
rect -2995 10605 -2955 10610
rect -2795 10640 -2755 10645
rect -2795 10610 -2790 10640
rect -2790 10610 -2760 10640
rect -2760 10610 -2755 10640
rect -2795 10605 -2755 10610
rect -2595 10640 -2555 10645
rect -2595 10610 -2590 10640
rect -2590 10610 -2560 10640
rect -2560 10610 -2555 10640
rect -2595 10605 -2555 10610
rect -2395 10640 -2355 10645
rect -2395 10610 -2390 10640
rect -2390 10610 -2360 10640
rect -2360 10610 -2355 10640
rect -2395 10605 -2355 10610
rect -2195 10640 -2155 10645
rect -2195 10610 -2190 10640
rect -2190 10610 -2160 10640
rect -2160 10610 -2155 10640
rect -2195 10605 -2155 10610
rect -1995 10640 -1955 10645
rect -1995 10610 -1990 10640
rect -1990 10610 -1960 10640
rect -1960 10610 -1955 10640
rect -1995 10605 -1955 10610
rect -1695 10640 -1655 10645
rect -1695 10610 -1690 10640
rect -1690 10610 -1660 10640
rect -1660 10610 -1655 10640
rect -1695 10605 -1655 10610
rect -2995 10590 -2955 10595
rect -2995 10560 -2990 10590
rect -2990 10560 -2960 10590
rect -2960 10560 -2955 10590
rect -2995 10555 -2955 10560
rect -2795 10590 -2755 10595
rect -2795 10560 -2790 10590
rect -2790 10560 -2760 10590
rect -2760 10560 -2755 10590
rect -2795 10555 -2755 10560
rect -2595 10590 -2555 10595
rect -2595 10560 -2590 10590
rect -2590 10560 -2560 10590
rect -2560 10560 -2555 10590
rect -2595 10555 -2555 10560
rect -2395 10590 -2355 10595
rect -2395 10560 -2390 10590
rect -2390 10560 -2360 10590
rect -2360 10560 -2355 10590
rect -2395 10555 -2355 10560
rect -2195 10590 -2155 10595
rect -2195 10560 -2190 10590
rect -2190 10560 -2160 10590
rect -2160 10560 -2155 10590
rect -2195 10555 -2155 10560
rect -1995 10590 -1955 10595
rect -1995 10560 -1990 10590
rect -1990 10560 -1960 10590
rect -1960 10560 -1955 10590
rect -1995 10555 -1955 10560
rect -1695 10590 -1655 10595
rect -1695 10560 -1690 10590
rect -1690 10560 -1660 10590
rect -1660 10560 -1655 10590
rect -1695 10555 -1655 10560
rect -2995 10540 -2955 10545
rect -2995 10510 -2990 10540
rect -2990 10510 -2960 10540
rect -2960 10510 -2955 10540
rect -2995 10505 -2955 10510
rect -2795 10540 -2755 10545
rect -2795 10510 -2790 10540
rect -2790 10510 -2760 10540
rect -2760 10510 -2755 10540
rect -2795 10505 -2755 10510
rect -2595 10540 -2555 10545
rect -2595 10510 -2590 10540
rect -2590 10510 -2560 10540
rect -2560 10510 -2555 10540
rect -2595 10505 -2555 10510
rect -2395 10540 -2355 10545
rect -2395 10510 -2390 10540
rect -2390 10510 -2360 10540
rect -2360 10510 -2355 10540
rect -2395 10505 -2355 10510
rect -2195 10540 -2155 10545
rect -2195 10510 -2190 10540
rect -2190 10510 -2160 10540
rect -2160 10510 -2155 10540
rect -2195 10505 -2155 10510
rect -1995 10540 -1955 10545
rect -1995 10510 -1990 10540
rect -1990 10510 -1960 10540
rect -1960 10510 -1955 10540
rect -1995 10505 -1955 10510
rect -1695 10540 -1655 10545
rect -1695 10510 -1690 10540
rect -1690 10510 -1660 10540
rect -1660 10510 -1655 10540
rect -1695 10505 -1655 10510
rect -1795 10205 -1755 10245
rect -1895 10105 -1855 10145
rect -2095 9705 -2055 9745
rect -2295 9505 -2255 9545
rect -2995 9340 -2955 9345
rect -2995 9310 -2990 9340
rect -2990 9310 -2960 9340
rect -2960 9310 -2955 9340
rect -2995 9305 -2955 9310
rect -2795 9340 -2755 9345
rect -2795 9310 -2790 9340
rect -2790 9310 -2760 9340
rect -2760 9310 -2755 9340
rect -2795 9305 -2755 9310
rect -2595 9340 -2555 9345
rect -2595 9310 -2590 9340
rect -2590 9310 -2560 9340
rect -2560 9310 -2555 9340
rect -2595 9305 -2555 9310
rect -2395 9340 -2355 9345
rect -2395 9310 -2390 9340
rect -2390 9310 -2360 9340
rect -2360 9310 -2355 9340
rect -2395 9305 -2355 9310
rect -2195 9340 -2155 9345
rect -2195 9310 -2190 9340
rect -2190 9310 -2160 9340
rect -2160 9310 -2155 9340
rect -2195 9305 -2155 9310
rect -1995 9340 -1955 9345
rect -1995 9310 -1990 9340
rect -1990 9310 -1960 9340
rect -1960 9310 -1955 9340
rect -1995 9305 -1955 9310
rect -1695 9340 -1655 9345
rect -1695 9310 -1690 9340
rect -1690 9310 -1660 9340
rect -1660 9310 -1655 9340
rect -1695 9305 -1655 9310
rect -2995 9290 -2955 9295
rect -2995 9260 -2990 9290
rect -2990 9260 -2960 9290
rect -2960 9260 -2955 9290
rect -2995 9255 -2955 9260
rect -2795 9290 -2755 9295
rect -2795 9260 -2790 9290
rect -2790 9260 -2760 9290
rect -2760 9260 -2755 9290
rect -2795 9255 -2755 9260
rect -2595 9290 -2555 9295
rect -2595 9260 -2590 9290
rect -2590 9260 -2560 9290
rect -2560 9260 -2555 9290
rect -2595 9255 -2555 9260
rect -2395 9290 -2355 9295
rect -2395 9260 -2390 9290
rect -2390 9260 -2360 9290
rect -2360 9260 -2355 9290
rect -2395 9255 -2355 9260
rect -2195 9290 -2155 9295
rect -2195 9260 -2190 9290
rect -2190 9260 -2160 9290
rect -2160 9260 -2155 9290
rect -2195 9255 -2155 9260
rect -1995 9290 -1955 9295
rect -1995 9260 -1990 9290
rect -1990 9260 -1960 9290
rect -1960 9260 -1955 9290
rect -1995 9255 -1955 9260
rect -1695 9290 -1655 9295
rect -1695 9260 -1690 9290
rect -1690 9260 -1660 9290
rect -1660 9260 -1655 9290
rect -1695 9255 -1655 9260
rect -2995 9240 -2955 9245
rect -2995 9210 -2990 9240
rect -2990 9210 -2960 9240
rect -2960 9210 -2955 9240
rect -2995 9205 -2955 9210
rect -2795 9240 -2755 9245
rect -2795 9210 -2790 9240
rect -2790 9210 -2760 9240
rect -2760 9210 -2755 9240
rect -2795 9205 -2755 9210
rect -2595 9240 -2555 9245
rect -2595 9210 -2590 9240
rect -2590 9210 -2560 9240
rect -2560 9210 -2555 9240
rect -2595 9205 -2555 9210
rect -2395 9240 -2355 9245
rect -2395 9210 -2390 9240
rect -2390 9210 -2360 9240
rect -2360 9210 -2355 9240
rect -2395 9205 -2355 9210
rect -2195 9240 -2155 9245
rect -2195 9210 -2190 9240
rect -2190 9210 -2160 9240
rect -2160 9210 -2155 9240
rect -2195 9205 -2155 9210
rect -1995 9240 -1955 9245
rect -1995 9210 -1990 9240
rect -1990 9210 -1960 9240
rect -1960 9210 -1955 9240
rect -1995 9205 -1955 9210
rect -1695 9240 -1655 9245
rect -1695 9210 -1690 9240
rect -1690 9210 -1660 9240
rect -1660 9210 -1655 9240
rect -1695 9205 -1655 9210
rect -2495 9005 -2455 9045
rect -2695 8805 -2655 8845
rect -2895 8405 -2855 8445
rect -2995 8040 -2955 8045
rect -2995 8010 -2990 8040
rect -2990 8010 -2960 8040
rect -2960 8010 -2955 8040
rect -2995 8005 -2955 8010
rect -2795 8040 -2755 8045
rect -2795 8010 -2790 8040
rect -2790 8010 -2760 8040
rect -2760 8010 -2755 8040
rect -2795 8005 -2755 8010
rect -2595 8040 -2555 8045
rect -2595 8010 -2590 8040
rect -2590 8010 -2560 8040
rect -2560 8010 -2555 8040
rect -2595 8005 -2555 8010
rect -2395 8040 -2355 8045
rect -2395 8010 -2390 8040
rect -2390 8010 -2360 8040
rect -2360 8010 -2355 8040
rect -2395 8005 -2355 8010
rect -2195 8040 -2155 8045
rect -2195 8010 -2190 8040
rect -2190 8010 -2160 8040
rect -2160 8010 -2155 8040
rect -2195 8005 -2155 8010
rect -1995 8040 -1955 8045
rect -1995 8010 -1990 8040
rect -1990 8010 -1960 8040
rect -1960 8010 -1955 8040
rect -1995 8005 -1955 8010
rect -1695 8040 -1655 8045
rect -1695 8010 -1690 8040
rect -1690 8010 -1660 8040
rect -1660 8010 -1655 8040
rect -1695 8005 -1655 8010
rect -2995 7990 -2955 7995
rect -2995 7960 -2990 7990
rect -2990 7960 -2960 7990
rect -2960 7960 -2955 7990
rect -2995 7955 -2955 7960
rect -2795 7990 -2755 7995
rect -2795 7960 -2790 7990
rect -2790 7960 -2760 7990
rect -2760 7960 -2755 7990
rect -2795 7955 -2755 7960
rect -2595 7990 -2555 7995
rect -2595 7960 -2590 7990
rect -2590 7960 -2560 7990
rect -2560 7960 -2555 7990
rect -2595 7955 -2555 7960
rect -2395 7990 -2355 7995
rect -2395 7960 -2390 7990
rect -2390 7960 -2360 7990
rect -2360 7960 -2355 7990
rect -2395 7955 -2355 7960
rect -2195 7990 -2155 7995
rect -2195 7960 -2190 7990
rect -2190 7960 -2160 7990
rect -2160 7960 -2155 7990
rect -2195 7955 -2155 7960
rect -1995 7990 -1955 7995
rect -1995 7960 -1990 7990
rect -1990 7960 -1960 7990
rect -1960 7960 -1955 7990
rect -1995 7955 -1955 7960
rect -1695 7990 -1655 7995
rect -1695 7960 -1690 7990
rect -1690 7960 -1660 7990
rect -1660 7960 -1655 7990
rect -1695 7955 -1655 7960
rect -2995 7940 -2955 7945
rect -2995 7910 -2990 7940
rect -2990 7910 -2960 7940
rect -2960 7910 -2955 7940
rect -2995 7905 -2955 7910
rect -2795 7940 -2755 7945
rect -2795 7910 -2790 7940
rect -2790 7910 -2760 7940
rect -2760 7910 -2755 7940
rect -2795 7905 -2755 7910
rect -2595 7940 -2555 7945
rect -2595 7910 -2590 7940
rect -2590 7910 -2560 7940
rect -2560 7910 -2555 7940
rect -2595 7905 -2555 7910
rect -2395 7940 -2355 7945
rect -2395 7910 -2390 7940
rect -2390 7910 -2360 7940
rect -2360 7910 -2355 7940
rect -2395 7905 -2355 7910
rect -2195 7940 -2155 7945
rect -2195 7910 -2190 7940
rect -2190 7910 -2160 7940
rect -2160 7910 -2155 7940
rect -2195 7905 -2155 7910
rect -1995 7940 -1955 7945
rect -1995 7910 -1990 7940
rect -1990 7910 -1960 7940
rect -1960 7910 -1955 7940
rect -1995 7905 -1955 7910
rect -1695 7940 -1655 7945
rect -1695 7910 -1690 7940
rect -1690 7910 -1660 7940
rect -1660 7910 -1655 7940
rect -1695 7905 -1655 7910
rect -2995 7740 -2955 7745
rect -2995 7710 -2990 7740
rect -2990 7710 -2960 7740
rect -2960 7710 -2955 7740
rect -2995 7705 -2955 7710
rect -2795 7740 -2755 7745
rect -2795 7710 -2790 7740
rect -2790 7710 -2760 7740
rect -2760 7710 -2755 7740
rect -2795 7705 -2755 7710
rect -2595 7740 -2555 7745
rect -2595 7710 -2590 7740
rect -2590 7710 -2560 7740
rect -2560 7710 -2555 7740
rect -2595 7705 -2555 7710
rect -2395 7740 -2355 7745
rect -2395 7710 -2390 7740
rect -2390 7710 -2360 7740
rect -2360 7710 -2355 7740
rect -2395 7705 -2355 7710
rect -2195 7740 -2155 7745
rect -2195 7710 -2190 7740
rect -2190 7710 -2160 7740
rect -2160 7710 -2155 7740
rect -2195 7705 -2155 7710
rect -1995 7740 -1955 7745
rect -1995 7710 -1990 7740
rect -1990 7710 -1960 7740
rect -1960 7710 -1955 7740
rect -1995 7705 -1955 7710
rect -1695 7740 -1655 7745
rect -1695 7710 -1690 7740
rect -1690 7710 -1660 7740
rect -1660 7710 -1655 7740
rect -1695 7705 -1655 7710
rect -2995 7690 -2955 7695
rect -2995 7660 -2990 7690
rect -2990 7660 -2960 7690
rect -2960 7660 -2955 7690
rect -2995 7655 -2955 7660
rect -2795 7690 -2755 7695
rect -2795 7660 -2790 7690
rect -2790 7660 -2760 7690
rect -2760 7660 -2755 7690
rect -2795 7655 -2755 7660
rect -2595 7690 -2555 7695
rect -2595 7660 -2590 7690
rect -2590 7660 -2560 7690
rect -2560 7660 -2555 7690
rect -2595 7655 -2555 7660
rect -2395 7690 -2355 7695
rect -2395 7660 -2390 7690
rect -2390 7660 -2360 7690
rect -2360 7660 -2355 7690
rect -2395 7655 -2355 7660
rect -2195 7690 -2155 7695
rect -2195 7660 -2190 7690
rect -2190 7660 -2160 7690
rect -2160 7660 -2155 7690
rect -2195 7655 -2155 7660
rect -1995 7690 -1955 7695
rect -1995 7660 -1990 7690
rect -1990 7660 -1960 7690
rect -1960 7660 -1955 7690
rect -1995 7655 -1955 7660
rect -1695 7690 -1655 7695
rect -1695 7660 -1690 7690
rect -1690 7660 -1660 7690
rect -1660 7660 -1655 7690
rect -1695 7655 -1655 7660
rect -2995 7640 -2955 7645
rect -2995 7610 -2990 7640
rect -2990 7610 -2960 7640
rect -2960 7610 -2955 7640
rect -2995 7605 -2955 7610
rect -2795 7640 -2755 7645
rect -2795 7610 -2790 7640
rect -2790 7610 -2760 7640
rect -2760 7610 -2755 7640
rect -2795 7605 -2755 7610
rect -2595 7640 -2555 7645
rect -2595 7610 -2590 7640
rect -2590 7610 -2560 7640
rect -2560 7610 -2555 7640
rect -2595 7605 -2555 7610
rect -2395 7640 -2355 7645
rect -2395 7610 -2390 7640
rect -2390 7610 -2360 7640
rect -2360 7610 -2355 7640
rect -2395 7605 -2355 7610
rect -2195 7640 -2155 7645
rect -2195 7610 -2190 7640
rect -2190 7610 -2160 7640
rect -2160 7610 -2155 7640
rect -2195 7605 -2155 7610
rect -1995 7640 -1955 7645
rect -1995 7610 -1990 7640
rect -1990 7610 -1960 7640
rect -1960 7610 -1955 7640
rect -1995 7605 -1955 7610
rect -1695 7640 -1655 7645
rect -1695 7610 -1690 7640
rect -1690 7610 -1660 7640
rect -1660 7610 -1655 7640
rect -1695 7605 -1655 7610
rect -2895 7205 -2855 7245
rect -2695 6805 -2655 6845
rect -2495 6605 -2455 6645
rect -2995 6440 -2955 6445
rect -2995 6410 -2990 6440
rect -2990 6410 -2960 6440
rect -2960 6410 -2955 6440
rect -2995 6405 -2955 6410
rect -2795 6440 -2755 6445
rect -2795 6410 -2790 6440
rect -2790 6410 -2760 6440
rect -2760 6410 -2755 6440
rect -2795 6405 -2755 6410
rect -2595 6440 -2555 6445
rect -2595 6410 -2590 6440
rect -2590 6410 -2560 6440
rect -2560 6410 -2555 6440
rect -2595 6405 -2555 6410
rect -2395 6440 -2355 6445
rect -2395 6410 -2390 6440
rect -2390 6410 -2360 6440
rect -2360 6410 -2355 6440
rect -2395 6405 -2355 6410
rect -2195 6440 -2155 6445
rect -2195 6410 -2190 6440
rect -2190 6410 -2160 6440
rect -2160 6410 -2155 6440
rect -2195 6405 -2155 6410
rect -1995 6440 -1955 6445
rect -1995 6410 -1990 6440
rect -1990 6410 -1960 6440
rect -1960 6410 -1955 6440
rect -1995 6405 -1955 6410
rect -1695 6440 -1655 6445
rect -1695 6410 -1690 6440
rect -1690 6410 -1660 6440
rect -1660 6410 -1655 6440
rect -1695 6405 -1655 6410
rect -2995 6390 -2955 6395
rect -2995 6360 -2990 6390
rect -2990 6360 -2960 6390
rect -2960 6360 -2955 6390
rect -2995 6355 -2955 6360
rect -2795 6390 -2755 6395
rect -2795 6360 -2790 6390
rect -2790 6360 -2760 6390
rect -2760 6360 -2755 6390
rect -2795 6355 -2755 6360
rect -2595 6390 -2555 6395
rect -2595 6360 -2590 6390
rect -2590 6360 -2560 6390
rect -2560 6360 -2555 6390
rect -2595 6355 -2555 6360
rect -2395 6390 -2355 6395
rect -2395 6360 -2390 6390
rect -2390 6360 -2360 6390
rect -2360 6360 -2355 6390
rect -2395 6355 -2355 6360
rect -2195 6390 -2155 6395
rect -2195 6360 -2190 6390
rect -2190 6360 -2160 6390
rect -2160 6360 -2155 6390
rect -2195 6355 -2155 6360
rect -1995 6390 -1955 6395
rect -1995 6360 -1990 6390
rect -1990 6360 -1960 6390
rect -1960 6360 -1955 6390
rect -1995 6355 -1955 6360
rect -1695 6390 -1655 6395
rect -1695 6360 -1690 6390
rect -1690 6360 -1660 6390
rect -1660 6360 -1655 6390
rect -1695 6355 -1655 6360
rect -2995 6340 -2955 6345
rect -2995 6310 -2990 6340
rect -2990 6310 -2960 6340
rect -2960 6310 -2955 6340
rect -2995 6305 -2955 6310
rect -2795 6340 -2755 6345
rect -2795 6310 -2790 6340
rect -2790 6310 -2760 6340
rect -2760 6310 -2755 6340
rect -2795 6305 -2755 6310
rect -2595 6340 -2555 6345
rect -2595 6310 -2590 6340
rect -2590 6310 -2560 6340
rect -2560 6310 -2555 6340
rect -2595 6305 -2555 6310
rect -2395 6340 -2355 6345
rect -2395 6310 -2390 6340
rect -2390 6310 -2360 6340
rect -2360 6310 -2355 6340
rect -2395 6305 -2355 6310
rect -2195 6340 -2155 6345
rect -2195 6310 -2190 6340
rect -2190 6310 -2160 6340
rect -2160 6310 -2155 6340
rect -2195 6305 -2155 6310
rect -1995 6340 -1955 6345
rect -1995 6310 -1990 6340
rect -1990 6310 -1960 6340
rect -1960 6310 -1955 6340
rect -1995 6305 -1955 6310
rect -1695 6340 -1655 6345
rect -1695 6310 -1690 6340
rect -1690 6310 -1660 6340
rect -1660 6310 -1655 6340
rect -1695 6305 -1655 6310
rect -2295 6105 -2255 6145
rect -2095 5905 -2055 5945
rect -1895 5505 -1855 5545
rect -1795 5405 -1755 5445
rect -2995 5140 -2955 5145
rect -2995 5110 -2990 5140
rect -2990 5110 -2960 5140
rect -2960 5110 -2955 5140
rect -2995 5105 -2955 5110
rect -2795 5140 -2755 5145
rect -2795 5110 -2790 5140
rect -2790 5110 -2760 5140
rect -2760 5110 -2755 5140
rect -2795 5105 -2755 5110
rect -2595 5140 -2555 5145
rect -2595 5110 -2590 5140
rect -2590 5110 -2560 5140
rect -2560 5110 -2555 5140
rect -2595 5105 -2555 5110
rect -2395 5140 -2355 5145
rect -2395 5110 -2390 5140
rect -2390 5110 -2360 5140
rect -2360 5110 -2355 5140
rect -2395 5105 -2355 5110
rect -2195 5140 -2155 5145
rect -2195 5110 -2190 5140
rect -2190 5110 -2160 5140
rect -2160 5110 -2155 5140
rect -2195 5105 -2155 5110
rect -1995 5140 -1955 5145
rect -1995 5110 -1990 5140
rect -1990 5110 -1960 5140
rect -1960 5110 -1955 5140
rect -1995 5105 -1955 5110
rect -1695 5140 -1655 5145
rect -1695 5110 -1690 5140
rect -1690 5110 -1660 5140
rect -1660 5110 -1655 5140
rect -1695 5105 -1655 5110
rect -2995 5090 -2955 5095
rect -2995 5060 -2990 5090
rect -2990 5060 -2960 5090
rect -2960 5060 -2955 5090
rect -2995 5055 -2955 5060
rect -2795 5090 -2755 5095
rect -2795 5060 -2790 5090
rect -2790 5060 -2760 5090
rect -2760 5060 -2755 5090
rect -2795 5055 -2755 5060
rect -2595 5090 -2555 5095
rect -2595 5060 -2590 5090
rect -2590 5060 -2560 5090
rect -2560 5060 -2555 5090
rect -2595 5055 -2555 5060
rect -2395 5090 -2355 5095
rect -2395 5060 -2390 5090
rect -2390 5060 -2360 5090
rect -2360 5060 -2355 5090
rect -2395 5055 -2355 5060
rect -2195 5090 -2155 5095
rect -2195 5060 -2190 5090
rect -2190 5060 -2160 5090
rect -2160 5060 -2155 5090
rect -2195 5055 -2155 5060
rect -1995 5090 -1955 5095
rect -1995 5060 -1990 5090
rect -1990 5060 -1960 5090
rect -1960 5060 -1955 5090
rect -1995 5055 -1955 5060
rect -1695 5090 -1655 5095
rect -1695 5060 -1690 5090
rect -1690 5060 -1660 5090
rect -1660 5060 -1655 5090
rect -1695 5055 -1655 5060
rect -2995 5040 -2955 5045
rect -2995 5010 -2990 5040
rect -2990 5010 -2960 5040
rect -2960 5010 -2955 5040
rect -2995 5005 -2955 5010
rect -2795 5040 -2755 5045
rect -2795 5010 -2790 5040
rect -2790 5010 -2760 5040
rect -2760 5010 -2755 5040
rect -2795 5005 -2755 5010
rect -2595 5040 -2555 5045
rect -2595 5010 -2590 5040
rect -2590 5010 -2560 5040
rect -2560 5010 -2555 5040
rect -2595 5005 -2555 5010
rect -2395 5040 -2355 5045
rect -2395 5010 -2390 5040
rect -2390 5010 -2360 5040
rect -2360 5010 -2355 5040
rect -2395 5005 -2355 5010
rect -2195 5040 -2155 5045
rect -2195 5010 -2190 5040
rect -2190 5010 -2160 5040
rect -2160 5010 -2155 5040
rect -2195 5005 -2155 5010
rect -1995 5040 -1955 5045
rect -1995 5010 -1990 5040
rect -1990 5010 -1960 5040
rect -1960 5010 -1955 5040
rect -1995 5005 -1955 5010
rect -1695 5040 -1655 5045
rect -1695 5010 -1690 5040
rect -1690 5010 -1660 5040
rect -1660 5010 -1655 5040
rect -1695 5005 -1655 5010
rect -3395 4805 -3355 4845
rect 39805 4740 39845 4745
rect 39805 4710 39810 4740
rect 39810 4710 39840 4740
rect 39840 4710 39845 4740
rect 39805 4705 39845 4710
rect 39905 4640 39945 4645
rect 39905 4610 39910 4640
rect 39910 4610 39940 4640
rect 39940 4610 39945 4640
rect 39905 4605 39945 4610
rect 39955 4640 39995 4645
rect 39955 4610 39960 4640
rect 39960 4610 39990 4640
rect 39990 4610 39995 4640
rect 39955 4605 39995 4610
rect 40005 4640 40045 4645
rect 40005 4610 40010 4640
rect 40010 4610 40040 4640
rect 40040 4610 40045 4640
rect 40005 4605 40045 4610
rect 40055 4640 40095 4645
rect 40055 4610 40060 4640
rect 40060 4610 40090 4640
rect 40090 4610 40095 4640
rect 40055 4605 40095 4610
rect 40105 4640 40145 4645
rect 40105 4610 40110 4640
rect 40110 4610 40140 4640
rect 40140 4610 40145 4640
rect 40105 4605 40145 4610
rect 40155 4640 40195 4645
rect 40155 4610 40160 4640
rect 40160 4610 40190 4640
rect 40190 4610 40195 4640
rect 40155 4605 40195 4610
rect 40205 4640 40245 4645
rect 40205 4610 40210 4640
rect 40210 4610 40240 4640
rect 40240 4610 40245 4640
rect 40205 4605 40245 4610
rect 40255 4640 40295 4645
rect 40255 4610 40260 4640
rect 40260 4610 40290 4640
rect 40290 4610 40295 4640
rect 40255 4605 40295 4610
rect 40305 4640 40345 4645
rect 40305 4610 40310 4640
rect 40310 4610 40340 4640
rect 40340 4610 40345 4640
rect 40305 4605 40345 4610
rect 40355 4640 40395 4645
rect 40355 4610 40360 4640
rect 40360 4610 40390 4640
rect 40390 4610 40395 4640
rect 40355 4605 40395 4610
rect 40405 4640 40445 4645
rect 40405 4610 40410 4640
rect 40410 4610 40440 4640
rect 40440 4610 40445 4640
rect 40405 4605 40445 4610
rect 40455 4640 40495 4645
rect 40455 4610 40460 4640
rect 40460 4610 40490 4640
rect 40490 4610 40495 4640
rect 40455 4605 40495 4610
rect 40505 4640 40545 4645
rect 40505 4610 40510 4640
rect 40510 4610 40540 4640
rect 40540 4610 40545 4640
rect 40505 4605 40545 4610
rect 40555 4640 40595 4645
rect 40555 4610 40560 4640
rect 40560 4610 40590 4640
rect 40590 4610 40595 4640
rect 40555 4605 40595 4610
rect 40605 4640 40645 4645
rect 40605 4610 40610 4640
rect 40610 4610 40640 4640
rect 40640 4610 40645 4640
rect 40605 4605 40645 4610
rect 40655 4640 40695 4645
rect 40655 4610 40660 4640
rect 40660 4610 40690 4640
rect 40690 4610 40695 4640
rect 40655 4605 40695 4610
rect 40705 4640 40745 4645
rect 40705 4610 40710 4640
rect 40710 4610 40740 4640
rect 40740 4610 40745 4640
rect 40705 4605 40745 4610
rect 40755 4640 40795 4645
rect 40755 4610 40760 4640
rect 40760 4610 40790 4640
rect 40790 4610 40795 4640
rect 40755 4605 40795 4610
rect 40805 4640 40845 4645
rect 40805 4610 40810 4640
rect 40810 4610 40840 4640
rect 40840 4610 40845 4640
rect 40805 4605 40845 4610
rect 40855 4640 40895 4645
rect 40855 4610 40860 4640
rect 40860 4610 40890 4640
rect 40890 4610 40895 4640
rect 40855 4605 40895 4610
rect 39905 4590 39945 4595
rect 39905 4560 39910 4590
rect 39910 4560 39940 4590
rect 39940 4560 39945 4590
rect 39905 4555 39945 4560
rect 39955 4590 39995 4595
rect 39955 4560 39960 4590
rect 39960 4560 39990 4590
rect 39990 4560 39995 4590
rect 39955 4555 39995 4560
rect 40005 4590 40045 4595
rect 40005 4560 40010 4590
rect 40010 4560 40040 4590
rect 40040 4560 40045 4590
rect 40005 4555 40045 4560
rect 40055 4590 40095 4595
rect 40055 4560 40060 4590
rect 40060 4560 40090 4590
rect 40090 4560 40095 4590
rect 40055 4555 40095 4560
rect 40105 4590 40145 4595
rect 40105 4560 40110 4590
rect 40110 4560 40140 4590
rect 40140 4560 40145 4590
rect 40105 4555 40145 4560
rect 40155 4590 40195 4595
rect 40155 4560 40160 4590
rect 40160 4560 40190 4590
rect 40190 4560 40195 4590
rect 40155 4555 40195 4560
rect 40205 4590 40245 4595
rect 40205 4560 40210 4590
rect 40210 4560 40240 4590
rect 40240 4560 40245 4590
rect 40205 4555 40245 4560
rect 40255 4590 40295 4595
rect 40255 4560 40260 4590
rect 40260 4560 40290 4590
rect 40290 4560 40295 4590
rect 40255 4555 40295 4560
rect 40305 4590 40345 4595
rect 40305 4560 40310 4590
rect 40310 4560 40340 4590
rect 40340 4560 40345 4590
rect 40305 4555 40345 4560
rect 40355 4590 40395 4595
rect 40355 4560 40360 4590
rect 40360 4560 40390 4590
rect 40390 4560 40395 4590
rect 40355 4555 40395 4560
rect 40405 4590 40445 4595
rect 40405 4560 40410 4590
rect 40410 4560 40440 4590
rect 40440 4560 40445 4590
rect 40405 4555 40445 4560
rect 40455 4590 40495 4595
rect 40455 4560 40460 4590
rect 40460 4560 40490 4590
rect 40490 4560 40495 4590
rect 40455 4555 40495 4560
rect 40505 4590 40545 4595
rect 40505 4560 40510 4590
rect 40510 4560 40540 4590
rect 40540 4560 40545 4590
rect 40505 4555 40545 4560
rect 40555 4590 40595 4595
rect 40555 4560 40560 4590
rect 40560 4560 40590 4590
rect 40590 4560 40595 4590
rect 40555 4555 40595 4560
rect 40605 4590 40645 4595
rect 40605 4560 40610 4590
rect 40610 4560 40640 4590
rect 40640 4560 40645 4590
rect 40605 4555 40645 4560
rect 40655 4590 40695 4595
rect 40655 4560 40660 4590
rect 40660 4560 40690 4590
rect 40690 4560 40695 4590
rect 40655 4555 40695 4560
rect 40705 4590 40745 4595
rect 40705 4560 40710 4590
rect 40710 4560 40740 4590
rect 40740 4560 40745 4590
rect 40705 4555 40745 4560
rect 40755 4590 40795 4595
rect 40755 4560 40760 4590
rect 40760 4560 40790 4590
rect 40790 4560 40795 4590
rect 40755 4555 40795 4560
rect 40805 4590 40845 4595
rect 40805 4560 40810 4590
rect 40810 4560 40840 4590
rect 40840 4560 40845 4590
rect 40805 4555 40845 4560
rect 40855 4590 40895 4595
rect 40855 4560 40860 4590
rect 40860 4560 40890 4590
rect 40890 4560 40895 4590
rect 40855 4555 40895 4560
rect 39905 4540 39945 4545
rect 39905 4510 39910 4540
rect 39910 4510 39940 4540
rect 39940 4510 39945 4540
rect 39905 4505 39945 4510
rect 39955 4540 39995 4545
rect 39955 4510 39960 4540
rect 39960 4510 39990 4540
rect 39990 4510 39995 4540
rect 39955 4505 39995 4510
rect 40005 4540 40045 4545
rect 40005 4510 40010 4540
rect 40010 4510 40040 4540
rect 40040 4510 40045 4540
rect 40005 4505 40045 4510
rect 40055 4540 40095 4545
rect 40055 4510 40060 4540
rect 40060 4510 40090 4540
rect 40090 4510 40095 4540
rect 40055 4505 40095 4510
rect 40105 4540 40145 4545
rect 40105 4510 40110 4540
rect 40110 4510 40140 4540
rect 40140 4510 40145 4540
rect 40105 4505 40145 4510
rect 40155 4540 40195 4545
rect 40155 4510 40160 4540
rect 40160 4510 40190 4540
rect 40190 4510 40195 4540
rect 40155 4505 40195 4510
rect 40205 4540 40245 4545
rect 40205 4510 40210 4540
rect 40210 4510 40240 4540
rect 40240 4510 40245 4540
rect 40205 4505 40245 4510
rect 40255 4540 40295 4545
rect 40255 4510 40260 4540
rect 40260 4510 40290 4540
rect 40290 4510 40295 4540
rect 40255 4505 40295 4510
rect 40305 4540 40345 4545
rect 40305 4510 40310 4540
rect 40310 4510 40340 4540
rect 40340 4510 40345 4540
rect 40305 4505 40345 4510
rect 40355 4540 40395 4545
rect 40355 4510 40360 4540
rect 40360 4510 40390 4540
rect 40390 4510 40395 4540
rect 40355 4505 40395 4510
rect 40405 4540 40445 4545
rect 40405 4510 40410 4540
rect 40410 4510 40440 4540
rect 40440 4510 40445 4540
rect 40405 4505 40445 4510
rect 40455 4540 40495 4545
rect 40455 4510 40460 4540
rect 40460 4510 40490 4540
rect 40490 4510 40495 4540
rect 40455 4505 40495 4510
rect 40505 4540 40545 4545
rect 40505 4510 40510 4540
rect 40510 4510 40540 4540
rect 40540 4510 40545 4540
rect 40505 4505 40545 4510
rect 40555 4540 40595 4545
rect 40555 4510 40560 4540
rect 40560 4510 40590 4540
rect 40590 4510 40595 4540
rect 40555 4505 40595 4510
rect 40605 4540 40645 4545
rect 40605 4510 40610 4540
rect 40610 4510 40640 4540
rect 40640 4510 40645 4540
rect 40605 4505 40645 4510
rect 40655 4540 40695 4545
rect 40655 4510 40660 4540
rect 40660 4510 40690 4540
rect 40690 4510 40695 4540
rect 40655 4505 40695 4510
rect 40705 4540 40745 4545
rect 40705 4510 40710 4540
rect 40710 4510 40740 4540
rect 40740 4510 40745 4540
rect 40705 4505 40745 4510
rect 40755 4540 40795 4545
rect 40755 4510 40760 4540
rect 40760 4510 40790 4540
rect 40790 4510 40795 4540
rect 40755 4505 40795 4510
rect 40805 4540 40845 4545
rect 40805 4510 40810 4540
rect 40810 4510 40840 4540
rect 40840 4510 40845 4540
rect 40805 4505 40845 4510
rect 40855 4540 40895 4545
rect 40855 4510 40860 4540
rect 40860 4510 40890 4540
rect 40890 4510 40895 4540
rect 40855 4505 40895 4510
rect 39905 4490 39945 4495
rect 39905 4460 39910 4490
rect 39910 4460 39940 4490
rect 39940 4460 39945 4490
rect 39905 4455 39945 4460
rect 39955 4490 39995 4495
rect 39955 4460 39960 4490
rect 39960 4460 39990 4490
rect 39990 4460 39995 4490
rect 39955 4455 39995 4460
rect 40005 4490 40045 4495
rect 40005 4460 40010 4490
rect 40010 4460 40040 4490
rect 40040 4460 40045 4490
rect 40005 4455 40045 4460
rect 40055 4490 40095 4495
rect 40055 4460 40060 4490
rect 40060 4460 40090 4490
rect 40090 4460 40095 4490
rect 40055 4455 40095 4460
rect 40105 4490 40145 4495
rect 40105 4460 40110 4490
rect 40110 4460 40140 4490
rect 40140 4460 40145 4490
rect 40105 4455 40145 4460
rect 40155 4490 40195 4495
rect 40155 4460 40160 4490
rect 40160 4460 40190 4490
rect 40190 4460 40195 4490
rect 40155 4455 40195 4460
rect 40205 4490 40245 4495
rect 40205 4460 40210 4490
rect 40210 4460 40240 4490
rect 40240 4460 40245 4490
rect 40205 4455 40245 4460
rect 40255 4490 40295 4495
rect 40255 4460 40260 4490
rect 40260 4460 40290 4490
rect 40290 4460 40295 4490
rect 40255 4455 40295 4460
rect 40305 4490 40345 4495
rect 40305 4460 40310 4490
rect 40310 4460 40340 4490
rect 40340 4460 40345 4490
rect 40305 4455 40345 4460
rect 40355 4490 40395 4495
rect 40355 4460 40360 4490
rect 40360 4460 40390 4490
rect 40390 4460 40395 4490
rect 40355 4455 40395 4460
rect 40405 4490 40445 4495
rect 40405 4460 40410 4490
rect 40410 4460 40440 4490
rect 40440 4460 40445 4490
rect 40405 4455 40445 4460
rect 40455 4490 40495 4495
rect 40455 4460 40460 4490
rect 40460 4460 40490 4490
rect 40490 4460 40495 4490
rect 40455 4455 40495 4460
rect 40505 4490 40545 4495
rect 40505 4460 40510 4490
rect 40510 4460 40540 4490
rect 40540 4460 40545 4490
rect 40505 4455 40545 4460
rect 40555 4490 40595 4495
rect 40555 4460 40560 4490
rect 40560 4460 40590 4490
rect 40590 4460 40595 4490
rect 40555 4455 40595 4460
rect 40605 4490 40645 4495
rect 40605 4460 40610 4490
rect 40610 4460 40640 4490
rect 40640 4460 40645 4490
rect 40605 4455 40645 4460
rect 40655 4490 40695 4495
rect 40655 4460 40660 4490
rect 40660 4460 40690 4490
rect 40690 4460 40695 4490
rect 40655 4455 40695 4460
rect 40705 4490 40745 4495
rect 40705 4460 40710 4490
rect 40710 4460 40740 4490
rect 40740 4460 40745 4490
rect 40705 4455 40745 4460
rect 40755 4490 40795 4495
rect 40755 4460 40760 4490
rect 40760 4460 40790 4490
rect 40790 4460 40795 4490
rect 40755 4455 40795 4460
rect 40805 4490 40845 4495
rect 40805 4460 40810 4490
rect 40810 4460 40840 4490
rect 40840 4460 40845 4490
rect 40805 4455 40845 4460
rect 40855 4490 40895 4495
rect 40855 4460 40860 4490
rect 40860 4460 40890 4490
rect 40890 4460 40895 4490
rect 40855 4455 40895 4460
rect 39905 4440 39945 4445
rect 39905 4410 39910 4440
rect 39910 4410 39940 4440
rect 39940 4410 39945 4440
rect 39905 4405 39945 4410
rect 39955 4440 39995 4445
rect 39955 4410 39960 4440
rect 39960 4410 39990 4440
rect 39990 4410 39995 4440
rect 39955 4405 39995 4410
rect 40005 4440 40045 4445
rect 40005 4410 40010 4440
rect 40010 4410 40040 4440
rect 40040 4410 40045 4440
rect 40005 4405 40045 4410
rect 40055 4440 40095 4445
rect 40055 4410 40060 4440
rect 40060 4410 40090 4440
rect 40090 4410 40095 4440
rect 40055 4405 40095 4410
rect 40105 4440 40145 4445
rect 40105 4410 40110 4440
rect 40110 4410 40140 4440
rect 40140 4410 40145 4440
rect 40105 4405 40145 4410
rect 40155 4440 40195 4445
rect 40155 4410 40160 4440
rect 40160 4410 40190 4440
rect 40190 4410 40195 4440
rect 40155 4405 40195 4410
rect 40205 4440 40245 4445
rect 40205 4410 40210 4440
rect 40210 4410 40240 4440
rect 40240 4410 40245 4440
rect 40205 4405 40245 4410
rect 40255 4440 40295 4445
rect 40255 4410 40260 4440
rect 40260 4410 40290 4440
rect 40290 4410 40295 4440
rect 40255 4405 40295 4410
rect 40305 4440 40345 4445
rect 40305 4410 40310 4440
rect 40310 4410 40340 4440
rect 40340 4410 40345 4440
rect 40305 4405 40345 4410
rect 40355 4440 40395 4445
rect 40355 4410 40360 4440
rect 40360 4410 40390 4440
rect 40390 4410 40395 4440
rect 40355 4405 40395 4410
rect 40405 4440 40445 4445
rect 40405 4410 40410 4440
rect 40410 4410 40440 4440
rect 40440 4410 40445 4440
rect 40405 4405 40445 4410
rect 40455 4440 40495 4445
rect 40455 4410 40460 4440
rect 40460 4410 40490 4440
rect 40490 4410 40495 4440
rect 40455 4405 40495 4410
rect 40505 4440 40545 4445
rect 40505 4410 40510 4440
rect 40510 4410 40540 4440
rect 40540 4410 40545 4440
rect 40505 4405 40545 4410
rect 40555 4440 40595 4445
rect 40555 4410 40560 4440
rect 40560 4410 40590 4440
rect 40590 4410 40595 4440
rect 40555 4405 40595 4410
rect 40605 4440 40645 4445
rect 40605 4410 40610 4440
rect 40610 4410 40640 4440
rect 40640 4410 40645 4440
rect 40605 4405 40645 4410
rect 40655 4440 40695 4445
rect 40655 4410 40660 4440
rect 40660 4410 40690 4440
rect 40690 4410 40695 4440
rect 40655 4405 40695 4410
rect 40705 4440 40745 4445
rect 40705 4410 40710 4440
rect 40710 4410 40740 4440
rect 40740 4410 40745 4440
rect 40705 4405 40745 4410
rect 40755 4440 40795 4445
rect 40755 4410 40760 4440
rect 40760 4410 40790 4440
rect 40790 4410 40795 4440
rect 40755 4405 40795 4410
rect 40805 4440 40845 4445
rect 40805 4410 40810 4440
rect 40810 4410 40840 4440
rect 40840 4410 40845 4440
rect 40805 4405 40845 4410
rect 40855 4440 40895 4445
rect 40855 4410 40860 4440
rect 40860 4410 40890 4440
rect 40890 4410 40895 4440
rect 40855 4405 40895 4410
rect 39805 4340 39845 4345
rect 39805 4310 39810 4340
rect 39810 4310 39840 4340
rect 39840 4310 39845 4340
rect 39805 4305 39845 4310
rect -3195 4205 -3155 4245
rect -3495 3840 -3455 3845
rect -3495 3810 -3490 3840
rect -3490 3810 -3460 3840
rect -3460 3810 -3455 3840
rect -3495 3805 -3455 3810
rect -3295 3840 -3255 3845
rect -3295 3810 -3290 3840
rect -3290 3810 -3260 3840
rect -3260 3810 -3255 3840
rect -3295 3805 -3255 3810
rect -3095 3840 -3055 3845
rect -3095 3810 -3090 3840
rect -3090 3810 -3060 3840
rect -3060 3810 -3055 3840
rect -3095 3805 -3055 3810
rect -1595 3840 -1555 3845
rect -1595 3810 -1590 3840
rect -1590 3810 -1560 3840
rect -1560 3810 -1555 3840
rect -1595 3805 -1555 3810
rect -1095 3840 -1055 3845
rect -1095 3810 -1090 3840
rect -1090 3810 -1060 3840
rect -1060 3810 -1055 3840
rect -1095 3805 -1055 3810
rect -895 3840 -855 3845
rect -895 3810 -890 3840
rect -890 3810 -860 3840
rect -860 3810 -855 3840
rect -895 3805 -855 3810
rect -695 3840 -655 3845
rect -695 3810 -690 3840
rect -690 3810 -660 3840
rect -660 3810 -655 3840
rect -695 3805 -655 3810
rect -495 3840 -455 3845
rect -495 3810 -490 3840
rect -490 3810 -460 3840
rect -460 3810 -455 3840
rect -495 3805 -455 3810
rect -295 3840 -255 3845
rect -295 3810 -290 3840
rect -290 3810 -260 3840
rect -260 3810 -255 3840
rect -295 3805 -255 3810
rect -95 3840 -55 3845
rect -95 3810 -90 3840
rect -90 3810 -60 3840
rect -60 3810 -55 3840
rect -95 3805 -55 3810
rect -3495 3790 -3455 3795
rect -3495 3760 -3490 3790
rect -3490 3760 -3460 3790
rect -3460 3760 -3455 3790
rect -3495 3755 -3455 3760
rect -3295 3790 -3255 3795
rect -3295 3760 -3290 3790
rect -3290 3760 -3260 3790
rect -3260 3760 -3255 3790
rect -3295 3755 -3255 3760
rect -3095 3790 -3055 3795
rect -3095 3760 -3090 3790
rect -3090 3760 -3060 3790
rect -3060 3760 -3055 3790
rect -3095 3755 -3055 3760
rect -1595 3790 -1555 3795
rect -1595 3760 -1590 3790
rect -1590 3760 -1560 3790
rect -1560 3760 -1555 3790
rect -1595 3755 -1555 3760
rect -1095 3790 -1055 3795
rect -1095 3760 -1090 3790
rect -1090 3760 -1060 3790
rect -1060 3760 -1055 3790
rect -1095 3755 -1055 3760
rect -895 3790 -855 3795
rect -895 3760 -890 3790
rect -890 3760 -860 3790
rect -860 3760 -855 3790
rect -895 3755 -855 3760
rect -695 3790 -655 3795
rect -695 3760 -690 3790
rect -690 3760 -660 3790
rect -660 3760 -655 3790
rect -695 3755 -655 3760
rect -495 3790 -455 3795
rect -495 3760 -490 3790
rect -490 3760 -460 3790
rect -460 3760 -455 3790
rect -495 3755 -455 3760
rect -295 3790 -255 3795
rect -295 3760 -290 3790
rect -290 3760 -260 3790
rect -260 3760 -255 3790
rect -295 3755 -255 3760
rect -95 3790 -55 3795
rect -95 3760 -90 3790
rect -90 3760 -60 3790
rect -60 3760 -55 3790
rect -95 3755 -55 3760
rect -3495 3740 -3455 3745
rect -3495 3710 -3490 3740
rect -3490 3710 -3460 3740
rect -3460 3710 -3455 3740
rect -3495 3705 -3455 3710
rect -3295 3740 -3255 3745
rect -3295 3710 -3290 3740
rect -3290 3710 -3260 3740
rect -3260 3710 -3255 3740
rect -3295 3705 -3255 3710
rect -3095 3740 -3055 3745
rect -3095 3710 -3090 3740
rect -3090 3710 -3060 3740
rect -3060 3710 -3055 3740
rect -3095 3705 -3055 3710
rect -1595 3740 -1555 3745
rect -1595 3710 -1590 3740
rect -1590 3710 -1560 3740
rect -1560 3710 -1555 3740
rect -1595 3705 -1555 3710
rect -1095 3740 -1055 3745
rect -1095 3710 -1090 3740
rect -1090 3710 -1060 3740
rect -1060 3710 -1055 3740
rect -1095 3705 -1055 3710
rect -895 3740 -855 3745
rect -895 3710 -890 3740
rect -890 3710 -860 3740
rect -860 3710 -855 3740
rect -895 3705 -855 3710
rect -695 3740 -655 3745
rect -695 3710 -690 3740
rect -690 3710 -660 3740
rect -660 3710 -655 3740
rect -695 3705 -655 3710
rect -495 3740 -455 3745
rect -495 3710 -490 3740
rect -490 3710 -460 3740
rect -460 3710 -455 3740
rect -495 3705 -455 3710
rect -295 3740 -255 3745
rect -295 3710 -290 3740
rect -290 3710 -260 3740
rect -260 3710 -255 3740
rect -295 3705 -255 3710
rect -95 3740 -55 3745
rect -95 3710 -90 3740
rect -90 3710 -60 3740
rect -60 3710 -55 3740
rect -95 3705 -55 3710
rect -1495 3405 -1455 3445
rect -1395 3305 -1355 3345
rect -1295 3205 -1255 3245
rect -1195 3105 -1155 3145
rect -995 2705 -955 2745
rect -795 2505 -755 2545
rect -3495 2140 -3455 2145
rect -3495 2110 -3490 2140
rect -3490 2110 -3460 2140
rect -3460 2110 -3455 2140
rect -3495 2105 -3455 2110
rect -3295 2140 -3255 2145
rect -3295 2110 -3290 2140
rect -3290 2110 -3260 2140
rect -3260 2110 -3255 2140
rect -3295 2105 -3255 2110
rect -3095 2140 -3055 2145
rect -3095 2110 -3090 2140
rect -3090 2110 -3060 2140
rect -3060 2110 -3055 2140
rect -3095 2105 -3055 2110
rect -1595 2140 -1555 2145
rect -1595 2110 -1590 2140
rect -1590 2110 -1560 2140
rect -1560 2110 -1555 2140
rect -1595 2105 -1555 2110
rect -1095 2140 -1055 2145
rect -1095 2110 -1090 2140
rect -1090 2110 -1060 2140
rect -1060 2110 -1055 2140
rect -1095 2105 -1055 2110
rect -895 2140 -855 2145
rect -895 2110 -890 2140
rect -890 2110 -860 2140
rect -860 2110 -855 2140
rect -895 2105 -855 2110
rect -695 2140 -655 2145
rect -695 2110 -690 2140
rect -690 2110 -660 2140
rect -660 2110 -655 2140
rect -695 2105 -655 2110
rect -495 2140 -455 2145
rect -495 2110 -490 2140
rect -490 2110 -460 2140
rect -460 2110 -455 2140
rect -495 2105 -455 2110
rect -295 2140 -255 2145
rect -295 2110 -290 2140
rect -290 2110 -260 2140
rect -260 2110 -255 2140
rect -295 2105 -255 2110
rect -95 2140 -55 2145
rect -95 2110 -90 2140
rect -90 2110 -60 2140
rect -60 2110 -55 2140
rect -95 2105 -55 2110
rect -3495 2090 -3455 2095
rect -3495 2060 -3490 2090
rect -3490 2060 -3460 2090
rect -3460 2060 -3455 2090
rect -3495 2055 -3455 2060
rect -3295 2090 -3255 2095
rect -3295 2060 -3290 2090
rect -3290 2060 -3260 2090
rect -3260 2060 -3255 2090
rect -3295 2055 -3255 2060
rect -3095 2090 -3055 2095
rect -3095 2060 -3090 2090
rect -3090 2060 -3060 2090
rect -3060 2060 -3055 2090
rect -3095 2055 -3055 2060
rect -1595 2090 -1555 2095
rect -1595 2060 -1590 2090
rect -1590 2060 -1560 2090
rect -1560 2060 -1555 2090
rect -1595 2055 -1555 2060
rect -1095 2090 -1055 2095
rect -1095 2060 -1090 2090
rect -1090 2060 -1060 2090
rect -1060 2060 -1055 2090
rect -1095 2055 -1055 2060
rect -895 2090 -855 2095
rect -895 2060 -890 2090
rect -890 2060 -860 2090
rect -860 2060 -855 2090
rect -895 2055 -855 2060
rect -695 2090 -655 2095
rect -695 2060 -690 2090
rect -690 2060 -660 2090
rect -660 2060 -655 2090
rect -695 2055 -655 2060
rect -495 2090 -455 2095
rect -495 2060 -490 2090
rect -490 2060 -460 2090
rect -460 2060 -455 2090
rect -495 2055 -455 2060
rect -295 2090 -255 2095
rect -295 2060 -290 2090
rect -290 2060 -260 2090
rect -260 2060 -255 2090
rect -295 2055 -255 2060
rect -95 2090 -55 2095
rect -95 2060 -90 2090
rect -90 2060 -60 2090
rect -60 2060 -55 2090
rect -95 2055 -55 2060
rect -3495 2040 -3455 2045
rect -3495 2010 -3490 2040
rect -3490 2010 -3460 2040
rect -3460 2010 -3455 2040
rect -3495 2005 -3455 2010
rect -3295 2040 -3255 2045
rect -3295 2010 -3290 2040
rect -3290 2010 -3260 2040
rect -3260 2010 -3255 2040
rect -3295 2005 -3255 2010
rect -3095 2040 -3055 2045
rect -3095 2010 -3090 2040
rect -3090 2010 -3060 2040
rect -3060 2010 -3055 2040
rect -3095 2005 -3055 2010
rect -1595 2040 -1555 2045
rect -1595 2010 -1590 2040
rect -1590 2010 -1560 2040
rect -1560 2010 -1555 2040
rect -1595 2005 -1555 2010
rect -1095 2040 -1055 2045
rect -1095 2010 -1090 2040
rect -1090 2010 -1060 2040
rect -1060 2010 -1055 2040
rect -1095 2005 -1055 2010
rect -895 2040 -855 2045
rect -895 2010 -890 2040
rect -890 2010 -860 2040
rect -860 2010 -855 2040
rect -895 2005 -855 2010
rect -695 2040 -655 2045
rect -695 2010 -690 2040
rect -690 2010 -660 2040
rect -660 2010 -655 2040
rect -695 2005 -655 2010
rect -495 2040 -455 2045
rect -495 2010 -490 2040
rect -490 2010 -460 2040
rect -460 2010 -455 2040
rect -495 2005 -455 2010
rect -295 2040 -255 2045
rect -295 2010 -290 2040
rect -290 2010 -260 2040
rect -260 2010 -255 2040
rect -295 2005 -255 2010
rect -95 2040 -55 2045
rect -95 2010 -90 2040
rect -90 2010 -60 2040
rect -60 2010 -55 2040
rect -95 2005 -55 2010
rect -595 1605 -555 1645
rect -395 1405 -355 1445
rect -195 1005 -155 1045
rect -3495 440 -3455 445
rect -3495 410 -3490 440
rect -3490 410 -3460 440
rect -3460 410 -3455 440
rect -3495 405 -3455 410
rect -3295 440 -3255 445
rect -3295 410 -3290 440
rect -3290 410 -3260 440
rect -3260 410 -3255 440
rect -3295 405 -3255 410
rect -3095 440 -3055 445
rect -3095 410 -3090 440
rect -3090 410 -3060 440
rect -3060 410 -3055 440
rect -3095 405 -3055 410
rect -1595 440 -1555 445
rect -1595 410 -1590 440
rect -1590 410 -1560 440
rect -1560 410 -1555 440
rect -1595 405 -1555 410
rect -1095 440 -1055 445
rect -1095 410 -1090 440
rect -1090 410 -1060 440
rect -1060 410 -1055 440
rect -1095 405 -1055 410
rect -895 440 -855 445
rect -895 410 -890 440
rect -890 410 -860 440
rect -860 410 -855 440
rect -895 405 -855 410
rect -695 440 -655 445
rect -695 410 -690 440
rect -690 410 -660 440
rect -660 410 -655 440
rect -695 405 -655 410
rect -495 440 -455 445
rect -495 410 -490 440
rect -490 410 -460 440
rect -460 410 -455 440
rect -495 405 -455 410
rect -295 440 -255 445
rect -295 410 -290 440
rect -290 410 -260 440
rect -260 410 -255 440
rect -295 405 -255 410
rect -95 440 -55 445
rect -95 410 -90 440
rect -90 410 -60 440
rect -60 410 -55 440
rect -95 405 -55 410
rect -3495 390 -3455 395
rect -3495 360 -3490 390
rect -3490 360 -3460 390
rect -3460 360 -3455 390
rect -3495 355 -3455 360
rect -3295 390 -3255 395
rect -3295 360 -3290 390
rect -3290 360 -3260 390
rect -3260 360 -3255 390
rect -3295 355 -3255 360
rect -3095 390 -3055 395
rect -3095 360 -3090 390
rect -3090 360 -3060 390
rect -3060 360 -3055 390
rect -3095 355 -3055 360
rect -1595 390 -1555 395
rect -1595 360 -1590 390
rect -1590 360 -1560 390
rect -1560 360 -1555 390
rect -1595 355 -1555 360
rect -1095 390 -1055 395
rect -1095 360 -1090 390
rect -1090 360 -1060 390
rect -1060 360 -1055 390
rect -1095 355 -1055 360
rect -895 390 -855 395
rect -895 360 -890 390
rect -890 360 -860 390
rect -860 360 -855 390
rect -895 355 -855 360
rect -695 390 -655 395
rect -695 360 -690 390
rect -690 360 -660 390
rect -660 360 -655 390
rect -695 355 -655 360
rect -495 390 -455 395
rect -495 360 -490 390
rect -490 360 -460 390
rect -460 360 -455 390
rect -495 355 -455 360
rect -295 390 -255 395
rect -295 360 -290 390
rect -290 360 -260 390
rect -260 360 -255 390
rect -295 355 -255 360
rect -95 390 -55 395
rect -95 360 -90 390
rect -90 360 -60 390
rect -60 360 -55 390
rect -95 355 -55 360
rect -3495 340 -3455 345
rect -3495 310 -3490 340
rect -3490 310 -3460 340
rect -3460 310 -3455 340
rect -3495 305 -3455 310
rect -3295 340 -3255 345
rect -3295 310 -3290 340
rect -3290 310 -3260 340
rect -3260 310 -3255 340
rect -3295 305 -3255 310
rect -3095 340 -3055 345
rect -3095 310 -3090 340
rect -3090 310 -3060 340
rect -3060 310 -3055 340
rect -3095 305 -3055 310
rect -1595 340 -1555 345
rect -1595 310 -1590 340
rect -1590 310 -1560 340
rect -1560 310 -1555 340
rect -1595 305 -1555 310
rect -1095 340 -1055 345
rect -1095 310 -1090 340
rect -1090 310 -1060 340
rect -1060 310 -1055 340
rect -1095 305 -1055 310
rect -895 340 -855 345
rect -895 310 -890 340
rect -890 310 -860 340
rect -860 310 -855 340
rect -895 305 -855 310
rect -695 340 -655 345
rect -695 310 -690 340
rect -690 310 -660 340
rect -660 310 -655 340
rect -695 305 -655 310
rect -495 340 -455 345
rect -495 310 -490 340
rect -490 310 -460 340
rect -460 310 -455 340
rect -495 305 -455 310
rect -295 340 -255 345
rect -295 310 -290 340
rect -290 310 -260 340
rect -260 310 -255 340
rect -295 305 -255 310
rect -95 340 -55 345
rect -95 310 -90 340
rect -90 310 -60 340
rect -60 310 -55 340
rect -95 305 -55 310
<< mimcap >>
rect 150 17850 3150 17900
rect 150 17200 200 17850
rect 3100 17200 3150 17850
rect 150 17150 3150 17200
rect 3400 17850 6400 17900
rect 3400 17200 3450 17850
rect 6350 17200 6400 17850
rect 3400 17150 6400 17200
rect 6650 17850 9650 17900
rect 6650 17200 6700 17850
rect 9600 17200 9650 17850
rect 6650 17150 9650 17200
rect 9900 17850 12900 17900
rect 9900 17200 9950 17850
rect 12850 17200 12900 17850
rect 9900 17150 12900 17200
rect 13150 17850 16150 17900
rect 13150 17200 13200 17850
rect 16100 17200 16150 17850
rect 13150 17150 16150 17200
rect 16400 17850 19400 17900
rect 16400 17200 16450 17850
rect 19350 17200 19400 17850
rect 16400 17150 19400 17200
rect 19650 17850 22650 17900
rect 19650 17200 19700 17850
rect 22600 17200 22650 17850
rect 19650 17150 22650 17200
rect 22900 17850 25900 17900
rect 22900 17200 22950 17850
rect 25850 17200 25900 17850
rect 22900 17150 25900 17200
rect 26150 17850 29150 17900
rect 26150 17200 26200 17850
rect 29100 17200 29150 17850
rect 26150 17150 29150 17200
rect 29400 17850 32400 17900
rect 29400 17200 29450 17850
rect 32350 17200 32400 17850
rect 29400 17150 32400 17200
rect 32650 17850 35650 17900
rect 32650 17200 32700 17850
rect 35600 17200 35650 17850
rect 32650 17150 35650 17200
rect 35900 17850 38900 17900
rect 35900 17200 35950 17850
rect 38850 17200 38900 17850
rect 35900 17150 38900 17200
rect 39150 17850 39700 17900
rect 39150 17200 39200 17850
rect 39650 17200 39700 17850
rect 39150 17150 39700 17200
rect 150 16650 3150 16700
rect 150 16000 200 16650
rect 3100 16000 3150 16650
rect 150 15950 3150 16000
rect 3400 16650 6400 16700
rect 3400 16000 3450 16650
rect 6350 16000 6400 16650
rect 3400 15950 6400 16000
rect 6650 16650 9650 16700
rect 6650 16000 6700 16650
rect 9600 16000 9650 16650
rect 6650 15950 9650 16000
rect 9900 16650 12900 16700
rect 9900 16000 9950 16650
rect 12850 16000 12900 16650
rect 9900 15950 12900 16000
rect 13150 16650 16150 16700
rect 13150 16000 13200 16650
rect 16100 16000 16150 16650
rect 13150 15950 16150 16000
rect 16400 16650 19400 16700
rect 16400 16000 16450 16650
rect 19350 16000 19400 16650
rect 16400 15950 19400 16000
rect 19650 16650 22650 16700
rect 19650 16000 19700 16650
rect 22600 16000 22650 16650
rect 19650 15950 22650 16000
rect 22900 16650 25900 16700
rect 22900 16000 22950 16650
rect 25850 16000 25900 16650
rect 22900 15950 25900 16000
rect 26150 16650 29150 16700
rect 26150 16000 26200 16650
rect 29100 16000 29150 16650
rect 26150 15950 29150 16000
rect 29400 16650 32400 16700
rect 29400 16000 29450 16650
rect 32350 16000 32400 16650
rect 29400 15950 32400 16000
rect 32650 16650 35650 16700
rect 32650 16000 32700 16650
rect 35600 16000 35650 16650
rect 32650 15950 35650 16000
rect 35900 16650 38900 16700
rect 35900 16000 35950 16650
rect 38850 16000 38900 16650
rect 35900 15950 38900 16000
rect 39150 16650 39700 16700
rect 39150 16000 39200 16650
rect 39650 16000 39700 16650
rect 39150 15950 39700 16000
<< mimcapcontact >>
rect 200 17200 3100 17850
rect 3450 17200 6350 17850
rect 6700 17200 9600 17850
rect 9950 17200 12850 17850
rect 13200 17200 16100 17850
rect 16450 17200 19350 17850
rect 19700 17200 22600 17850
rect 22950 17200 25850 17850
rect 26200 17200 29100 17850
rect 29450 17200 32350 17850
rect 32700 17200 35600 17850
rect 35950 17200 38850 17850
rect 39200 17200 39650 17850
rect 200 16000 3100 16650
rect 3450 16000 6350 16650
rect 6700 16000 9600 16650
rect 9950 16000 12850 16650
rect 13200 16000 16100 16650
rect 16450 16000 19350 16650
rect 19700 16000 22600 16650
rect 22950 16000 25850 16650
rect 26200 16000 29100 16650
rect 29450 16000 32350 16650
rect 32700 16000 35600 16650
rect 35950 16000 38850 16650
rect 39200 16000 39650 16650
<< metal4 >>
rect -3500 16945 -3450 18150
rect -3500 16905 -3495 16945
rect -3455 16905 -3450 16945
rect -3500 15745 -3450 16905
rect -3500 15705 -3495 15745
rect -3455 15705 -3450 15745
rect -3500 15345 -3450 15705
rect -3500 15305 -3495 15345
rect -3455 15305 -3450 15345
rect -3500 15295 -3450 15305
rect -3500 15255 -3495 15295
rect -3455 15255 -3450 15295
rect -3500 15245 -3450 15255
rect -3500 15205 -3495 15245
rect -3455 15205 -3450 15245
rect -3500 13645 -3450 15205
rect -3500 13605 -3495 13645
rect -3455 13605 -3450 13645
rect -3500 13595 -3450 13605
rect -3500 13555 -3495 13595
rect -3455 13555 -3450 13595
rect -3500 13545 -3450 13555
rect -3500 13505 -3495 13545
rect -3455 13505 -3450 13545
rect -3500 11945 -3450 13505
rect -3500 11905 -3495 11945
rect -3455 11905 -3450 11945
rect -3500 11895 -3450 11905
rect -3500 11855 -3495 11895
rect -3455 11855 -3450 11895
rect -3500 11845 -3450 11855
rect -3500 11805 -3495 11845
rect -3455 11805 -3450 11845
rect -3500 3845 -3450 11805
rect -3500 3805 -3495 3845
rect -3455 3805 -3450 3845
rect -3500 3795 -3450 3805
rect -3500 3755 -3495 3795
rect -3455 3755 -3450 3795
rect -3500 3745 -3450 3755
rect -3500 3705 -3495 3745
rect -3455 3705 -3450 3745
rect -3500 2145 -3450 3705
rect -3500 2105 -3495 2145
rect -3455 2105 -3450 2145
rect -3500 2095 -3450 2105
rect -3500 2055 -3495 2095
rect -3455 2055 -3450 2095
rect -3500 2045 -3450 2055
rect -3500 2005 -3495 2045
rect -3455 2005 -3450 2045
rect -3500 445 -3450 2005
rect -3500 405 -3495 445
rect -3455 405 -3450 445
rect -3500 395 -3450 405
rect -3500 355 -3495 395
rect -3455 355 -3450 395
rect -3500 345 -3450 355
rect -3500 305 -3495 345
rect -3455 305 -3450 345
rect -3500 0 -3450 305
rect -3400 10845 -3350 18150
rect -3400 10805 -3395 10845
rect -3355 10805 -3350 10845
rect -3400 4845 -3350 10805
rect -3400 4805 -3395 4845
rect -3355 4805 -3350 4845
rect -3400 0 -3350 4805
rect -3300 16945 -3250 18150
rect -3300 16905 -3295 16945
rect -3255 16905 -3250 16945
rect -3300 15745 -3250 16905
rect -3300 15705 -3295 15745
rect -3255 15705 -3250 15745
rect -3300 15345 -3250 15705
rect -3300 15305 -3295 15345
rect -3255 15305 -3250 15345
rect -3300 15295 -3250 15305
rect -3300 15255 -3295 15295
rect -3255 15255 -3250 15295
rect -3300 15245 -3250 15255
rect -3300 15205 -3295 15245
rect -3255 15205 -3250 15245
rect -3300 13645 -3250 15205
rect -3300 13605 -3295 13645
rect -3255 13605 -3250 13645
rect -3300 13595 -3250 13605
rect -3300 13555 -3295 13595
rect -3255 13555 -3250 13595
rect -3300 13545 -3250 13555
rect -3300 13505 -3295 13545
rect -3255 13505 -3250 13545
rect -3300 11945 -3250 13505
rect -3300 11905 -3295 11945
rect -3255 11905 -3250 11945
rect -3300 11895 -3250 11905
rect -3300 11855 -3295 11895
rect -3255 11855 -3250 11895
rect -3300 11845 -3250 11855
rect -3300 11805 -3295 11845
rect -3255 11805 -3250 11845
rect -3300 3845 -3250 11805
rect -3300 3805 -3295 3845
rect -3255 3805 -3250 3845
rect -3300 3795 -3250 3805
rect -3300 3755 -3295 3795
rect -3255 3755 -3250 3795
rect -3300 3745 -3250 3755
rect -3300 3705 -3295 3745
rect -3255 3705 -3250 3745
rect -3300 2145 -3250 3705
rect -3300 2105 -3295 2145
rect -3255 2105 -3250 2145
rect -3300 2095 -3250 2105
rect -3300 2055 -3295 2095
rect -3255 2055 -3250 2095
rect -3300 2045 -3250 2055
rect -3300 2005 -3295 2045
rect -3255 2005 -3250 2045
rect -3300 445 -3250 2005
rect -3300 405 -3295 445
rect -3255 405 -3250 445
rect -3300 395 -3250 405
rect -3300 355 -3295 395
rect -3255 355 -3250 395
rect -3300 345 -3250 355
rect -3300 305 -3295 345
rect -3255 305 -3250 345
rect -3300 0 -3250 305
rect -3200 11445 -3150 18150
rect -3200 11405 -3195 11445
rect -3155 11405 -3150 11445
rect -3200 4245 -3150 11405
rect -3200 4205 -3195 4245
rect -3155 4205 -3150 4245
rect -3200 0 -3150 4205
rect -3100 16945 -3050 18150
rect -3100 16905 -3095 16945
rect -3055 16905 -3050 16945
rect -3100 15745 -3050 16905
rect -3100 15705 -3095 15745
rect -3055 15705 -3050 15745
rect -3100 15345 -3050 15705
rect -3100 15305 -3095 15345
rect -3055 15305 -3050 15345
rect -3100 15295 -3050 15305
rect -3100 15255 -3095 15295
rect -3055 15255 -3050 15295
rect -3100 15245 -3050 15255
rect -3100 15205 -3095 15245
rect -3055 15205 -3050 15245
rect -3100 13645 -3050 15205
rect -3100 13605 -3095 13645
rect -3055 13605 -3050 13645
rect -3100 13595 -3050 13605
rect -3100 13555 -3095 13595
rect -3055 13555 -3050 13595
rect -3100 13545 -3050 13555
rect -3100 13505 -3095 13545
rect -3055 13505 -3050 13545
rect -3100 11945 -3050 13505
rect -3100 11905 -3095 11945
rect -3055 11905 -3050 11945
rect -3100 11895 -3050 11905
rect -3100 11855 -3095 11895
rect -3055 11855 -3050 11895
rect -3100 11845 -3050 11855
rect -3100 11805 -3095 11845
rect -3055 11805 -3050 11845
rect -3100 3845 -3050 11805
rect -3100 3805 -3095 3845
rect -3055 3805 -3050 3845
rect -3100 3795 -3050 3805
rect -3100 3755 -3095 3795
rect -3055 3755 -3050 3795
rect -3100 3745 -3050 3755
rect -3100 3705 -3095 3745
rect -3055 3705 -3050 3745
rect -3100 2145 -3050 3705
rect -3100 2105 -3095 2145
rect -3055 2105 -3050 2145
rect -3100 2095 -3050 2105
rect -3100 2055 -3095 2095
rect -3055 2055 -3050 2095
rect -3100 2045 -3050 2055
rect -3100 2005 -3095 2045
rect -3055 2005 -3050 2045
rect -3100 445 -3050 2005
rect -3100 405 -3095 445
rect -3055 405 -3050 445
rect -3100 395 -3050 405
rect -3100 355 -3095 395
rect -3055 355 -3050 395
rect -3100 345 -3050 355
rect -3100 305 -3095 345
rect -3055 305 -3050 345
rect -3100 0 -3050 305
rect -3000 18100 -1650 18150
rect -3000 17150 -2950 18100
rect -2900 17150 -2850 18100
rect -2800 17150 -2750 18100
rect -2700 17150 -2650 18100
rect -2600 17150 -2550 18100
rect -2500 17150 -2450 18100
rect -2400 17150 -2350 18100
rect -2300 17150 -2250 18100
rect -2200 17150 -2150 18100
rect -2100 17150 -2050 18100
rect -2000 17150 -1950 18100
rect -1900 17150 -1850 18100
rect -1800 17150 -1750 18100
rect -1700 17150 -1650 18100
rect -3000 17100 -1650 17150
rect -3000 15750 -2950 17100
rect -2900 15750 -2850 17100
rect -2800 15750 -2750 17100
rect -3000 15700 -2750 15750
rect -3000 10645 -2950 15700
rect -3000 10605 -2995 10645
rect -2955 10605 -2950 10645
rect -3000 10595 -2950 10605
rect -3000 10555 -2995 10595
rect -2955 10555 -2950 10595
rect -3000 10545 -2950 10555
rect -3000 10505 -2995 10545
rect -2955 10505 -2950 10545
rect -3000 9345 -2950 10505
rect -3000 9305 -2995 9345
rect -2955 9305 -2950 9345
rect -3000 9295 -2950 9305
rect -3000 9255 -2995 9295
rect -2955 9255 -2950 9295
rect -3000 9245 -2950 9255
rect -3000 9205 -2995 9245
rect -2955 9205 -2950 9245
rect -3000 8045 -2950 9205
rect -3000 8005 -2995 8045
rect -2955 8005 -2950 8045
rect -3000 7995 -2950 8005
rect -3000 7955 -2995 7995
rect -2955 7955 -2950 7995
rect -3000 7945 -2950 7955
rect -3000 7905 -2995 7945
rect -2955 7905 -2950 7945
rect -3000 7745 -2950 7905
rect -3000 7705 -2995 7745
rect -2955 7705 -2950 7745
rect -3000 7695 -2950 7705
rect -3000 7655 -2995 7695
rect -2955 7655 -2950 7695
rect -3000 7645 -2950 7655
rect -3000 7605 -2995 7645
rect -2955 7605 -2950 7645
rect -3000 6445 -2950 7605
rect -3000 6405 -2995 6445
rect -2955 6405 -2950 6445
rect -3000 6395 -2950 6405
rect -3000 6355 -2995 6395
rect -2955 6355 -2950 6395
rect -3000 6345 -2950 6355
rect -3000 6305 -2995 6345
rect -2955 6305 -2950 6345
rect -3000 5145 -2950 6305
rect -3000 5105 -2995 5145
rect -2955 5105 -2950 5145
rect -3000 5095 -2950 5105
rect -3000 5055 -2995 5095
rect -2955 5055 -2950 5095
rect -3000 5045 -2950 5055
rect -3000 5005 -2995 5045
rect -2955 5005 -2950 5045
rect -3000 0 -2950 5005
rect -2900 8445 -2850 15650
rect -2900 8405 -2895 8445
rect -2855 8405 -2850 8445
rect -2900 7245 -2850 8405
rect -2900 7205 -2895 7245
rect -2855 7205 -2850 7245
rect -2900 0 -2850 7205
rect -2800 10645 -2750 15700
rect -2800 10605 -2795 10645
rect -2755 10605 -2750 10645
rect -2800 10595 -2750 10605
rect -2800 10555 -2795 10595
rect -2755 10555 -2750 10595
rect -2800 10545 -2750 10555
rect -2800 10505 -2795 10545
rect -2755 10505 -2750 10545
rect -2800 9345 -2750 10505
rect -2800 9305 -2795 9345
rect -2755 9305 -2750 9345
rect -2800 9295 -2750 9305
rect -2800 9255 -2795 9295
rect -2755 9255 -2750 9295
rect -2800 9245 -2750 9255
rect -2800 9205 -2795 9245
rect -2755 9205 -2750 9245
rect -2800 8045 -2750 9205
rect -2800 8005 -2795 8045
rect -2755 8005 -2750 8045
rect -2800 7995 -2750 8005
rect -2800 7955 -2795 7995
rect -2755 7955 -2750 7995
rect -2800 7945 -2750 7955
rect -2800 7905 -2795 7945
rect -2755 7905 -2750 7945
rect -2800 7745 -2750 7905
rect -2800 7705 -2795 7745
rect -2755 7705 -2750 7745
rect -2800 7695 -2750 7705
rect -2800 7655 -2795 7695
rect -2755 7655 -2750 7695
rect -2800 7645 -2750 7655
rect -2800 7605 -2795 7645
rect -2755 7605 -2750 7645
rect -2800 6445 -2750 7605
rect -2800 6405 -2795 6445
rect -2755 6405 -2750 6445
rect -2800 6395 -2750 6405
rect -2800 6355 -2795 6395
rect -2755 6355 -2750 6395
rect -2800 6345 -2750 6355
rect -2800 6305 -2795 6345
rect -2755 6305 -2750 6345
rect -2800 5145 -2750 6305
rect -2800 5105 -2795 5145
rect -2755 5105 -2750 5145
rect -2800 5095 -2750 5105
rect -2800 5055 -2795 5095
rect -2755 5055 -2750 5095
rect -2800 5045 -2750 5055
rect -2800 5005 -2795 5045
rect -2755 5005 -2750 5045
rect -2800 0 -2750 5005
rect -2700 17045 -2650 17050
rect -2700 17005 -2695 17045
rect -2655 17005 -2650 17045
rect -2700 8845 -2650 17005
rect -2700 8805 -2695 8845
rect -2655 8805 -2650 8845
rect -2700 6845 -2650 8805
rect -2700 6805 -2695 6845
rect -2655 6805 -2650 6845
rect -2700 0 -2650 6805
rect -2600 15750 -2550 17100
rect -2500 15750 -2450 17100
rect -2400 15750 -2350 17100
rect -2300 15750 -2250 17100
rect -2200 15750 -2150 17100
rect -2100 15750 -2050 17100
rect -2000 15750 -1950 17100
rect -1900 15750 -1850 17100
rect -1800 15750 -1750 17100
rect -1700 15750 -1650 17100
rect -2600 15700 -1650 15750
rect -2600 10645 -2550 15700
rect -2600 10605 -2595 10645
rect -2555 10605 -2550 10645
rect -2600 10595 -2550 10605
rect -2600 10555 -2595 10595
rect -2555 10555 -2550 10595
rect -2600 10545 -2550 10555
rect -2600 10505 -2595 10545
rect -2555 10505 -2550 10545
rect -2600 9345 -2550 10505
rect -2600 9305 -2595 9345
rect -2555 9305 -2550 9345
rect -2600 9295 -2550 9305
rect -2600 9255 -2595 9295
rect -2555 9255 -2550 9295
rect -2600 9245 -2550 9255
rect -2600 9205 -2595 9245
rect -2555 9205 -2550 9245
rect -2600 8045 -2550 9205
rect -2600 8005 -2595 8045
rect -2555 8005 -2550 8045
rect -2600 7995 -2550 8005
rect -2600 7955 -2595 7995
rect -2555 7955 -2550 7995
rect -2600 7945 -2550 7955
rect -2600 7905 -2595 7945
rect -2555 7905 -2550 7945
rect -2600 7745 -2550 7905
rect -2600 7705 -2595 7745
rect -2555 7705 -2550 7745
rect -2600 7695 -2550 7705
rect -2600 7655 -2595 7695
rect -2555 7655 -2550 7695
rect -2600 7645 -2550 7655
rect -2600 7605 -2595 7645
rect -2555 7605 -2550 7645
rect -2600 6445 -2550 7605
rect -2600 6405 -2595 6445
rect -2555 6405 -2550 6445
rect -2600 6395 -2550 6405
rect -2600 6355 -2595 6395
rect -2555 6355 -2550 6395
rect -2600 6345 -2550 6355
rect -2600 6305 -2595 6345
rect -2555 6305 -2550 6345
rect -2600 5145 -2550 6305
rect -2600 5105 -2595 5145
rect -2555 5105 -2550 5145
rect -2600 5095 -2550 5105
rect -2600 5055 -2595 5095
rect -2555 5055 -2550 5095
rect -2600 5045 -2550 5055
rect -2600 5005 -2595 5045
rect -2555 5005 -2550 5045
rect -2600 0 -2550 5005
rect -2500 9045 -2450 15650
rect -2500 9005 -2495 9045
rect -2455 9005 -2450 9045
rect -2500 6645 -2450 9005
rect -2500 6605 -2495 6645
rect -2455 6605 -2450 6645
rect -2500 0 -2450 6605
rect -2400 10645 -2350 15700
rect -2400 10605 -2395 10645
rect -2355 10605 -2350 10645
rect -2400 10595 -2350 10605
rect -2400 10555 -2395 10595
rect -2355 10555 -2350 10595
rect -2400 10545 -2350 10555
rect -2400 10505 -2395 10545
rect -2355 10505 -2350 10545
rect -2400 9345 -2350 10505
rect -2400 9305 -2395 9345
rect -2355 9305 -2350 9345
rect -2400 9295 -2350 9305
rect -2400 9255 -2395 9295
rect -2355 9255 -2350 9295
rect -2400 9245 -2350 9255
rect -2400 9205 -2395 9245
rect -2355 9205 -2350 9245
rect -2400 8045 -2350 9205
rect -2400 8005 -2395 8045
rect -2355 8005 -2350 8045
rect -2400 7995 -2350 8005
rect -2400 7955 -2395 7995
rect -2355 7955 -2350 7995
rect -2400 7945 -2350 7955
rect -2400 7905 -2395 7945
rect -2355 7905 -2350 7945
rect -2400 7745 -2350 7905
rect -2400 7705 -2395 7745
rect -2355 7705 -2350 7745
rect -2400 7695 -2350 7705
rect -2400 7655 -2395 7695
rect -2355 7655 -2350 7695
rect -2400 7645 -2350 7655
rect -2400 7605 -2395 7645
rect -2355 7605 -2350 7645
rect -2400 6445 -2350 7605
rect -2400 6405 -2395 6445
rect -2355 6405 -2350 6445
rect -2400 6395 -2350 6405
rect -2400 6355 -2395 6395
rect -2355 6355 -2350 6395
rect -2400 6345 -2350 6355
rect -2400 6305 -2395 6345
rect -2355 6305 -2350 6345
rect -2400 5145 -2350 6305
rect -2400 5105 -2395 5145
rect -2355 5105 -2350 5145
rect -2400 5095 -2350 5105
rect -2400 5055 -2395 5095
rect -2355 5055 -2350 5095
rect -2400 5045 -2350 5055
rect -2400 5005 -2395 5045
rect -2355 5005 -2350 5045
rect -2400 0 -2350 5005
rect -2300 9545 -2250 15650
rect -2300 9505 -2295 9545
rect -2255 9505 -2250 9545
rect -2300 6145 -2250 9505
rect -2300 6105 -2295 6145
rect -2255 6105 -2250 6145
rect -2300 0 -2250 6105
rect -2200 10645 -2150 15700
rect -2200 10605 -2195 10645
rect -2155 10605 -2150 10645
rect -2200 10595 -2150 10605
rect -2200 10555 -2195 10595
rect -2155 10555 -2150 10595
rect -2200 10545 -2150 10555
rect -2200 10505 -2195 10545
rect -2155 10505 -2150 10545
rect -2200 9345 -2150 10505
rect -2200 9305 -2195 9345
rect -2155 9305 -2150 9345
rect -2200 9295 -2150 9305
rect -2200 9255 -2195 9295
rect -2155 9255 -2150 9295
rect -2200 9245 -2150 9255
rect -2200 9205 -2195 9245
rect -2155 9205 -2150 9245
rect -2200 8045 -2150 9205
rect -2200 8005 -2195 8045
rect -2155 8005 -2150 8045
rect -2200 7995 -2150 8005
rect -2200 7955 -2195 7995
rect -2155 7955 -2150 7995
rect -2200 7945 -2150 7955
rect -2200 7905 -2195 7945
rect -2155 7905 -2150 7945
rect -2200 7745 -2150 7905
rect -2200 7705 -2195 7745
rect -2155 7705 -2150 7745
rect -2200 7695 -2150 7705
rect -2200 7655 -2195 7695
rect -2155 7655 -2150 7695
rect -2200 7645 -2150 7655
rect -2200 7605 -2195 7645
rect -2155 7605 -2150 7645
rect -2200 6445 -2150 7605
rect -2200 6405 -2195 6445
rect -2155 6405 -2150 6445
rect -2200 6395 -2150 6405
rect -2200 6355 -2195 6395
rect -2155 6355 -2150 6395
rect -2200 6345 -2150 6355
rect -2200 6305 -2195 6345
rect -2155 6305 -2150 6345
rect -2200 5145 -2150 6305
rect -2200 5105 -2195 5145
rect -2155 5105 -2150 5145
rect -2200 5095 -2150 5105
rect -2200 5055 -2195 5095
rect -2155 5055 -2150 5095
rect -2200 5045 -2150 5055
rect -2200 5005 -2195 5045
rect -2155 5005 -2150 5045
rect -2200 0 -2150 5005
rect -2100 9745 -2050 15650
rect -2100 9705 -2095 9745
rect -2055 9705 -2050 9745
rect -2100 5945 -2050 9705
rect -2100 5905 -2095 5945
rect -2055 5905 -2050 5945
rect -2100 0 -2050 5905
rect -2000 10645 -1950 15700
rect -2000 10605 -1995 10645
rect -1955 10605 -1950 10645
rect -2000 10595 -1950 10605
rect -2000 10555 -1995 10595
rect -1955 10555 -1950 10595
rect -2000 10545 -1950 10555
rect -2000 10505 -1995 10545
rect -1955 10505 -1950 10545
rect -2000 9345 -1950 10505
rect -2000 9305 -1995 9345
rect -1955 9305 -1950 9345
rect -2000 9295 -1950 9305
rect -2000 9255 -1995 9295
rect -1955 9255 -1950 9295
rect -2000 9245 -1950 9255
rect -2000 9205 -1995 9245
rect -1955 9205 -1950 9245
rect -2000 8045 -1950 9205
rect -2000 8005 -1995 8045
rect -1955 8005 -1950 8045
rect -2000 7995 -1950 8005
rect -2000 7955 -1995 7995
rect -1955 7955 -1950 7995
rect -2000 7945 -1950 7955
rect -2000 7905 -1995 7945
rect -1955 7905 -1950 7945
rect -2000 7745 -1950 7905
rect -2000 7705 -1995 7745
rect -1955 7705 -1950 7745
rect -2000 7695 -1950 7705
rect -2000 7655 -1995 7695
rect -1955 7655 -1950 7695
rect -2000 7645 -1950 7655
rect -2000 7605 -1995 7645
rect -1955 7605 -1950 7645
rect -2000 6445 -1950 7605
rect -2000 6405 -1995 6445
rect -1955 6405 -1950 6445
rect -2000 6395 -1950 6405
rect -2000 6355 -1995 6395
rect -1955 6355 -1950 6395
rect -2000 6345 -1950 6355
rect -2000 6305 -1995 6345
rect -1955 6305 -1950 6345
rect -2000 5145 -1950 6305
rect -2000 5105 -1995 5145
rect -1955 5105 -1950 5145
rect -2000 5095 -1950 5105
rect -2000 5055 -1995 5095
rect -1955 5055 -1950 5095
rect -2000 5045 -1950 5055
rect -2000 5005 -1995 5045
rect -1955 5005 -1950 5045
rect -2000 0 -1950 5005
rect -1900 10145 -1850 15650
rect -1900 10105 -1895 10145
rect -1855 10105 -1850 10145
rect -1900 5545 -1850 10105
rect -1900 5505 -1895 5545
rect -1855 5505 -1850 5545
rect -1900 0 -1850 5505
rect -1800 10245 -1750 15650
rect -1800 10205 -1795 10245
rect -1755 10205 -1750 10245
rect -1800 5445 -1750 10205
rect -1800 5405 -1795 5445
rect -1755 5405 -1750 5445
rect -1800 0 -1750 5405
rect -1700 10645 -1650 15700
rect -1700 10605 -1695 10645
rect -1655 10605 -1650 10645
rect -1700 10595 -1650 10605
rect -1700 10555 -1695 10595
rect -1655 10555 -1650 10595
rect -1700 10545 -1650 10555
rect -1700 10505 -1695 10545
rect -1655 10505 -1650 10545
rect -1700 9345 -1650 10505
rect -1700 9305 -1695 9345
rect -1655 9305 -1650 9345
rect -1700 9295 -1650 9305
rect -1700 9255 -1695 9295
rect -1655 9255 -1650 9295
rect -1700 9245 -1650 9255
rect -1700 9205 -1695 9245
rect -1655 9205 -1650 9245
rect -1700 8045 -1650 9205
rect -1700 8005 -1695 8045
rect -1655 8005 -1650 8045
rect -1700 7995 -1650 8005
rect -1700 7955 -1695 7995
rect -1655 7955 -1650 7995
rect -1700 7945 -1650 7955
rect -1700 7905 -1695 7945
rect -1655 7905 -1650 7945
rect -1700 7745 -1650 7905
rect -1700 7705 -1695 7745
rect -1655 7705 -1650 7745
rect -1700 7695 -1650 7705
rect -1700 7655 -1695 7695
rect -1655 7655 -1650 7695
rect -1700 7645 -1650 7655
rect -1700 7605 -1695 7645
rect -1655 7605 -1650 7645
rect -1700 6445 -1650 7605
rect -1700 6405 -1695 6445
rect -1655 6405 -1650 6445
rect -1700 6395 -1650 6405
rect -1700 6355 -1695 6395
rect -1655 6355 -1650 6395
rect -1700 6345 -1650 6355
rect -1700 6305 -1695 6345
rect -1655 6305 -1650 6345
rect -1700 5145 -1650 6305
rect -1700 5105 -1695 5145
rect -1655 5105 -1650 5145
rect -1700 5095 -1650 5105
rect -1700 5055 -1695 5095
rect -1655 5055 -1650 5095
rect -1700 5045 -1650 5055
rect -1700 5005 -1695 5045
rect -1655 5005 -1650 5045
rect -1700 0 -1650 5005
rect -1600 16945 -1550 18150
rect -1600 16905 -1595 16945
rect -1555 16905 -1550 16945
rect -1600 15745 -1550 16905
rect -1600 15705 -1595 15745
rect -1555 15705 -1550 15745
rect -1600 15345 -1550 15705
rect -1600 15305 -1595 15345
rect -1555 15305 -1550 15345
rect -1600 15295 -1550 15305
rect -1600 15255 -1595 15295
rect -1555 15255 -1550 15295
rect -1600 15245 -1550 15255
rect -1600 15205 -1595 15245
rect -1555 15205 -1550 15245
rect -1600 13645 -1550 15205
rect -1600 13605 -1595 13645
rect -1555 13605 -1550 13645
rect -1600 13595 -1550 13605
rect -1600 13555 -1595 13595
rect -1555 13555 -1550 13595
rect -1600 13545 -1550 13555
rect -1600 13505 -1595 13545
rect -1555 13505 -1550 13545
rect -1600 11945 -1550 13505
rect -1600 11905 -1595 11945
rect -1555 11905 -1550 11945
rect -1600 11895 -1550 11905
rect -1600 11855 -1595 11895
rect -1555 11855 -1550 11895
rect -1600 11845 -1550 11855
rect -1600 11805 -1595 11845
rect -1555 11805 -1550 11845
rect -1600 3845 -1550 11805
rect -1600 3805 -1595 3845
rect -1555 3805 -1550 3845
rect -1600 3795 -1550 3805
rect -1600 3755 -1595 3795
rect -1555 3755 -1550 3795
rect -1600 3745 -1550 3755
rect -1600 3705 -1595 3745
rect -1555 3705 -1550 3745
rect -1600 2145 -1550 3705
rect -1600 2105 -1595 2145
rect -1555 2105 -1550 2145
rect -1600 2095 -1550 2105
rect -1600 2055 -1595 2095
rect -1555 2055 -1550 2095
rect -1600 2045 -1550 2055
rect -1600 2005 -1595 2045
rect -1555 2005 -1550 2045
rect -1600 445 -1550 2005
rect -1600 405 -1595 445
rect -1555 405 -1550 445
rect -1600 395 -1550 405
rect -1600 355 -1595 395
rect -1555 355 -1550 395
rect -1600 345 -1550 355
rect -1600 305 -1595 345
rect -1555 305 -1550 345
rect -1600 0 -1550 305
rect -1500 12245 -1450 18150
rect -1500 12205 -1495 12245
rect -1455 12205 -1450 12245
rect -1500 3445 -1450 12205
rect -1500 3405 -1495 3445
rect -1455 3405 -1450 3445
rect -1500 0 -1450 3405
rect -1400 12345 -1350 18150
rect -1400 12305 -1395 12345
rect -1355 12305 -1350 12345
rect -1400 3345 -1350 12305
rect -1400 3305 -1395 3345
rect -1355 3305 -1350 3345
rect -1400 0 -1350 3305
rect -1300 18100 -1250 18150
rect -1300 12445 -1250 18050
rect -1200 18100 -50 18150
rect -1200 16950 -1150 18100
rect -1100 16950 -1050 18100
rect -1000 16950 -950 18100
rect -900 16950 -850 18100
rect -800 16950 -750 18100
rect -700 16950 -650 18100
rect -600 16950 -550 18100
rect -500 16950 -450 18100
rect -400 16950 -350 18100
rect -300 16950 -250 18100
rect -200 16950 -150 18100
rect -100 16950 -50 18100
rect -1200 16945 -50 16950
rect -1200 16905 -1195 16945
rect -1155 16905 -1095 16945
rect -1055 16905 -995 16945
rect -955 16905 -895 16945
rect -855 16905 -795 16945
rect -755 16905 -695 16945
rect -655 16905 -595 16945
rect -555 16905 -495 16945
rect -455 16905 -395 16945
rect -355 16905 -295 16945
rect -255 16905 -195 16945
rect -155 16905 -95 16945
rect -55 16905 -50 16945
rect -1200 16900 -50 16905
rect -1200 15750 -1150 16900
rect -1100 15750 -1050 16900
rect -1000 15750 -950 16900
rect -900 15750 -850 16900
rect -800 15750 -750 16900
rect -700 15750 -650 16900
rect -600 15750 -550 16900
rect -500 15750 -450 16900
rect -1200 15745 -450 15750
rect -1200 15705 -1195 15745
rect -1155 15705 -1095 15745
rect -1055 15705 -995 15745
rect -955 15705 -895 15745
rect -855 15705 -695 15745
rect -655 15705 -595 15745
rect -555 15705 -495 15745
rect -455 15705 -450 15745
rect -1200 15700 -450 15705
rect -1300 12405 -1295 12445
rect -1255 12405 -1250 12445
rect -1300 3245 -1250 12405
rect -1300 3205 -1295 3245
rect -1255 3205 -1250 3245
rect -1300 0 -1250 3205
rect -1200 12545 -1150 15650
rect -1200 12505 -1195 12545
rect -1155 12505 -1150 12545
rect -1200 3145 -1150 12505
rect -1200 3105 -1195 3145
rect -1155 3105 -1150 3145
rect -1200 0 -1150 3105
rect -1100 15345 -1050 15700
rect -1100 15305 -1095 15345
rect -1055 15305 -1050 15345
rect -1100 15295 -1050 15305
rect -1100 15255 -1095 15295
rect -1055 15255 -1050 15295
rect -1100 15245 -1050 15255
rect -1100 15205 -1095 15245
rect -1055 15205 -1050 15245
rect -1100 13645 -1050 15205
rect -1100 13605 -1095 13645
rect -1055 13605 -1050 13645
rect -1100 13595 -1050 13605
rect -1100 13555 -1095 13595
rect -1055 13555 -1050 13595
rect -1100 13545 -1050 13555
rect -1100 13505 -1095 13545
rect -1055 13505 -1050 13545
rect -1100 11945 -1050 13505
rect -1100 11905 -1095 11945
rect -1055 11905 -1050 11945
rect -1100 11895 -1050 11905
rect -1100 11855 -1095 11895
rect -1055 11855 -1050 11895
rect -1100 11845 -1050 11855
rect -1100 11805 -1095 11845
rect -1055 11805 -1050 11845
rect -1100 3845 -1050 11805
rect -1100 3805 -1095 3845
rect -1055 3805 -1050 3845
rect -1100 3795 -1050 3805
rect -1100 3755 -1095 3795
rect -1055 3755 -1050 3795
rect -1100 3745 -1050 3755
rect -1100 3705 -1095 3745
rect -1055 3705 -1050 3745
rect -1100 2145 -1050 3705
rect -1100 2105 -1095 2145
rect -1055 2105 -1050 2145
rect -1100 2095 -1050 2105
rect -1100 2055 -1095 2095
rect -1055 2055 -1050 2095
rect -1100 2045 -1050 2055
rect -1100 2005 -1095 2045
rect -1055 2005 -1050 2045
rect -1100 445 -1050 2005
rect -1100 405 -1095 445
rect -1055 405 -1050 445
rect -1100 395 -1050 405
rect -1100 355 -1095 395
rect -1055 355 -1050 395
rect -1100 345 -1050 355
rect -1100 305 -1095 345
rect -1055 305 -1050 345
rect -1100 0 -1050 305
rect -1000 12945 -950 15650
rect -1000 12905 -995 12945
rect -955 12905 -950 12945
rect -1000 2745 -950 12905
rect -1000 2705 -995 2745
rect -955 2705 -950 2745
rect -1000 0 -950 2705
rect -900 15345 -850 15700
rect -900 15305 -895 15345
rect -855 15305 -850 15345
rect -900 15295 -850 15305
rect -900 15255 -895 15295
rect -855 15255 -850 15295
rect -900 15245 -850 15255
rect -900 15205 -895 15245
rect -855 15205 -850 15245
rect -900 13645 -850 15205
rect -900 13605 -895 13645
rect -855 13605 -850 13645
rect -900 13595 -850 13605
rect -900 13555 -895 13595
rect -855 13555 -850 13595
rect -900 13545 -850 13555
rect -900 13505 -895 13545
rect -855 13505 -850 13545
rect -900 11945 -850 13505
rect -900 11905 -895 11945
rect -855 11905 -850 11945
rect -900 11895 -850 11905
rect -900 11855 -895 11895
rect -855 11855 -850 11895
rect -900 11845 -850 11855
rect -900 11805 -895 11845
rect -855 11805 -850 11845
rect -900 3845 -850 11805
rect -900 3805 -895 3845
rect -855 3805 -850 3845
rect -900 3795 -850 3805
rect -900 3755 -895 3795
rect -855 3755 -850 3795
rect -900 3745 -850 3755
rect -900 3705 -895 3745
rect -855 3705 -850 3745
rect -900 2145 -850 3705
rect -900 2105 -895 2145
rect -855 2105 -850 2145
rect -900 2095 -850 2105
rect -900 2055 -895 2095
rect -855 2055 -850 2095
rect -900 2045 -850 2055
rect -900 2005 -895 2045
rect -855 2005 -850 2045
rect -900 445 -850 2005
rect -900 405 -895 445
rect -855 405 -850 445
rect -900 395 -850 405
rect -900 355 -895 395
rect -855 355 -850 395
rect -900 345 -850 355
rect -900 305 -895 345
rect -855 305 -850 345
rect -900 0 -850 305
rect -800 13145 -750 15650
rect -800 13105 -795 13145
rect -755 13105 -750 13145
rect -800 2545 -750 13105
rect -800 2505 -795 2545
rect -755 2505 -750 2545
rect -800 0 -750 2505
rect -700 15345 -650 15700
rect -700 15305 -695 15345
rect -655 15305 -650 15345
rect -700 15295 -650 15305
rect -700 15255 -695 15295
rect -655 15255 -650 15295
rect -700 15245 -650 15255
rect -700 15205 -695 15245
rect -655 15205 -650 15245
rect -700 13645 -650 15205
rect -700 13605 -695 13645
rect -655 13605 -650 13645
rect -700 13595 -650 13605
rect -700 13555 -695 13595
rect -655 13555 -650 13595
rect -700 13545 -650 13555
rect -700 13505 -695 13545
rect -655 13505 -650 13545
rect -700 11945 -650 13505
rect -700 11905 -695 11945
rect -655 11905 -650 11945
rect -700 11895 -650 11905
rect -700 11855 -695 11895
rect -655 11855 -650 11895
rect -700 11845 -650 11855
rect -700 11805 -695 11845
rect -655 11805 -650 11845
rect -700 3845 -650 11805
rect -700 3805 -695 3845
rect -655 3805 -650 3845
rect -700 3795 -650 3805
rect -700 3755 -695 3795
rect -655 3755 -650 3795
rect -700 3745 -650 3755
rect -700 3705 -695 3745
rect -655 3705 -650 3745
rect -700 2145 -650 3705
rect -700 2105 -695 2145
rect -655 2105 -650 2145
rect -700 2095 -650 2105
rect -700 2055 -695 2095
rect -655 2055 -650 2095
rect -700 2045 -650 2055
rect -700 2005 -695 2045
rect -655 2005 -650 2045
rect -700 445 -650 2005
rect -700 405 -695 445
rect -655 405 -650 445
rect -700 395 -650 405
rect -700 355 -695 395
rect -655 355 -650 395
rect -700 345 -650 355
rect -700 305 -695 345
rect -655 305 -650 345
rect -700 0 -650 305
rect -600 14045 -550 15650
rect -600 14005 -595 14045
rect -555 14005 -550 14045
rect -600 1645 -550 14005
rect -600 1605 -595 1645
rect -555 1605 -550 1645
rect -600 0 -550 1605
rect -500 15345 -450 15700
rect -500 15305 -495 15345
rect -455 15305 -450 15345
rect -500 15295 -450 15305
rect -500 15255 -495 15295
rect -455 15255 -450 15295
rect -500 15245 -450 15255
rect -500 15205 -495 15245
rect -455 15205 -450 15245
rect -500 13645 -450 15205
rect -500 13605 -495 13645
rect -455 13605 -450 13645
rect -500 13595 -450 13605
rect -500 13555 -495 13595
rect -455 13555 -450 13595
rect -500 13545 -450 13555
rect -500 13505 -495 13545
rect -455 13505 -450 13545
rect -500 11945 -450 13505
rect -500 11905 -495 11945
rect -455 11905 -450 11945
rect -500 11895 -450 11905
rect -500 11855 -495 11895
rect -455 11855 -450 11895
rect -500 11845 -450 11855
rect -500 11805 -495 11845
rect -455 11805 -450 11845
rect -500 3845 -450 11805
rect -500 3805 -495 3845
rect -455 3805 -450 3845
rect -500 3795 -450 3805
rect -500 3755 -495 3795
rect -455 3755 -450 3795
rect -500 3745 -450 3755
rect -500 3705 -495 3745
rect -455 3705 -450 3745
rect -500 2145 -450 3705
rect -500 2105 -495 2145
rect -455 2105 -450 2145
rect -500 2095 -450 2105
rect -500 2055 -495 2095
rect -455 2055 -450 2095
rect -500 2045 -450 2055
rect -500 2005 -495 2045
rect -455 2005 -450 2045
rect -500 445 -450 2005
rect -500 405 -495 445
rect -455 405 -450 445
rect -500 395 -450 405
rect -500 355 -495 395
rect -455 355 -450 395
rect -500 345 -450 355
rect -500 305 -495 345
rect -455 305 -450 345
rect -500 0 -450 305
rect -400 16845 -350 16850
rect -400 16805 -395 16845
rect -355 16805 -350 16845
rect -400 14245 -350 16805
rect -400 14205 -395 14245
rect -355 14205 -350 14245
rect -400 1445 -350 14205
rect -400 1405 -395 1445
rect -355 1405 -350 1445
rect -400 0 -350 1405
rect -300 15750 -250 16900
rect -200 15750 -150 16900
rect -100 15750 -50 16900
rect -300 15745 -50 15750
rect -300 15705 -295 15745
rect -255 15705 -195 15745
rect -155 15705 -95 15745
rect -55 15705 -50 15745
rect -300 15700 -50 15705
rect 0 18145 39750 18150
rect 0 18105 5 18145
rect 45 18105 55 18145
rect 95 18105 105 18145
rect 145 18105 155 18145
rect 195 18105 205 18145
rect 245 18105 255 18145
rect 295 18105 305 18145
rect 345 18105 355 18145
rect 395 18105 405 18145
rect 445 18105 455 18145
rect 495 18105 505 18145
rect 545 18105 555 18145
rect 595 18105 605 18145
rect 645 18105 655 18145
rect 695 18105 705 18145
rect 745 18105 755 18145
rect 795 18105 805 18145
rect 845 18105 855 18145
rect 895 18105 905 18145
rect 945 18105 955 18145
rect 995 18105 1005 18145
rect 1045 18105 1055 18145
rect 1095 18105 1105 18145
rect 1145 18105 1155 18145
rect 1195 18105 1205 18145
rect 1245 18105 1255 18145
rect 1295 18105 1305 18145
rect 1345 18105 1355 18145
rect 1395 18105 1405 18145
rect 1445 18105 1455 18145
rect 1495 18105 1505 18145
rect 1545 18105 1555 18145
rect 1595 18105 1605 18145
rect 1645 18105 1655 18145
rect 1695 18105 1705 18145
rect 1745 18105 1755 18145
rect 1795 18105 1805 18145
rect 1845 18105 1855 18145
rect 1895 18105 1905 18145
rect 1945 18105 1955 18145
rect 1995 18105 2005 18145
rect 2045 18105 2055 18145
rect 2095 18105 2105 18145
rect 2145 18105 2155 18145
rect 2195 18105 2205 18145
rect 2245 18105 2255 18145
rect 2295 18105 2305 18145
rect 2345 18105 2355 18145
rect 2395 18105 2405 18145
rect 2445 18105 2455 18145
rect 2495 18105 2505 18145
rect 2545 18105 2555 18145
rect 2595 18105 2605 18145
rect 2645 18105 2655 18145
rect 2695 18105 2705 18145
rect 2745 18105 2755 18145
rect 2795 18105 2805 18145
rect 2845 18105 2855 18145
rect 2895 18105 2905 18145
rect 2945 18105 2955 18145
rect 2995 18105 3005 18145
rect 3045 18105 3055 18145
rect 3095 18105 3105 18145
rect 3145 18105 3155 18145
rect 3195 18105 3205 18145
rect 3245 18105 3255 18145
rect 3295 18105 3305 18145
rect 3345 18105 3355 18145
rect 3395 18105 3405 18145
rect 3445 18105 3455 18145
rect 3495 18105 3505 18145
rect 3545 18105 3555 18145
rect 3595 18105 3605 18145
rect 3645 18105 3655 18145
rect 3695 18105 3705 18145
rect 3745 18105 3755 18145
rect 3795 18105 3805 18145
rect 3845 18105 3855 18145
rect 3895 18105 3905 18145
rect 3945 18105 3955 18145
rect 3995 18105 4005 18145
rect 4045 18105 4055 18145
rect 4095 18105 4105 18145
rect 4145 18105 4155 18145
rect 4195 18105 4205 18145
rect 4245 18105 4255 18145
rect 4295 18105 4305 18145
rect 4345 18105 4355 18145
rect 4395 18105 4405 18145
rect 4445 18105 4455 18145
rect 4495 18105 4505 18145
rect 4545 18105 4555 18145
rect 4595 18105 4605 18145
rect 4645 18105 4655 18145
rect 4695 18105 4705 18145
rect 4745 18105 4755 18145
rect 4795 18105 4805 18145
rect 4845 18105 4855 18145
rect 4895 18105 4905 18145
rect 4945 18105 4955 18145
rect 4995 18105 5005 18145
rect 5045 18105 5055 18145
rect 5095 18105 5105 18145
rect 5145 18105 5155 18145
rect 5195 18105 5205 18145
rect 5245 18105 5255 18145
rect 5295 18105 5305 18145
rect 5345 18105 5355 18145
rect 5395 18105 5405 18145
rect 5445 18105 5455 18145
rect 5495 18105 5505 18145
rect 5545 18105 5555 18145
rect 5595 18105 5605 18145
rect 5645 18105 5655 18145
rect 5695 18105 5705 18145
rect 5745 18105 5755 18145
rect 5795 18105 5805 18145
rect 5845 18105 5855 18145
rect 5895 18105 5905 18145
rect 5945 18105 5955 18145
rect 5995 18105 6005 18145
rect 6045 18105 6055 18145
rect 6095 18105 6105 18145
rect 6145 18105 6155 18145
rect 6195 18105 6205 18145
rect 6245 18105 6255 18145
rect 6295 18105 6305 18145
rect 6345 18105 6355 18145
rect 6395 18105 6405 18145
rect 6445 18105 6455 18145
rect 6495 18105 6505 18145
rect 6545 18105 6555 18145
rect 6595 18105 6605 18145
rect 6645 18105 6655 18145
rect 6695 18105 6705 18145
rect 6745 18105 6755 18145
rect 6795 18105 6805 18145
rect 6845 18105 6855 18145
rect 6895 18105 6905 18145
rect 6945 18105 6955 18145
rect 6995 18105 7005 18145
rect 7045 18105 7055 18145
rect 7095 18105 7105 18145
rect 7145 18105 7155 18145
rect 7195 18105 7205 18145
rect 7245 18105 7255 18145
rect 7295 18105 7305 18145
rect 7345 18105 7355 18145
rect 7395 18105 7405 18145
rect 7445 18105 7455 18145
rect 7495 18105 7505 18145
rect 7545 18105 7555 18145
rect 7595 18105 7605 18145
rect 7645 18105 7655 18145
rect 7695 18105 7705 18145
rect 7745 18105 7755 18145
rect 7795 18105 7805 18145
rect 7845 18105 7855 18145
rect 7895 18105 7905 18145
rect 7945 18105 7955 18145
rect 7995 18105 8005 18145
rect 8045 18105 8055 18145
rect 8095 18105 8105 18145
rect 8145 18105 8155 18145
rect 8195 18105 8205 18145
rect 8245 18105 8255 18145
rect 8295 18105 8305 18145
rect 8345 18105 8355 18145
rect 8395 18105 8405 18145
rect 8445 18105 8455 18145
rect 8495 18105 8505 18145
rect 8545 18105 8555 18145
rect 8595 18105 8605 18145
rect 8645 18105 8655 18145
rect 8695 18105 8705 18145
rect 8745 18105 8755 18145
rect 8795 18105 8805 18145
rect 8845 18105 8855 18145
rect 8895 18105 8905 18145
rect 8945 18105 8955 18145
rect 8995 18105 9005 18145
rect 9045 18105 9055 18145
rect 9095 18105 9105 18145
rect 9145 18105 9155 18145
rect 9195 18105 9205 18145
rect 9245 18105 9255 18145
rect 9295 18105 9305 18145
rect 9345 18105 9355 18145
rect 9395 18105 9405 18145
rect 9445 18105 9455 18145
rect 9495 18105 9505 18145
rect 9545 18105 9555 18145
rect 9595 18105 9605 18145
rect 9645 18105 9655 18145
rect 9695 18105 9705 18145
rect 9745 18105 9755 18145
rect 9795 18105 9805 18145
rect 9845 18105 9855 18145
rect 9895 18105 9905 18145
rect 9945 18105 9955 18145
rect 9995 18105 10005 18145
rect 10045 18105 10055 18145
rect 10095 18105 10105 18145
rect 10145 18105 10155 18145
rect 10195 18105 10205 18145
rect 10245 18105 10255 18145
rect 10295 18105 10305 18145
rect 10345 18105 10355 18145
rect 10395 18105 10405 18145
rect 10445 18105 10455 18145
rect 10495 18105 10505 18145
rect 10545 18105 10555 18145
rect 10595 18105 10605 18145
rect 10645 18105 10655 18145
rect 10695 18105 10705 18145
rect 10745 18105 10755 18145
rect 10795 18105 10805 18145
rect 10845 18105 10855 18145
rect 10895 18105 10905 18145
rect 10945 18105 10955 18145
rect 10995 18105 11005 18145
rect 11045 18105 11055 18145
rect 11095 18105 11105 18145
rect 11145 18105 11155 18145
rect 11195 18105 11205 18145
rect 11245 18105 11255 18145
rect 11295 18105 11305 18145
rect 11345 18105 11355 18145
rect 11395 18105 11405 18145
rect 11445 18105 11455 18145
rect 11495 18105 11505 18145
rect 11545 18105 11555 18145
rect 11595 18105 11605 18145
rect 11645 18105 11655 18145
rect 11695 18105 11705 18145
rect 11745 18105 11755 18145
rect 11795 18105 11805 18145
rect 11845 18105 11855 18145
rect 11895 18105 11905 18145
rect 11945 18105 11955 18145
rect 11995 18105 12005 18145
rect 12045 18105 12055 18145
rect 12095 18105 12105 18145
rect 12145 18105 12155 18145
rect 12195 18105 12205 18145
rect 12245 18105 12255 18145
rect 12295 18105 12305 18145
rect 12345 18105 12355 18145
rect 12395 18105 12405 18145
rect 12445 18105 12455 18145
rect 12495 18105 12505 18145
rect 12545 18105 12555 18145
rect 12595 18105 12605 18145
rect 12645 18105 12655 18145
rect 12695 18105 12705 18145
rect 12745 18105 12755 18145
rect 12795 18105 12805 18145
rect 12845 18105 12855 18145
rect 12895 18105 12905 18145
rect 12945 18105 12955 18145
rect 12995 18105 13005 18145
rect 13045 18105 13055 18145
rect 13095 18105 13105 18145
rect 13145 18105 13155 18145
rect 13195 18105 13205 18145
rect 13245 18105 13255 18145
rect 13295 18105 13305 18145
rect 13345 18105 13355 18145
rect 13395 18105 13405 18145
rect 13445 18105 13455 18145
rect 13495 18105 13505 18145
rect 13545 18105 13555 18145
rect 13595 18105 13605 18145
rect 13645 18105 13655 18145
rect 13695 18105 13705 18145
rect 13745 18105 13755 18145
rect 13795 18105 13805 18145
rect 13845 18105 13855 18145
rect 13895 18105 13905 18145
rect 13945 18105 13955 18145
rect 13995 18105 14005 18145
rect 14045 18105 14055 18145
rect 14095 18105 14105 18145
rect 14145 18105 14155 18145
rect 14195 18105 14205 18145
rect 14245 18105 14255 18145
rect 14295 18105 14305 18145
rect 14345 18105 14355 18145
rect 14395 18105 14405 18145
rect 14445 18105 14455 18145
rect 14495 18105 14505 18145
rect 14545 18105 14555 18145
rect 14595 18105 14605 18145
rect 14645 18105 14655 18145
rect 14695 18105 14705 18145
rect 14745 18105 14755 18145
rect 14795 18105 14805 18145
rect 14845 18105 14855 18145
rect 14895 18105 14905 18145
rect 14945 18105 14955 18145
rect 14995 18105 15005 18145
rect 15045 18105 15055 18145
rect 15095 18105 15105 18145
rect 15145 18105 15155 18145
rect 15195 18105 15205 18145
rect 15245 18105 15255 18145
rect 15295 18105 15305 18145
rect 15345 18105 15355 18145
rect 15395 18105 15405 18145
rect 15445 18105 15455 18145
rect 15495 18105 15505 18145
rect 15545 18105 15555 18145
rect 15595 18105 15605 18145
rect 15645 18105 15655 18145
rect 15695 18105 15705 18145
rect 15745 18105 15755 18145
rect 15795 18105 15805 18145
rect 15845 18105 15855 18145
rect 15895 18105 15905 18145
rect 15945 18105 15955 18145
rect 15995 18105 16005 18145
rect 16045 18105 16055 18145
rect 16095 18105 16105 18145
rect 16145 18105 16155 18145
rect 16195 18105 16205 18145
rect 16245 18105 16255 18145
rect 16295 18105 16305 18145
rect 16345 18105 16355 18145
rect 16395 18105 16405 18145
rect 16445 18105 16455 18145
rect 16495 18105 16505 18145
rect 16545 18105 16555 18145
rect 16595 18105 16605 18145
rect 16645 18105 16655 18145
rect 16695 18105 16705 18145
rect 16745 18105 16755 18145
rect 16795 18105 16805 18145
rect 16845 18105 16855 18145
rect 16895 18105 16905 18145
rect 16945 18105 16955 18145
rect 16995 18105 17005 18145
rect 17045 18105 17055 18145
rect 17095 18105 17105 18145
rect 17145 18105 17155 18145
rect 17195 18105 17205 18145
rect 17245 18105 17255 18145
rect 17295 18105 17305 18145
rect 17345 18105 17355 18145
rect 17395 18105 17405 18145
rect 17445 18105 17455 18145
rect 17495 18105 17505 18145
rect 17545 18105 17555 18145
rect 17595 18105 17605 18145
rect 17645 18105 17655 18145
rect 17695 18105 17705 18145
rect 17745 18105 17755 18145
rect 17795 18105 17805 18145
rect 17845 18105 17855 18145
rect 17895 18105 17905 18145
rect 17945 18105 17955 18145
rect 17995 18105 18005 18145
rect 18045 18105 18055 18145
rect 18095 18105 18105 18145
rect 18145 18105 18155 18145
rect 18195 18105 18205 18145
rect 18245 18105 18255 18145
rect 18295 18105 18305 18145
rect 18345 18105 18355 18145
rect 18395 18105 18405 18145
rect 18445 18105 18455 18145
rect 18495 18105 18505 18145
rect 18545 18105 18555 18145
rect 18595 18105 18605 18145
rect 18645 18105 18655 18145
rect 18695 18105 18705 18145
rect 18745 18105 18755 18145
rect 18795 18105 18805 18145
rect 18845 18105 18855 18145
rect 18895 18105 18905 18145
rect 18945 18105 18955 18145
rect 18995 18105 19005 18145
rect 19045 18105 19055 18145
rect 19095 18105 19105 18145
rect 19145 18105 19155 18145
rect 19195 18105 19205 18145
rect 19245 18105 19255 18145
rect 19295 18105 19305 18145
rect 19345 18105 19355 18145
rect 19395 18105 19405 18145
rect 19445 18105 19455 18145
rect 19495 18105 19505 18145
rect 19545 18105 19555 18145
rect 19595 18105 19605 18145
rect 19645 18105 19655 18145
rect 19695 18105 19705 18145
rect 19745 18105 19755 18145
rect 19795 18105 19805 18145
rect 19845 18105 19855 18145
rect 19895 18105 19905 18145
rect 19945 18105 19955 18145
rect 19995 18105 20005 18145
rect 20045 18105 20055 18145
rect 20095 18105 20105 18145
rect 20145 18105 20155 18145
rect 20195 18105 20205 18145
rect 20245 18105 20255 18145
rect 20295 18105 20305 18145
rect 20345 18105 20355 18145
rect 20395 18105 20405 18145
rect 20445 18105 20455 18145
rect 20495 18105 20505 18145
rect 20545 18105 20555 18145
rect 20595 18105 20605 18145
rect 20645 18105 20655 18145
rect 20695 18105 20705 18145
rect 20745 18105 20755 18145
rect 20795 18105 20805 18145
rect 20845 18105 20855 18145
rect 20895 18105 20905 18145
rect 20945 18105 20955 18145
rect 20995 18105 21005 18145
rect 21045 18105 21055 18145
rect 21095 18105 21105 18145
rect 21145 18105 21155 18145
rect 21195 18105 21205 18145
rect 21245 18105 21255 18145
rect 21295 18105 21305 18145
rect 21345 18105 21355 18145
rect 21395 18105 21405 18145
rect 21445 18105 21455 18145
rect 21495 18105 21505 18145
rect 21545 18105 21555 18145
rect 21595 18105 21605 18145
rect 21645 18105 21655 18145
rect 21695 18105 21705 18145
rect 21745 18105 21755 18145
rect 21795 18105 21805 18145
rect 21845 18105 21855 18145
rect 21895 18105 21905 18145
rect 21945 18105 21955 18145
rect 21995 18105 22005 18145
rect 22045 18105 22055 18145
rect 22095 18105 22105 18145
rect 22145 18105 22155 18145
rect 22195 18105 22205 18145
rect 22245 18105 22255 18145
rect 22295 18105 22305 18145
rect 22345 18105 22355 18145
rect 22395 18105 22405 18145
rect 22445 18105 22455 18145
rect 22495 18105 22505 18145
rect 22545 18105 22555 18145
rect 22595 18105 22605 18145
rect 22645 18105 22655 18145
rect 22695 18105 22705 18145
rect 22745 18105 22755 18145
rect 22795 18105 22805 18145
rect 22845 18105 22855 18145
rect 22895 18105 22905 18145
rect 22945 18105 22955 18145
rect 22995 18105 23005 18145
rect 23045 18105 23055 18145
rect 23095 18105 23105 18145
rect 23145 18105 23155 18145
rect 23195 18105 23205 18145
rect 23245 18105 23255 18145
rect 23295 18105 23305 18145
rect 23345 18105 23355 18145
rect 23395 18105 23405 18145
rect 23445 18105 23455 18145
rect 23495 18105 23505 18145
rect 23545 18105 23555 18145
rect 23595 18105 23605 18145
rect 23645 18105 23655 18145
rect 23695 18105 23705 18145
rect 23745 18105 23755 18145
rect 23795 18105 23805 18145
rect 23845 18105 23855 18145
rect 23895 18105 23905 18145
rect 23945 18105 23955 18145
rect 23995 18105 24005 18145
rect 24045 18105 24055 18145
rect 24095 18105 24105 18145
rect 24145 18105 24155 18145
rect 24195 18105 24205 18145
rect 24245 18105 24255 18145
rect 24295 18105 24305 18145
rect 24345 18105 24355 18145
rect 24395 18105 24405 18145
rect 24445 18105 24455 18145
rect 24495 18105 24505 18145
rect 24545 18105 24555 18145
rect 24595 18105 24605 18145
rect 24645 18105 24655 18145
rect 24695 18105 24705 18145
rect 24745 18105 24755 18145
rect 24795 18105 24805 18145
rect 24845 18105 24855 18145
rect 24895 18105 24905 18145
rect 24945 18105 24955 18145
rect 24995 18105 25005 18145
rect 25045 18105 25055 18145
rect 25095 18105 25105 18145
rect 25145 18105 25155 18145
rect 25195 18105 25205 18145
rect 25245 18105 25255 18145
rect 25295 18105 25305 18145
rect 25345 18105 25355 18145
rect 25395 18105 25405 18145
rect 25445 18105 25455 18145
rect 25495 18105 25505 18145
rect 25545 18105 25555 18145
rect 25595 18105 25605 18145
rect 25645 18105 25655 18145
rect 25695 18105 25705 18145
rect 25745 18105 25755 18145
rect 25795 18105 25805 18145
rect 25845 18105 25855 18145
rect 25895 18105 25905 18145
rect 25945 18105 25955 18145
rect 25995 18105 26005 18145
rect 26045 18105 26055 18145
rect 26095 18105 26105 18145
rect 26145 18105 26155 18145
rect 26195 18105 26205 18145
rect 26245 18105 26255 18145
rect 26295 18105 26305 18145
rect 26345 18105 26355 18145
rect 26395 18105 26405 18145
rect 26445 18105 26455 18145
rect 26495 18105 26505 18145
rect 26545 18105 26555 18145
rect 26595 18105 26605 18145
rect 26645 18105 26655 18145
rect 26695 18105 26705 18145
rect 26745 18105 26755 18145
rect 26795 18105 26805 18145
rect 26845 18105 26855 18145
rect 26895 18105 26905 18145
rect 26945 18105 26955 18145
rect 26995 18105 27005 18145
rect 27045 18105 27055 18145
rect 27095 18105 27105 18145
rect 27145 18105 27155 18145
rect 27195 18105 27205 18145
rect 27245 18105 27255 18145
rect 27295 18105 27305 18145
rect 27345 18105 27355 18145
rect 27395 18105 27405 18145
rect 27445 18105 27455 18145
rect 27495 18105 27505 18145
rect 27545 18105 27555 18145
rect 27595 18105 27605 18145
rect 27645 18105 27655 18145
rect 27695 18105 27705 18145
rect 27745 18105 27755 18145
rect 27795 18105 27805 18145
rect 27845 18105 27855 18145
rect 27895 18105 27905 18145
rect 27945 18105 27955 18145
rect 27995 18105 28005 18145
rect 28045 18105 28055 18145
rect 28095 18105 28105 18145
rect 28145 18105 28155 18145
rect 28195 18105 28205 18145
rect 28245 18105 28255 18145
rect 28295 18105 28305 18145
rect 28345 18105 28355 18145
rect 28395 18105 28405 18145
rect 28445 18105 28455 18145
rect 28495 18105 28505 18145
rect 28545 18105 28555 18145
rect 28595 18105 28605 18145
rect 28645 18105 28655 18145
rect 28695 18105 28705 18145
rect 28745 18105 28755 18145
rect 28795 18105 28805 18145
rect 28845 18105 28855 18145
rect 28895 18105 28905 18145
rect 28945 18105 28955 18145
rect 28995 18105 29005 18145
rect 29045 18105 29055 18145
rect 29095 18105 29105 18145
rect 29145 18105 29155 18145
rect 29195 18105 29205 18145
rect 29245 18105 29255 18145
rect 29295 18105 29305 18145
rect 29345 18105 29355 18145
rect 29395 18105 29405 18145
rect 29445 18105 29455 18145
rect 29495 18105 29505 18145
rect 29545 18105 29555 18145
rect 29595 18105 29605 18145
rect 29645 18105 29655 18145
rect 29695 18105 29705 18145
rect 29745 18105 29755 18145
rect 29795 18105 29805 18145
rect 29845 18105 29855 18145
rect 29895 18105 29905 18145
rect 29945 18105 29955 18145
rect 29995 18105 30005 18145
rect 30045 18105 30055 18145
rect 30095 18105 30105 18145
rect 30145 18105 30155 18145
rect 30195 18105 30205 18145
rect 30245 18105 30255 18145
rect 30295 18105 30305 18145
rect 30345 18105 30355 18145
rect 30395 18105 30405 18145
rect 30445 18105 30455 18145
rect 30495 18105 30505 18145
rect 30545 18105 30555 18145
rect 30595 18105 30605 18145
rect 30645 18105 30655 18145
rect 30695 18105 30705 18145
rect 30745 18105 30755 18145
rect 30795 18105 30805 18145
rect 30845 18105 30855 18145
rect 30895 18105 30905 18145
rect 30945 18105 30955 18145
rect 30995 18105 31005 18145
rect 31045 18105 31055 18145
rect 31095 18105 31105 18145
rect 31145 18105 31155 18145
rect 31195 18105 31205 18145
rect 31245 18105 31255 18145
rect 31295 18105 31305 18145
rect 31345 18105 31355 18145
rect 31395 18105 31405 18145
rect 31445 18105 31455 18145
rect 31495 18105 31505 18145
rect 31545 18105 31555 18145
rect 31595 18105 31605 18145
rect 31645 18105 31655 18145
rect 31695 18105 31705 18145
rect 31745 18105 31755 18145
rect 31795 18105 31805 18145
rect 31845 18105 31855 18145
rect 31895 18105 31905 18145
rect 31945 18105 31955 18145
rect 31995 18105 32005 18145
rect 32045 18105 32055 18145
rect 32095 18105 32105 18145
rect 32145 18105 32155 18145
rect 32195 18105 32205 18145
rect 32245 18105 32255 18145
rect 32295 18105 32305 18145
rect 32345 18105 32355 18145
rect 32395 18105 32405 18145
rect 32445 18105 32455 18145
rect 32495 18105 32505 18145
rect 32545 18105 32555 18145
rect 32595 18105 32605 18145
rect 32645 18105 32655 18145
rect 32695 18105 32705 18145
rect 32745 18105 32755 18145
rect 32795 18105 32805 18145
rect 32845 18105 32855 18145
rect 32895 18105 32905 18145
rect 32945 18105 32955 18145
rect 32995 18105 33005 18145
rect 33045 18105 33055 18145
rect 33095 18105 33105 18145
rect 33145 18105 33155 18145
rect 33195 18105 33205 18145
rect 33245 18105 33255 18145
rect 33295 18105 33305 18145
rect 33345 18105 33355 18145
rect 33395 18105 33405 18145
rect 33445 18105 33455 18145
rect 33495 18105 33505 18145
rect 33545 18105 33555 18145
rect 33595 18105 33605 18145
rect 33645 18105 33655 18145
rect 33695 18105 33705 18145
rect 33745 18105 33755 18145
rect 33795 18105 33805 18145
rect 33845 18105 33855 18145
rect 33895 18105 33905 18145
rect 33945 18105 33955 18145
rect 33995 18105 34005 18145
rect 34045 18105 34055 18145
rect 34095 18105 34105 18145
rect 34145 18105 34155 18145
rect 34195 18105 34205 18145
rect 34245 18105 34255 18145
rect 34295 18105 34305 18145
rect 34345 18105 34355 18145
rect 34395 18105 34405 18145
rect 34445 18105 34455 18145
rect 34495 18105 34505 18145
rect 34545 18105 34555 18145
rect 34595 18105 34605 18145
rect 34645 18105 34655 18145
rect 34695 18105 34705 18145
rect 34745 18105 34755 18145
rect 34795 18105 34805 18145
rect 34845 18105 34855 18145
rect 34895 18105 34905 18145
rect 34945 18105 34955 18145
rect 34995 18105 35005 18145
rect 35045 18105 35055 18145
rect 35095 18105 35105 18145
rect 35145 18105 35155 18145
rect 35195 18105 35205 18145
rect 35245 18105 35255 18145
rect 35295 18105 35305 18145
rect 35345 18105 35355 18145
rect 35395 18105 35405 18145
rect 35445 18105 35455 18145
rect 35495 18105 35505 18145
rect 35545 18105 35555 18145
rect 35595 18105 35605 18145
rect 35645 18105 35655 18145
rect 35695 18105 35705 18145
rect 35745 18105 35755 18145
rect 35795 18105 35805 18145
rect 35845 18105 35855 18145
rect 35895 18105 35905 18145
rect 35945 18105 35955 18145
rect 35995 18105 36005 18145
rect 36045 18105 36055 18145
rect 36095 18105 36105 18145
rect 36145 18105 36155 18145
rect 36195 18105 36205 18145
rect 36245 18105 36255 18145
rect 36295 18105 36305 18145
rect 36345 18105 36355 18145
rect 36395 18105 36405 18145
rect 36445 18105 36455 18145
rect 36495 18105 36505 18145
rect 36545 18105 36555 18145
rect 36595 18105 36605 18145
rect 36645 18105 36655 18145
rect 36695 18105 36705 18145
rect 36745 18105 36755 18145
rect 36795 18105 36805 18145
rect 36845 18105 36855 18145
rect 36895 18105 36905 18145
rect 36945 18105 36955 18145
rect 36995 18105 37005 18145
rect 37045 18105 37055 18145
rect 37095 18105 37105 18145
rect 37145 18105 37155 18145
rect 37195 18105 37205 18145
rect 37245 18105 37255 18145
rect 37295 18105 37305 18145
rect 37345 18105 37355 18145
rect 37395 18105 37405 18145
rect 37445 18105 37455 18145
rect 37495 18105 37505 18145
rect 37545 18105 37555 18145
rect 37595 18105 37605 18145
rect 37645 18105 37655 18145
rect 37695 18105 37705 18145
rect 37745 18105 37755 18145
rect 37795 18105 37805 18145
rect 37845 18105 37855 18145
rect 37895 18105 37905 18145
rect 37945 18105 37955 18145
rect 37995 18105 38005 18145
rect 38045 18105 38055 18145
rect 38095 18105 38105 18145
rect 38145 18105 38155 18145
rect 38195 18105 38205 18145
rect 38245 18105 38255 18145
rect 38295 18105 38305 18145
rect 38345 18105 38355 18145
rect 38395 18105 38405 18145
rect 38445 18105 38455 18145
rect 38495 18105 38505 18145
rect 38545 18105 38555 18145
rect 38595 18105 38605 18145
rect 38645 18105 38655 18145
rect 38695 18105 38705 18145
rect 38745 18105 38755 18145
rect 38795 18105 38805 18145
rect 38845 18105 38855 18145
rect 38895 18105 38905 18145
rect 38945 18105 38955 18145
rect 38995 18105 39005 18145
rect 39045 18105 39055 18145
rect 39095 18105 39105 18145
rect 39145 18105 39155 18145
rect 39195 18105 39205 18145
rect 39245 18105 39255 18145
rect 39295 18105 39305 18145
rect 39345 18105 39355 18145
rect 39395 18105 39405 18145
rect 39445 18105 39455 18145
rect 39495 18105 39505 18145
rect 39545 18105 39555 18145
rect 39595 18105 39605 18145
rect 39645 18105 39655 18145
rect 39695 18105 39705 18145
rect 39745 18105 39750 18145
rect 0 18045 39750 18105
rect 0 18005 5 18045
rect 45 18005 55 18045
rect 95 18005 105 18045
rect 145 18005 155 18045
rect 195 18005 205 18045
rect 245 18005 255 18045
rect 295 18005 305 18045
rect 345 18005 355 18045
rect 395 18005 405 18045
rect 445 18005 455 18045
rect 495 18005 505 18045
rect 545 18005 555 18045
rect 595 18005 605 18045
rect 645 18005 655 18045
rect 695 18005 705 18045
rect 745 18005 755 18045
rect 795 18005 805 18045
rect 845 18005 855 18045
rect 895 18005 905 18045
rect 945 18005 955 18045
rect 995 18005 1005 18045
rect 1045 18005 1055 18045
rect 1095 18005 1105 18045
rect 1145 18005 1155 18045
rect 1195 18005 1205 18045
rect 1245 18005 1255 18045
rect 1295 18005 1305 18045
rect 1345 18005 1355 18045
rect 1395 18005 1405 18045
rect 1445 18005 1455 18045
rect 1495 18005 1505 18045
rect 1545 18005 1555 18045
rect 1595 18005 1605 18045
rect 1645 18005 1655 18045
rect 1695 18005 1705 18045
rect 1745 18005 1755 18045
rect 1795 18005 1805 18045
rect 1845 18005 1855 18045
rect 1895 18005 1905 18045
rect 1945 18005 1955 18045
rect 1995 18005 2005 18045
rect 2045 18005 2055 18045
rect 2095 18005 2105 18045
rect 2145 18005 2155 18045
rect 2195 18005 2205 18045
rect 2245 18005 2255 18045
rect 2295 18005 2305 18045
rect 2345 18005 2355 18045
rect 2395 18005 2405 18045
rect 2445 18005 2455 18045
rect 2495 18005 2505 18045
rect 2545 18005 2555 18045
rect 2595 18005 2605 18045
rect 2645 18005 2655 18045
rect 2695 18005 2705 18045
rect 2745 18005 2755 18045
rect 2795 18005 2805 18045
rect 2845 18005 2855 18045
rect 2895 18005 2905 18045
rect 2945 18005 2955 18045
rect 2995 18005 3005 18045
rect 3045 18005 3055 18045
rect 3095 18005 3105 18045
rect 3145 18005 3155 18045
rect 3195 18005 3205 18045
rect 3245 18005 3255 18045
rect 3295 18005 3305 18045
rect 3345 18005 3355 18045
rect 3395 18005 3405 18045
rect 3445 18005 3455 18045
rect 3495 18005 3505 18045
rect 3545 18005 3555 18045
rect 3595 18005 3605 18045
rect 3645 18005 3655 18045
rect 3695 18005 3705 18045
rect 3745 18005 3755 18045
rect 3795 18005 3805 18045
rect 3845 18005 3855 18045
rect 3895 18005 3905 18045
rect 3945 18005 3955 18045
rect 3995 18005 4005 18045
rect 4045 18005 4055 18045
rect 4095 18005 4105 18045
rect 4145 18005 4155 18045
rect 4195 18005 4205 18045
rect 4245 18005 4255 18045
rect 4295 18005 4305 18045
rect 4345 18005 4355 18045
rect 4395 18005 4405 18045
rect 4445 18005 4455 18045
rect 4495 18005 4505 18045
rect 4545 18005 4555 18045
rect 4595 18005 4605 18045
rect 4645 18005 4655 18045
rect 4695 18005 4705 18045
rect 4745 18005 4755 18045
rect 4795 18005 4805 18045
rect 4845 18005 4855 18045
rect 4895 18005 4905 18045
rect 4945 18005 4955 18045
rect 4995 18005 5005 18045
rect 5045 18005 5055 18045
rect 5095 18005 5105 18045
rect 5145 18005 5155 18045
rect 5195 18005 5205 18045
rect 5245 18005 5255 18045
rect 5295 18005 5305 18045
rect 5345 18005 5355 18045
rect 5395 18005 5405 18045
rect 5445 18005 5455 18045
rect 5495 18005 5505 18045
rect 5545 18005 5555 18045
rect 5595 18005 5605 18045
rect 5645 18005 5655 18045
rect 5695 18005 5705 18045
rect 5745 18005 5755 18045
rect 5795 18005 5805 18045
rect 5845 18005 5855 18045
rect 5895 18005 5905 18045
rect 5945 18005 5955 18045
rect 5995 18005 6005 18045
rect 6045 18005 6055 18045
rect 6095 18005 6105 18045
rect 6145 18005 6155 18045
rect 6195 18005 6205 18045
rect 6245 18005 6255 18045
rect 6295 18005 6305 18045
rect 6345 18005 6355 18045
rect 6395 18005 6405 18045
rect 6445 18005 6455 18045
rect 6495 18005 6505 18045
rect 6545 18005 6555 18045
rect 6595 18005 6605 18045
rect 6645 18005 6655 18045
rect 6695 18005 6705 18045
rect 6745 18005 6755 18045
rect 6795 18005 6805 18045
rect 6845 18005 6855 18045
rect 6895 18005 6905 18045
rect 6945 18005 6955 18045
rect 6995 18005 7005 18045
rect 7045 18005 7055 18045
rect 7095 18005 7105 18045
rect 7145 18005 7155 18045
rect 7195 18005 7205 18045
rect 7245 18005 7255 18045
rect 7295 18005 7305 18045
rect 7345 18005 7355 18045
rect 7395 18005 7405 18045
rect 7445 18005 7455 18045
rect 7495 18005 7505 18045
rect 7545 18005 7555 18045
rect 7595 18005 7605 18045
rect 7645 18005 7655 18045
rect 7695 18005 7705 18045
rect 7745 18005 7755 18045
rect 7795 18005 7805 18045
rect 7845 18005 7855 18045
rect 7895 18005 7905 18045
rect 7945 18005 7955 18045
rect 7995 18005 8005 18045
rect 8045 18005 8055 18045
rect 8095 18005 8105 18045
rect 8145 18005 8155 18045
rect 8195 18005 8205 18045
rect 8245 18005 8255 18045
rect 8295 18005 8305 18045
rect 8345 18005 8355 18045
rect 8395 18005 8405 18045
rect 8445 18005 8455 18045
rect 8495 18005 8505 18045
rect 8545 18005 8555 18045
rect 8595 18005 8605 18045
rect 8645 18005 8655 18045
rect 8695 18005 8705 18045
rect 8745 18005 8755 18045
rect 8795 18005 8805 18045
rect 8845 18005 8855 18045
rect 8895 18005 8905 18045
rect 8945 18005 8955 18045
rect 8995 18005 9005 18045
rect 9045 18005 9055 18045
rect 9095 18005 9105 18045
rect 9145 18005 9155 18045
rect 9195 18005 9205 18045
rect 9245 18005 9255 18045
rect 9295 18005 9305 18045
rect 9345 18005 9355 18045
rect 9395 18005 9405 18045
rect 9445 18005 9455 18045
rect 9495 18005 9505 18045
rect 9545 18005 9555 18045
rect 9595 18005 9605 18045
rect 9645 18005 9655 18045
rect 9695 18005 9705 18045
rect 9745 18005 9755 18045
rect 9795 18005 9805 18045
rect 9845 18005 9855 18045
rect 9895 18005 9905 18045
rect 9945 18005 9955 18045
rect 9995 18005 10005 18045
rect 10045 18005 10055 18045
rect 10095 18005 10105 18045
rect 10145 18005 10155 18045
rect 10195 18005 10205 18045
rect 10245 18005 10255 18045
rect 10295 18005 10305 18045
rect 10345 18005 10355 18045
rect 10395 18005 10405 18045
rect 10445 18005 10455 18045
rect 10495 18005 10505 18045
rect 10545 18005 10555 18045
rect 10595 18005 10605 18045
rect 10645 18005 10655 18045
rect 10695 18005 10705 18045
rect 10745 18005 10755 18045
rect 10795 18005 10805 18045
rect 10845 18005 10855 18045
rect 10895 18005 10905 18045
rect 10945 18005 10955 18045
rect 10995 18005 11005 18045
rect 11045 18005 11055 18045
rect 11095 18005 11105 18045
rect 11145 18005 11155 18045
rect 11195 18005 11205 18045
rect 11245 18005 11255 18045
rect 11295 18005 11305 18045
rect 11345 18005 11355 18045
rect 11395 18005 11405 18045
rect 11445 18005 11455 18045
rect 11495 18005 11505 18045
rect 11545 18005 11555 18045
rect 11595 18005 11605 18045
rect 11645 18005 11655 18045
rect 11695 18005 11705 18045
rect 11745 18005 11755 18045
rect 11795 18005 11805 18045
rect 11845 18005 11855 18045
rect 11895 18005 11905 18045
rect 11945 18005 11955 18045
rect 11995 18005 12005 18045
rect 12045 18005 12055 18045
rect 12095 18005 12105 18045
rect 12145 18005 12155 18045
rect 12195 18005 12205 18045
rect 12245 18005 12255 18045
rect 12295 18005 12305 18045
rect 12345 18005 12355 18045
rect 12395 18005 12405 18045
rect 12445 18005 12455 18045
rect 12495 18005 12505 18045
rect 12545 18005 12555 18045
rect 12595 18005 12605 18045
rect 12645 18005 12655 18045
rect 12695 18005 12705 18045
rect 12745 18005 12755 18045
rect 12795 18005 12805 18045
rect 12845 18005 12855 18045
rect 12895 18005 12905 18045
rect 12945 18005 12955 18045
rect 12995 18005 13005 18045
rect 13045 18005 13055 18045
rect 13095 18005 13105 18045
rect 13145 18005 13155 18045
rect 13195 18005 13205 18045
rect 13245 18005 13255 18045
rect 13295 18005 13305 18045
rect 13345 18005 13355 18045
rect 13395 18005 13405 18045
rect 13445 18005 13455 18045
rect 13495 18005 13505 18045
rect 13545 18005 13555 18045
rect 13595 18005 13605 18045
rect 13645 18005 13655 18045
rect 13695 18005 13705 18045
rect 13745 18005 13755 18045
rect 13795 18005 13805 18045
rect 13845 18005 13855 18045
rect 13895 18005 13905 18045
rect 13945 18005 13955 18045
rect 13995 18005 14005 18045
rect 14045 18005 14055 18045
rect 14095 18005 14105 18045
rect 14145 18005 14155 18045
rect 14195 18005 14205 18045
rect 14245 18005 14255 18045
rect 14295 18005 14305 18045
rect 14345 18005 14355 18045
rect 14395 18005 14405 18045
rect 14445 18005 14455 18045
rect 14495 18005 14505 18045
rect 14545 18005 14555 18045
rect 14595 18005 14605 18045
rect 14645 18005 14655 18045
rect 14695 18005 14705 18045
rect 14745 18005 14755 18045
rect 14795 18005 14805 18045
rect 14845 18005 14855 18045
rect 14895 18005 14905 18045
rect 14945 18005 14955 18045
rect 14995 18005 15005 18045
rect 15045 18005 15055 18045
rect 15095 18005 15105 18045
rect 15145 18005 15155 18045
rect 15195 18005 15205 18045
rect 15245 18005 15255 18045
rect 15295 18005 15305 18045
rect 15345 18005 15355 18045
rect 15395 18005 15405 18045
rect 15445 18005 15455 18045
rect 15495 18005 15505 18045
rect 15545 18005 15555 18045
rect 15595 18005 15605 18045
rect 15645 18005 15655 18045
rect 15695 18005 15705 18045
rect 15745 18005 15755 18045
rect 15795 18005 15805 18045
rect 15845 18005 15855 18045
rect 15895 18005 15905 18045
rect 15945 18005 15955 18045
rect 15995 18005 16005 18045
rect 16045 18005 16055 18045
rect 16095 18005 16105 18045
rect 16145 18005 16155 18045
rect 16195 18005 16205 18045
rect 16245 18005 16255 18045
rect 16295 18005 16305 18045
rect 16345 18005 16355 18045
rect 16395 18005 16405 18045
rect 16445 18005 16455 18045
rect 16495 18005 16505 18045
rect 16545 18005 16555 18045
rect 16595 18005 16605 18045
rect 16645 18005 16655 18045
rect 16695 18005 16705 18045
rect 16745 18005 16755 18045
rect 16795 18005 16805 18045
rect 16845 18005 16855 18045
rect 16895 18005 16905 18045
rect 16945 18005 16955 18045
rect 16995 18005 17005 18045
rect 17045 18005 17055 18045
rect 17095 18005 17105 18045
rect 17145 18005 17155 18045
rect 17195 18005 17205 18045
rect 17245 18005 17255 18045
rect 17295 18005 17305 18045
rect 17345 18005 17355 18045
rect 17395 18005 17405 18045
rect 17445 18005 17455 18045
rect 17495 18005 17505 18045
rect 17545 18005 17555 18045
rect 17595 18005 17605 18045
rect 17645 18005 17655 18045
rect 17695 18005 17705 18045
rect 17745 18005 17755 18045
rect 17795 18005 17805 18045
rect 17845 18005 17855 18045
rect 17895 18005 17905 18045
rect 17945 18005 17955 18045
rect 17995 18005 18005 18045
rect 18045 18005 18055 18045
rect 18095 18005 18105 18045
rect 18145 18005 18155 18045
rect 18195 18005 18205 18045
rect 18245 18005 18255 18045
rect 18295 18005 18305 18045
rect 18345 18005 18355 18045
rect 18395 18005 18405 18045
rect 18445 18005 18455 18045
rect 18495 18005 18505 18045
rect 18545 18005 18555 18045
rect 18595 18005 18605 18045
rect 18645 18005 18655 18045
rect 18695 18005 18705 18045
rect 18745 18005 18755 18045
rect 18795 18005 18805 18045
rect 18845 18005 18855 18045
rect 18895 18005 18905 18045
rect 18945 18005 18955 18045
rect 18995 18005 19005 18045
rect 19045 18005 19055 18045
rect 19095 18005 19105 18045
rect 19145 18005 19155 18045
rect 19195 18005 19205 18045
rect 19245 18005 19255 18045
rect 19295 18005 19305 18045
rect 19345 18005 19355 18045
rect 19395 18005 19405 18045
rect 19445 18005 19455 18045
rect 19495 18005 19505 18045
rect 19545 18005 19555 18045
rect 19595 18005 19605 18045
rect 19645 18005 19655 18045
rect 19695 18005 19705 18045
rect 19745 18005 19755 18045
rect 19795 18005 19805 18045
rect 19845 18005 19855 18045
rect 19895 18005 19905 18045
rect 19945 18005 19955 18045
rect 19995 18005 20005 18045
rect 20045 18005 20055 18045
rect 20095 18005 20105 18045
rect 20145 18005 20155 18045
rect 20195 18005 20205 18045
rect 20245 18005 20255 18045
rect 20295 18005 20305 18045
rect 20345 18005 20355 18045
rect 20395 18005 20405 18045
rect 20445 18005 20455 18045
rect 20495 18005 20505 18045
rect 20545 18005 20555 18045
rect 20595 18005 20605 18045
rect 20645 18005 20655 18045
rect 20695 18005 20705 18045
rect 20745 18005 20755 18045
rect 20795 18005 20805 18045
rect 20845 18005 20855 18045
rect 20895 18005 20905 18045
rect 20945 18005 20955 18045
rect 20995 18005 21005 18045
rect 21045 18005 21055 18045
rect 21095 18005 21105 18045
rect 21145 18005 21155 18045
rect 21195 18005 21205 18045
rect 21245 18005 21255 18045
rect 21295 18005 21305 18045
rect 21345 18005 21355 18045
rect 21395 18005 21405 18045
rect 21445 18005 21455 18045
rect 21495 18005 21505 18045
rect 21545 18005 21555 18045
rect 21595 18005 21605 18045
rect 21645 18005 21655 18045
rect 21695 18005 21705 18045
rect 21745 18005 21755 18045
rect 21795 18005 21805 18045
rect 21845 18005 21855 18045
rect 21895 18005 21905 18045
rect 21945 18005 21955 18045
rect 21995 18005 22005 18045
rect 22045 18005 22055 18045
rect 22095 18005 22105 18045
rect 22145 18005 22155 18045
rect 22195 18005 22205 18045
rect 22245 18005 22255 18045
rect 22295 18005 22305 18045
rect 22345 18005 22355 18045
rect 22395 18005 22405 18045
rect 22445 18005 22455 18045
rect 22495 18005 22505 18045
rect 22545 18005 22555 18045
rect 22595 18005 22605 18045
rect 22645 18005 22655 18045
rect 22695 18005 22705 18045
rect 22745 18005 22755 18045
rect 22795 18005 22805 18045
rect 22845 18005 22855 18045
rect 22895 18005 22905 18045
rect 22945 18005 22955 18045
rect 22995 18005 23005 18045
rect 23045 18005 23055 18045
rect 23095 18005 23105 18045
rect 23145 18005 23155 18045
rect 23195 18005 23205 18045
rect 23245 18005 23255 18045
rect 23295 18005 23305 18045
rect 23345 18005 23355 18045
rect 23395 18005 23405 18045
rect 23445 18005 23455 18045
rect 23495 18005 23505 18045
rect 23545 18005 23555 18045
rect 23595 18005 23605 18045
rect 23645 18005 23655 18045
rect 23695 18005 23705 18045
rect 23745 18005 23755 18045
rect 23795 18005 23805 18045
rect 23845 18005 23855 18045
rect 23895 18005 23905 18045
rect 23945 18005 23955 18045
rect 23995 18005 24005 18045
rect 24045 18005 24055 18045
rect 24095 18005 24105 18045
rect 24145 18005 24155 18045
rect 24195 18005 24205 18045
rect 24245 18005 24255 18045
rect 24295 18005 24305 18045
rect 24345 18005 24355 18045
rect 24395 18005 24405 18045
rect 24445 18005 24455 18045
rect 24495 18005 24505 18045
rect 24545 18005 24555 18045
rect 24595 18005 24605 18045
rect 24645 18005 24655 18045
rect 24695 18005 24705 18045
rect 24745 18005 24755 18045
rect 24795 18005 24805 18045
rect 24845 18005 24855 18045
rect 24895 18005 24905 18045
rect 24945 18005 24955 18045
rect 24995 18005 25005 18045
rect 25045 18005 25055 18045
rect 25095 18005 25105 18045
rect 25145 18005 25155 18045
rect 25195 18005 25205 18045
rect 25245 18005 25255 18045
rect 25295 18005 25305 18045
rect 25345 18005 25355 18045
rect 25395 18005 25405 18045
rect 25445 18005 25455 18045
rect 25495 18005 25505 18045
rect 25545 18005 25555 18045
rect 25595 18005 25605 18045
rect 25645 18005 25655 18045
rect 25695 18005 25705 18045
rect 25745 18005 25755 18045
rect 25795 18005 25805 18045
rect 25845 18005 25855 18045
rect 25895 18005 25905 18045
rect 25945 18005 25955 18045
rect 25995 18005 26005 18045
rect 26045 18005 26055 18045
rect 26095 18005 26105 18045
rect 26145 18005 26155 18045
rect 26195 18005 26205 18045
rect 26245 18005 26255 18045
rect 26295 18005 26305 18045
rect 26345 18005 26355 18045
rect 26395 18005 26405 18045
rect 26445 18005 26455 18045
rect 26495 18005 26505 18045
rect 26545 18005 26555 18045
rect 26595 18005 26605 18045
rect 26645 18005 26655 18045
rect 26695 18005 26705 18045
rect 26745 18005 26755 18045
rect 26795 18005 26805 18045
rect 26845 18005 26855 18045
rect 26895 18005 26905 18045
rect 26945 18005 26955 18045
rect 26995 18005 27005 18045
rect 27045 18005 27055 18045
rect 27095 18005 27105 18045
rect 27145 18005 27155 18045
rect 27195 18005 27205 18045
rect 27245 18005 27255 18045
rect 27295 18005 27305 18045
rect 27345 18005 27355 18045
rect 27395 18005 27405 18045
rect 27445 18005 27455 18045
rect 27495 18005 27505 18045
rect 27545 18005 27555 18045
rect 27595 18005 27605 18045
rect 27645 18005 27655 18045
rect 27695 18005 27705 18045
rect 27745 18005 27755 18045
rect 27795 18005 27805 18045
rect 27845 18005 27855 18045
rect 27895 18005 27905 18045
rect 27945 18005 27955 18045
rect 27995 18005 28005 18045
rect 28045 18005 28055 18045
rect 28095 18005 28105 18045
rect 28145 18005 28155 18045
rect 28195 18005 28205 18045
rect 28245 18005 28255 18045
rect 28295 18005 28305 18045
rect 28345 18005 28355 18045
rect 28395 18005 28405 18045
rect 28445 18005 28455 18045
rect 28495 18005 28505 18045
rect 28545 18005 28555 18045
rect 28595 18005 28605 18045
rect 28645 18005 28655 18045
rect 28695 18005 28705 18045
rect 28745 18005 28755 18045
rect 28795 18005 28805 18045
rect 28845 18005 28855 18045
rect 28895 18005 28905 18045
rect 28945 18005 28955 18045
rect 28995 18005 29005 18045
rect 29045 18005 29055 18045
rect 29095 18005 29105 18045
rect 29145 18005 29155 18045
rect 29195 18005 29205 18045
rect 29245 18005 29255 18045
rect 29295 18005 29305 18045
rect 29345 18005 29355 18045
rect 29395 18005 29405 18045
rect 29445 18005 29455 18045
rect 29495 18005 29505 18045
rect 29545 18005 29555 18045
rect 29595 18005 29605 18045
rect 29645 18005 29655 18045
rect 29695 18005 29705 18045
rect 29745 18005 29755 18045
rect 29795 18005 29805 18045
rect 29845 18005 29855 18045
rect 29895 18005 29905 18045
rect 29945 18005 29955 18045
rect 29995 18005 30005 18045
rect 30045 18005 30055 18045
rect 30095 18005 30105 18045
rect 30145 18005 30155 18045
rect 30195 18005 30205 18045
rect 30245 18005 30255 18045
rect 30295 18005 30305 18045
rect 30345 18005 30355 18045
rect 30395 18005 30405 18045
rect 30445 18005 30455 18045
rect 30495 18005 30505 18045
rect 30545 18005 30555 18045
rect 30595 18005 30605 18045
rect 30645 18005 30655 18045
rect 30695 18005 30705 18045
rect 30745 18005 30755 18045
rect 30795 18005 30805 18045
rect 30845 18005 30855 18045
rect 30895 18005 30905 18045
rect 30945 18005 30955 18045
rect 30995 18005 31005 18045
rect 31045 18005 31055 18045
rect 31095 18005 31105 18045
rect 31145 18005 31155 18045
rect 31195 18005 31205 18045
rect 31245 18005 31255 18045
rect 31295 18005 31305 18045
rect 31345 18005 31355 18045
rect 31395 18005 31405 18045
rect 31445 18005 31455 18045
rect 31495 18005 31505 18045
rect 31545 18005 31555 18045
rect 31595 18005 31605 18045
rect 31645 18005 31655 18045
rect 31695 18005 31705 18045
rect 31745 18005 31755 18045
rect 31795 18005 31805 18045
rect 31845 18005 31855 18045
rect 31895 18005 31905 18045
rect 31945 18005 31955 18045
rect 31995 18005 32005 18045
rect 32045 18005 32055 18045
rect 32095 18005 32105 18045
rect 32145 18005 32155 18045
rect 32195 18005 32205 18045
rect 32245 18005 32255 18045
rect 32295 18005 32305 18045
rect 32345 18005 32355 18045
rect 32395 18005 32405 18045
rect 32445 18005 32455 18045
rect 32495 18005 32505 18045
rect 32545 18005 32555 18045
rect 32595 18005 32605 18045
rect 32645 18005 32655 18045
rect 32695 18005 32705 18045
rect 32745 18005 32755 18045
rect 32795 18005 32805 18045
rect 32845 18005 32855 18045
rect 32895 18005 32905 18045
rect 32945 18005 32955 18045
rect 32995 18005 33005 18045
rect 33045 18005 33055 18045
rect 33095 18005 33105 18045
rect 33145 18005 33155 18045
rect 33195 18005 33205 18045
rect 33245 18005 33255 18045
rect 33295 18005 33305 18045
rect 33345 18005 33355 18045
rect 33395 18005 33405 18045
rect 33445 18005 33455 18045
rect 33495 18005 33505 18045
rect 33545 18005 33555 18045
rect 33595 18005 33605 18045
rect 33645 18005 33655 18045
rect 33695 18005 33705 18045
rect 33745 18005 33755 18045
rect 33795 18005 33805 18045
rect 33845 18005 33855 18045
rect 33895 18005 33905 18045
rect 33945 18005 33955 18045
rect 33995 18005 34005 18045
rect 34045 18005 34055 18045
rect 34095 18005 34105 18045
rect 34145 18005 34155 18045
rect 34195 18005 34205 18045
rect 34245 18005 34255 18045
rect 34295 18005 34305 18045
rect 34345 18005 34355 18045
rect 34395 18005 34405 18045
rect 34445 18005 34455 18045
rect 34495 18005 34505 18045
rect 34545 18005 34555 18045
rect 34595 18005 34605 18045
rect 34645 18005 34655 18045
rect 34695 18005 34705 18045
rect 34745 18005 34755 18045
rect 34795 18005 34805 18045
rect 34845 18005 34855 18045
rect 34895 18005 34905 18045
rect 34945 18005 34955 18045
rect 34995 18005 35005 18045
rect 35045 18005 35055 18045
rect 35095 18005 35105 18045
rect 35145 18005 35155 18045
rect 35195 18005 35205 18045
rect 35245 18005 35255 18045
rect 35295 18005 35305 18045
rect 35345 18005 35355 18045
rect 35395 18005 35405 18045
rect 35445 18005 35455 18045
rect 35495 18005 35505 18045
rect 35545 18005 35555 18045
rect 35595 18005 35605 18045
rect 35645 18005 35655 18045
rect 35695 18005 35705 18045
rect 35745 18005 35755 18045
rect 35795 18005 35805 18045
rect 35845 18005 35855 18045
rect 35895 18005 35905 18045
rect 35945 18005 35955 18045
rect 35995 18005 36005 18045
rect 36045 18005 36055 18045
rect 36095 18005 36105 18045
rect 36145 18005 36155 18045
rect 36195 18005 36205 18045
rect 36245 18005 36255 18045
rect 36295 18005 36305 18045
rect 36345 18005 36355 18045
rect 36395 18005 36405 18045
rect 36445 18005 36455 18045
rect 36495 18005 36505 18045
rect 36545 18005 36555 18045
rect 36595 18005 36605 18045
rect 36645 18005 36655 18045
rect 36695 18005 36705 18045
rect 36745 18005 36755 18045
rect 36795 18005 36805 18045
rect 36845 18005 36855 18045
rect 36895 18005 36905 18045
rect 36945 18005 36955 18045
rect 36995 18005 37005 18045
rect 37045 18005 37055 18045
rect 37095 18005 37105 18045
rect 37145 18005 37155 18045
rect 37195 18005 37205 18045
rect 37245 18005 37255 18045
rect 37295 18005 37305 18045
rect 37345 18005 37355 18045
rect 37395 18005 37405 18045
rect 37445 18005 37455 18045
rect 37495 18005 37505 18045
rect 37545 18005 37555 18045
rect 37595 18005 37605 18045
rect 37645 18005 37655 18045
rect 37695 18005 37705 18045
rect 37745 18005 37755 18045
rect 37795 18005 37805 18045
rect 37845 18005 37855 18045
rect 37895 18005 37905 18045
rect 37945 18005 37955 18045
rect 37995 18005 38005 18045
rect 38045 18005 38055 18045
rect 38095 18005 38105 18045
rect 38145 18005 38155 18045
rect 38195 18005 38205 18045
rect 38245 18005 38255 18045
rect 38295 18005 38305 18045
rect 38345 18005 38355 18045
rect 38395 18005 38405 18045
rect 38445 18005 38455 18045
rect 38495 18005 38505 18045
rect 38545 18005 38555 18045
rect 38595 18005 38605 18045
rect 38645 18005 38655 18045
rect 38695 18005 38705 18045
rect 38745 18005 38755 18045
rect 38795 18005 38805 18045
rect 38845 18005 38855 18045
rect 38895 18005 38905 18045
rect 38945 18005 38955 18045
rect 38995 18005 39005 18045
rect 39045 18005 39055 18045
rect 39095 18005 39105 18045
rect 39145 18005 39155 18045
rect 39195 18005 39205 18045
rect 39245 18005 39255 18045
rect 39295 18005 39305 18045
rect 39345 18005 39355 18045
rect 39395 18005 39405 18045
rect 39445 18005 39455 18045
rect 39495 18005 39505 18045
rect 39545 18005 39555 18045
rect 39595 18005 39605 18045
rect 39645 18005 39655 18045
rect 39695 18005 39705 18045
rect 39745 18005 39750 18045
rect 0 18000 39750 18005
rect 0 16950 50 18000
rect 100 17850 3200 17950
rect 100 17200 200 17850
rect 3100 17200 3200 17850
rect 100 17050 3200 17200
rect 3350 17850 6450 17950
rect 3350 17200 3450 17850
rect 6350 17200 6450 17850
rect 3350 17050 6450 17200
rect 6600 17850 9700 17950
rect 6600 17200 6700 17850
rect 9600 17200 9700 17850
rect 6600 17050 9700 17200
rect 9850 17850 12950 17950
rect 9850 17200 9950 17850
rect 12850 17200 12950 17850
rect 9850 17050 12950 17200
rect 13100 17850 16200 17950
rect 13100 17200 13200 17850
rect 16100 17200 16200 17850
rect 13100 17050 16200 17200
rect 16350 17850 19450 17950
rect 16350 17200 16450 17850
rect 19350 17200 19450 17850
rect 16350 17050 19450 17200
rect 19600 17850 22700 17950
rect 19600 17200 19700 17850
rect 22600 17200 22700 17850
rect 19600 17050 22700 17200
rect 22850 17850 25950 17950
rect 22850 17200 22950 17850
rect 25850 17200 25950 17850
rect 22850 17050 25950 17200
rect 26100 17850 29200 17950
rect 26100 17200 26200 17850
rect 29100 17200 29200 17850
rect 26100 17050 29200 17200
rect 29350 17850 32450 17950
rect 29350 17200 29450 17850
rect 32350 17200 32450 17850
rect 29350 17050 32450 17200
rect 32600 17850 35700 17950
rect 32600 17200 32700 17850
rect 35600 17200 35700 17850
rect 32600 17050 35700 17200
rect 35850 17850 38950 17950
rect 35850 17200 35950 17850
rect 38850 17200 38950 17850
rect 35850 17050 38950 17200
rect 39100 17850 39750 17950
rect 39100 17200 39200 17850
rect 39650 17200 39750 17850
rect 39100 17050 39750 17200
rect 100 17045 39750 17050
rect 100 17005 105 17045
rect 145 17005 155 17045
rect 195 17005 205 17045
rect 245 17005 255 17045
rect 295 17005 305 17045
rect 345 17005 355 17045
rect 395 17005 405 17045
rect 445 17005 455 17045
rect 495 17005 505 17045
rect 545 17005 555 17045
rect 595 17005 605 17045
rect 645 17005 655 17045
rect 695 17005 705 17045
rect 745 17005 755 17045
rect 795 17005 805 17045
rect 845 17005 855 17045
rect 895 17005 905 17045
rect 945 17005 955 17045
rect 995 17005 1005 17045
rect 1045 17005 1055 17045
rect 1095 17005 1105 17045
rect 1145 17005 1155 17045
rect 1195 17005 1205 17045
rect 1245 17005 1255 17045
rect 1295 17005 1305 17045
rect 1345 17005 1355 17045
rect 1395 17005 1405 17045
rect 1445 17005 1455 17045
rect 1495 17005 1505 17045
rect 1545 17005 1555 17045
rect 1595 17005 1605 17045
rect 1645 17005 1655 17045
rect 1695 17005 1705 17045
rect 1745 17005 1755 17045
rect 1795 17005 1805 17045
rect 1845 17005 1855 17045
rect 1895 17005 1905 17045
rect 1945 17005 1955 17045
rect 1995 17005 2005 17045
rect 2045 17005 2055 17045
rect 2095 17005 2105 17045
rect 2145 17005 2155 17045
rect 2195 17005 2205 17045
rect 2245 17005 2255 17045
rect 2295 17005 2305 17045
rect 2345 17005 2355 17045
rect 2395 17005 2405 17045
rect 2445 17005 2455 17045
rect 2495 17005 2505 17045
rect 2545 17005 2555 17045
rect 2595 17005 2605 17045
rect 2645 17005 2655 17045
rect 2695 17005 2705 17045
rect 2745 17005 2755 17045
rect 2795 17005 2805 17045
rect 2845 17005 2855 17045
rect 2895 17005 2905 17045
rect 2945 17005 2955 17045
rect 2995 17005 3005 17045
rect 3045 17005 3055 17045
rect 3095 17005 3105 17045
rect 3145 17005 3155 17045
rect 3195 17005 3205 17045
rect 3245 17005 3255 17045
rect 3295 17005 3305 17045
rect 3345 17005 3355 17045
rect 3395 17005 3405 17045
rect 3445 17005 3455 17045
rect 3495 17005 3505 17045
rect 3545 17005 3555 17045
rect 3595 17005 3605 17045
rect 3645 17005 3655 17045
rect 3695 17005 3705 17045
rect 3745 17005 3755 17045
rect 3795 17005 3805 17045
rect 3845 17005 3855 17045
rect 3895 17005 3905 17045
rect 3945 17005 3955 17045
rect 3995 17005 4005 17045
rect 4045 17005 4055 17045
rect 4095 17005 4105 17045
rect 4145 17005 4155 17045
rect 4195 17005 4205 17045
rect 4245 17005 4255 17045
rect 4295 17005 4305 17045
rect 4345 17005 4355 17045
rect 4395 17005 4405 17045
rect 4445 17005 4455 17045
rect 4495 17005 4505 17045
rect 4545 17005 4555 17045
rect 4595 17005 4605 17045
rect 4645 17005 4655 17045
rect 4695 17005 4705 17045
rect 4745 17005 4755 17045
rect 4795 17005 4805 17045
rect 4845 17005 4855 17045
rect 4895 17005 4905 17045
rect 4945 17005 4955 17045
rect 4995 17005 5005 17045
rect 5045 17005 5055 17045
rect 5095 17005 5105 17045
rect 5145 17005 5155 17045
rect 5195 17005 5205 17045
rect 5245 17005 5255 17045
rect 5295 17005 5305 17045
rect 5345 17005 5355 17045
rect 5395 17005 5405 17045
rect 5445 17005 5455 17045
rect 5495 17005 5505 17045
rect 5545 17005 5555 17045
rect 5595 17005 5605 17045
rect 5645 17005 5655 17045
rect 5695 17005 5705 17045
rect 5745 17005 5755 17045
rect 5795 17005 5805 17045
rect 5845 17005 5855 17045
rect 5895 17005 5905 17045
rect 5945 17005 5955 17045
rect 5995 17005 6005 17045
rect 6045 17005 6055 17045
rect 6095 17005 6105 17045
rect 6145 17005 6155 17045
rect 6195 17005 6205 17045
rect 6245 17005 6255 17045
rect 6295 17005 6305 17045
rect 6345 17005 6355 17045
rect 6395 17005 6405 17045
rect 6445 17005 6455 17045
rect 6495 17005 6505 17045
rect 6545 17005 6555 17045
rect 6595 17005 6605 17045
rect 6645 17005 6655 17045
rect 6695 17005 6705 17045
rect 6745 17005 6755 17045
rect 6795 17005 6805 17045
rect 6845 17005 6855 17045
rect 6895 17005 6905 17045
rect 6945 17005 6955 17045
rect 6995 17005 7005 17045
rect 7045 17005 7055 17045
rect 7095 17005 7105 17045
rect 7145 17005 7155 17045
rect 7195 17005 7205 17045
rect 7245 17005 7255 17045
rect 7295 17005 7305 17045
rect 7345 17005 7355 17045
rect 7395 17005 7405 17045
rect 7445 17005 7455 17045
rect 7495 17005 7505 17045
rect 7545 17005 7555 17045
rect 7595 17005 7605 17045
rect 7645 17005 7655 17045
rect 7695 17005 7705 17045
rect 7745 17005 7755 17045
rect 7795 17005 7805 17045
rect 7845 17005 7855 17045
rect 7895 17005 7905 17045
rect 7945 17005 7955 17045
rect 7995 17005 8005 17045
rect 8045 17005 8055 17045
rect 8095 17005 8105 17045
rect 8145 17005 8155 17045
rect 8195 17005 8205 17045
rect 8245 17005 8255 17045
rect 8295 17005 8305 17045
rect 8345 17005 8355 17045
rect 8395 17005 8405 17045
rect 8445 17005 8455 17045
rect 8495 17005 8505 17045
rect 8545 17005 8555 17045
rect 8595 17005 8605 17045
rect 8645 17005 8655 17045
rect 8695 17005 8705 17045
rect 8745 17005 8755 17045
rect 8795 17005 8805 17045
rect 8845 17005 8855 17045
rect 8895 17005 8905 17045
rect 8945 17005 8955 17045
rect 8995 17005 9005 17045
rect 9045 17005 9055 17045
rect 9095 17005 9105 17045
rect 9145 17005 9155 17045
rect 9195 17005 9205 17045
rect 9245 17005 9255 17045
rect 9295 17005 9305 17045
rect 9345 17005 9355 17045
rect 9395 17005 9405 17045
rect 9445 17005 9455 17045
rect 9495 17005 9505 17045
rect 9545 17005 9555 17045
rect 9595 17005 9605 17045
rect 9645 17005 9655 17045
rect 9695 17005 9705 17045
rect 9745 17005 9755 17045
rect 9795 17005 9805 17045
rect 9845 17005 9855 17045
rect 9895 17005 9905 17045
rect 9945 17005 9955 17045
rect 9995 17005 10005 17045
rect 10045 17005 10055 17045
rect 10095 17005 10105 17045
rect 10145 17005 10155 17045
rect 10195 17005 10205 17045
rect 10245 17005 10255 17045
rect 10295 17005 10305 17045
rect 10345 17005 10355 17045
rect 10395 17005 10405 17045
rect 10445 17005 10455 17045
rect 10495 17005 10505 17045
rect 10545 17005 10555 17045
rect 10595 17005 10605 17045
rect 10645 17005 10655 17045
rect 10695 17005 10705 17045
rect 10745 17005 10755 17045
rect 10795 17005 10805 17045
rect 10845 17005 10855 17045
rect 10895 17005 10905 17045
rect 10945 17005 10955 17045
rect 10995 17005 11005 17045
rect 11045 17005 11055 17045
rect 11095 17005 11105 17045
rect 11145 17005 11155 17045
rect 11195 17005 11205 17045
rect 11245 17005 11255 17045
rect 11295 17005 11305 17045
rect 11345 17005 11355 17045
rect 11395 17005 11405 17045
rect 11445 17005 11455 17045
rect 11495 17005 11505 17045
rect 11545 17005 11555 17045
rect 11595 17005 11605 17045
rect 11645 17005 11655 17045
rect 11695 17005 11705 17045
rect 11745 17005 11755 17045
rect 11795 17005 11805 17045
rect 11845 17005 11855 17045
rect 11895 17005 11905 17045
rect 11945 17005 11955 17045
rect 11995 17005 12005 17045
rect 12045 17005 12055 17045
rect 12095 17005 12105 17045
rect 12145 17005 12155 17045
rect 12195 17005 12205 17045
rect 12245 17005 12255 17045
rect 12295 17005 12305 17045
rect 12345 17005 12355 17045
rect 12395 17005 12405 17045
rect 12445 17005 12455 17045
rect 12495 17005 12505 17045
rect 12545 17005 12555 17045
rect 12595 17005 12605 17045
rect 12645 17005 12655 17045
rect 12695 17005 12705 17045
rect 12745 17005 12755 17045
rect 12795 17005 12805 17045
rect 12845 17005 12855 17045
rect 12895 17005 12905 17045
rect 12945 17005 12955 17045
rect 12995 17005 13005 17045
rect 13045 17005 13055 17045
rect 13095 17005 13105 17045
rect 13145 17005 13155 17045
rect 13195 17005 13205 17045
rect 13245 17005 13255 17045
rect 13295 17005 13305 17045
rect 13345 17005 13355 17045
rect 13395 17005 13405 17045
rect 13445 17005 13455 17045
rect 13495 17005 13505 17045
rect 13545 17005 13555 17045
rect 13595 17005 13605 17045
rect 13645 17005 13655 17045
rect 13695 17005 13705 17045
rect 13745 17005 13755 17045
rect 13795 17005 13805 17045
rect 13845 17005 13855 17045
rect 13895 17005 13905 17045
rect 13945 17005 13955 17045
rect 13995 17005 14005 17045
rect 14045 17005 14055 17045
rect 14095 17005 14105 17045
rect 14145 17005 14155 17045
rect 14195 17005 14205 17045
rect 14245 17005 14255 17045
rect 14295 17005 14305 17045
rect 14345 17005 14355 17045
rect 14395 17005 14405 17045
rect 14445 17005 14455 17045
rect 14495 17005 14505 17045
rect 14545 17005 14555 17045
rect 14595 17005 14605 17045
rect 14645 17005 14655 17045
rect 14695 17005 14705 17045
rect 14745 17005 14755 17045
rect 14795 17005 14805 17045
rect 14845 17005 14855 17045
rect 14895 17005 14905 17045
rect 14945 17005 14955 17045
rect 14995 17005 15005 17045
rect 15045 17005 15055 17045
rect 15095 17005 15105 17045
rect 15145 17005 15155 17045
rect 15195 17005 15205 17045
rect 15245 17005 15255 17045
rect 15295 17005 15305 17045
rect 15345 17005 15355 17045
rect 15395 17005 15405 17045
rect 15445 17005 15455 17045
rect 15495 17005 15505 17045
rect 15545 17005 15555 17045
rect 15595 17005 15605 17045
rect 15645 17005 15655 17045
rect 15695 17005 15705 17045
rect 15745 17005 15755 17045
rect 15795 17005 15805 17045
rect 15845 17005 15855 17045
rect 15895 17005 15905 17045
rect 15945 17005 15955 17045
rect 15995 17005 16005 17045
rect 16045 17005 16055 17045
rect 16095 17005 16105 17045
rect 16145 17005 16155 17045
rect 16195 17005 16205 17045
rect 16245 17005 16255 17045
rect 16295 17005 16305 17045
rect 16345 17005 16355 17045
rect 16395 17005 16405 17045
rect 16445 17005 16455 17045
rect 16495 17005 16505 17045
rect 16545 17005 16555 17045
rect 16595 17005 16605 17045
rect 16645 17005 16655 17045
rect 16695 17005 16705 17045
rect 16745 17005 16755 17045
rect 16795 17005 16805 17045
rect 16845 17005 16855 17045
rect 16895 17005 16905 17045
rect 16945 17005 16955 17045
rect 16995 17005 17005 17045
rect 17045 17005 17055 17045
rect 17095 17005 17105 17045
rect 17145 17005 17155 17045
rect 17195 17005 17205 17045
rect 17245 17005 17255 17045
rect 17295 17005 17305 17045
rect 17345 17005 17355 17045
rect 17395 17005 17405 17045
rect 17445 17005 17455 17045
rect 17495 17005 17505 17045
rect 17545 17005 17555 17045
rect 17595 17005 17605 17045
rect 17645 17005 17655 17045
rect 17695 17005 17705 17045
rect 17745 17005 17755 17045
rect 17795 17005 17805 17045
rect 17845 17005 17855 17045
rect 17895 17005 17905 17045
rect 17945 17005 17955 17045
rect 17995 17005 18005 17045
rect 18045 17005 18055 17045
rect 18095 17005 18105 17045
rect 18145 17005 18155 17045
rect 18195 17005 18205 17045
rect 18245 17005 18255 17045
rect 18295 17005 18305 17045
rect 18345 17005 18355 17045
rect 18395 17005 18405 17045
rect 18445 17005 18455 17045
rect 18495 17005 18505 17045
rect 18545 17005 18555 17045
rect 18595 17005 18605 17045
rect 18645 17005 18655 17045
rect 18695 17005 18705 17045
rect 18745 17005 18755 17045
rect 18795 17005 18805 17045
rect 18845 17005 18855 17045
rect 18895 17005 18905 17045
rect 18945 17005 18955 17045
rect 18995 17005 19005 17045
rect 19045 17005 19055 17045
rect 19095 17005 19105 17045
rect 19145 17005 19155 17045
rect 19195 17005 19205 17045
rect 19245 17005 19255 17045
rect 19295 17005 19305 17045
rect 19345 17005 19355 17045
rect 19395 17005 19405 17045
rect 19445 17005 19455 17045
rect 19495 17005 19505 17045
rect 19545 17005 19555 17045
rect 19595 17005 19605 17045
rect 19645 17005 19655 17045
rect 19695 17005 19705 17045
rect 19745 17005 19755 17045
rect 19795 17005 19805 17045
rect 19845 17005 19855 17045
rect 19895 17005 19905 17045
rect 19945 17005 19955 17045
rect 19995 17005 20005 17045
rect 20045 17005 20055 17045
rect 20095 17005 20105 17045
rect 20145 17005 20155 17045
rect 20195 17005 20205 17045
rect 20245 17005 20255 17045
rect 20295 17005 20305 17045
rect 20345 17005 20355 17045
rect 20395 17005 20405 17045
rect 20445 17005 20455 17045
rect 20495 17005 20505 17045
rect 20545 17005 20555 17045
rect 20595 17005 20605 17045
rect 20645 17005 20655 17045
rect 20695 17005 20705 17045
rect 20745 17005 20755 17045
rect 20795 17005 20805 17045
rect 20845 17005 20855 17045
rect 20895 17005 20905 17045
rect 20945 17005 20955 17045
rect 20995 17005 21005 17045
rect 21045 17005 21055 17045
rect 21095 17005 21105 17045
rect 21145 17005 21155 17045
rect 21195 17005 21205 17045
rect 21245 17005 21255 17045
rect 21295 17005 21305 17045
rect 21345 17005 21355 17045
rect 21395 17005 21405 17045
rect 21445 17005 21455 17045
rect 21495 17005 21505 17045
rect 21545 17005 21555 17045
rect 21595 17005 21605 17045
rect 21645 17005 21655 17045
rect 21695 17005 21705 17045
rect 21745 17005 21755 17045
rect 21795 17005 21805 17045
rect 21845 17005 21855 17045
rect 21895 17005 21905 17045
rect 21945 17005 21955 17045
rect 21995 17005 22005 17045
rect 22045 17005 22055 17045
rect 22095 17005 22105 17045
rect 22145 17005 22155 17045
rect 22195 17005 22205 17045
rect 22245 17005 22255 17045
rect 22295 17005 22305 17045
rect 22345 17005 22355 17045
rect 22395 17005 22405 17045
rect 22445 17005 22455 17045
rect 22495 17005 22505 17045
rect 22545 17005 22555 17045
rect 22595 17005 22605 17045
rect 22645 17005 22655 17045
rect 22695 17005 22705 17045
rect 22745 17005 22755 17045
rect 22795 17005 22805 17045
rect 22845 17005 22855 17045
rect 22895 17005 22905 17045
rect 22945 17005 22955 17045
rect 22995 17005 23005 17045
rect 23045 17005 23055 17045
rect 23095 17005 23105 17045
rect 23145 17005 23155 17045
rect 23195 17005 23205 17045
rect 23245 17005 23255 17045
rect 23295 17005 23305 17045
rect 23345 17005 23355 17045
rect 23395 17005 23405 17045
rect 23445 17005 23455 17045
rect 23495 17005 23505 17045
rect 23545 17005 23555 17045
rect 23595 17005 23605 17045
rect 23645 17005 23655 17045
rect 23695 17005 23705 17045
rect 23745 17005 23755 17045
rect 23795 17005 23805 17045
rect 23845 17005 23855 17045
rect 23895 17005 23905 17045
rect 23945 17005 23955 17045
rect 23995 17005 24005 17045
rect 24045 17005 24055 17045
rect 24095 17005 24105 17045
rect 24145 17005 24155 17045
rect 24195 17005 24205 17045
rect 24245 17005 24255 17045
rect 24295 17005 24305 17045
rect 24345 17005 24355 17045
rect 24395 17005 24405 17045
rect 24445 17005 24455 17045
rect 24495 17005 24505 17045
rect 24545 17005 24555 17045
rect 24595 17005 24605 17045
rect 24645 17005 24655 17045
rect 24695 17005 24705 17045
rect 24745 17005 24755 17045
rect 24795 17005 24805 17045
rect 24845 17005 24855 17045
rect 24895 17005 24905 17045
rect 24945 17005 24955 17045
rect 24995 17005 25005 17045
rect 25045 17005 25055 17045
rect 25095 17005 25105 17045
rect 25145 17005 25155 17045
rect 25195 17005 25205 17045
rect 25245 17005 25255 17045
rect 25295 17005 25305 17045
rect 25345 17005 25355 17045
rect 25395 17005 25405 17045
rect 25445 17005 25455 17045
rect 25495 17005 25505 17045
rect 25545 17005 25555 17045
rect 25595 17005 25605 17045
rect 25645 17005 25655 17045
rect 25695 17005 25705 17045
rect 25745 17005 25755 17045
rect 25795 17005 25805 17045
rect 25845 17005 25855 17045
rect 25895 17005 25905 17045
rect 25945 17005 25955 17045
rect 25995 17005 26005 17045
rect 26045 17005 26055 17045
rect 26095 17005 26105 17045
rect 26145 17005 26155 17045
rect 26195 17005 26205 17045
rect 26245 17005 26255 17045
rect 26295 17005 26305 17045
rect 26345 17005 26355 17045
rect 26395 17005 26405 17045
rect 26445 17005 26455 17045
rect 26495 17005 26505 17045
rect 26545 17005 26555 17045
rect 26595 17005 26605 17045
rect 26645 17005 26655 17045
rect 26695 17005 26705 17045
rect 26745 17005 26755 17045
rect 26795 17005 26805 17045
rect 26845 17005 26855 17045
rect 26895 17005 26905 17045
rect 26945 17005 26955 17045
rect 26995 17005 27005 17045
rect 27045 17005 27055 17045
rect 27095 17005 27105 17045
rect 27145 17005 27155 17045
rect 27195 17005 27205 17045
rect 27245 17005 27255 17045
rect 27295 17005 27305 17045
rect 27345 17005 27355 17045
rect 27395 17005 27405 17045
rect 27445 17005 27455 17045
rect 27495 17005 27505 17045
rect 27545 17005 27555 17045
rect 27595 17005 27605 17045
rect 27645 17005 27655 17045
rect 27695 17005 27705 17045
rect 27745 17005 27755 17045
rect 27795 17005 27805 17045
rect 27845 17005 27855 17045
rect 27895 17005 27905 17045
rect 27945 17005 27955 17045
rect 27995 17005 28005 17045
rect 28045 17005 28055 17045
rect 28095 17005 28105 17045
rect 28145 17005 28155 17045
rect 28195 17005 28205 17045
rect 28245 17005 28255 17045
rect 28295 17005 28305 17045
rect 28345 17005 28355 17045
rect 28395 17005 28405 17045
rect 28445 17005 28455 17045
rect 28495 17005 28505 17045
rect 28545 17005 28555 17045
rect 28595 17005 28605 17045
rect 28645 17005 28655 17045
rect 28695 17005 28705 17045
rect 28745 17005 28755 17045
rect 28795 17005 28805 17045
rect 28845 17005 28855 17045
rect 28895 17005 28905 17045
rect 28945 17005 28955 17045
rect 28995 17005 29005 17045
rect 29045 17005 29055 17045
rect 29095 17005 29105 17045
rect 29145 17005 29155 17045
rect 29195 17005 29205 17045
rect 29245 17005 29255 17045
rect 29295 17005 29305 17045
rect 29345 17005 29355 17045
rect 29395 17005 29405 17045
rect 29445 17005 29455 17045
rect 29495 17005 29505 17045
rect 29545 17005 29555 17045
rect 29595 17005 29605 17045
rect 29645 17005 29655 17045
rect 29695 17005 29705 17045
rect 29745 17005 29755 17045
rect 29795 17005 29805 17045
rect 29845 17005 29855 17045
rect 29895 17005 29905 17045
rect 29945 17005 29955 17045
rect 29995 17005 30005 17045
rect 30045 17005 30055 17045
rect 30095 17005 30105 17045
rect 30145 17005 30155 17045
rect 30195 17005 30205 17045
rect 30245 17005 30255 17045
rect 30295 17005 30305 17045
rect 30345 17005 30355 17045
rect 30395 17005 30405 17045
rect 30445 17005 30455 17045
rect 30495 17005 30505 17045
rect 30545 17005 30555 17045
rect 30595 17005 30605 17045
rect 30645 17005 30655 17045
rect 30695 17005 30705 17045
rect 30745 17005 30755 17045
rect 30795 17005 30805 17045
rect 30845 17005 30855 17045
rect 30895 17005 30905 17045
rect 30945 17005 30955 17045
rect 30995 17005 31005 17045
rect 31045 17005 31055 17045
rect 31095 17005 31105 17045
rect 31145 17005 31155 17045
rect 31195 17005 31205 17045
rect 31245 17005 31255 17045
rect 31295 17005 31305 17045
rect 31345 17005 31355 17045
rect 31395 17005 31405 17045
rect 31445 17005 31455 17045
rect 31495 17005 31505 17045
rect 31545 17005 31555 17045
rect 31595 17005 31605 17045
rect 31645 17005 31655 17045
rect 31695 17005 31705 17045
rect 31745 17005 31755 17045
rect 31795 17005 31805 17045
rect 31845 17005 31855 17045
rect 31895 17005 31905 17045
rect 31945 17005 31955 17045
rect 31995 17005 32005 17045
rect 32045 17005 32055 17045
rect 32095 17005 32105 17045
rect 32145 17005 32155 17045
rect 32195 17005 32205 17045
rect 32245 17005 32255 17045
rect 32295 17005 32305 17045
rect 32345 17005 32355 17045
rect 32395 17005 32405 17045
rect 32445 17005 32455 17045
rect 32495 17005 32505 17045
rect 32545 17005 32555 17045
rect 32595 17005 32605 17045
rect 32645 17005 32655 17045
rect 32695 17005 32705 17045
rect 32745 17005 32755 17045
rect 32795 17005 32805 17045
rect 32845 17005 32855 17045
rect 32895 17005 32905 17045
rect 32945 17005 32955 17045
rect 32995 17005 33005 17045
rect 33045 17005 33055 17045
rect 33095 17005 33105 17045
rect 33145 17005 33155 17045
rect 33195 17005 33205 17045
rect 33245 17005 33255 17045
rect 33295 17005 33305 17045
rect 33345 17005 33355 17045
rect 33395 17005 33405 17045
rect 33445 17005 33455 17045
rect 33495 17005 33505 17045
rect 33545 17005 33555 17045
rect 33595 17005 33605 17045
rect 33645 17005 33655 17045
rect 33695 17005 33705 17045
rect 33745 17005 33755 17045
rect 33795 17005 33805 17045
rect 33845 17005 33855 17045
rect 33895 17005 33905 17045
rect 33945 17005 33955 17045
rect 33995 17005 34005 17045
rect 34045 17005 34055 17045
rect 34095 17005 34105 17045
rect 34145 17005 34155 17045
rect 34195 17005 34205 17045
rect 34245 17005 34255 17045
rect 34295 17005 34305 17045
rect 34345 17005 34355 17045
rect 34395 17005 34405 17045
rect 34445 17005 34455 17045
rect 34495 17005 34505 17045
rect 34545 17005 34555 17045
rect 34595 17005 34605 17045
rect 34645 17005 34655 17045
rect 34695 17005 34705 17045
rect 34745 17005 34755 17045
rect 34795 17005 34805 17045
rect 34845 17005 34855 17045
rect 34895 17005 34905 17045
rect 34945 17005 34955 17045
rect 34995 17005 35005 17045
rect 35045 17005 35055 17045
rect 35095 17005 35105 17045
rect 35145 17005 35155 17045
rect 35195 17005 35205 17045
rect 35245 17005 35255 17045
rect 35295 17005 35305 17045
rect 35345 17005 35355 17045
rect 35395 17005 35405 17045
rect 35445 17005 35455 17045
rect 35495 17005 35505 17045
rect 35545 17005 35555 17045
rect 35595 17005 35605 17045
rect 35645 17005 35655 17045
rect 35695 17005 35705 17045
rect 35745 17005 35755 17045
rect 35795 17005 35805 17045
rect 35845 17005 35855 17045
rect 35895 17005 35905 17045
rect 35945 17005 35955 17045
rect 35995 17005 36005 17045
rect 36045 17005 36055 17045
rect 36095 17005 36105 17045
rect 36145 17005 36155 17045
rect 36195 17005 36205 17045
rect 36245 17005 36255 17045
rect 36295 17005 36305 17045
rect 36345 17005 36355 17045
rect 36395 17005 36405 17045
rect 36445 17005 36455 17045
rect 36495 17005 36505 17045
rect 36545 17005 36555 17045
rect 36595 17005 36605 17045
rect 36645 17005 36655 17045
rect 36695 17005 36705 17045
rect 36745 17005 36755 17045
rect 36795 17005 36805 17045
rect 36845 17005 36855 17045
rect 36895 17005 36905 17045
rect 36945 17005 36955 17045
rect 36995 17005 37005 17045
rect 37045 17005 37055 17045
rect 37095 17005 37105 17045
rect 37145 17005 37155 17045
rect 37195 17005 37205 17045
rect 37245 17005 37255 17045
rect 37295 17005 37305 17045
rect 37345 17005 37355 17045
rect 37395 17005 37405 17045
rect 37445 17005 37455 17045
rect 37495 17005 37505 17045
rect 37545 17005 37555 17045
rect 37595 17005 37605 17045
rect 37645 17005 37655 17045
rect 37695 17005 37705 17045
rect 37745 17005 37755 17045
rect 37795 17005 37805 17045
rect 37845 17005 37855 17045
rect 37895 17005 37905 17045
rect 37945 17005 37955 17045
rect 37995 17005 38005 17045
rect 38045 17005 38055 17045
rect 38095 17005 38105 17045
rect 38145 17005 38155 17045
rect 38195 17005 38205 17045
rect 38245 17005 38255 17045
rect 38295 17005 38305 17045
rect 38345 17005 38355 17045
rect 38395 17005 38405 17045
rect 38445 17005 38455 17045
rect 38495 17005 38505 17045
rect 38545 17005 38555 17045
rect 38595 17005 38605 17045
rect 38645 17005 38655 17045
rect 38695 17005 38705 17045
rect 38745 17005 38755 17045
rect 38795 17005 38805 17045
rect 38845 17005 38855 17045
rect 38895 17005 38905 17045
rect 38945 17005 38955 17045
rect 38995 17005 39005 17045
rect 39045 17005 39055 17045
rect 39095 17005 39105 17045
rect 39145 17005 39155 17045
rect 39195 17005 39205 17045
rect 39245 17005 39255 17045
rect 39295 17005 39305 17045
rect 39345 17005 39355 17045
rect 39395 17005 39405 17045
rect 39445 17005 39455 17045
rect 39495 17005 39505 17045
rect 39545 17005 39555 17045
rect 39595 17005 39605 17045
rect 39645 17005 39655 17045
rect 39695 17005 39705 17045
rect 39745 17005 39750 17045
rect 100 17000 39750 17005
rect 0 16945 39750 16950
rect 0 16905 5 16945
rect 45 16905 55 16945
rect 95 16905 105 16945
rect 145 16905 155 16945
rect 195 16905 205 16945
rect 245 16905 255 16945
rect 295 16905 305 16945
rect 345 16905 355 16945
rect 395 16905 405 16945
rect 445 16905 455 16945
rect 495 16905 505 16945
rect 545 16905 555 16945
rect 595 16905 605 16945
rect 645 16905 655 16945
rect 695 16905 705 16945
rect 745 16905 755 16945
rect 795 16905 805 16945
rect 845 16905 855 16945
rect 895 16905 905 16945
rect 945 16905 955 16945
rect 995 16905 1005 16945
rect 1045 16905 1055 16945
rect 1095 16905 1105 16945
rect 1145 16905 1155 16945
rect 1195 16905 1205 16945
rect 1245 16905 1255 16945
rect 1295 16905 1305 16945
rect 1345 16905 1355 16945
rect 1395 16905 1405 16945
rect 1445 16905 1455 16945
rect 1495 16905 1505 16945
rect 1545 16905 1555 16945
rect 1595 16905 1605 16945
rect 1645 16905 1655 16945
rect 1695 16905 1705 16945
rect 1745 16905 1755 16945
rect 1795 16905 1805 16945
rect 1845 16905 1855 16945
rect 1895 16905 1905 16945
rect 1945 16905 1955 16945
rect 1995 16905 2005 16945
rect 2045 16905 2055 16945
rect 2095 16905 2105 16945
rect 2145 16905 2155 16945
rect 2195 16905 2205 16945
rect 2245 16905 2255 16945
rect 2295 16905 2305 16945
rect 2345 16905 2355 16945
rect 2395 16905 2405 16945
rect 2445 16905 2455 16945
rect 2495 16905 2505 16945
rect 2545 16905 2555 16945
rect 2595 16905 2605 16945
rect 2645 16905 2655 16945
rect 2695 16905 2705 16945
rect 2745 16905 2755 16945
rect 2795 16905 2805 16945
rect 2845 16905 2855 16945
rect 2895 16905 2905 16945
rect 2945 16905 2955 16945
rect 2995 16905 3005 16945
rect 3045 16905 3055 16945
rect 3095 16905 3105 16945
rect 3145 16905 3155 16945
rect 3195 16905 3205 16945
rect 3245 16905 3255 16945
rect 3295 16905 3305 16945
rect 3345 16905 3355 16945
rect 3395 16905 3405 16945
rect 3445 16905 3455 16945
rect 3495 16905 3505 16945
rect 3545 16905 3555 16945
rect 3595 16905 3605 16945
rect 3645 16905 3655 16945
rect 3695 16905 3705 16945
rect 3745 16905 3755 16945
rect 3795 16905 3805 16945
rect 3845 16905 3855 16945
rect 3895 16905 3905 16945
rect 3945 16905 3955 16945
rect 3995 16905 4005 16945
rect 4045 16905 4055 16945
rect 4095 16905 4105 16945
rect 4145 16905 4155 16945
rect 4195 16905 4205 16945
rect 4245 16905 4255 16945
rect 4295 16905 4305 16945
rect 4345 16905 4355 16945
rect 4395 16905 4405 16945
rect 4445 16905 4455 16945
rect 4495 16905 4505 16945
rect 4545 16905 4555 16945
rect 4595 16905 4605 16945
rect 4645 16905 4655 16945
rect 4695 16905 4705 16945
rect 4745 16905 4755 16945
rect 4795 16905 4805 16945
rect 4845 16905 4855 16945
rect 4895 16905 4905 16945
rect 4945 16905 4955 16945
rect 4995 16905 5005 16945
rect 5045 16905 5055 16945
rect 5095 16905 5105 16945
rect 5145 16905 5155 16945
rect 5195 16905 5205 16945
rect 5245 16905 5255 16945
rect 5295 16905 5305 16945
rect 5345 16905 5355 16945
rect 5395 16905 5405 16945
rect 5445 16905 5455 16945
rect 5495 16905 5505 16945
rect 5545 16905 5555 16945
rect 5595 16905 5605 16945
rect 5645 16905 5655 16945
rect 5695 16905 5705 16945
rect 5745 16905 5755 16945
rect 5795 16905 5805 16945
rect 5845 16905 5855 16945
rect 5895 16905 5905 16945
rect 5945 16905 5955 16945
rect 5995 16905 6005 16945
rect 6045 16905 6055 16945
rect 6095 16905 6105 16945
rect 6145 16905 6155 16945
rect 6195 16905 6205 16945
rect 6245 16905 6255 16945
rect 6295 16905 6305 16945
rect 6345 16905 6355 16945
rect 6395 16905 6405 16945
rect 6445 16905 6455 16945
rect 6495 16905 6505 16945
rect 6545 16905 6555 16945
rect 6595 16905 6605 16945
rect 6645 16905 6655 16945
rect 6695 16905 6705 16945
rect 6745 16905 6755 16945
rect 6795 16905 6805 16945
rect 6845 16905 6855 16945
rect 6895 16905 6905 16945
rect 6945 16905 6955 16945
rect 6995 16905 7005 16945
rect 7045 16905 7055 16945
rect 7095 16905 7105 16945
rect 7145 16905 7155 16945
rect 7195 16905 7205 16945
rect 7245 16905 7255 16945
rect 7295 16905 7305 16945
rect 7345 16905 7355 16945
rect 7395 16905 7405 16945
rect 7445 16905 7455 16945
rect 7495 16905 7505 16945
rect 7545 16905 7555 16945
rect 7595 16905 7605 16945
rect 7645 16905 7655 16945
rect 7695 16905 7705 16945
rect 7745 16905 7755 16945
rect 7795 16905 7805 16945
rect 7845 16905 7855 16945
rect 7895 16905 7905 16945
rect 7945 16905 7955 16945
rect 7995 16905 8005 16945
rect 8045 16905 8055 16945
rect 8095 16905 8105 16945
rect 8145 16905 8155 16945
rect 8195 16905 8205 16945
rect 8245 16905 8255 16945
rect 8295 16905 8305 16945
rect 8345 16905 8355 16945
rect 8395 16905 8405 16945
rect 8445 16905 8455 16945
rect 8495 16905 8505 16945
rect 8545 16905 8555 16945
rect 8595 16905 8605 16945
rect 8645 16905 8655 16945
rect 8695 16905 8705 16945
rect 8745 16905 8755 16945
rect 8795 16905 8805 16945
rect 8845 16905 8855 16945
rect 8895 16905 8905 16945
rect 8945 16905 8955 16945
rect 8995 16905 9005 16945
rect 9045 16905 9055 16945
rect 9095 16905 9105 16945
rect 9145 16905 9155 16945
rect 9195 16905 9205 16945
rect 9245 16905 9255 16945
rect 9295 16905 9305 16945
rect 9345 16905 9355 16945
rect 9395 16905 9405 16945
rect 9445 16905 9455 16945
rect 9495 16905 9505 16945
rect 9545 16905 9555 16945
rect 9595 16905 9605 16945
rect 9645 16905 9655 16945
rect 9695 16905 9705 16945
rect 9745 16905 9755 16945
rect 9795 16905 9805 16945
rect 9845 16905 9855 16945
rect 9895 16905 9905 16945
rect 9945 16905 9955 16945
rect 9995 16905 10005 16945
rect 10045 16905 10055 16945
rect 10095 16905 10105 16945
rect 10145 16905 10155 16945
rect 10195 16905 10205 16945
rect 10245 16905 10255 16945
rect 10295 16905 10305 16945
rect 10345 16905 10355 16945
rect 10395 16905 10405 16945
rect 10445 16905 10455 16945
rect 10495 16905 10505 16945
rect 10545 16905 10555 16945
rect 10595 16905 10605 16945
rect 10645 16905 10655 16945
rect 10695 16905 10705 16945
rect 10745 16905 10755 16945
rect 10795 16905 10805 16945
rect 10845 16905 10855 16945
rect 10895 16905 10905 16945
rect 10945 16905 10955 16945
rect 10995 16905 11005 16945
rect 11045 16905 11055 16945
rect 11095 16905 11105 16945
rect 11145 16905 11155 16945
rect 11195 16905 11205 16945
rect 11245 16905 11255 16945
rect 11295 16905 11305 16945
rect 11345 16905 11355 16945
rect 11395 16905 11405 16945
rect 11445 16905 11455 16945
rect 11495 16905 11505 16945
rect 11545 16905 11555 16945
rect 11595 16905 11605 16945
rect 11645 16905 11655 16945
rect 11695 16905 11705 16945
rect 11745 16905 11755 16945
rect 11795 16905 11805 16945
rect 11845 16905 11855 16945
rect 11895 16905 11905 16945
rect 11945 16905 11955 16945
rect 11995 16905 12005 16945
rect 12045 16905 12055 16945
rect 12095 16905 12105 16945
rect 12145 16905 12155 16945
rect 12195 16905 12205 16945
rect 12245 16905 12255 16945
rect 12295 16905 12305 16945
rect 12345 16905 12355 16945
rect 12395 16905 12405 16945
rect 12445 16905 12455 16945
rect 12495 16905 12505 16945
rect 12545 16905 12555 16945
rect 12595 16905 12605 16945
rect 12645 16905 12655 16945
rect 12695 16905 12705 16945
rect 12745 16905 12755 16945
rect 12795 16905 12805 16945
rect 12845 16905 12855 16945
rect 12895 16905 12905 16945
rect 12945 16905 12955 16945
rect 12995 16905 13005 16945
rect 13045 16905 13055 16945
rect 13095 16905 13105 16945
rect 13145 16905 13155 16945
rect 13195 16905 13205 16945
rect 13245 16905 13255 16945
rect 13295 16905 13305 16945
rect 13345 16905 13355 16945
rect 13395 16905 13405 16945
rect 13445 16905 13455 16945
rect 13495 16905 13505 16945
rect 13545 16905 13555 16945
rect 13595 16905 13605 16945
rect 13645 16905 13655 16945
rect 13695 16905 13705 16945
rect 13745 16905 13755 16945
rect 13795 16905 13805 16945
rect 13845 16905 13855 16945
rect 13895 16905 13905 16945
rect 13945 16905 13955 16945
rect 13995 16905 14005 16945
rect 14045 16905 14055 16945
rect 14095 16905 14105 16945
rect 14145 16905 14155 16945
rect 14195 16905 14205 16945
rect 14245 16905 14255 16945
rect 14295 16905 14305 16945
rect 14345 16905 14355 16945
rect 14395 16905 14405 16945
rect 14445 16905 14455 16945
rect 14495 16905 14505 16945
rect 14545 16905 14555 16945
rect 14595 16905 14605 16945
rect 14645 16905 14655 16945
rect 14695 16905 14705 16945
rect 14745 16905 14755 16945
rect 14795 16905 14805 16945
rect 14845 16905 14855 16945
rect 14895 16905 14905 16945
rect 14945 16905 14955 16945
rect 14995 16905 15005 16945
rect 15045 16905 15055 16945
rect 15095 16905 15105 16945
rect 15145 16905 15155 16945
rect 15195 16905 15205 16945
rect 15245 16905 15255 16945
rect 15295 16905 15305 16945
rect 15345 16905 15355 16945
rect 15395 16905 15405 16945
rect 15445 16905 15455 16945
rect 15495 16905 15505 16945
rect 15545 16905 15555 16945
rect 15595 16905 15605 16945
rect 15645 16905 15655 16945
rect 15695 16905 15705 16945
rect 15745 16905 15755 16945
rect 15795 16905 15805 16945
rect 15845 16905 15855 16945
rect 15895 16905 15905 16945
rect 15945 16905 15955 16945
rect 15995 16905 16005 16945
rect 16045 16905 16055 16945
rect 16095 16905 16105 16945
rect 16145 16905 16155 16945
rect 16195 16905 16205 16945
rect 16245 16905 16255 16945
rect 16295 16905 16305 16945
rect 16345 16905 16355 16945
rect 16395 16905 16405 16945
rect 16445 16905 16455 16945
rect 16495 16905 16505 16945
rect 16545 16905 16555 16945
rect 16595 16905 16605 16945
rect 16645 16905 16655 16945
rect 16695 16905 16705 16945
rect 16745 16905 16755 16945
rect 16795 16905 16805 16945
rect 16845 16905 16855 16945
rect 16895 16905 16905 16945
rect 16945 16905 16955 16945
rect 16995 16905 17005 16945
rect 17045 16905 17055 16945
rect 17095 16905 17105 16945
rect 17145 16905 17155 16945
rect 17195 16905 17205 16945
rect 17245 16905 17255 16945
rect 17295 16905 17305 16945
rect 17345 16905 17355 16945
rect 17395 16905 17405 16945
rect 17445 16905 17455 16945
rect 17495 16905 17505 16945
rect 17545 16905 17555 16945
rect 17595 16905 17605 16945
rect 17645 16905 17655 16945
rect 17695 16905 17705 16945
rect 17745 16905 17755 16945
rect 17795 16905 17805 16945
rect 17845 16905 17855 16945
rect 17895 16905 17905 16945
rect 17945 16905 17955 16945
rect 17995 16905 18005 16945
rect 18045 16905 18055 16945
rect 18095 16905 18105 16945
rect 18145 16905 18155 16945
rect 18195 16905 18205 16945
rect 18245 16905 18255 16945
rect 18295 16905 18305 16945
rect 18345 16905 18355 16945
rect 18395 16905 18405 16945
rect 18445 16905 18455 16945
rect 18495 16905 18505 16945
rect 18545 16905 18555 16945
rect 18595 16905 18605 16945
rect 18645 16905 18655 16945
rect 18695 16905 18705 16945
rect 18745 16905 18755 16945
rect 18795 16905 18805 16945
rect 18845 16905 18855 16945
rect 18895 16905 18905 16945
rect 18945 16905 18955 16945
rect 18995 16905 19005 16945
rect 19045 16905 19055 16945
rect 19095 16905 19105 16945
rect 19145 16905 19155 16945
rect 19195 16905 19205 16945
rect 19245 16905 19255 16945
rect 19295 16905 19305 16945
rect 19345 16905 19355 16945
rect 19395 16905 19405 16945
rect 19445 16905 19455 16945
rect 19495 16905 19505 16945
rect 19545 16905 19555 16945
rect 19595 16905 19605 16945
rect 19645 16905 19655 16945
rect 19695 16905 19705 16945
rect 19745 16905 19755 16945
rect 19795 16905 19805 16945
rect 19845 16905 19855 16945
rect 19895 16905 19905 16945
rect 19945 16905 19955 16945
rect 19995 16905 20005 16945
rect 20045 16905 20055 16945
rect 20095 16905 20105 16945
rect 20145 16905 20155 16945
rect 20195 16905 20205 16945
rect 20245 16905 20255 16945
rect 20295 16905 20305 16945
rect 20345 16905 20355 16945
rect 20395 16905 20405 16945
rect 20445 16905 20455 16945
rect 20495 16905 20505 16945
rect 20545 16905 20555 16945
rect 20595 16905 20605 16945
rect 20645 16905 20655 16945
rect 20695 16905 20705 16945
rect 20745 16905 20755 16945
rect 20795 16905 20805 16945
rect 20845 16905 20855 16945
rect 20895 16905 20905 16945
rect 20945 16905 20955 16945
rect 20995 16905 21005 16945
rect 21045 16905 21055 16945
rect 21095 16905 21105 16945
rect 21145 16905 21155 16945
rect 21195 16905 21205 16945
rect 21245 16905 21255 16945
rect 21295 16905 21305 16945
rect 21345 16905 21355 16945
rect 21395 16905 21405 16945
rect 21445 16905 21455 16945
rect 21495 16905 21505 16945
rect 21545 16905 21555 16945
rect 21595 16905 21605 16945
rect 21645 16905 21655 16945
rect 21695 16905 21705 16945
rect 21745 16905 21755 16945
rect 21795 16905 21805 16945
rect 21845 16905 21855 16945
rect 21895 16905 21905 16945
rect 21945 16905 21955 16945
rect 21995 16905 22005 16945
rect 22045 16905 22055 16945
rect 22095 16905 22105 16945
rect 22145 16905 22155 16945
rect 22195 16905 22205 16945
rect 22245 16905 22255 16945
rect 22295 16905 22305 16945
rect 22345 16905 22355 16945
rect 22395 16905 22405 16945
rect 22445 16905 22455 16945
rect 22495 16905 22505 16945
rect 22545 16905 22555 16945
rect 22595 16905 22605 16945
rect 22645 16905 22655 16945
rect 22695 16905 22705 16945
rect 22745 16905 22755 16945
rect 22795 16905 22805 16945
rect 22845 16905 22855 16945
rect 22895 16905 22905 16945
rect 22945 16905 22955 16945
rect 22995 16905 23005 16945
rect 23045 16905 23055 16945
rect 23095 16905 23105 16945
rect 23145 16905 23155 16945
rect 23195 16905 23205 16945
rect 23245 16905 23255 16945
rect 23295 16905 23305 16945
rect 23345 16905 23355 16945
rect 23395 16905 23405 16945
rect 23445 16905 23455 16945
rect 23495 16905 23505 16945
rect 23545 16905 23555 16945
rect 23595 16905 23605 16945
rect 23645 16905 23655 16945
rect 23695 16905 23705 16945
rect 23745 16905 23755 16945
rect 23795 16905 23805 16945
rect 23845 16905 23855 16945
rect 23895 16905 23905 16945
rect 23945 16905 23955 16945
rect 23995 16905 24005 16945
rect 24045 16905 24055 16945
rect 24095 16905 24105 16945
rect 24145 16905 24155 16945
rect 24195 16905 24205 16945
rect 24245 16905 24255 16945
rect 24295 16905 24305 16945
rect 24345 16905 24355 16945
rect 24395 16905 24405 16945
rect 24445 16905 24455 16945
rect 24495 16905 24505 16945
rect 24545 16905 24555 16945
rect 24595 16905 24605 16945
rect 24645 16905 24655 16945
rect 24695 16905 24705 16945
rect 24745 16905 24755 16945
rect 24795 16905 24805 16945
rect 24845 16905 24855 16945
rect 24895 16905 24905 16945
rect 24945 16905 24955 16945
rect 24995 16905 25005 16945
rect 25045 16905 25055 16945
rect 25095 16905 25105 16945
rect 25145 16905 25155 16945
rect 25195 16905 25205 16945
rect 25245 16905 25255 16945
rect 25295 16905 25305 16945
rect 25345 16905 25355 16945
rect 25395 16905 25405 16945
rect 25445 16905 25455 16945
rect 25495 16905 25505 16945
rect 25545 16905 25555 16945
rect 25595 16905 25605 16945
rect 25645 16905 25655 16945
rect 25695 16905 25705 16945
rect 25745 16905 25755 16945
rect 25795 16905 25805 16945
rect 25845 16905 25855 16945
rect 25895 16905 25905 16945
rect 25945 16905 25955 16945
rect 25995 16905 26005 16945
rect 26045 16905 26055 16945
rect 26095 16905 26105 16945
rect 26145 16905 26155 16945
rect 26195 16905 26205 16945
rect 26245 16905 26255 16945
rect 26295 16905 26305 16945
rect 26345 16905 26355 16945
rect 26395 16905 26405 16945
rect 26445 16905 26455 16945
rect 26495 16905 26505 16945
rect 26545 16905 26555 16945
rect 26595 16905 26605 16945
rect 26645 16905 26655 16945
rect 26695 16905 26705 16945
rect 26745 16905 26755 16945
rect 26795 16905 26805 16945
rect 26845 16905 26855 16945
rect 26895 16905 26905 16945
rect 26945 16905 26955 16945
rect 26995 16905 27005 16945
rect 27045 16905 27055 16945
rect 27095 16905 27105 16945
rect 27145 16905 27155 16945
rect 27195 16905 27205 16945
rect 27245 16905 27255 16945
rect 27295 16905 27305 16945
rect 27345 16905 27355 16945
rect 27395 16905 27405 16945
rect 27445 16905 27455 16945
rect 27495 16905 27505 16945
rect 27545 16905 27555 16945
rect 27595 16905 27605 16945
rect 27645 16905 27655 16945
rect 27695 16905 27705 16945
rect 27745 16905 27755 16945
rect 27795 16905 27805 16945
rect 27845 16905 27855 16945
rect 27895 16905 27905 16945
rect 27945 16905 27955 16945
rect 27995 16905 28005 16945
rect 28045 16905 28055 16945
rect 28095 16905 28105 16945
rect 28145 16905 28155 16945
rect 28195 16905 28205 16945
rect 28245 16905 28255 16945
rect 28295 16905 28305 16945
rect 28345 16905 28355 16945
rect 28395 16905 28405 16945
rect 28445 16905 28455 16945
rect 28495 16905 28505 16945
rect 28545 16905 28555 16945
rect 28595 16905 28605 16945
rect 28645 16905 28655 16945
rect 28695 16905 28705 16945
rect 28745 16905 28755 16945
rect 28795 16905 28805 16945
rect 28845 16905 28855 16945
rect 28895 16905 28905 16945
rect 28945 16905 28955 16945
rect 28995 16905 29005 16945
rect 29045 16905 29055 16945
rect 29095 16905 29105 16945
rect 29145 16905 29155 16945
rect 29195 16905 29205 16945
rect 29245 16905 29255 16945
rect 29295 16905 29305 16945
rect 29345 16905 29355 16945
rect 29395 16905 29405 16945
rect 29445 16905 29455 16945
rect 29495 16905 29505 16945
rect 29545 16905 29555 16945
rect 29595 16905 29605 16945
rect 29645 16905 29655 16945
rect 29695 16905 29705 16945
rect 29745 16905 29755 16945
rect 29795 16905 29805 16945
rect 29845 16905 29855 16945
rect 29895 16905 29905 16945
rect 29945 16905 29955 16945
rect 29995 16905 30005 16945
rect 30045 16905 30055 16945
rect 30095 16905 30105 16945
rect 30145 16905 30155 16945
rect 30195 16905 30205 16945
rect 30245 16905 30255 16945
rect 30295 16905 30305 16945
rect 30345 16905 30355 16945
rect 30395 16905 30405 16945
rect 30445 16905 30455 16945
rect 30495 16905 30505 16945
rect 30545 16905 30555 16945
rect 30595 16905 30605 16945
rect 30645 16905 30655 16945
rect 30695 16905 30705 16945
rect 30745 16905 30755 16945
rect 30795 16905 30805 16945
rect 30845 16905 30855 16945
rect 30895 16905 30905 16945
rect 30945 16905 30955 16945
rect 30995 16905 31005 16945
rect 31045 16905 31055 16945
rect 31095 16905 31105 16945
rect 31145 16905 31155 16945
rect 31195 16905 31205 16945
rect 31245 16905 31255 16945
rect 31295 16905 31305 16945
rect 31345 16905 31355 16945
rect 31395 16905 31405 16945
rect 31445 16905 31455 16945
rect 31495 16905 31505 16945
rect 31545 16905 31555 16945
rect 31595 16905 31605 16945
rect 31645 16905 31655 16945
rect 31695 16905 31705 16945
rect 31745 16905 31755 16945
rect 31795 16905 31805 16945
rect 31845 16905 31855 16945
rect 31895 16905 31905 16945
rect 31945 16905 31955 16945
rect 31995 16905 32005 16945
rect 32045 16905 32055 16945
rect 32095 16905 32105 16945
rect 32145 16905 32155 16945
rect 32195 16905 32205 16945
rect 32245 16905 32255 16945
rect 32295 16905 32305 16945
rect 32345 16905 32355 16945
rect 32395 16905 32405 16945
rect 32445 16905 32455 16945
rect 32495 16905 32505 16945
rect 32545 16905 32555 16945
rect 32595 16905 32605 16945
rect 32645 16905 32655 16945
rect 32695 16905 32705 16945
rect 32745 16905 32755 16945
rect 32795 16905 32805 16945
rect 32845 16905 32855 16945
rect 32895 16905 32905 16945
rect 32945 16905 32955 16945
rect 32995 16905 33005 16945
rect 33045 16905 33055 16945
rect 33095 16905 33105 16945
rect 33145 16905 33155 16945
rect 33195 16905 33205 16945
rect 33245 16905 33255 16945
rect 33295 16905 33305 16945
rect 33345 16905 33355 16945
rect 33395 16905 33405 16945
rect 33445 16905 33455 16945
rect 33495 16905 33505 16945
rect 33545 16905 33555 16945
rect 33595 16905 33605 16945
rect 33645 16905 33655 16945
rect 33695 16905 33705 16945
rect 33745 16905 33755 16945
rect 33795 16905 33805 16945
rect 33845 16905 33855 16945
rect 33895 16905 33905 16945
rect 33945 16905 33955 16945
rect 33995 16905 34005 16945
rect 34045 16905 34055 16945
rect 34095 16905 34105 16945
rect 34145 16905 34155 16945
rect 34195 16905 34205 16945
rect 34245 16905 34255 16945
rect 34295 16905 34305 16945
rect 34345 16905 34355 16945
rect 34395 16905 34405 16945
rect 34445 16905 34455 16945
rect 34495 16905 34505 16945
rect 34545 16905 34555 16945
rect 34595 16905 34605 16945
rect 34645 16905 34655 16945
rect 34695 16905 34705 16945
rect 34745 16905 34755 16945
rect 34795 16905 34805 16945
rect 34845 16905 34855 16945
rect 34895 16905 34905 16945
rect 34945 16905 34955 16945
rect 34995 16905 35005 16945
rect 35045 16905 35055 16945
rect 35095 16905 35105 16945
rect 35145 16905 35155 16945
rect 35195 16905 35205 16945
rect 35245 16905 35255 16945
rect 35295 16905 35305 16945
rect 35345 16905 35355 16945
rect 35395 16905 35405 16945
rect 35445 16905 35455 16945
rect 35495 16905 35505 16945
rect 35545 16905 35555 16945
rect 35595 16905 35605 16945
rect 35645 16905 35655 16945
rect 35695 16905 35705 16945
rect 35745 16905 35755 16945
rect 35795 16905 35805 16945
rect 35845 16905 35855 16945
rect 35895 16905 35905 16945
rect 35945 16905 35955 16945
rect 35995 16905 36005 16945
rect 36045 16905 36055 16945
rect 36095 16905 36105 16945
rect 36145 16905 36155 16945
rect 36195 16905 36205 16945
rect 36245 16905 36255 16945
rect 36295 16905 36305 16945
rect 36345 16905 36355 16945
rect 36395 16905 36405 16945
rect 36445 16905 36455 16945
rect 36495 16905 36505 16945
rect 36545 16905 36555 16945
rect 36595 16905 36605 16945
rect 36645 16905 36655 16945
rect 36695 16905 36705 16945
rect 36745 16905 36755 16945
rect 36795 16905 36805 16945
rect 36845 16905 36855 16945
rect 36895 16905 36905 16945
rect 36945 16905 36955 16945
rect 36995 16905 37005 16945
rect 37045 16905 37055 16945
rect 37095 16905 37105 16945
rect 37145 16905 37155 16945
rect 37195 16905 37205 16945
rect 37245 16905 37255 16945
rect 37295 16905 37305 16945
rect 37345 16905 37355 16945
rect 37395 16905 37405 16945
rect 37445 16905 37455 16945
rect 37495 16905 37505 16945
rect 37545 16905 37555 16945
rect 37595 16905 37605 16945
rect 37645 16905 37655 16945
rect 37695 16905 37705 16945
rect 37745 16905 37755 16945
rect 37795 16905 37805 16945
rect 37845 16905 37855 16945
rect 37895 16905 37905 16945
rect 37945 16905 37955 16945
rect 37995 16905 38005 16945
rect 38045 16905 38055 16945
rect 38095 16905 38105 16945
rect 38145 16905 38155 16945
rect 38195 16905 38205 16945
rect 38245 16905 38255 16945
rect 38295 16905 38305 16945
rect 38345 16905 38355 16945
rect 38395 16905 38405 16945
rect 38445 16905 38455 16945
rect 38495 16905 38505 16945
rect 38545 16905 38555 16945
rect 38595 16905 38605 16945
rect 38645 16905 38655 16945
rect 38695 16905 38705 16945
rect 38745 16905 38755 16945
rect 38795 16905 38805 16945
rect 38845 16905 38855 16945
rect 38895 16905 38905 16945
rect 38945 16905 38955 16945
rect 38995 16905 39005 16945
rect 39045 16905 39055 16945
rect 39095 16905 39105 16945
rect 39145 16905 39155 16945
rect 39195 16905 39205 16945
rect 39245 16905 39255 16945
rect 39295 16905 39305 16945
rect 39345 16905 39355 16945
rect 39395 16905 39405 16945
rect 39445 16905 39455 16945
rect 39495 16905 39505 16945
rect 39545 16905 39555 16945
rect 39595 16905 39605 16945
rect 39645 16905 39655 16945
rect 39695 16905 39705 16945
rect 39745 16905 39750 16945
rect 0 16900 39750 16905
rect 0 15850 50 16900
rect 100 16845 39750 16850
rect 100 16805 105 16845
rect 145 16805 155 16845
rect 195 16805 205 16845
rect 245 16805 255 16845
rect 295 16805 305 16845
rect 345 16805 355 16845
rect 395 16805 405 16845
rect 445 16805 455 16845
rect 495 16805 505 16845
rect 545 16805 555 16845
rect 595 16805 605 16845
rect 645 16805 655 16845
rect 695 16805 705 16845
rect 745 16805 755 16845
rect 795 16805 805 16845
rect 845 16805 855 16845
rect 895 16805 905 16845
rect 945 16805 955 16845
rect 995 16805 1005 16845
rect 1045 16805 1055 16845
rect 1095 16805 1105 16845
rect 1145 16805 1155 16845
rect 1195 16805 1205 16845
rect 1245 16805 1255 16845
rect 1295 16805 1305 16845
rect 1345 16805 1355 16845
rect 1395 16805 1405 16845
rect 1445 16805 1455 16845
rect 1495 16805 1505 16845
rect 1545 16805 1555 16845
rect 1595 16805 1605 16845
rect 1645 16805 1655 16845
rect 1695 16805 1705 16845
rect 1745 16805 1755 16845
rect 1795 16805 1805 16845
rect 1845 16805 1855 16845
rect 1895 16805 1905 16845
rect 1945 16805 1955 16845
rect 1995 16805 2005 16845
rect 2045 16805 2055 16845
rect 2095 16805 2105 16845
rect 2145 16805 2155 16845
rect 2195 16805 2205 16845
rect 2245 16805 2255 16845
rect 2295 16805 2305 16845
rect 2345 16805 2355 16845
rect 2395 16805 2405 16845
rect 2445 16805 2455 16845
rect 2495 16805 2505 16845
rect 2545 16805 2555 16845
rect 2595 16805 2605 16845
rect 2645 16805 2655 16845
rect 2695 16805 2705 16845
rect 2745 16805 2755 16845
rect 2795 16805 2805 16845
rect 2845 16805 2855 16845
rect 2895 16805 2905 16845
rect 2945 16805 2955 16845
rect 2995 16805 3005 16845
rect 3045 16805 3055 16845
rect 3095 16805 3105 16845
rect 3145 16805 3155 16845
rect 3195 16805 3205 16845
rect 3245 16805 3255 16845
rect 3295 16805 3305 16845
rect 3345 16805 3355 16845
rect 3395 16805 3405 16845
rect 3445 16805 3455 16845
rect 3495 16805 3505 16845
rect 3545 16805 3555 16845
rect 3595 16805 3605 16845
rect 3645 16805 3655 16845
rect 3695 16805 3705 16845
rect 3745 16805 3755 16845
rect 3795 16805 3805 16845
rect 3845 16805 3855 16845
rect 3895 16805 3905 16845
rect 3945 16805 3955 16845
rect 3995 16805 4005 16845
rect 4045 16805 4055 16845
rect 4095 16805 4105 16845
rect 4145 16805 4155 16845
rect 4195 16805 4205 16845
rect 4245 16805 4255 16845
rect 4295 16805 4305 16845
rect 4345 16805 4355 16845
rect 4395 16805 4405 16845
rect 4445 16805 4455 16845
rect 4495 16805 4505 16845
rect 4545 16805 4555 16845
rect 4595 16805 4605 16845
rect 4645 16805 4655 16845
rect 4695 16805 4705 16845
rect 4745 16805 4755 16845
rect 4795 16805 4805 16845
rect 4845 16805 4855 16845
rect 4895 16805 4905 16845
rect 4945 16805 4955 16845
rect 4995 16805 5005 16845
rect 5045 16805 5055 16845
rect 5095 16805 5105 16845
rect 5145 16805 5155 16845
rect 5195 16805 5205 16845
rect 5245 16805 5255 16845
rect 5295 16805 5305 16845
rect 5345 16805 5355 16845
rect 5395 16805 5405 16845
rect 5445 16805 5455 16845
rect 5495 16805 5505 16845
rect 5545 16805 5555 16845
rect 5595 16805 5605 16845
rect 5645 16805 5655 16845
rect 5695 16805 5705 16845
rect 5745 16805 5755 16845
rect 5795 16805 5805 16845
rect 5845 16805 5855 16845
rect 5895 16805 5905 16845
rect 5945 16805 5955 16845
rect 5995 16805 6005 16845
rect 6045 16805 6055 16845
rect 6095 16805 6105 16845
rect 6145 16805 6155 16845
rect 6195 16805 6205 16845
rect 6245 16805 6255 16845
rect 6295 16805 6305 16845
rect 6345 16805 6355 16845
rect 6395 16805 6405 16845
rect 6445 16805 6455 16845
rect 6495 16805 6505 16845
rect 6545 16805 6555 16845
rect 6595 16805 6605 16845
rect 6645 16805 6655 16845
rect 6695 16805 6705 16845
rect 6745 16805 6755 16845
rect 6795 16805 6805 16845
rect 6845 16805 6855 16845
rect 6895 16805 6905 16845
rect 6945 16805 6955 16845
rect 6995 16805 7005 16845
rect 7045 16805 7055 16845
rect 7095 16805 7105 16845
rect 7145 16805 7155 16845
rect 7195 16805 7205 16845
rect 7245 16805 7255 16845
rect 7295 16805 7305 16845
rect 7345 16805 7355 16845
rect 7395 16805 7405 16845
rect 7445 16805 7455 16845
rect 7495 16805 7505 16845
rect 7545 16805 7555 16845
rect 7595 16805 7605 16845
rect 7645 16805 7655 16845
rect 7695 16805 7705 16845
rect 7745 16805 7755 16845
rect 7795 16805 7805 16845
rect 7845 16805 7855 16845
rect 7895 16805 7905 16845
rect 7945 16805 7955 16845
rect 7995 16805 8005 16845
rect 8045 16805 8055 16845
rect 8095 16805 8105 16845
rect 8145 16805 8155 16845
rect 8195 16805 8205 16845
rect 8245 16805 8255 16845
rect 8295 16805 8305 16845
rect 8345 16805 8355 16845
rect 8395 16805 8405 16845
rect 8445 16805 8455 16845
rect 8495 16805 8505 16845
rect 8545 16805 8555 16845
rect 8595 16805 8605 16845
rect 8645 16805 8655 16845
rect 8695 16805 8705 16845
rect 8745 16805 8755 16845
rect 8795 16805 8805 16845
rect 8845 16805 8855 16845
rect 8895 16805 8905 16845
rect 8945 16805 8955 16845
rect 8995 16805 9005 16845
rect 9045 16805 9055 16845
rect 9095 16805 9105 16845
rect 9145 16805 9155 16845
rect 9195 16805 9205 16845
rect 9245 16805 9255 16845
rect 9295 16805 9305 16845
rect 9345 16805 9355 16845
rect 9395 16805 9405 16845
rect 9445 16805 9455 16845
rect 9495 16805 9505 16845
rect 9545 16805 9555 16845
rect 9595 16805 9605 16845
rect 9645 16805 9655 16845
rect 9695 16805 9705 16845
rect 9745 16805 9755 16845
rect 9795 16805 9805 16845
rect 9845 16805 9855 16845
rect 9895 16805 9905 16845
rect 9945 16805 9955 16845
rect 9995 16805 10005 16845
rect 10045 16805 10055 16845
rect 10095 16805 10105 16845
rect 10145 16805 10155 16845
rect 10195 16805 10205 16845
rect 10245 16805 10255 16845
rect 10295 16805 10305 16845
rect 10345 16805 10355 16845
rect 10395 16805 10405 16845
rect 10445 16805 10455 16845
rect 10495 16805 10505 16845
rect 10545 16805 10555 16845
rect 10595 16805 10605 16845
rect 10645 16805 10655 16845
rect 10695 16805 10705 16845
rect 10745 16805 10755 16845
rect 10795 16805 10805 16845
rect 10845 16805 10855 16845
rect 10895 16805 10905 16845
rect 10945 16805 10955 16845
rect 10995 16805 11005 16845
rect 11045 16805 11055 16845
rect 11095 16805 11105 16845
rect 11145 16805 11155 16845
rect 11195 16805 11205 16845
rect 11245 16805 11255 16845
rect 11295 16805 11305 16845
rect 11345 16805 11355 16845
rect 11395 16805 11405 16845
rect 11445 16805 11455 16845
rect 11495 16805 11505 16845
rect 11545 16805 11555 16845
rect 11595 16805 11605 16845
rect 11645 16805 11655 16845
rect 11695 16805 11705 16845
rect 11745 16805 11755 16845
rect 11795 16805 11805 16845
rect 11845 16805 11855 16845
rect 11895 16805 11905 16845
rect 11945 16805 11955 16845
rect 11995 16805 12005 16845
rect 12045 16805 12055 16845
rect 12095 16805 12105 16845
rect 12145 16805 12155 16845
rect 12195 16805 12205 16845
rect 12245 16805 12255 16845
rect 12295 16805 12305 16845
rect 12345 16805 12355 16845
rect 12395 16805 12405 16845
rect 12445 16805 12455 16845
rect 12495 16805 12505 16845
rect 12545 16805 12555 16845
rect 12595 16805 12605 16845
rect 12645 16805 12655 16845
rect 12695 16805 12705 16845
rect 12745 16805 12755 16845
rect 12795 16805 12805 16845
rect 12845 16805 12855 16845
rect 12895 16805 12905 16845
rect 12945 16805 12955 16845
rect 12995 16805 13005 16845
rect 13045 16805 13055 16845
rect 13095 16805 13105 16845
rect 13145 16805 13155 16845
rect 13195 16805 13205 16845
rect 13245 16805 13255 16845
rect 13295 16805 13305 16845
rect 13345 16805 13355 16845
rect 13395 16805 13405 16845
rect 13445 16805 13455 16845
rect 13495 16805 13505 16845
rect 13545 16805 13555 16845
rect 13595 16805 13605 16845
rect 13645 16805 13655 16845
rect 13695 16805 13705 16845
rect 13745 16805 13755 16845
rect 13795 16805 13805 16845
rect 13845 16805 13855 16845
rect 13895 16805 13905 16845
rect 13945 16805 13955 16845
rect 13995 16805 14005 16845
rect 14045 16805 14055 16845
rect 14095 16805 14105 16845
rect 14145 16805 14155 16845
rect 14195 16805 14205 16845
rect 14245 16805 14255 16845
rect 14295 16805 14305 16845
rect 14345 16805 14355 16845
rect 14395 16805 14405 16845
rect 14445 16805 14455 16845
rect 14495 16805 14505 16845
rect 14545 16805 14555 16845
rect 14595 16805 14605 16845
rect 14645 16805 14655 16845
rect 14695 16805 14705 16845
rect 14745 16805 14755 16845
rect 14795 16805 14805 16845
rect 14845 16805 14855 16845
rect 14895 16805 14905 16845
rect 14945 16805 14955 16845
rect 14995 16805 15005 16845
rect 15045 16805 15055 16845
rect 15095 16805 15105 16845
rect 15145 16805 15155 16845
rect 15195 16805 15205 16845
rect 15245 16805 15255 16845
rect 15295 16805 15305 16845
rect 15345 16805 15355 16845
rect 15395 16805 15405 16845
rect 15445 16805 15455 16845
rect 15495 16805 15505 16845
rect 15545 16805 15555 16845
rect 15595 16805 15605 16845
rect 15645 16805 15655 16845
rect 15695 16805 15705 16845
rect 15745 16805 15755 16845
rect 15795 16805 15805 16845
rect 15845 16805 15855 16845
rect 15895 16805 15905 16845
rect 15945 16805 15955 16845
rect 15995 16805 16005 16845
rect 16045 16805 16055 16845
rect 16095 16805 16105 16845
rect 16145 16805 16155 16845
rect 16195 16805 16205 16845
rect 16245 16805 16255 16845
rect 16295 16805 16305 16845
rect 16345 16805 16355 16845
rect 16395 16805 16405 16845
rect 16445 16805 16455 16845
rect 16495 16805 16505 16845
rect 16545 16805 16555 16845
rect 16595 16805 16605 16845
rect 16645 16805 16655 16845
rect 16695 16805 16705 16845
rect 16745 16805 16755 16845
rect 16795 16805 16805 16845
rect 16845 16805 16855 16845
rect 16895 16805 16905 16845
rect 16945 16805 16955 16845
rect 16995 16805 17005 16845
rect 17045 16805 17055 16845
rect 17095 16805 17105 16845
rect 17145 16805 17155 16845
rect 17195 16805 17205 16845
rect 17245 16805 17255 16845
rect 17295 16805 17305 16845
rect 17345 16805 17355 16845
rect 17395 16805 17405 16845
rect 17445 16805 17455 16845
rect 17495 16805 17505 16845
rect 17545 16805 17555 16845
rect 17595 16805 17605 16845
rect 17645 16805 17655 16845
rect 17695 16805 17705 16845
rect 17745 16805 17755 16845
rect 17795 16805 17805 16845
rect 17845 16805 17855 16845
rect 17895 16805 17905 16845
rect 17945 16805 17955 16845
rect 17995 16805 18005 16845
rect 18045 16805 18055 16845
rect 18095 16805 18105 16845
rect 18145 16805 18155 16845
rect 18195 16805 18205 16845
rect 18245 16805 18255 16845
rect 18295 16805 18305 16845
rect 18345 16805 18355 16845
rect 18395 16805 18405 16845
rect 18445 16805 18455 16845
rect 18495 16805 18505 16845
rect 18545 16805 18555 16845
rect 18595 16805 18605 16845
rect 18645 16805 18655 16845
rect 18695 16805 18705 16845
rect 18745 16805 18755 16845
rect 18795 16805 18805 16845
rect 18845 16805 18855 16845
rect 18895 16805 18905 16845
rect 18945 16805 18955 16845
rect 18995 16805 19005 16845
rect 19045 16805 19055 16845
rect 19095 16805 19105 16845
rect 19145 16805 19155 16845
rect 19195 16805 19205 16845
rect 19245 16805 19255 16845
rect 19295 16805 19305 16845
rect 19345 16805 19355 16845
rect 19395 16805 19405 16845
rect 19445 16805 19455 16845
rect 19495 16805 19505 16845
rect 19545 16805 19555 16845
rect 19595 16805 19605 16845
rect 19645 16805 19655 16845
rect 19695 16805 19705 16845
rect 19745 16805 19755 16845
rect 19795 16805 19805 16845
rect 19845 16805 19855 16845
rect 19895 16805 19905 16845
rect 19945 16805 19955 16845
rect 19995 16805 20005 16845
rect 20045 16805 20055 16845
rect 20095 16805 20105 16845
rect 20145 16805 20155 16845
rect 20195 16805 20205 16845
rect 20245 16805 20255 16845
rect 20295 16805 20305 16845
rect 20345 16805 20355 16845
rect 20395 16805 20405 16845
rect 20445 16805 20455 16845
rect 20495 16805 20505 16845
rect 20545 16805 20555 16845
rect 20595 16805 20605 16845
rect 20645 16805 20655 16845
rect 20695 16805 20705 16845
rect 20745 16805 20755 16845
rect 20795 16805 20805 16845
rect 20845 16805 20855 16845
rect 20895 16805 20905 16845
rect 20945 16805 20955 16845
rect 20995 16805 21005 16845
rect 21045 16805 21055 16845
rect 21095 16805 21105 16845
rect 21145 16805 21155 16845
rect 21195 16805 21205 16845
rect 21245 16805 21255 16845
rect 21295 16805 21305 16845
rect 21345 16805 21355 16845
rect 21395 16805 21405 16845
rect 21445 16805 21455 16845
rect 21495 16805 21505 16845
rect 21545 16805 21555 16845
rect 21595 16805 21605 16845
rect 21645 16805 21655 16845
rect 21695 16805 21705 16845
rect 21745 16805 21755 16845
rect 21795 16805 21805 16845
rect 21845 16805 21855 16845
rect 21895 16805 21905 16845
rect 21945 16805 21955 16845
rect 21995 16805 22005 16845
rect 22045 16805 22055 16845
rect 22095 16805 22105 16845
rect 22145 16805 22155 16845
rect 22195 16805 22205 16845
rect 22245 16805 22255 16845
rect 22295 16805 22305 16845
rect 22345 16805 22355 16845
rect 22395 16805 22405 16845
rect 22445 16805 22455 16845
rect 22495 16805 22505 16845
rect 22545 16805 22555 16845
rect 22595 16805 22605 16845
rect 22645 16805 22655 16845
rect 22695 16805 22705 16845
rect 22745 16805 22755 16845
rect 22795 16805 22805 16845
rect 22845 16805 22855 16845
rect 22895 16805 22905 16845
rect 22945 16805 22955 16845
rect 22995 16805 23005 16845
rect 23045 16805 23055 16845
rect 23095 16805 23105 16845
rect 23145 16805 23155 16845
rect 23195 16805 23205 16845
rect 23245 16805 23255 16845
rect 23295 16805 23305 16845
rect 23345 16805 23355 16845
rect 23395 16805 23405 16845
rect 23445 16805 23455 16845
rect 23495 16805 23505 16845
rect 23545 16805 23555 16845
rect 23595 16805 23605 16845
rect 23645 16805 23655 16845
rect 23695 16805 23705 16845
rect 23745 16805 23755 16845
rect 23795 16805 23805 16845
rect 23845 16805 23855 16845
rect 23895 16805 23905 16845
rect 23945 16805 23955 16845
rect 23995 16805 24005 16845
rect 24045 16805 24055 16845
rect 24095 16805 24105 16845
rect 24145 16805 24155 16845
rect 24195 16805 24205 16845
rect 24245 16805 24255 16845
rect 24295 16805 24305 16845
rect 24345 16805 24355 16845
rect 24395 16805 24405 16845
rect 24445 16805 24455 16845
rect 24495 16805 24505 16845
rect 24545 16805 24555 16845
rect 24595 16805 24605 16845
rect 24645 16805 24655 16845
rect 24695 16805 24705 16845
rect 24745 16805 24755 16845
rect 24795 16805 24805 16845
rect 24845 16805 24855 16845
rect 24895 16805 24905 16845
rect 24945 16805 24955 16845
rect 24995 16805 25005 16845
rect 25045 16805 25055 16845
rect 25095 16805 25105 16845
rect 25145 16805 25155 16845
rect 25195 16805 25205 16845
rect 25245 16805 25255 16845
rect 25295 16805 25305 16845
rect 25345 16805 25355 16845
rect 25395 16805 25405 16845
rect 25445 16805 25455 16845
rect 25495 16805 25505 16845
rect 25545 16805 25555 16845
rect 25595 16805 25605 16845
rect 25645 16805 25655 16845
rect 25695 16805 25705 16845
rect 25745 16805 25755 16845
rect 25795 16805 25805 16845
rect 25845 16805 25855 16845
rect 25895 16805 25905 16845
rect 25945 16805 25955 16845
rect 25995 16805 26005 16845
rect 26045 16805 26055 16845
rect 26095 16805 26105 16845
rect 26145 16805 26155 16845
rect 26195 16805 26205 16845
rect 26245 16805 26255 16845
rect 26295 16805 26305 16845
rect 26345 16805 26355 16845
rect 26395 16805 26405 16845
rect 26445 16805 26455 16845
rect 26495 16805 26505 16845
rect 26545 16805 26555 16845
rect 26595 16805 26605 16845
rect 26645 16805 26655 16845
rect 26695 16805 26705 16845
rect 26745 16805 26755 16845
rect 26795 16805 26805 16845
rect 26845 16805 26855 16845
rect 26895 16805 26905 16845
rect 26945 16805 26955 16845
rect 26995 16805 27005 16845
rect 27045 16805 27055 16845
rect 27095 16805 27105 16845
rect 27145 16805 27155 16845
rect 27195 16805 27205 16845
rect 27245 16805 27255 16845
rect 27295 16805 27305 16845
rect 27345 16805 27355 16845
rect 27395 16805 27405 16845
rect 27445 16805 27455 16845
rect 27495 16805 27505 16845
rect 27545 16805 27555 16845
rect 27595 16805 27605 16845
rect 27645 16805 27655 16845
rect 27695 16805 27705 16845
rect 27745 16805 27755 16845
rect 27795 16805 27805 16845
rect 27845 16805 27855 16845
rect 27895 16805 27905 16845
rect 27945 16805 27955 16845
rect 27995 16805 28005 16845
rect 28045 16805 28055 16845
rect 28095 16805 28105 16845
rect 28145 16805 28155 16845
rect 28195 16805 28205 16845
rect 28245 16805 28255 16845
rect 28295 16805 28305 16845
rect 28345 16805 28355 16845
rect 28395 16805 28405 16845
rect 28445 16805 28455 16845
rect 28495 16805 28505 16845
rect 28545 16805 28555 16845
rect 28595 16805 28605 16845
rect 28645 16805 28655 16845
rect 28695 16805 28705 16845
rect 28745 16805 28755 16845
rect 28795 16805 28805 16845
rect 28845 16805 28855 16845
rect 28895 16805 28905 16845
rect 28945 16805 28955 16845
rect 28995 16805 29005 16845
rect 29045 16805 29055 16845
rect 29095 16805 29105 16845
rect 29145 16805 29155 16845
rect 29195 16805 29205 16845
rect 29245 16805 29255 16845
rect 29295 16805 29305 16845
rect 29345 16805 29355 16845
rect 29395 16805 29405 16845
rect 29445 16805 29455 16845
rect 29495 16805 29505 16845
rect 29545 16805 29555 16845
rect 29595 16805 29605 16845
rect 29645 16805 29655 16845
rect 29695 16805 29705 16845
rect 29745 16805 29755 16845
rect 29795 16805 29805 16845
rect 29845 16805 29855 16845
rect 29895 16805 29905 16845
rect 29945 16805 29955 16845
rect 29995 16805 30005 16845
rect 30045 16805 30055 16845
rect 30095 16805 30105 16845
rect 30145 16805 30155 16845
rect 30195 16805 30205 16845
rect 30245 16805 30255 16845
rect 30295 16805 30305 16845
rect 30345 16805 30355 16845
rect 30395 16805 30405 16845
rect 30445 16805 30455 16845
rect 30495 16805 30505 16845
rect 30545 16805 30555 16845
rect 30595 16805 30605 16845
rect 30645 16805 30655 16845
rect 30695 16805 30705 16845
rect 30745 16805 30755 16845
rect 30795 16805 30805 16845
rect 30845 16805 30855 16845
rect 30895 16805 30905 16845
rect 30945 16805 30955 16845
rect 30995 16805 31005 16845
rect 31045 16805 31055 16845
rect 31095 16805 31105 16845
rect 31145 16805 31155 16845
rect 31195 16805 31205 16845
rect 31245 16805 31255 16845
rect 31295 16805 31305 16845
rect 31345 16805 31355 16845
rect 31395 16805 31405 16845
rect 31445 16805 31455 16845
rect 31495 16805 31505 16845
rect 31545 16805 31555 16845
rect 31595 16805 31605 16845
rect 31645 16805 31655 16845
rect 31695 16805 31705 16845
rect 31745 16805 31755 16845
rect 31795 16805 31805 16845
rect 31845 16805 31855 16845
rect 31895 16805 31905 16845
rect 31945 16805 31955 16845
rect 31995 16805 32005 16845
rect 32045 16805 32055 16845
rect 32095 16805 32105 16845
rect 32145 16805 32155 16845
rect 32195 16805 32205 16845
rect 32245 16805 32255 16845
rect 32295 16805 32305 16845
rect 32345 16805 32355 16845
rect 32395 16805 32405 16845
rect 32445 16805 32455 16845
rect 32495 16805 32505 16845
rect 32545 16805 32555 16845
rect 32595 16805 32605 16845
rect 32645 16805 32655 16845
rect 32695 16805 32705 16845
rect 32745 16805 32755 16845
rect 32795 16805 32805 16845
rect 32845 16805 32855 16845
rect 32895 16805 32905 16845
rect 32945 16805 32955 16845
rect 32995 16805 33005 16845
rect 33045 16805 33055 16845
rect 33095 16805 33105 16845
rect 33145 16805 33155 16845
rect 33195 16805 33205 16845
rect 33245 16805 33255 16845
rect 33295 16805 33305 16845
rect 33345 16805 33355 16845
rect 33395 16805 33405 16845
rect 33445 16805 33455 16845
rect 33495 16805 33505 16845
rect 33545 16805 33555 16845
rect 33595 16805 33605 16845
rect 33645 16805 33655 16845
rect 33695 16805 33705 16845
rect 33745 16805 33755 16845
rect 33795 16805 33805 16845
rect 33845 16805 33855 16845
rect 33895 16805 33905 16845
rect 33945 16805 33955 16845
rect 33995 16805 34005 16845
rect 34045 16805 34055 16845
rect 34095 16805 34105 16845
rect 34145 16805 34155 16845
rect 34195 16805 34205 16845
rect 34245 16805 34255 16845
rect 34295 16805 34305 16845
rect 34345 16805 34355 16845
rect 34395 16805 34405 16845
rect 34445 16805 34455 16845
rect 34495 16805 34505 16845
rect 34545 16805 34555 16845
rect 34595 16805 34605 16845
rect 34645 16805 34655 16845
rect 34695 16805 34705 16845
rect 34745 16805 34755 16845
rect 34795 16805 34805 16845
rect 34845 16805 34855 16845
rect 34895 16805 34905 16845
rect 34945 16805 34955 16845
rect 34995 16805 35005 16845
rect 35045 16805 35055 16845
rect 35095 16805 35105 16845
rect 35145 16805 35155 16845
rect 35195 16805 35205 16845
rect 35245 16805 35255 16845
rect 35295 16805 35305 16845
rect 35345 16805 35355 16845
rect 35395 16805 35405 16845
rect 35445 16805 35455 16845
rect 35495 16805 35505 16845
rect 35545 16805 35555 16845
rect 35595 16805 35605 16845
rect 35645 16805 35655 16845
rect 35695 16805 35705 16845
rect 35745 16805 35755 16845
rect 35795 16805 35805 16845
rect 35845 16805 35855 16845
rect 35895 16805 35905 16845
rect 35945 16805 35955 16845
rect 35995 16805 36005 16845
rect 36045 16805 36055 16845
rect 36095 16805 36105 16845
rect 36145 16805 36155 16845
rect 36195 16805 36205 16845
rect 36245 16805 36255 16845
rect 36295 16805 36305 16845
rect 36345 16805 36355 16845
rect 36395 16805 36405 16845
rect 36445 16805 36455 16845
rect 36495 16805 36505 16845
rect 36545 16805 36555 16845
rect 36595 16805 36605 16845
rect 36645 16805 36655 16845
rect 36695 16805 36705 16845
rect 36745 16805 36755 16845
rect 36795 16805 36805 16845
rect 36845 16805 36855 16845
rect 36895 16805 36905 16845
rect 36945 16805 36955 16845
rect 36995 16805 37005 16845
rect 37045 16805 37055 16845
rect 37095 16805 37105 16845
rect 37145 16805 37155 16845
rect 37195 16805 37205 16845
rect 37245 16805 37255 16845
rect 37295 16805 37305 16845
rect 37345 16805 37355 16845
rect 37395 16805 37405 16845
rect 37445 16805 37455 16845
rect 37495 16805 37505 16845
rect 37545 16805 37555 16845
rect 37595 16805 37605 16845
rect 37645 16805 37655 16845
rect 37695 16805 37705 16845
rect 37745 16805 37755 16845
rect 37795 16805 37805 16845
rect 37845 16805 37855 16845
rect 37895 16805 37905 16845
rect 37945 16805 37955 16845
rect 37995 16805 38005 16845
rect 38045 16805 38055 16845
rect 38095 16805 38105 16845
rect 38145 16805 38155 16845
rect 38195 16805 38205 16845
rect 38245 16805 38255 16845
rect 38295 16805 38305 16845
rect 38345 16805 38355 16845
rect 38395 16805 38405 16845
rect 38445 16805 38455 16845
rect 38495 16805 38505 16845
rect 38545 16805 38555 16845
rect 38595 16805 38605 16845
rect 38645 16805 38655 16845
rect 38695 16805 38705 16845
rect 38745 16805 38755 16845
rect 38795 16805 38805 16845
rect 38845 16805 38855 16845
rect 38895 16805 38905 16845
rect 38945 16805 38955 16845
rect 38995 16805 39005 16845
rect 39045 16805 39055 16845
rect 39095 16805 39105 16845
rect 39145 16805 39155 16845
rect 39195 16805 39205 16845
rect 39245 16805 39255 16845
rect 39295 16805 39305 16845
rect 39345 16805 39355 16845
rect 39395 16805 39405 16845
rect 39445 16805 39455 16845
rect 39495 16805 39505 16845
rect 39545 16805 39555 16845
rect 39595 16805 39605 16845
rect 39645 16805 39655 16845
rect 39695 16805 39705 16845
rect 39745 16805 39750 16845
rect 100 16800 39750 16805
rect 100 16650 3200 16800
rect 100 16000 200 16650
rect 3100 16000 3200 16650
rect 100 15900 3200 16000
rect 3350 16650 6450 16800
rect 3350 16000 3450 16650
rect 6350 16000 6450 16650
rect 3350 15900 6450 16000
rect 6600 16650 9700 16800
rect 6600 16000 6700 16650
rect 9600 16000 9700 16650
rect 6600 15900 9700 16000
rect 9850 16650 12950 16800
rect 9850 16000 9950 16650
rect 12850 16000 12950 16650
rect 9850 15900 12950 16000
rect 13100 16650 16200 16800
rect 13100 16000 13200 16650
rect 16100 16000 16200 16650
rect 13100 15900 16200 16000
rect 16350 16650 19450 16800
rect 16350 16000 16450 16650
rect 19350 16000 19450 16650
rect 16350 15900 19450 16000
rect 19600 16650 22700 16800
rect 19600 16000 19700 16650
rect 22600 16000 22700 16650
rect 19600 15900 22700 16000
rect 22850 16650 25950 16800
rect 22850 16000 22950 16650
rect 25850 16000 25950 16650
rect 22850 15900 25950 16000
rect 26100 16650 29200 16800
rect 26100 16000 26200 16650
rect 29100 16000 29200 16650
rect 26100 15900 29200 16000
rect 29350 16650 32450 16800
rect 29350 16000 29450 16650
rect 32350 16000 32450 16650
rect 29350 15900 32450 16000
rect 32600 16650 35700 16800
rect 32600 16000 32700 16650
rect 35600 16000 35700 16650
rect 32600 15900 35700 16000
rect 35850 16650 38950 16800
rect 35850 16000 35950 16650
rect 38850 16000 38950 16650
rect 35850 15900 38950 16000
rect 39100 16650 39750 16800
rect 39100 16000 39200 16650
rect 39650 16000 39750 16650
rect 39100 15900 39750 16000
rect 0 15845 39750 15850
rect 0 15805 5 15845
rect 45 15805 55 15845
rect 95 15805 105 15845
rect 145 15805 155 15845
rect 195 15805 205 15845
rect 245 15805 255 15845
rect 295 15805 305 15845
rect 345 15805 355 15845
rect 395 15805 405 15845
rect 445 15805 455 15845
rect 495 15805 505 15845
rect 545 15805 555 15845
rect 595 15805 605 15845
rect 645 15805 655 15845
rect 695 15805 705 15845
rect 745 15805 755 15845
rect 795 15805 805 15845
rect 845 15805 855 15845
rect 895 15805 905 15845
rect 945 15805 955 15845
rect 995 15805 1005 15845
rect 1045 15805 1055 15845
rect 1095 15805 1105 15845
rect 1145 15805 1155 15845
rect 1195 15805 1205 15845
rect 1245 15805 1255 15845
rect 1295 15805 1305 15845
rect 1345 15805 1355 15845
rect 1395 15805 1405 15845
rect 1445 15805 1455 15845
rect 1495 15805 1505 15845
rect 1545 15805 1555 15845
rect 1595 15805 1605 15845
rect 1645 15805 1655 15845
rect 1695 15805 1705 15845
rect 1745 15805 1755 15845
rect 1795 15805 1805 15845
rect 1845 15805 1855 15845
rect 1895 15805 1905 15845
rect 1945 15805 1955 15845
rect 1995 15805 2005 15845
rect 2045 15805 2055 15845
rect 2095 15805 2105 15845
rect 2145 15805 2155 15845
rect 2195 15805 2205 15845
rect 2245 15805 2255 15845
rect 2295 15805 2305 15845
rect 2345 15805 2355 15845
rect 2395 15805 2405 15845
rect 2445 15805 2455 15845
rect 2495 15805 2505 15845
rect 2545 15805 2555 15845
rect 2595 15805 2605 15845
rect 2645 15805 2655 15845
rect 2695 15805 2705 15845
rect 2745 15805 2755 15845
rect 2795 15805 2805 15845
rect 2845 15805 2855 15845
rect 2895 15805 2905 15845
rect 2945 15805 2955 15845
rect 2995 15805 3005 15845
rect 3045 15805 3055 15845
rect 3095 15805 3105 15845
rect 3145 15805 3155 15845
rect 3195 15805 3205 15845
rect 3245 15805 3255 15845
rect 3295 15805 3305 15845
rect 3345 15805 3355 15845
rect 3395 15805 3405 15845
rect 3445 15805 3455 15845
rect 3495 15805 3505 15845
rect 3545 15805 3555 15845
rect 3595 15805 3605 15845
rect 3645 15805 3655 15845
rect 3695 15805 3705 15845
rect 3745 15805 3755 15845
rect 3795 15805 3805 15845
rect 3845 15805 3855 15845
rect 3895 15805 3905 15845
rect 3945 15805 3955 15845
rect 3995 15805 4005 15845
rect 4045 15805 4055 15845
rect 4095 15805 4105 15845
rect 4145 15805 4155 15845
rect 4195 15805 4205 15845
rect 4245 15805 4255 15845
rect 4295 15805 4305 15845
rect 4345 15805 4355 15845
rect 4395 15805 4405 15845
rect 4445 15805 4455 15845
rect 4495 15805 4505 15845
rect 4545 15805 4555 15845
rect 4595 15805 4605 15845
rect 4645 15805 4655 15845
rect 4695 15805 4705 15845
rect 4745 15805 4755 15845
rect 4795 15805 4805 15845
rect 4845 15805 4855 15845
rect 4895 15805 4905 15845
rect 4945 15805 4955 15845
rect 4995 15805 5005 15845
rect 5045 15805 5055 15845
rect 5095 15805 5105 15845
rect 5145 15805 5155 15845
rect 5195 15805 5205 15845
rect 5245 15805 5255 15845
rect 5295 15805 5305 15845
rect 5345 15805 5355 15845
rect 5395 15805 5405 15845
rect 5445 15805 5455 15845
rect 5495 15805 5505 15845
rect 5545 15805 5555 15845
rect 5595 15805 5605 15845
rect 5645 15805 5655 15845
rect 5695 15805 5705 15845
rect 5745 15805 5755 15845
rect 5795 15805 5805 15845
rect 5845 15805 5855 15845
rect 5895 15805 5905 15845
rect 5945 15805 5955 15845
rect 5995 15805 6005 15845
rect 6045 15805 6055 15845
rect 6095 15805 6105 15845
rect 6145 15805 6155 15845
rect 6195 15805 6205 15845
rect 6245 15805 6255 15845
rect 6295 15805 6305 15845
rect 6345 15805 6355 15845
rect 6395 15805 6405 15845
rect 6445 15805 6455 15845
rect 6495 15805 6505 15845
rect 6545 15805 6555 15845
rect 6595 15805 6605 15845
rect 6645 15805 6655 15845
rect 6695 15805 6705 15845
rect 6745 15805 6755 15845
rect 6795 15805 6805 15845
rect 6845 15805 6855 15845
rect 6895 15805 6905 15845
rect 6945 15805 6955 15845
rect 6995 15805 7005 15845
rect 7045 15805 7055 15845
rect 7095 15805 7105 15845
rect 7145 15805 7155 15845
rect 7195 15805 7205 15845
rect 7245 15805 7255 15845
rect 7295 15805 7305 15845
rect 7345 15805 7355 15845
rect 7395 15805 7405 15845
rect 7445 15805 7455 15845
rect 7495 15805 7505 15845
rect 7545 15805 7555 15845
rect 7595 15805 7605 15845
rect 7645 15805 7655 15845
rect 7695 15805 7705 15845
rect 7745 15805 7755 15845
rect 7795 15805 7805 15845
rect 7845 15805 7855 15845
rect 7895 15805 7905 15845
rect 7945 15805 7955 15845
rect 7995 15805 8005 15845
rect 8045 15805 8055 15845
rect 8095 15805 8105 15845
rect 8145 15805 8155 15845
rect 8195 15805 8205 15845
rect 8245 15805 8255 15845
rect 8295 15805 8305 15845
rect 8345 15805 8355 15845
rect 8395 15805 8405 15845
rect 8445 15805 8455 15845
rect 8495 15805 8505 15845
rect 8545 15805 8555 15845
rect 8595 15805 8605 15845
rect 8645 15805 8655 15845
rect 8695 15805 8705 15845
rect 8745 15805 8755 15845
rect 8795 15805 8805 15845
rect 8845 15805 8855 15845
rect 8895 15805 8905 15845
rect 8945 15805 8955 15845
rect 8995 15805 9005 15845
rect 9045 15805 9055 15845
rect 9095 15805 9105 15845
rect 9145 15805 9155 15845
rect 9195 15805 9205 15845
rect 9245 15805 9255 15845
rect 9295 15805 9305 15845
rect 9345 15805 9355 15845
rect 9395 15805 9405 15845
rect 9445 15805 9455 15845
rect 9495 15805 9505 15845
rect 9545 15805 9555 15845
rect 9595 15805 9605 15845
rect 9645 15805 9655 15845
rect 9695 15805 9705 15845
rect 9745 15805 9755 15845
rect 9795 15805 9805 15845
rect 9845 15805 9855 15845
rect 9895 15805 9905 15845
rect 9945 15805 9955 15845
rect 9995 15805 10005 15845
rect 10045 15805 10055 15845
rect 10095 15805 10105 15845
rect 10145 15805 10155 15845
rect 10195 15805 10205 15845
rect 10245 15805 10255 15845
rect 10295 15805 10305 15845
rect 10345 15805 10355 15845
rect 10395 15805 10405 15845
rect 10445 15805 10455 15845
rect 10495 15805 10505 15845
rect 10545 15805 10555 15845
rect 10595 15805 10605 15845
rect 10645 15805 10655 15845
rect 10695 15805 10705 15845
rect 10745 15805 10755 15845
rect 10795 15805 10805 15845
rect 10845 15805 10855 15845
rect 10895 15805 10905 15845
rect 10945 15805 10955 15845
rect 10995 15805 11005 15845
rect 11045 15805 11055 15845
rect 11095 15805 11105 15845
rect 11145 15805 11155 15845
rect 11195 15805 11205 15845
rect 11245 15805 11255 15845
rect 11295 15805 11305 15845
rect 11345 15805 11355 15845
rect 11395 15805 11405 15845
rect 11445 15805 11455 15845
rect 11495 15805 11505 15845
rect 11545 15805 11555 15845
rect 11595 15805 11605 15845
rect 11645 15805 11655 15845
rect 11695 15805 11705 15845
rect 11745 15805 11755 15845
rect 11795 15805 11805 15845
rect 11845 15805 11855 15845
rect 11895 15805 11905 15845
rect 11945 15805 11955 15845
rect 11995 15805 12005 15845
rect 12045 15805 12055 15845
rect 12095 15805 12105 15845
rect 12145 15805 12155 15845
rect 12195 15805 12205 15845
rect 12245 15805 12255 15845
rect 12295 15805 12305 15845
rect 12345 15805 12355 15845
rect 12395 15805 12405 15845
rect 12445 15805 12455 15845
rect 12495 15805 12505 15845
rect 12545 15805 12555 15845
rect 12595 15805 12605 15845
rect 12645 15805 12655 15845
rect 12695 15805 12705 15845
rect 12745 15805 12755 15845
rect 12795 15805 12805 15845
rect 12845 15805 12855 15845
rect 12895 15805 12905 15845
rect 12945 15805 12955 15845
rect 12995 15805 13005 15845
rect 13045 15805 13055 15845
rect 13095 15805 13105 15845
rect 13145 15805 13155 15845
rect 13195 15805 13205 15845
rect 13245 15805 13255 15845
rect 13295 15805 13305 15845
rect 13345 15805 13355 15845
rect 13395 15805 13405 15845
rect 13445 15805 13455 15845
rect 13495 15805 13505 15845
rect 13545 15805 13555 15845
rect 13595 15805 13605 15845
rect 13645 15805 13655 15845
rect 13695 15805 13705 15845
rect 13745 15805 13755 15845
rect 13795 15805 13805 15845
rect 13845 15805 13855 15845
rect 13895 15805 13905 15845
rect 13945 15805 13955 15845
rect 13995 15805 14005 15845
rect 14045 15805 14055 15845
rect 14095 15805 14105 15845
rect 14145 15805 14155 15845
rect 14195 15805 14205 15845
rect 14245 15805 14255 15845
rect 14295 15805 14305 15845
rect 14345 15805 14355 15845
rect 14395 15805 14405 15845
rect 14445 15805 14455 15845
rect 14495 15805 14505 15845
rect 14545 15805 14555 15845
rect 14595 15805 14605 15845
rect 14645 15805 14655 15845
rect 14695 15805 14705 15845
rect 14745 15805 14755 15845
rect 14795 15805 14805 15845
rect 14845 15805 14855 15845
rect 14895 15805 14905 15845
rect 14945 15805 14955 15845
rect 14995 15805 15005 15845
rect 15045 15805 15055 15845
rect 15095 15805 15105 15845
rect 15145 15805 15155 15845
rect 15195 15805 15205 15845
rect 15245 15805 15255 15845
rect 15295 15805 15305 15845
rect 15345 15805 15355 15845
rect 15395 15805 15405 15845
rect 15445 15805 15455 15845
rect 15495 15805 15505 15845
rect 15545 15805 15555 15845
rect 15595 15805 15605 15845
rect 15645 15805 15655 15845
rect 15695 15805 15705 15845
rect 15745 15805 15755 15845
rect 15795 15805 15805 15845
rect 15845 15805 15855 15845
rect 15895 15805 15905 15845
rect 15945 15805 15955 15845
rect 15995 15805 16005 15845
rect 16045 15805 16055 15845
rect 16095 15805 16105 15845
rect 16145 15805 16155 15845
rect 16195 15805 16205 15845
rect 16245 15805 16255 15845
rect 16295 15805 16305 15845
rect 16345 15805 16355 15845
rect 16395 15805 16405 15845
rect 16445 15805 16455 15845
rect 16495 15805 16505 15845
rect 16545 15805 16555 15845
rect 16595 15805 16605 15845
rect 16645 15805 16655 15845
rect 16695 15805 16705 15845
rect 16745 15805 16755 15845
rect 16795 15805 16805 15845
rect 16845 15805 16855 15845
rect 16895 15805 16905 15845
rect 16945 15805 16955 15845
rect 16995 15805 17005 15845
rect 17045 15805 17055 15845
rect 17095 15805 17105 15845
rect 17145 15805 17155 15845
rect 17195 15805 17205 15845
rect 17245 15805 17255 15845
rect 17295 15805 17305 15845
rect 17345 15805 17355 15845
rect 17395 15805 17405 15845
rect 17445 15805 17455 15845
rect 17495 15805 17505 15845
rect 17545 15805 17555 15845
rect 17595 15805 17605 15845
rect 17645 15805 17655 15845
rect 17695 15805 17705 15845
rect 17745 15805 17755 15845
rect 17795 15805 17805 15845
rect 17845 15805 17855 15845
rect 17895 15805 17905 15845
rect 17945 15805 17955 15845
rect 17995 15805 18005 15845
rect 18045 15805 18055 15845
rect 18095 15805 18105 15845
rect 18145 15805 18155 15845
rect 18195 15805 18205 15845
rect 18245 15805 18255 15845
rect 18295 15805 18305 15845
rect 18345 15805 18355 15845
rect 18395 15805 18405 15845
rect 18445 15805 18455 15845
rect 18495 15805 18505 15845
rect 18545 15805 18555 15845
rect 18595 15805 18605 15845
rect 18645 15805 18655 15845
rect 18695 15805 18705 15845
rect 18745 15805 18755 15845
rect 18795 15805 18805 15845
rect 18845 15805 18855 15845
rect 18895 15805 18905 15845
rect 18945 15805 18955 15845
rect 18995 15805 19005 15845
rect 19045 15805 19055 15845
rect 19095 15805 19105 15845
rect 19145 15805 19155 15845
rect 19195 15805 19205 15845
rect 19245 15805 19255 15845
rect 19295 15805 19305 15845
rect 19345 15805 19355 15845
rect 19395 15805 19405 15845
rect 19445 15805 19455 15845
rect 19495 15805 19505 15845
rect 19545 15805 19555 15845
rect 19595 15805 19605 15845
rect 19645 15805 19655 15845
rect 19695 15805 19705 15845
rect 19745 15805 19755 15845
rect 19795 15805 19805 15845
rect 19845 15805 19855 15845
rect 19895 15805 19905 15845
rect 19945 15805 19955 15845
rect 19995 15805 20005 15845
rect 20045 15805 20055 15845
rect 20095 15805 20105 15845
rect 20145 15805 20155 15845
rect 20195 15805 20205 15845
rect 20245 15805 20255 15845
rect 20295 15805 20305 15845
rect 20345 15805 20355 15845
rect 20395 15805 20405 15845
rect 20445 15805 20455 15845
rect 20495 15805 20505 15845
rect 20545 15805 20555 15845
rect 20595 15805 20605 15845
rect 20645 15805 20655 15845
rect 20695 15805 20705 15845
rect 20745 15805 20755 15845
rect 20795 15805 20805 15845
rect 20845 15805 20855 15845
rect 20895 15805 20905 15845
rect 20945 15805 20955 15845
rect 20995 15805 21005 15845
rect 21045 15805 21055 15845
rect 21095 15805 21105 15845
rect 21145 15805 21155 15845
rect 21195 15805 21205 15845
rect 21245 15805 21255 15845
rect 21295 15805 21305 15845
rect 21345 15805 21355 15845
rect 21395 15805 21405 15845
rect 21445 15805 21455 15845
rect 21495 15805 21505 15845
rect 21545 15805 21555 15845
rect 21595 15805 21605 15845
rect 21645 15805 21655 15845
rect 21695 15805 21705 15845
rect 21745 15805 21755 15845
rect 21795 15805 21805 15845
rect 21845 15805 21855 15845
rect 21895 15805 21905 15845
rect 21945 15805 21955 15845
rect 21995 15805 22005 15845
rect 22045 15805 22055 15845
rect 22095 15805 22105 15845
rect 22145 15805 22155 15845
rect 22195 15805 22205 15845
rect 22245 15805 22255 15845
rect 22295 15805 22305 15845
rect 22345 15805 22355 15845
rect 22395 15805 22405 15845
rect 22445 15805 22455 15845
rect 22495 15805 22505 15845
rect 22545 15805 22555 15845
rect 22595 15805 22605 15845
rect 22645 15805 22655 15845
rect 22695 15805 22705 15845
rect 22745 15805 22755 15845
rect 22795 15805 22805 15845
rect 22845 15805 22855 15845
rect 22895 15805 22905 15845
rect 22945 15805 22955 15845
rect 22995 15805 23005 15845
rect 23045 15805 23055 15845
rect 23095 15805 23105 15845
rect 23145 15805 23155 15845
rect 23195 15805 23205 15845
rect 23245 15805 23255 15845
rect 23295 15805 23305 15845
rect 23345 15805 23355 15845
rect 23395 15805 23405 15845
rect 23445 15805 23455 15845
rect 23495 15805 23505 15845
rect 23545 15805 23555 15845
rect 23595 15805 23605 15845
rect 23645 15805 23655 15845
rect 23695 15805 23705 15845
rect 23745 15805 23755 15845
rect 23795 15805 23805 15845
rect 23845 15805 23855 15845
rect 23895 15805 23905 15845
rect 23945 15805 23955 15845
rect 23995 15805 24005 15845
rect 24045 15805 24055 15845
rect 24095 15805 24105 15845
rect 24145 15805 24155 15845
rect 24195 15805 24205 15845
rect 24245 15805 24255 15845
rect 24295 15805 24305 15845
rect 24345 15805 24355 15845
rect 24395 15805 24405 15845
rect 24445 15805 24455 15845
rect 24495 15805 24505 15845
rect 24545 15805 24555 15845
rect 24595 15805 24605 15845
rect 24645 15805 24655 15845
rect 24695 15805 24705 15845
rect 24745 15805 24755 15845
rect 24795 15805 24805 15845
rect 24845 15805 24855 15845
rect 24895 15805 24905 15845
rect 24945 15805 24955 15845
rect 24995 15805 25005 15845
rect 25045 15805 25055 15845
rect 25095 15805 25105 15845
rect 25145 15805 25155 15845
rect 25195 15805 25205 15845
rect 25245 15805 25255 15845
rect 25295 15805 25305 15845
rect 25345 15805 25355 15845
rect 25395 15805 25405 15845
rect 25445 15805 25455 15845
rect 25495 15805 25505 15845
rect 25545 15805 25555 15845
rect 25595 15805 25605 15845
rect 25645 15805 25655 15845
rect 25695 15805 25705 15845
rect 25745 15805 25755 15845
rect 25795 15805 25805 15845
rect 25845 15805 25855 15845
rect 25895 15805 25905 15845
rect 25945 15805 25955 15845
rect 25995 15805 26005 15845
rect 26045 15805 26055 15845
rect 26095 15805 26105 15845
rect 26145 15805 26155 15845
rect 26195 15805 26205 15845
rect 26245 15805 26255 15845
rect 26295 15805 26305 15845
rect 26345 15805 26355 15845
rect 26395 15805 26405 15845
rect 26445 15805 26455 15845
rect 26495 15805 26505 15845
rect 26545 15805 26555 15845
rect 26595 15805 26605 15845
rect 26645 15805 26655 15845
rect 26695 15805 26705 15845
rect 26745 15805 26755 15845
rect 26795 15805 26805 15845
rect 26845 15805 26855 15845
rect 26895 15805 26905 15845
rect 26945 15805 26955 15845
rect 26995 15805 27005 15845
rect 27045 15805 27055 15845
rect 27095 15805 27105 15845
rect 27145 15805 27155 15845
rect 27195 15805 27205 15845
rect 27245 15805 27255 15845
rect 27295 15805 27305 15845
rect 27345 15805 27355 15845
rect 27395 15805 27405 15845
rect 27445 15805 27455 15845
rect 27495 15805 27505 15845
rect 27545 15805 27555 15845
rect 27595 15805 27605 15845
rect 27645 15805 27655 15845
rect 27695 15805 27705 15845
rect 27745 15805 27755 15845
rect 27795 15805 27805 15845
rect 27845 15805 27855 15845
rect 27895 15805 27905 15845
rect 27945 15805 27955 15845
rect 27995 15805 28005 15845
rect 28045 15805 28055 15845
rect 28095 15805 28105 15845
rect 28145 15805 28155 15845
rect 28195 15805 28205 15845
rect 28245 15805 28255 15845
rect 28295 15805 28305 15845
rect 28345 15805 28355 15845
rect 28395 15805 28405 15845
rect 28445 15805 28455 15845
rect 28495 15805 28505 15845
rect 28545 15805 28555 15845
rect 28595 15805 28605 15845
rect 28645 15805 28655 15845
rect 28695 15805 28705 15845
rect 28745 15805 28755 15845
rect 28795 15805 28805 15845
rect 28845 15805 28855 15845
rect 28895 15805 28905 15845
rect 28945 15805 28955 15845
rect 28995 15805 29005 15845
rect 29045 15805 29055 15845
rect 29095 15805 29105 15845
rect 29145 15805 29155 15845
rect 29195 15805 29205 15845
rect 29245 15805 29255 15845
rect 29295 15805 29305 15845
rect 29345 15805 29355 15845
rect 29395 15805 29405 15845
rect 29445 15805 29455 15845
rect 29495 15805 29505 15845
rect 29545 15805 29555 15845
rect 29595 15805 29605 15845
rect 29645 15805 29655 15845
rect 29695 15805 29705 15845
rect 29745 15805 29755 15845
rect 29795 15805 29805 15845
rect 29845 15805 29855 15845
rect 29895 15805 29905 15845
rect 29945 15805 29955 15845
rect 29995 15805 30005 15845
rect 30045 15805 30055 15845
rect 30095 15805 30105 15845
rect 30145 15805 30155 15845
rect 30195 15805 30205 15845
rect 30245 15805 30255 15845
rect 30295 15805 30305 15845
rect 30345 15805 30355 15845
rect 30395 15805 30405 15845
rect 30445 15805 30455 15845
rect 30495 15805 30505 15845
rect 30545 15805 30555 15845
rect 30595 15805 30605 15845
rect 30645 15805 30655 15845
rect 30695 15805 30705 15845
rect 30745 15805 30755 15845
rect 30795 15805 30805 15845
rect 30845 15805 30855 15845
rect 30895 15805 30905 15845
rect 30945 15805 30955 15845
rect 30995 15805 31005 15845
rect 31045 15805 31055 15845
rect 31095 15805 31105 15845
rect 31145 15805 31155 15845
rect 31195 15805 31205 15845
rect 31245 15805 31255 15845
rect 31295 15805 31305 15845
rect 31345 15805 31355 15845
rect 31395 15805 31405 15845
rect 31445 15805 31455 15845
rect 31495 15805 31505 15845
rect 31545 15805 31555 15845
rect 31595 15805 31605 15845
rect 31645 15805 31655 15845
rect 31695 15805 31705 15845
rect 31745 15805 31755 15845
rect 31795 15805 31805 15845
rect 31845 15805 31855 15845
rect 31895 15805 31905 15845
rect 31945 15805 31955 15845
rect 31995 15805 32005 15845
rect 32045 15805 32055 15845
rect 32095 15805 32105 15845
rect 32145 15805 32155 15845
rect 32195 15805 32205 15845
rect 32245 15805 32255 15845
rect 32295 15805 32305 15845
rect 32345 15805 32355 15845
rect 32395 15805 32405 15845
rect 32445 15805 32455 15845
rect 32495 15805 32505 15845
rect 32545 15805 32555 15845
rect 32595 15805 32605 15845
rect 32645 15805 32655 15845
rect 32695 15805 32705 15845
rect 32745 15805 32755 15845
rect 32795 15805 32805 15845
rect 32845 15805 32855 15845
rect 32895 15805 32905 15845
rect 32945 15805 32955 15845
rect 32995 15805 33005 15845
rect 33045 15805 33055 15845
rect 33095 15805 33105 15845
rect 33145 15805 33155 15845
rect 33195 15805 33205 15845
rect 33245 15805 33255 15845
rect 33295 15805 33305 15845
rect 33345 15805 33355 15845
rect 33395 15805 33405 15845
rect 33445 15805 33455 15845
rect 33495 15805 33505 15845
rect 33545 15805 33555 15845
rect 33595 15805 33605 15845
rect 33645 15805 33655 15845
rect 33695 15805 33705 15845
rect 33745 15805 33755 15845
rect 33795 15805 33805 15845
rect 33845 15805 33855 15845
rect 33895 15805 33905 15845
rect 33945 15805 33955 15845
rect 33995 15805 34005 15845
rect 34045 15805 34055 15845
rect 34095 15805 34105 15845
rect 34145 15805 34155 15845
rect 34195 15805 34205 15845
rect 34245 15805 34255 15845
rect 34295 15805 34305 15845
rect 34345 15805 34355 15845
rect 34395 15805 34405 15845
rect 34445 15805 34455 15845
rect 34495 15805 34505 15845
rect 34545 15805 34555 15845
rect 34595 15805 34605 15845
rect 34645 15805 34655 15845
rect 34695 15805 34705 15845
rect 34745 15805 34755 15845
rect 34795 15805 34805 15845
rect 34845 15805 34855 15845
rect 34895 15805 34905 15845
rect 34945 15805 34955 15845
rect 34995 15805 35005 15845
rect 35045 15805 35055 15845
rect 35095 15805 35105 15845
rect 35145 15805 35155 15845
rect 35195 15805 35205 15845
rect 35245 15805 35255 15845
rect 35295 15805 35305 15845
rect 35345 15805 35355 15845
rect 35395 15805 35405 15845
rect 35445 15805 35455 15845
rect 35495 15805 35505 15845
rect 35545 15805 35555 15845
rect 35595 15805 35605 15845
rect 35645 15805 35655 15845
rect 35695 15805 35705 15845
rect 35745 15805 35755 15845
rect 35795 15805 35805 15845
rect 35845 15805 35855 15845
rect 35895 15805 35905 15845
rect 35945 15805 35955 15845
rect 35995 15805 36005 15845
rect 36045 15805 36055 15845
rect 36095 15805 36105 15845
rect 36145 15805 36155 15845
rect 36195 15805 36205 15845
rect 36245 15805 36255 15845
rect 36295 15805 36305 15845
rect 36345 15805 36355 15845
rect 36395 15805 36405 15845
rect 36445 15805 36455 15845
rect 36495 15805 36505 15845
rect 36545 15805 36555 15845
rect 36595 15805 36605 15845
rect 36645 15805 36655 15845
rect 36695 15805 36705 15845
rect 36745 15805 36755 15845
rect 36795 15805 36805 15845
rect 36845 15805 36855 15845
rect 36895 15805 36905 15845
rect 36945 15805 36955 15845
rect 36995 15805 37005 15845
rect 37045 15805 37055 15845
rect 37095 15805 37105 15845
rect 37145 15805 37155 15845
rect 37195 15805 37205 15845
rect 37245 15805 37255 15845
rect 37295 15805 37305 15845
rect 37345 15805 37355 15845
rect 37395 15805 37405 15845
rect 37445 15805 37455 15845
rect 37495 15805 37505 15845
rect 37545 15805 37555 15845
rect 37595 15805 37605 15845
rect 37645 15805 37655 15845
rect 37695 15805 37705 15845
rect 37745 15805 37755 15845
rect 37795 15805 37805 15845
rect 37845 15805 37855 15845
rect 37895 15805 37905 15845
rect 37945 15805 37955 15845
rect 37995 15805 38005 15845
rect 38045 15805 38055 15845
rect 38095 15805 38105 15845
rect 38145 15805 38155 15845
rect 38195 15805 38205 15845
rect 38245 15805 38255 15845
rect 38295 15805 38305 15845
rect 38345 15805 38355 15845
rect 38395 15805 38405 15845
rect 38445 15805 38455 15845
rect 38495 15805 38505 15845
rect 38545 15805 38555 15845
rect 38595 15805 38605 15845
rect 38645 15805 38655 15845
rect 38695 15805 38705 15845
rect 38745 15805 38755 15845
rect 38795 15805 38805 15845
rect 38845 15805 38855 15845
rect 38895 15805 38905 15845
rect 38945 15805 38955 15845
rect 38995 15805 39005 15845
rect 39045 15805 39055 15845
rect 39095 15805 39105 15845
rect 39145 15805 39155 15845
rect 39195 15805 39205 15845
rect 39245 15805 39255 15845
rect 39295 15805 39305 15845
rect 39345 15805 39355 15845
rect 39395 15805 39405 15845
rect 39445 15805 39455 15845
rect 39495 15805 39505 15845
rect 39545 15805 39555 15845
rect 39595 15805 39605 15845
rect 39645 15805 39655 15845
rect 39695 15805 39705 15845
rect 39745 15805 39750 15845
rect 0 15745 39750 15805
rect 0 15705 5 15745
rect 45 15705 55 15745
rect 95 15705 105 15745
rect 145 15705 155 15745
rect 195 15705 205 15745
rect 245 15705 255 15745
rect 295 15705 305 15745
rect 345 15705 355 15745
rect 395 15705 405 15745
rect 445 15705 455 15745
rect 495 15705 505 15745
rect 545 15705 555 15745
rect 595 15705 605 15745
rect 645 15705 655 15745
rect 695 15705 705 15745
rect 745 15705 755 15745
rect 795 15705 805 15745
rect 845 15705 855 15745
rect 895 15705 905 15745
rect 945 15705 955 15745
rect 995 15705 1005 15745
rect 1045 15705 1055 15745
rect 1095 15705 1105 15745
rect 1145 15705 1155 15745
rect 1195 15705 1205 15745
rect 1245 15705 1255 15745
rect 1295 15705 1305 15745
rect 1345 15705 1355 15745
rect 1395 15705 1405 15745
rect 1445 15705 1455 15745
rect 1495 15705 1505 15745
rect 1545 15705 1555 15745
rect 1595 15705 1605 15745
rect 1645 15705 1655 15745
rect 1695 15705 1705 15745
rect 1745 15705 1755 15745
rect 1795 15705 1805 15745
rect 1845 15705 1855 15745
rect 1895 15705 1905 15745
rect 1945 15705 1955 15745
rect 1995 15705 2005 15745
rect 2045 15705 2055 15745
rect 2095 15705 2105 15745
rect 2145 15705 2155 15745
rect 2195 15705 2205 15745
rect 2245 15705 2255 15745
rect 2295 15705 2305 15745
rect 2345 15705 2355 15745
rect 2395 15705 2405 15745
rect 2445 15705 2455 15745
rect 2495 15705 2505 15745
rect 2545 15705 2555 15745
rect 2595 15705 2605 15745
rect 2645 15705 2655 15745
rect 2695 15705 2705 15745
rect 2745 15705 2755 15745
rect 2795 15705 2805 15745
rect 2845 15705 2855 15745
rect 2895 15705 2905 15745
rect 2945 15705 2955 15745
rect 2995 15705 3005 15745
rect 3045 15705 3055 15745
rect 3095 15705 3105 15745
rect 3145 15705 3155 15745
rect 3195 15705 3205 15745
rect 3245 15705 3255 15745
rect 3295 15705 3305 15745
rect 3345 15705 3355 15745
rect 3395 15705 3405 15745
rect 3445 15705 3455 15745
rect 3495 15705 3505 15745
rect 3545 15705 3555 15745
rect 3595 15705 3605 15745
rect 3645 15705 3655 15745
rect 3695 15705 3705 15745
rect 3745 15705 3755 15745
rect 3795 15705 3805 15745
rect 3845 15705 3855 15745
rect 3895 15705 3905 15745
rect 3945 15705 3955 15745
rect 3995 15705 4005 15745
rect 4045 15705 4055 15745
rect 4095 15705 4105 15745
rect 4145 15705 4155 15745
rect 4195 15705 4205 15745
rect 4245 15705 4255 15745
rect 4295 15705 4305 15745
rect 4345 15705 4355 15745
rect 4395 15705 4405 15745
rect 4445 15705 4455 15745
rect 4495 15705 4505 15745
rect 4545 15705 4555 15745
rect 4595 15705 4605 15745
rect 4645 15705 4655 15745
rect 4695 15705 4705 15745
rect 4745 15705 4755 15745
rect 4795 15705 4805 15745
rect 4845 15705 4855 15745
rect 4895 15705 4905 15745
rect 4945 15705 4955 15745
rect 4995 15705 5005 15745
rect 5045 15705 5055 15745
rect 5095 15705 5105 15745
rect 5145 15705 5155 15745
rect 5195 15705 5205 15745
rect 5245 15705 5255 15745
rect 5295 15705 5305 15745
rect 5345 15705 5355 15745
rect 5395 15705 5405 15745
rect 5445 15705 5455 15745
rect 5495 15705 5505 15745
rect 5545 15705 5555 15745
rect 5595 15705 5605 15745
rect 5645 15705 5655 15745
rect 5695 15705 5705 15745
rect 5745 15705 5755 15745
rect 5795 15705 5805 15745
rect 5845 15705 5855 15745
rect 5895 15705 5905 15745
rect 5945 15705 5955 15745
rect 5995 15705 6005 15745
rect 6045 15705 6055 15745
rect 6095 15705 6105 15745
rect 6145 15705 6155 15745
rect 6195 15705 6205 15745
rect 6245 15705 6255 15745
rect 6295 15705 6305 15745
rect 6345 15705 6355 15745
rect 6395 15705 6405 15745
rect 6445 15705 6455 15745
rect 6495 15705 6505 15745
rect 6545 15705 6555 15745
rect 6595 15705 6605 15745
rect 6645 15705 6655 15745
rect 6695 15705 6705 15745
rect 6745 15705 6755 15745
rect 6795 15705 6805 15745
rect 6845 15705 6855 15745
rect 6895 15705 6905 15745
rect 6945 15705 6955 15745
rect 6995 15705 7005 15745
rect 7045 15705 7055 15745
rect 7095 15705 7105 15745
rect 7145 15705 7155 15745
rect 7195 15705 7205 15745
rect 7245 15705 7255 15745
rect 7295 15705 7305 15745
rect 7345 15705 7355 15745
rect 7395 15705 7405 15745
rect 7445 15705 7455 15745
rect 7495 15705 7505 15745
rect 7545 15705 7555 15745
rect 7595 15705 7605 15745
rect 7645 15705 7655 15745
rect 7695 15705 7705 15745
rect 7745 15705 7755 15745
rect 7795 15705 7805 15745
rect 7845 15705 7855 15745
rect 7895 15705 7905 15745
rect 7945 15705 7955 15745
rect 7995 15705 8005 15745
rect 8045 15705 8055 15745
rect 8095 15705 8105 15745
rect 8145 15705 8155 15745
rect 8195 15705 8205 15745
rect 8245 15705 8255 15745
rect 8295 15705 8305 15745
rect 8345 15705 8355 15745
rect 8395 15705 8405 15745
rect 8445 15705 8455 15745
rect 8495 15705 8505 15745
rect 8545 15705 8555 15745
rect 8595 15705 8605 15745
rect 8645 15705 8655 15745
rect 8695 15705 8705 15745
rect 8745 15705 8755 15745
rect 8795 15705 8805 15745
rect 8845 15705 8855 15745
rect 8895 15705 8905 15745
rect 8945 15705 8955 15745
rect 8995 15705 9005 15745
rect 9045 15705 9055 15745
rect 9095 15705 9105 15745
rect 9145 15705 9155 15745
rect 9195 15705 9205 15745
rect 9245 15705 9255 15745
rect 9295 15705 9305 15745
rect 9345 15705 9355 15745
rect 9395 15705 9405 15745
rect 9445 15705 9455 15745
rect 9495 15705 9505 15745
rect 9545 15705 9555 15745
rect 9595 15705 9605 15745
rect 9645 15705 9655 15745
rect 9695 15705 9705 15745
rect 9745 15705 9755 15745
rect 9795 15705 9805 15745
rect 9845 15705 9855 15745
rect 9895 15705 9905 15745
rect 9945 15705 9955 15745
rect 9995 15705 10005 15745
rect 10045 15705 10055 15745
rect 10095 15705 10105 15745
rect 10145 15705 10155 15745
rect 10195 15705 10205 15745
rect 10245 15705 10255 15745
rect 10295 15705 10305 15745
rect 10345 15705 10355 15745
rect 10395 15705 10405 15745
rect 10445 15705 10455 15745
rect 10495 15705 10505 15745
rect 10545 15705 10555 15745
rect 10595 15705 10605 15745
rect 10645 15705 10655 15745
rect 10695 15705 10705 15745
rect 10745 15705 10755 15745
rect 10795 15705 10805 15745
rect 10845 15705 10855 15745
rect 10895 15705 10905 15745
rect 10945 15705 10955 15745
rect 10995 15705 11005 15745
rect 11045 15705 11055 15745
rect 11095 15705 11105 15745
rect 11145 15705 11155 15745
rect 11195 15705 11205 15745
rect 11245 15705 11255 15745
rect 11295 15705 11305 15745
rect 11345 15705 11355 15745
rect 11395 15705 11405 15745
rect 11445 15705 11455 15745
rect 11495 15705 11505 15745
rect 11545 15705 11555 15745
rect 11595 15705 11605 15745
rect 11645 15705 11655 15745
rect 11695 15705 11705 15745
rect 11745 15705 11755 15745
rect 11795 15705 11805 15745
rect 11845 15705 11855 15745
rect 11895 15705 11905 15745
rect 11945 15705 11955 15745
rect 11995 15705 12005 15745
rect 12045 15705 12055 15745
rect 12095 15705 12105 15745
rect 12145 15705 12155 15745
rect 12195 15705 12205 15745
rect 12245 15705 12255 15745
rect 12295 15705 12305 15745
rect 12345 15705 12355 15745
rect 12395 15705 12405 15745
rect 12445 15705 12455 15745
rect 12495 15705 12505 15745
rect 12545 15705 12555 15745
rect 12595 15705 12605 15745
rect 12645 15705 12655 15745
rect 12695 15705 12705 15745
rect 12745 15705 12755 15745
rect 12795 15705 12805 15745
rect 12845 15705 12855 15745
rect 12895 15705 12905 15745
rect 12945 15705 12955 15745
rect 12995 15705 13005 15745
rect 13045 15705 13055 15745
rect 13095 15705 13105 15745
rect 13145 15705 13155 15745
rect 13195 15705 13205 15745
rect 13245 15705 13255 15745
rect 13295 15705 13305 15745
rect 13345 15705 13355 15745
rect 13395 15705 13405 15745
rect 13445 15705 13455 15745
rect 13495 15705 13505 15745
rect 13545 15705 13555 15745
rect 13595 15705 13605 15745
rect 13645 15705 13655 15745
rect 13695 15705 13705 15745
rect 13745 15705 13755 15745
rect 13795 15705 13805 15745
rect 13845 15705 13855 15745
rect 13895 15705 13905 15745
rect 13945 15705 13955 15745
rect 13995 15705 14005 15745
rect 14045 15705 14055 15745
rect 14095 15705 14105 15745
rect 14145 15705 14155 15745
rect 14195 15705 14205 15745
rect 14245 15705 14255 15745
rect 14295 15705 14305 15745
rect 14345 15705 14355 15745
rect 14395 15705 14405 15745
rect 14445 15705 14455 15745
rect 14495 15705 14505 15745
rect 14545 15705 14555 15745
rect 14595 15705 14605 15745
rect 14645 15705 14655 15745
rect 14695 15705 14705 15745
rect 14745 15705 14755 15745
rect 14795 15705 14805 15745
rect 14845 15705 14855 15745
rect 14895 15705 14905 15745
rect 14945 15705 14955 15745
rect 14995 15705 15005 15745
rect 15045 15705 15055 15745
rect 15095 15705 15105 15745
rect 15145 15705 15155 15745
rect 15195 15705 15205 15745
rect 15245 15705 15255 15745
rect 15295 15705 15305 15745
rect 15345 15705 15355 15745
rect 15395 15705 15405 15745
rect 15445 15705 15455 15745
rect 15495 15705 15505 15745
rect 15545 15705 15555 15745
rect 15595 15705 15605 15745
rect 15645 15705 15655 15745
rect 15695 15705 15705 15745
rect 15745 15705 15755 15745
rect 15795 15705 15805 15745
rect 15845 15705 15855 15745
rect 15895 15705 15905 15745
rect 15945 15705 15955 15745
rect 15995 15705 16005 15745
rect 16045 15705 16055 15745
rect 16095 15705 16105 15745
rect 16145 15705 16155 15745
rect 16195 15705 16205 15745
rect 16245 15705 16255 15745
rect 16295 15705 16305 15745
rect 16345 15705 16355 15745
rect 16395 15705 16405 15745
rect 16445 15705 16455 15745
rect 16495 15705 16505 15745
rect 16545 15705 16555 15745
rect 16595 15705 16605 15745
rect 16645 15705 16655 15745
rect 16695 15705 16705 15745
rect 16745 15705 16755 15745
rect 16795 15705 16805 15745
rect 16845 15705 16855 15745
rect 16895 15705 16905 15745
rect 16945 15705 16955 15745
rect 16995 15705 17005 15745
rect 17045 15705 17055 15745
rect 17095 15705 17105 15745
rect 17145 15705 17155 15745
rect 17195 15705 17205 15745
rect 17245 15705 17255 15745
rect 17295 15705 17305 15745
rect 17345 15705 17355 15745
rect 17395 15705 17405 15745
rect 17445 15705 17455 15745
rect 17495 15705 17505 15745
rect 17545 15705 17555 15745
rect 17595 15705 17605 15745
rect 17645 15705 17655 15745
rect 17695 15705 17705 15745
rect 17745 15705 17755 15745
rect 17795 15705 17805 15745
rect 17845 15705 17855 15745
rect 17895 15705 17905 15745
rect 17945 15705 17955 15745
rect 17995 15705 18005 15745
rect 18045 15705 18055 15745
rect 18095 15705 18105 15745
rect 18145 15705 18155 15745
rect 18195 15705 18205 15745
rect 18245 15705 18255 15745
rect 18295 15705 18305 15745
rect 18345 15705 18355 15745
rect 18395 15705 18405 15745
rect 18445 15705 18455 15745
rect 18495 15705 18505 15745
rect 18545 15705 18555 15745
rect 18595 15705 18605 15745
rect 18645 15705 18655 15745
rect 18695 15705 18705 15745
rect 18745 15705 18755 15745
rect 18795 15705 18805 15745
rect 18845 15705 18855 15745
rect 18895 15705 18905 15745
rect 18945 15705 18955 15745
rect 18995 15705 19005 15745
rect 19045 15705 19055 15745
rect 19095 15705 19105 15745
rect 19145 15705 19155 15745
rect 19195 15705 19205 15745
rect 19245 15705 19255 15745
rect 19295 15705 19305 15745
rect 19345 15705 19355 15745
rect 19395 15705 19405 15745
rect 19445 15705 19455 15745
rect 19495 15705 19505 15745
rect 19545 15705 19555 15745
rect 19595 15705 19605 15745
rect 19645 15705 19655 15745
rect 19695 15705 19705 15745
rect 19745 15705 19755 15745
rect 19795 15705 19805 15745
rect 19845 15705 19855 15745
rect 19895 15705 19905 15745
rect 19945 15705 19955 15745
rect 19995 15705 20005 15745
rect 20045 15705 20055 15745
rect 20095 15705 20105 15745
rect 20145 15705 20155 15745
rect 20195 15705 20205 15745
rect 20245 15705 20255 15745
rect 20295 15705 20305 15745
rect 20345 15705 20355 15745
rect 20395 15705 20405 15745
rect 20445 15705 20455 15745
rect 20495 15705 20505 15745
rect 20545 15705 20555 15745
rect 20595 15705 20605 15745
rect 20645 15705 20655 15745
rect 20695 15705 20705 15745
rect 20745 15705 20755 15745
rect 20795 15705 20805 15745
rect 20845 15705 20855 15745
rect 20895 15705 20905 15745
rect 20945 15705 20955 15745
rect 20995 15705 21005 15745
rect 21045 15705 21055 15745
rect 21095 15705 21105 15745
rect 21145 15705 21155 15745
rect 21195 15705 21205 15745
rect 21245 15705 21255 15745
rect 21295 15705 21305 15745
rect 21345 15705 21355 15745
rect 21395 15705 21405 15745
rect 21445 15705 21455 15745
rect 21495 15705 21505 15745
rect 21545 15705 21555 15745
rect 21595 15705 21605 15745
rect 21645 15705 21655 15745
rect 21695 15705 21705 15745
rect 21745 15705 21755 15745
rect 21795 15705 21805 15745
rect 21845 15705 21855 15745
rect 21895 15705 21905 15745
rect 21945 15705 21955 15745
rect 21995 15705 22005 15745
rect 22045 15705 22055 15745
rect 22095 15705 22105 15745
rect 22145 15705 22155 15745
rect 22195 15705 22205 15745
rect 22245 15705 22255 15745
rect 22295 15705 22305 15745
rect 22345 15705 22355 15745
rect 22395 15705 22405 15745
rect 22445 15705 22455 15745
rect 22495 15705 22505 15745
rect 22545 15705 22555 15745
rect 22595 15705 22605 15745
rect 22645 15705 22655 15745
rect 22695 15705 22705 15745
rect 22745 15705 22755 15745
rect 22795 15705 22805 15745
rect 22845 15705 22855 15745
rect 22895 15705 22905 15745
rect 22945 15705 22955 15745
rect 22995 15705 23005 15745
rect 23045 15705 23055 15745
rect 23095 15705 23105 15745
rect 23145 15705 23155 15745
rect 23195 15705 23205 15745
rect 23245 15705 23255 15745
rect 23295 15705 23305 15745
rect 23345 15705 23355 15745
rect 23395 15705 23405 15745
rect 23445 15705 23455 15745
rect 23495 15705 23505 15745
rect 23545 15705 23555 15745
rect 23595 15705 23605 15745
rect 23645 15705 23655 15745
rect 23695 15705 23705 15745
rect 23745 15705 23755 15745
rect 23795 15705 23805 15745
rect 23845 15705 23855 15745
rect 23895 15705 23905 15745
rect 23945 15705 23955 15745
rect 23995 15705 24005 15745
rect 24045 15705 24055 15745
rect 24095 15705 24105 15745
rect 24145 15705 24155 15745
rect 24195 15705 24205 15745
rect 24245 15705 24255 15745
rect 24295 15705 24305 15745
rect 24345 15705 24355 15745
rect 24395 15705 24405 15745
rect 24445 15705 24455 15745
rect 24495 15705 24505 15745
rect 24545 15705 24555 15745
rect 24595 15705 24605 15745
rect 24645 15705 24655 15745
rect 24695 15705 24705 15745
rect 24745 15705 24755 15745
rect 24795 15705 24805 15745
rect 24845 15705 24855 15745
rect 24895 15705 24905 15745
rect 24945 15705 24955 15745
rect 24995 15705 25005 15745
rect 25045 15705 25055 15745
rect 25095 15705 25105 15745
rect 25145 15705 25155 15745
rect 25195 15705 25205 15745
rect 25245 15705 25255 15745
rect 25295 15705 25305 15745
rect 25345 15705 25355 15745
rect 25395 15705 25405 15745
rect 25445 15705 25455 15745
rect 25495 15705 25505 15745
rect 25545 15705 25555 15745
rect 25595 15705 25605 15745
rect 25645 15705 25655 15745
rect 25695 15705 25705 15745
rect 25745 15705 25755 15745
rect 25795 15705 25805 15745
rect 25845 15705 25855 15745
rect 25895 15705 25905 15745
rect 25945 15705 25955 15745
rect 25995 15705 26005 15745
rect 26045 15705 26055 15745
rect 26095 15705 26105 15745
rect 26145 15705 26155 15745
rect 26195 15705 26205 15745
rect 26245 15705 26255 15745
rect 26295 15705 26305 15745
rect 26345 15705 26355 15745
rect 26395 15705 26405 15745
rect 26445 15705 26455 15745
rect 26495 15705 26505 15745
rect 26545 15705 26555 15745
rect 26595 15705 26605 15745
rect 26645 15705 26655 15745
rect 26695 15705 26705 15745
rect 26745 15705 26755 15745
rect 26795 15705 26805 15745
rect 26845 15705 26855 15745
rect 26895 15705 26905 15745
rect 26945 15705 26955 15745
rect 26995 15705 27005 15745
rect 27045 15705 27055 15745
rect 27095 15705 27105 15745
rect 27145 15705 27155 15745
rect 27195 15705 27205 15745
rect 27245 15705 27255 15745
rect 27295 15705 27305 15745
rect 27345 15705 27355 15745
rect 27395 15705 27405 15745
rect 27445 15705 27455 15745
rect 27495 15705 27505 15745
rect 27545 15705 27555 15745
rect 27595 15705 27605 15745
rect 27645 15705 27655 15745
rect 27695 15705 27705 15745
rect 27745 15705 27755 15745
rect 27795 15705 27805 15745
rect 27845 15705 27855 15745
rect 27895 15705 27905 15745
rect 27945 15705 27955 15745
rect 27995 15705 28005 15745
rect 28045 15705 28055 15745
rect 28095 15705 28105 15745
rect 28145 15705 28155 15745
rect 28195 15705 28205 15745
rect 28245 15705 28255 15745
rect 28295 15705 28305 15745
rect 28345 15705 28355 15745
rect 28395 15705 28405 15745
rect 28445 15705 28455 15745
rect 28495 15705 28505 15745
rect 28545 15705 28555 15745
rect 28595 15705 28605 15745
rect 28645 15705 28655 15745
rect 28695 15705 28705 15745
rect 28745 15705 28755 15745
rect 28795 15705 28805 15745
rect 28845 15705 28855 15745
rect 28895 15705 28905 15745
rect 28945 15705 28955 15745
rect 28995 15705 29005 15745
rect 29045 15705 29055 15745
rect 29095 15705 29105 15745
rect 29145 15705 29155 15745
rect 29195 15705 29205 15745
rect 29245 15705 29255 15745
rect 29295 15705 29305 15745
rect 29345 15705 29355 15745
rect 29395 15705 29405 15745
rect 29445 15705 29455 15745
rect 29495 15705 29505 15745
rect 29545 15705 29555 15745
rect 29595 15705 29605 15745
rect 29645 15705 29655 15745
rect 29695 15705 29705 15745
rect 29745 15705 29755 15745
rect 29795 15705 29805 15745
rect 29845 15705 29855 15745
rect 29895 15705 29905 15745
rect 29945 15705 29955 15745
rect 29995 15705 30005 15745
rect 30045 15705 30055 15745
rect 30095 15705 30105 15745
rect 30145 15705 30155 15745
rect 30195 15705 30205 15745
rect 30245 15705 30255 15745
rect 30295 15705 30305 15745
rect 30345 15705 30355 15745
rect 30395 15705 30405 15745
rect 30445 15705 30455 15745
rect 30495 15705 30505 15745
rect 30545 15705 30555 15745
rect 30595 15705 30605 15745
rect 30645 15705 30655 15745
rect 30695 15705 30705 15745
rect 30745 15705 30755 15745
rect 30795 15705 30805 15745
rect 30845 15705 30855 15745
rect 30895 15705 30905 15745
rect 30945 15705 30955 15745
rect 30995 15705 31005 15745
rect 31045 15705 31055 15745
rect 31095 15705 31105 15745
rect 31145 15705 31155 15745
rect 31195 15705 31205 15745
rect 31245 15705 31255 15745
rect 31295 15705 31305 15745
rect 31345 15705 31355 15745
rect 31395 15705 31405 15745
rect 31445 15705 31455 15745
rect 31495 15705 31505 15745
rect 31545 15705 31555 15745
rect 31595 15705 31605 15745
rect 31645 15705 31655 15745
rect 31695 15705 31705 15745
rect 31745 15705 31755 15745
rect 31795 15705 31805 15745
rect 31845 15705 31855 15745
rect 31895 15705 31905 15745
rect 31945 15705 31955 15745
rect 31995 15705 32005 15745
rect 32045 15705 32055 15745
rect 32095 15705 32105 15745
rect 32145 15705 32155 15745
rect 32195 15705 32205 15745
rect 32245 15705 32255 15745
rect 32295 15705 32305 15745
rect 32345 15705 32355 15745
rect 32395 15705 32405 15745
rect 32445 15705 32455 15745
rect 32495 15705 32505 15745
rect 32545 15705 32555 15745
rect 32595 15705 32605 15745
rect 32645 15705 32655 15745
rect 32695 15705 32705 15745
rect 32745 15705 32755 15745
rect 32795 15705 32805 15745
rect 32845 15705 32855 15745
rect 32895 15705 32905 15745
rect 32945 15705 32955 15745
rect 32995 15705 33005 15745
rect 33045 15705 33055 15745
rect 33095 15705 33105 15745
rect 33145 15705 33155 15745
rect 33195 15705 33205 15745
rect 33245 15705 33255 15745
rect 33295 15705 33305 15745
rect 33345 15705 33355 15745
rect 33395 15705 33405 15745
rect 33445 15705 33455 15745
rect 33495 15705 33505 15745
rect 33545 15705 33555 15745
rect 33595 15705 33605 15745
rect 33645 15705 33655 15745
rect 33695 15705 33705 15745
rect 33745 15705 33755 15745
rect 33795 15705 33805 15745
rect 33845 15705 33855 15745
rect 33895 15705 33905 15745
rect 33945 15705 33955 15745
rect 33995 15705 34005 15745
rect 34045 15705 34055 15745
rect 34095 15705 34105 15745
rect 34145 15705 34155 15745
rect 34195 15705 34205 15745
rect 34245 15705 34255 15745
rect 34295 15705 34305 15745
rect 34345 15705 34355 15745
rect 34395 15705 34405 15745
rect 34445 15705 34455 15745
rect 34495 15705 34505 15745
rect 34545 15705 34555 15745
rect 34595 15705 34605 15745
rect 34645 15705 34655 15745
rect 34695 15705 34705 15745
rect 34745 15705 34755 15745
rect 34795 15705 34805 15745
rect 34845 15705 34855 15745
rect 34895 15705 34905 15745
rect 34945 15705 34955 15745
rect 34995 15705 35005 15745
rect 35045 15705 35055 15745
rect 35095 15705 35105 15745
rect 35145 15705 35155 15745
rect 35195 15705 35205 15745
rect 35245 15705 35255 15745
rect 35295 15705 35305 15745
rect 35345 15705 35355 15745
rect 35395 15705 35405 15745
rect 35445 15705 35455 15745
rect 35495 15705 35505 15745
rect 35545 15705 35555 15745
rect 35595 15705 35605 15745
rect 35645 15705 35655 15745
rect 35695 15705 35705 15745
rect 35745 15705 35755 15745
rect 35795 15705 35805 15745
rect 35845 15705 35855 15745
rect 35895 15705 35905 15745
rect 35945 15705 35955 15745
rect 35995 15705 36005 15745
rect 36045 15705 36055 15745
rect 36095 15705 36105 15745
rect 36145 15705 36155 15745
rect 36195 15705 36205 15745
rect 36245 15705 36255 15745
rect 36295 15705 36305 15745
rect 36345 15705 36355 15745
rect 36395 15705 36405 15745
rect 36445 15705 36455 15745
rect 36495 15705 36505 15745
rect 36545 15705 36555 15745
rect 36595 15705 36605 15745
rect 36645 15705 36655 15745
rect 36695 15705 36705 15745
rect 36745 15705 36755 15745
rect 36795 15705 36805 15745
rect 36845 15705 36855 15745
rect 36895 15705 36905 15745
rect 36945 15705 36955 15745
rect 36995 15705 37005 15745
rect 37045 15705 37055 15745
rect 37095 15705 37105 15745
rect 37145 15705 37155 15745
rect 37195 15705 37205 15745
rect 37245 15705 37255 15745
rect 37295 15705 37305 15745
rect 37345 15705 37355 15745
rect 37395 15705 37405 15745
rect 37445 15705 37455 15745
rect 37495 15705 37505 15745
rect 37545 15705 37555 15745
rect 37595 15705 37605 15745
rect 37645 15705 37655 15745
rect 37695 15705 37705 15745
rect 37745 15705 37755 15745
rect 37795 15705 37805 15745
rect 37845 15705 37855 15745
rect 37895 15705 37905 15745
rect 37945 15705 37955 15745
rect 37995 15705 38005 15745
rect 38045 15705 38055 15745
rect 38095 15705 38105 15745
rect 38145 15705 38155 15745
rect 38195 15705 38205 15745
rect 38245 15705 38255 15745
rect 38295 15705 38305 15745
rect 38345 15705 38355 15745
rect 38395 15705 38405 15745
rect 38445 15705 38455 15745
rect 38495 15705 38505 15745
rect 38545 15705 38555 15745
rect 38595 15705 38605 15745
rect 38645 15705 38655 15745
rect 38695 15705 38705 15745
rect 38745 15705 38755 15745
rect 38795 15705 38805 15745
rect 38845 15705 38855 15745
rect 38895 15705 38905 15745
rect 38945 15705 38955 15745
rect 38995 15705 39005 15745
rect 39045 15705 39055 15745
rect 39095 15705 39105 15745
rect 39145 15705 39155 15745
rect 39195 15705 39205 15745
rect 39245 15705 39255 15745
rect 39295 15705 39305 15745
rect 39345 15705 39355 15745
rect 39395 15705 39405 15745
rect 39445 15705 39455 15745
rect 39495 15705 39505 15745
rect 39545 15705 39555 15745
rect 39595 15705 39605 15745
rect 39645 15705 39655 15745
rect 39695 15705 39705 15745
rect 39745 15705 39750 15745
rect 0 15700 39750 15705
rect -300 15345 -250 15700
rect -300 15305 -295 15345
rect -255 15305 -250 15345
rect -300 15295 -250 15305
rect -300 15255 -295 15295
rect -255 15255 -250 15295
rect -300 15245 -250 15255
rect -300 15205 -295 15245
rect -255 15205 -250 15245
rect -300 13645 -250 15205
rect -300 13605 -295 13645
rect -255 13605 -250 13645
rect -300 13595 -250 13605
rect -300 13555 -295 13595
rect -255 13555 -250 13595
rect -300 13545 -250 13555
rect -300 13505 -295 13545
rect -255 13505 -250 13545
rect -300 11945 -250 13505
rect -300 11905 -295 11945
rect -255 11905 -250 11945
rect -300 11895 -250 11905
rect -300 11855 -295 11895
rect -255 11855 -250 11895
rect -300 11845 -250 11855
rect -300 11805 -295 11845
rect -255 11805 -250 11845
rect -300 3845 -250 11805
rect -300 3805 -295 3845
rect -255 3805 -250 3845
rect -300 3795 -250 3805
rect -300 3755 -295 3795
rect -255 3755 -250 3795
rect -300 3745 -250 3755
rect -300 3705 -295 3745
rect -255 3705 -250 3745
rect -300 2145 -250 3705
rect -300 2105 -295 2145
rect -255 2105 -250 2145
rect -300 2095 -250 2105
rect -300 2055 -295 2095
rect -255 2055 -250 2095
rect -300 2045 -250 2055
rect -300 2005 -295 2045
rect -255 2005 -250 2045
rect -300 445 -250 2005
rect -300 405 -295 445
rect -255 405 -250 445
rect -300 395 -250 405
rect -300 355 -295 395
rect -255 355 -250 395
rect -300 345 -250 355
rect -300 305 -295 345
rect -255 305 -250 345
rect -300 0 -250 305
rect -200 14645 -150 15650
rect -200 14605 -195 14645
rect -155 14605 -150 14645
rect -200 1045 -150 14605
rect -200 1005 -195 1045
rect -155 1005 -150 1045
rect -200 0 -150 1005
rect -100 15345 -50 15700
rect -100 15305 -95 15345
rect -55 15305 -50 15345
rect -100 15295 -50 15305
rect -100 15255 -95 15295
rect -55 15255 -50 15295
rect -100 15245 -50 15255
rect -100 15205 -95 15245
rect -55 15205 -50 15245
rect -100 13645 -50 15205
rect -100 13605 -95 13645
rect -55 13605 -50 13645
rect -100 13595 -50 13605
rect -100 13555 -95 13595
rect -55 13555 -50 13595
rect -100 13545 -50 13555
rect -100 13505 -95 13545
rect -55 13505 -50 13545
rect -100 11945 -50 13505
rect -100 11905 -95 11945
rect -55 11905 -50 11945
rect -100 11895 -50 11905
rect -100 11855 -95 11895
rect -55 11855 -50 11895
rect -100 11845 -50 11855
rect -100 11805 -95 11845
rect -55 11805 -50 11845
rect -100 3845 -50 11805
rect -100 3805 -95 3845
rect -55 3805 -50 3845
rect -100 3795 -50 3805
rect -100 3755 -95 3795
rect -55 3755 -50 3795
rect -100 3745 -50 3755
rect -100 3705 -95 3745
rect -55 3705 -50 3745
rect -100 2145 -50 3705
rect -100 2105 -95 2145
rect -55 2105 -50 2145
rect -100 2095 -50 2105
rect -100 2055 -95 2095
rect -55 2055 -50 2095
rect -100 2045 -50 2055
rect -100 2005 -95 2045
rect -55 2005 -50 2045
rect -100 445 -50 2005
rect -100 405 -95 445
rect -55 405 -50 445
rect -100 395 -50 405
rect -100 355 -95 395
rect -55 355 -50 395
rect -100 345 -50 355
rect -100 305 -95 345
rect -55 305 -50 345
rect -100 0 -50 305
rect 39800 11345 39850 18150
rect 39800 11305 39805 11345
rect 39845 11305 39850 11345
rect 39800 10945 39850 11305
rect 39800 10905 39805 10945
rect 39845 10905 39850 10945
rect 39800 4745 39850 10905
rect 39800 4705 39805 4745
rect 39845 4705 39850 4745
rect 39800 4345 39850 4705
rect 39800 4305 39805 4345
rect 39845 4305 39850 4345
rect 39800 0 39850 4305
rect 39900 18145 40900 18150
rect 39900 18105 39905 18145
rect 39945 18105 39955 18145
rect 39995 18105 40005 18145
rect 40045 18105 40055 18145
rect 40095 18105 40105 18145
rect 40145 18105 40155 18145
rect 40195 18105 40205 18145
rect 40245 18105 40255 18145
rect 40295 18105 40305 18145
rect 40345 18105 40355 18145
rect 40395 18105 40405 18145
rect 40445 18105 40455 18145
rect 40495 18105 40505 18145
rect 40545 18105 40555 18145
rect 40595 18105 40605 18145
rect 40645 18105 40655 18145
rect 40695 18105 40705 18145
rect 40745 18105 40755 18145
rect 40795 18105 40805 18145
rect 40845 18105 40855 18145
rect 40895 18105 40900 18145
rect 39900 16945 40900 18105
rect 39900 16905 39905 16945
rect 39945 16905 39955 16945
rect 39995 16905 40005 16945
rect 40045 16905 40055 16945
rect 40095 16905 40105 16945
rect 40145 16905 40155 16945
rect 40195 16905 40205 16945
rect 40245 16905 40255 16945
rect 40295 16905 40305 16945
rect 40345 16905 40355 16945
rect 40395 16905 40405 16945
rect 40445 16905 40455 16945
rect 40495 16905 40505 16945
rect 40545 16905 40555 16945
rect 40595 16905 40605 16945
rect 40645 16905 40655 16945
rect 40695 16905 40705 16945
rect 40745 16905 40755 16945
rect 40795 16905 40805 16945
rect 40845 16905 40855 16945
rect 40895 16905 40900 16945
rect 39900 15745 40900 16905
rect 39900 15705 39905 15745
rect 39945 15705 39955 15745
rect 39995 15705 40005 15745
rect 40045 15705 40055 15745
rect 40095 15705 40105 15745
rect 40145 15705 40155 15745
rect 40195 15705 40205 15745
rect 40245 15705 40255 15745
rect 40295 15705 40305 15745
rect 40345 15705 40355 15745
rect 40395 15705 40405 15745
rect 40445 15705 40455 15745
rect 40495 15705 40505 15745
rect 40545 15705 40555 15745
rect 40595 15705 40605 15745
rect 40645 15705 40655 15745
rect 40695 15705 40705 15745
rect 40745 15705 40755 15745
rect 40795 15705 40805 15745
rect 40845 15705 40855 15745
rect 40895 15705 40900 15745
rect 39900 11245 40900 15705
rect 39900 11205 39905 11245
rect 39945 11205 39955 11245
rect 39995 11205 40005 11245
rect 40045 11205 40055 11245
rect 40095 11205 40105 11245
rect 40145 11205 40155 11245
rect 40195 11205 40205 11245
rect 40245 11205 40255 11245
rect 40295 11205 40305 11245
rect 40345 11205 40355 11245
rect 40395 11205 40405 11245
rect 40445 11205 40455 11245
rect 40495 11205 40505 11245
rect 40545 11205 40555 11245
rect 40595 11205 40605 11245
rect 40645 11205 40655 11245
rect 40695 11205 40705 11245
rect 40745 11205 40755 11245
rect 40795 11205 40805 11245
rect 40845 11205 40855 11245
rect 40895 11205 40900 11245
rect 39900 11195 40900 11205
rect 39900 11155 39905 11195
rect 39945 11155 39955 11195
rect 39995 11155 40005 11195
rect 40045 11155 40055 11195
rect 40095 11155 40105 11195
rect 40145 11155 40155 11195
rect 40195 11155 40205 11195
rect 40245 11155 40255 11195
rect 40295 11155 40305 11195
rect 40345 11155 40355 11195
rect 40395 11155 40405 11195
rect 40445 11155 40455 11195
rect 40495 11155 40505 11195
rect 40545 11155 40555 11195
rect 40595 11155 40605 11195
rect 40645 11155 40655 11195
rect 40695 11155 40705 11195
rect 40745 11155 40755 11195
rect 40795 11155 40805 11195
rect 40845 11155 40855 11195
rect 40895 11155 40900 11195
rect 39900 11145 40900 11155
rect 39900 11105 39905 11145
rect 39945 11105 39955 11145
rect 39995 11105 40005 11145
rect 40045 11105 40055 11145
rect 40095 11105 40105 11145
rect 40145 11105 40155 11145
rect 40195 11105 40205 11145
rect 40245 11105 40255 11145
rect 40295 11105 40305 11145
rect 40345 11105 40355 11145
rect 40395 11105 40405 11145
rect 40445 11105 40455 11145
rect 40495 11105 40505 11145
rect 40545 11105 40555 11145
rect 40595 11105 40605 11145
rect 40645 11105 40655 11145
rect 40695 11105 40705 11145
rect 40745 11105 40755 11145
rect 40795 11105 40805 11145
rect 40845 11105 40855 11145
rect 40895 11105 40900 11145
rect 39900 11095 40900 11105
rect 39900 11055 39905 11095
rect 39945 11055 39955 11095
rect 39995 11055 40005 11095
rect 40045 11055 40055 11095
rect 40095 11055 40105 11095
rect 40145 11055 40155 11095
rect 40195 11055 40205 11095
rect 40245 11055 40255 11095
rect 40295 11055 40305 11095
rect 40345 11055 40355 11095
rect 40395 11055 40405 11095
rect 40445 11055 40455 11095
rect 40495 11055 40505 11095
rect 40545 11055 40555 11095
rect 40595 11055 40605 11095
rect 40645 11055 40655 11095
rect 40695 11055 40705 11095
rect 40745 11055 40755 11095
rect 40795 11055 40805 11095
rect 40845 11055 40855 11095
rect 40895 11055 40900 11095
rect 39900 11045 40900 11055
rect 39900 11005 39905 11045
rect 39945 11005 39955 11045
rect 39995 11005 40005 11045
rect 40045 11005 40055 11045
rect 40095 11005 40105 11045
rect 40145 11005 40155 11045
rect 40195 11005 40205 11045
rect 40245 11005 40255 11045
rect 40295 11005 40305 11045
rect 40345 11005 40355 11045
rect 40395 11005 40405 11045
rect 40445 11005 40455 11045
rect 40495 11005 40505 11045
rect 40545 11005 40555 11045
rect 40595 11005 40605 11045
rect 40645 11005 40655 11045
rect 40695 11005 40705 11045
rect 40745 11005 40755 11045
rect 40795 11005 40805 11045
rect 40845 11005 40855 11045
rect 40895 11005 40900 11045
rect 39900 4645 40900 11005
rect 39900 4605 39905 4645
rect 39945 4605 39955 4645
rect 39995 4605 40005 4645
rect 40045 4605 40055 4645
rect 40095 4605 40105 4645
rect 40145 4605 40155 4645
rect 40195 4605 40205 4645
rect 40245 4605 40255 4645
rect 40295 4605 40305 4645
rect 40345 4605 40355 4645
rect 40395 4605 40405 4645
rect 40445 4605 40455 4645
rect 40495 4605 40505 4645
rect 40545 4605 40555 4645
rect 40595 4605 40605 4645
rect 40645 4605 40655 4645
rect 40695 4605 40705 4645
rect 40745 4605 40755 4645
rect 40795 4605 40805 4645
rect 40845 4605 40855 4645
rect 40895 4605 40900 4645
rect 39900 4595 40900 4605
rect 39900 4555 39905 4595
rect 39945 4555 39955 4595
rect 39995 4555 40005 4595
rect 40045 4555 40055 4595
rect 40095 4555 40105 4595
rect 40145 4555 40155 4595
rect 40195 4555 40205 4595
rect 40245 4555 40255 4595
rect 40295 4555 40305 4595
rect 40345 4555 40355 4595
rect 40395 4555 40405 4595
rect 40445 4555 40455 4595
rect 40495 4555 40505 4595
rect 40545 4555 40555 4595
rect 40595 4555 40605 4595
rect 40645 4555 40655 4595
rect 40695 4555 40705 4595
rect 40745 4555 40755 4595
rect 40795 4555 40805 4595
rect 40845 4555 40855 4595
rect 40895 4555 40900 4595
rect 39900 4545 40900 4555
rect 39900 4505 39905 4545
rect 39945 4505 39955 4545
rect 39995 4505 40005 4545
rect 40045 4505 40055 4545
rect 40095 4505 40105 4545
rect 40145 4505 40155 4545
rect 40195 4505 40205 4545
rect 40245 4505 40255 4545
rect 40295 4505 40305 4545
rect 40345 4505 40355 4545
rect 40395 4505 40405 4545
rect 40445 4505 40455 4545
rect 40495 4505 40505 4545
rect 40545 4505 40555 4545
rect 40595 4505 40605 4545
rect 40645 4505 40655 4545
rect 40695 4505 40705 4545
rect 40745 4505 40755 4545
rect 40795 4505 40805 4545
rect 40845 4505 40855 4545
rect 40895 4505 40900 4545
rect 39900 4495 40900 4505
rect 39900 4455 39905 4495
rect 39945 4455 39955 4495
rect 39995 4455 40005 4495
rect 40045 4455 40055 4495
rect 40095 4455 40105 4495
rect 40145 4455 40155 4495
rect 40195 4455 40205 4495
rect 40245 4455 40255 4495
rect 40295 4455 40305 4495
rect 40345 4455 40355 4495
rect 40395 4455 40405 4495
rect 40445 4455 40455 4495
rect 40495 4455 40505 4495
rect 40545 4455 40555 4495
rect 40595 4455 40605 4495
rect 40645 4455 40655 4495
rect 40695 4455 40705 4495
rect 40745 4455 40755 4495
rect 40795 4455 40805 4495
rect 40845 4455 40855 4495
rect 40895 4455 40900 4495
rect 39900 4445 40900 4455
rect 39900 4405 39905 4445
rect 39945 4405 39955 4445
rect 39995 4405 40005 4445
rect 40045 4405 40055 4445
rect 40095 4405 40105 4445
rect 40145 4405 40155 4445
rect 40195 4405 40205 4445
rect 40245 4405 40255 4445
rect 40295 4405 40305 4445
rect 40345 4405 40355 4445
rect 40395 4405 40405 4445
rect 40445 4405 40455 4445
rect 40495 4405 40505 4445
rect 40545 4405 40555 4445
rect 40595 4405 40605 4445
rect 40645 4405 40655 4445
rect 40695 4405 40705 4445
rect 40745 4405 40755 4445
rect 40795 4405 40805 4445
rect 40845 4405 40855 4445
rect 40895 4405 40900 4445
rect 39900 0 40900 4405
<< rmetal4 >>
rect -1300 18050 -1250 18100
use lpopamp_slice  slice0
timestamp 1713022628
transform -1 0 38750 0 -1 13550
box -1000 -2100 38750 5750
use lpopamp_slice  slice1
timestamp 1713022628
transform 1 0 1000 0 1 2100
box -1000 -2100 38750 5750
<< labels >>
rlabel metal3 -50 1000 0 1050 0 xn
rlabel metal3 -50 1400 0 1450 0 ynm
rlabel metal3 -50 1600 0 1650 0 ynp
rlabel metal3 -50 2500 0 2550 0 znm
rlabel metal3 -50 2700 0 2750 0 znp
rlabel metal3 -50 3100 0 3150 0 bna
rlabel metal3 -50 3200 0 3250 0 bnb
rlabel metal3 -50 5400 0 5450 0 bpb
rlabel metal3 -50 5500 0 5550 0 bpa
rlabel metal3 -50 5900 0 5950 0 zpp
rlabel metal3 -50 6100 0 6150 0 zpm
rlabel metal3 -50 6800 0 6850 0 ypm
rlabel metal3 -50 7200 0 7250 0 xp
rlabel metal3 -50 6600 0 6650 0 ypp
rlabel locali 0 0 50 50 0 vsub
port 9 nsew
rlabel metal4 -3400 18100 -3350 18150 0 im
port 1 nsew
rlabel metal4 -3200 18100 -3150 18150 0 ip
port 2 nsew
rlabel metal4 39900 18100 40900 18150 0 o
port 3 nsew
rlabel metal4 -1300 18100 -1250 18150 0 ib
port 4 nsew
rlabel metal4 -1400 18100 -1350 18150 0 en
port 5 nsew
rlabel metal4 -1500 18100 -1450 18150 0 enb
port 6 nsew
rlabel metal4 -3000 18100 -1650 18150 0 avdd
port 7 nsew
rlabel metal4 -1200 18100 -50 18150 0 avss
port 8 nsew
<< end >>
